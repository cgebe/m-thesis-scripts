MUNTLIG FRÅGA H-0108/09
till frågestunden under sammanträdesperioden i mars I 2009
i enlighet med artikel 109 i arbetsordningen
från
Konstantinos Droutsas
till rådet
Angående: Krav på omedelbart frigivande av fem kubanska fångar i Förenta staterna
Det har nu gått mer än tio år sedan de fem kubanska patrioterna Gerardo Hernández, Antonio Guerrero, Ramón Labañino, Fernando González och René González greps på falska och ogrundade anklagelser.
Ett nytt internationellt initiativ är på gång för att omedelbart få de fem fångarna fria, och ett krav om detta har hittills undertecknats av mer än 500 framstående konstnärer och intellektuella från hela världen.
Fördömer rådet det fortsatta, olagliga kvarhållandet av de fem kubanerna?
Hur ställer sig rådet till appellerna från nationella parlament och från internationella och nationella organisationer och personligheter om ett omedelbart frigivande av de fem fängslade kubanska patrioterna?
MUNTLIG FRÅGA H-0287/09
till frågestunden under sammanträdesperioden i september 2009
i enlighet med artikel 116 i arbetsordningen
från
Athanasios Pafilis
till rådet
Angående: Kriminalisering av kommunistisk ideologi i Litauen
Den 9 juni antog Litauens parlament ändringar till strafflagen som innebär att det blir brottsligt – med straff på upp till tre års fängelse – att sprida propaganda om och förneka eller rättfärdiga kommunismens och fascismens folkmord eller att offentligt förtala medlemmar i Litauens frihetsrörelse som kämpade mot den sovjetiska ockupationen mellan 1944 och 1953.
Dessa bestämmelser är ett försök att med straffrättsliga åtgärder förfalska historien och jämställa kommunismen med fascismen.
Vad anser rådet om återupprättandet av fascismen och nazismen – i synnerhet genom hot om straffrättsliga åtgärder mot oliktänkande – och om förbudet mot yttrandefrihet och kriminaliseringen av kommunistisk ideologi i ett flertal EU-medlemsstater, särskilt i Baltikum, där kommunistpartiet är förbjudet och där dess medlemmar och andra antifascistiska demokrater förföljs?
MUNTLIG FRÅGA H-0321/09
till frågestunden under sammanträdesperioden i oktober 2009
i enlighet med artikel 116 i arbetsordningen
från
Maria Badia i Cutchet
till kommissionen
Angående: Utbildning inom den nya europeiska politiska strategin
I samband med den aktuella ekonomiska recesionen har man på flera håll efterlyst en ny europeisk strategi för sysselsättning och en hållbar och smart tillväxt.
Flera rekommendationer har gjorts på vitt skilda områden, men det finns inga indikationer om detta på utbildningsområdet, och det verkar inte heller ha tagits några konkreta initiativ från kommissionens eller medlemsstaternas sida.
MUNTLIG FRÅGA H-0369/09
till frågestunden under sammanträdesperioden i november 2009
i enlighet med artikel 116 i arbetsordningen
från
Chris Davies
till rådet
Angående: Associeringsavtalet mellan EU och Israel
Vilka åtgärder har rådet vidtagit för att trygga respekten för människorättsklausulerna i associeringsavtalet mellan EU och Israel?
MUNTLIG FRÅGA H-0392/09
till frågestunden under sammanträdesperioden i november 2009
i enlighet med artikel 116 i arbetsordningen
från
Justas Vincas Paleckis
till rådet
Angående: Ratificeringen av energistadgan
Ryssland undertecknade 1994 tillsammans med 50 andra länder fördraget om energistadgan och tillhörande dokument, men regeringen i Moskva har ännu inte ratificerat stadgan.
I augusti vägrade Ryssland officiellt att ratificera fördraget och dess protokoll om energieffektivitet och de därtill hörande miljöaspekterna.
Inte heller Vitryssland eller Norge har ratificerat energistadgan.
Sedan år 2000 försöker EU förgäves förmå Ryssland att ratificera stadgan samt att göra de nödvändiga investeringarna i utvecklingen av energiteknik, avmonopolisera energidistributionen och liberalisera energimarknadsrelaterade investeringar.
På EU-nivå har man på nytt bekräftat energistadgefördragets betydelse, liksom det faktum att alla länder som undertecknat det måste uppfylla sina förpliktelser.
Vilka ytterligare åtgärder bör man enligt rådets uppfattning vidta för att se till att dessa bestämmelser omsätts i praktiken?
MUNTLIG FRÅGA H-0457/09
till frågestunden under sammanträdesperioden i december 2009
i enlighet med artikel 116 i arbetsordningen
från
Kathleen Van Brempt
till kommissionen
Angående: Billiga leksakers säkerhet
En ny undersökning som har genomförts av kvalitetskontrollorganet TÜV visar att två av tre undersökta leksaker inte uppfyller dagens kvalitetskrav.
En tredjedel av dem innehåller till och med förbjudna mjukgörare (ftalater).
Eftersom testet var specifikt inriktat på billiga leksaker finns det även en viktig social dimension på detta problem.
Är kommissionen väl insatt i problemet?
Hur tänker kommissionen se till att de hårdare kraven i det nya leksaksdirektivet följs, när man uppenbarligen inte ens kan åstadkomma en efterlevnad av det tidigare direktivet?
Vilka åtgärder kommer kommissionen att vidta för att alla barn ska kunna växa upp med säkra leksaker?
MUNTLIG FRÅGA H-0008/10
till frågestunden under sammanträdesperioden i februari 2010
i enlighet med artikel 116 i arbetsordningen
från
Zigmantas Balčytis
till rådet
Angående: En gemensam inre energimarknad
Spanien, Belgien och Ungern, ordförandeskapstrion, säger i sin överenskommelse och långsiktiga strategi att en av de politiska prioriteringarna kommer att vara att skapa en gemensam inre energimarknad.
Eftersom projekten i fråga är mellanstatliga är ett lyckosamt genomförande inte bara beroende av att tillräckliga ekonomiska medel ställs till förfogande, utan också av den politiska viljan och intentionen hos de medlemsstater som deltar i projekten.
Gemenskapen har lovat att tala med en röst i samband med att man skapar en inre energimarknad.
MUNTLIG FRÅGA H-0046/10
till frågestunden under sammanträdesperioden i februari 2010
i enlighet med artikel 116 i arbetsordningen
från
Laima Liucija Andrikienė
till kommissionen
Angående: "Bananavtalets" konsekvenser för EU:s inhemska bananproducenter
EU ingick nyligen ett historiskt avtal inom ramen för Världshandelsorganisationen (WTO) med länderna i Latinamerika om lägre tullavgifter för import av bananer från denna region.
Detta historiska avtal kommer emellertid att få negativa konsekvenser för EU:s egna bananproducenter, som kommer att utsättas för hård konkurrens från de latinamerikanska bananproducenterna.
Tänker kommissionen ta fram mekanismer för att skydda de europeiska bananproducenterna i områden som till exempel Kanarieöarna eller Madeira?
MUNTLIG FRÅGA H-0202/10
till frågestunden under sammanträdesperioden i maj 2010
i enlighet med artikel 116 i arbetsordningen
från
Jean-Luc Bennahmias
till kommissionen
Angående: Ett europeiskt organ för kontroll av idrottsverksamhet
Under denna period av året då transferfönstret öppnas väcks många frågor om bristen på insyn i dessa spelarövergångar, bland annat i spelaragenternas ersättning.
Anser kommissionen att det är lämpligt att EU föreslår att det inrättas ett oberoende europeiskt organ för kontroll av denna verksamhet, grundat på den modell som används inom den franska organisationen Direction Nationale du Contrôle de Gestion (som har till uppgift att kontrollera professionella franska fotbollsklubbars konton) eller inom World Anti-Doping Agency (ett internationellt samarbetsorgan för bekämpning av dopning inom idrotten)?
Stödjer kommissionen inrättandet av ett organ som även är öppet för Europarådets medlemsstater och som skulle ha till uppgift att kontrollera den finansiella öppenheten i syfte att förhindra avvikelser och orättvisa villkor som leder till en snedvriden konkurrens mellan klubbarna?
Fråga till frågestunden H-0311/2010
till kommissionen
Sammanträdesperiod: juli 2010
Artikel 116 i arbetsordningen
Marian Harkin
(ALDE) Angående: Handelsförhandlingar
Kan kommissionen mot bakgrund av att så många som nio medlemsstater redan har uttryckt oro över återupptagandet av Mercosur-förhandlingarna klargöra när dessa förhandlingar kommer att inledas?
Fråga till frågestunden H-0435/2010
till kommissionen
Sammanträdesperiod: september II 2010
Artikel 116 i arbetsordningen
Baroness
Sarah Ludford
(ALDE) Angående: Diabetesforskning
Diabetes är en allvarlig kronisk sjukdom som drabbar mer än 30 miljoner personer i EU:s medlemsstater.
Det är alarmerande att sjukdomen ökar i alla åldersgrupper, och särskilt tragiskt bland ungdomar.
En intensiv och samordnad forskning krävs för att stävja denna epidemi samt finna ett botemedel och effektiva metoder för att förebygga den.
Kan kommissionen tala om hur GD Forskning ämnar se till att EU intar en framträdande roll i den globala diabetesforskningen?
Vilka åtgärder ämnar kommissionen mer specifikt vidta för att möjliggöra bättre samordning och kontinuerlig finansiering för diabetesforskningen i enlighet med den strategi som skisseras i det nyligen avslutade FP7 DIAMAP-projektet?
Fråga till frågestunden H-0478/2010
till kommissionen
Sammanträdesperiod: oktober 2010
Artikel 116 i arbetsordningen
Andrew Henry William Brons
(NI) Angående: Malis president
Jag skulle vilja veta hur kommissionen ser på det tal som Malis president höll inför Europaparlamentet förra veckan.
Presidenten klagade över att Mali förlorar kvalificerad arbetskraft till den industrialiserade delen av världen.
Han berättade att nästan 35 procent av Malis akademiker arbetar utomlands och att en hög men inte närmare angiven andel personer som är verksamma inom sjukvården arbetar i andra länder.
Anser kommissionen att det är moraliskt försvarbart att länder i den industrialiserade delen av världen lockar till sig sjukvårdspersonal från länder i tredje världen, som dessa länder har finansierat utbildningen för med mycket begränsade medel?
Fråga till frågestunden H-0506/2010
till rådet
Sammanträdesperiod: oktober 2010
Artikel 116 i arbetsordningen
Laima Liucija Andrikienė
(PPE) Angående: Om EU:s representation i FN och andra internationella organ
Vad har rådet för strategi för att åstadkomma att Europeiska unionens nyligen utsedda höga företrädare som Europeiska rådets ordförande, Herman Van Rompuy, och den höga representanten för utrikes frågor och säkerhetspolitik, Catherine Ashton, kan tala inför FN:s generalförsamling på EU:s vägnar?
Efter att Lissabonfördraget trätt i kraft bör det vara Europeiska rådets ordförande, inte företrädare för det land som leder Europeiska rådets roterande ordförandeskap, som företräder EU på stats- och regeringschefsnivå i internationella sammanhang.
Vilka åtgärder bör vidtas för att genomföra dessa bestämmelser i Lissabonfördraget i internationella organ som FN?
Fråga till frågestunden H-0517/2010
till kommissionen
Sammanträdesperiod: november 2010
Artikel 116 i arbetsordningen
Georgios Koumoutsakos
(PPE) Angående: Tullunionen mellan EU och Turkiet och snedvridning av konkurrensen
Ett stort problem för handelsförbindelserna mellan EU och Turkiet är emellertid förfalskade produkter och bristfälligt immaterialrättsligt skydd, något som avsevärt snedvrider konkurrensen även på den europeiska marknaden.
Jag vill mot bakgrund av detta fråga följande: Vilka åtgärder tänker kommissionen vidta, och inom vilken tidsram, för att bekämpa denna företeelse, som är det mest karakteristiska uttrycket för det allmänna och hela tiden växande problemet med förfalskning och piratkopiering?
Fråga till frågestunden H-0624/2010
till rådet
Sammanträdesperiod: januari 2011
Artikel 116 i arbetsordningen
Vilija Blinkevičiūtė
(S&D) Angående: Skydd av barnoffer
Stockholmsprogrammet som antagits av rådet innehåller viktiga förebyggande åtgärder och åtgärder för skydd av offren och tillvaratagande av deras rättigheter i kampen mot människohandeln.
Skyddet av barn bör uppmärksammas särskilt och eftersom barnen är den svagaste länken i samhället måste enorma resurser satsas på detta område.
Barn säljs för att utföra tvångsarbete och för att delta i olaglig verksamhet.
Dessutom är de offer för den illegala organhandeln.
För att lättare kunna samordna EU-politiken när det gäller kampen mot människohandeln har rådet bestämt att utse en EU-samordnare för kampen mot människohandel.
Kan rådet tala om huruvida EU:s samordnare för kampen mot människohandel också kommer att vara ansvarig för kampen mot barnhandel?
Vilka konkreta åtgärder har den samordnare som utses för skydd av barnoffer tänkt att vidta?
Fråga till frågestunden H-0641/2010
till kommissionen
Sammanträdesperiod: januari 2011
Artikel 116 i arbetsordningen
Andreas Schwab
(PPE) Angående: EU-stöd till statliga kinesiska byggkoncerner
I Polen pågår just nu bygget av en sammanlagt 50 km lång delsträcka av motorvägen A2 mellan Warszawa och Lodz.
Bygget av denna delsträcka finansieras av EU-medel (EU:s strukturfonder) samt med hjälp av ett lån från EIB.
Uppdraget att bygga delsträckan gav det polska generaldirektoratet för nationella lands- och motorvägar till ett konsortium av statliga kinesiska byggkoncerner med namnet Covec.
I konkurrens med europeiska byggföretag låg anbudspriserna från den kinesiska anbudsgivaren mer än 50 procent under de upphandlande myndigheternas kostnadsuppskattning och en tredjedel under anbuden från anbudsgivaren med det näst lägsta anbudet.
Kinesiska företag fick delta i denna upphandling, trots att europeiska företag för det mesta inte får delta i upphandlingar i Kina.
Den kinesiska marknaden förblir stängd för så gott som all konkurrens inom byggindustrin.
Kommer kommissionen att vidta de rättsliga åtgärder som ges genom det avtal om offentlig upphandling som EU har tecknat med vissa tredjeländer?
Anser kommissionen att Kina, som inte har undertecknat avtalet om offentlig upphandling, borde behandlas som om man hade gjort det?
Vad gör kommissionen för att övertala Kina att ansluta sig till avtalet om offentlig upphandling?
Fråga till frågestunden H-000004/2011
till rådet
Sammanträdesperiod: januari 2011
Artikel 116 i arbetsordningen
Georgios Toussas
(GUE/NGL) Angående: Europeiska unionen godkänner ett erkännande av nazisterna
Den 21 december 2010 – för andra året i följd – antog FN:s generalförsamling en resolution som fördömer hjälteförklarandet av dem som deltog i de fascistiska legionerna från Waffen SS, allmänna förklaringar som rättfärdigar det nazistiska förgångna och nazismen, resandet av minnesmärken över nazister och deras kollaboratörer, skändandet och rivandet av hedersmonument över dem som kämpat mot fascismen och nazismen, olaglig uppgrävning av kroppar och flyttning av kvarlevor av dem som föll offer för fascisterna och deras brutalitet.
Resolutionen godkändes med en förkrossande majoritet av FN:s medlemsstater (129 medlemsstater för) medan Förenta staterna för andra gången i rad röstade mot och fick stöd av EU:s samtliga medlemsstater, vilka avstod från att rösta.
Ska EU-ländernas nedlagda röster uppfattas som ett godkännande eller ett tyst stöd för den glorifiering och det återupprättand av hedern för kollaboratörerna till de nazistiska krigsförbrytarna, något som öppet pågår i en rad av EU:s medlemsstater, samtidigt som förföljelserna av veteraner som deltog i den antifascistiska kampen tilltar, liksom av kommunister och kommunistiska partier?
Hänger EU:s vägran att fördöma denna vämjeliga förvrängning och förfalskning av vår historia samman med försöken att jämställa nazismen med kommunismen, försök som saknar historisk grund?
Fråga till frågestunden H-000022/2011/ändr.2
till kommissionen
Sammanträdesperiod: februari 2011
Artikel 116 i arbetsordningen
Nikolaos Chountis
(GUE/NGL) Angående: Tillväxtpolitik, Greklands samförståndsavtal och kommissionens skyldigheter
Greklands ekonomiska politik bestäms helt och hållet av ”samförståndsavtalet”, som undertecknats av den grekiska regeringen tillsammans med IMF och kommissionen.
Till och med samförståndsavtalets tillskyndare erkänner att det inte utvecklats någon plan för ekonomisk tillväxt vare sig inom ramen för avtalet eller parallellt med detta.
Detta faktum förvärrar de finansiella problemen samt orsakar stagnation och missmod på den inhemska marknaden.
Kan kommissionen åtminstone tänka sig att se över reglerna så att medlemsstatens andel i samfinansierade program sänks?
Överväger kommissionen en gemensam politik, exempelvis avseende turism och stöd till småföretag, eller sociala åtgärder, för att gynna medlemsstaterna och medborgarna i södra Europa, som är de som drabbats hårdast av krisen?
Fråga till frågestunden H-000056/2011
till rådet
Sammanträdesperiod: februari 2011
Artikel 116 i arbetsordningen
Marian Harkin
(ALDE) Angående: Räddningsfond för euroområdet
Vad anser det ungerska ordförandeskapet om möjliga reformer av räddningsfonden för euroområdet, särskilt när det gäller återköp av förmånstagarnas statspapper och lägre räntor på räddningslån?
Fråga till frågestunden H-000139/2011
till kommissionen
Sammanträdesperiod: april 2011
Artikel 116 i arbetsordningen
Sandrine Bélier
(Verts/ALE) Angående: EU:s strategi för biologisk mångfald
en obligatorisk miljökomponent när det gäller jordbruksföretag inom den första pelaren; komponenten skulle bestå av samlad god lantbrukspraxis, till exempel växtföljd och grön infrastruktur,
bestämmelser inom den första pelaren som är särskilt avpassade för lantbrukare på Natura 2000-områden och för driften av ekologiska jordbruk och betes- eller ängsmark som drivs på ett intensivt sätt,
en andra pelare som har tydlig målinriktning och som förses med tillräckliga resurser, bland annat effektiva, frivilliga och fleråriga planer för att stödja de bönder som går längre än att tillämpa god grundläggande praxis och som bidrar till förverkligandet av EU:s mål när det gäller klimatförändringar, biologisk mångfald och vatten?
Fråga till frågestunden H-000203/2011
till kommissionen
Sammanträdesperiod: juni 2011
Artikel 116 i arbetsordningen
Vilija Blinkevičiūtė
(S&D) Angående: Ändring av rådets förordning (EEG) nr 1612/68 om arbetskraftens fria rörlighet inom gemenskapen
Rådets förordning (EEG) nr 1612/68 om arbetskraftens fria rörlighet inom gemenskapen utgör referensram för den fria rörligheten för arbetstagare och har redan ändrats ett antal gånger.
Europaparlamentet utarbetar för närvarande ett betänkande om främjandet av den yrkesmässiga rörligheten i EU.
Kommissionens företrädare, som deltog vid ett sammanträde i utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor, förklarade den 19 april 2011 att kommissionen skulle ändra förordningen för att förbättra den.
När tror kommissionen att detta arbete kommer att inledas?
MUNTLIG FRÅGA MED DEBATT O-0057/04
i enlighet med artikel 108 i arbetsordningen
från
Philippe Morillon
för Fiskeriutskottet
till kommissionen
Angående: Fiskenäringen och bränslepriset
Priset på bränsle som används inom fiskenäringen har ökat mycket under de åtta senaste åren, med en ökning på 82 procent mellan 1996 och 2004 (från 0,17 euro/liter till 0,31 euro/liter).
Bränslepriset inverkar i hög grad på driftskostnaderna.
Driftsförlusterna för till exempel en trålare i kategorin 16–20 meter kan variera mellan -2,5 procent och -42,1 procent på grundval av siffrorna för 2003.
Under denna period har dieselbränslet uppnått sin högsta prisnivå flera gånger (2000, 2002, 2004).
Följderna av detta är desto påtagligare och leder till en krissituation, på grund av flera sammanfallande faktorer: bränslepriset, lägre priser och minskat stöd.
Detta var situationen sommaren 2004.
Den tidigare krisen under 1993–1994, som var ännu allvarligare till följd av det varaktiga kursfallet med anledning av rederiernas skuldsättning, hade en dominoeffekt: krisen ledde till uppläggning av fartyg (ibland de nyaste), skrotning av fartyg och omstrukturering av rederier, fiskeriverksamhetens kollapsande i flera hamnar, förlorade arbetsplatser inom fisket och följderna därav på ekonomin i närbelägna små regioner, minskat antal studerande i utbildningsanstalter inom sjöfartssektorn och minskat antal unga sjömän, misskrediterande av fiskaryrket, försvagade förvaltningsstrukturer och mindre finansiering till fiskesektorn.
Diskussionen inom EU, som nästan enbart riktar sig på en hållbar förvaltning av fiskeresurserna i syfte att bevara de kommande generationernas intressen, är så gott som frånvarande i krissituationer.
Fiskesektorn förhåller sig misstroende till EU-institutionerna, vilket kan konstaterats vid varje val (och vilket naturligtvis accentueras under svåra perioder).
Situationen är verkligen paradoxal eftersom hela fiskeregioner skulle ha försvunnit från kartan utan den gemensamma fiskeripolitiken.
Åtar sig kommissionen att vidta åtgärder till förmån för de mest utsatta regionerna?
Kommer kommissionen att lägga fram förslag för att göra det möjligt för europeiska fiskerifonden, eller någon annan metod, att ingripa vid krisperioder och sålunda trygga framtiden för regioner utan verkliga alternativ?
MUNTLIG FRÅGA MED DEBATT O-0063/04
i enlighet med artikel 108 i arbetsordningen
från
Ilda Figueiredo
och
Marco Rizzo
för GUE/NGL -gruppen
till kommissionen
Angående: Rådets politiska överenskommelse om förslaget till direktiv om patentbarhet för datorrelaterade uppfinningar
Förslaget till direktiv om patentbarhet för datorrelaterade uppfinningar svarar inte upp mot de ekonomiska, forskningsrelaterade och kulturella utmaningar som programvaruindustrin står inför, och heller inte behovet av att främja uppfinningar och teknisk utveckling eller de särskilda behov som finns i små och medelstora företag.
Detta förslag till direktiv syftar till att öppna möjligheten att ta patent på människors kunnande, vilket tjänar de multinationella programvaruföretagens intresse av marknadsdominans och vinstintresse.
Den 18 maj 2004 nådde rådet om konkurrensfrågor en politisk överenskommelse om förslaget till direktiv om patentbarhet för datorrelaterade uppfinningar som öppnar dörren för patent på programvara.
Denna politiska överenskommelse ingicks genom kvalificerad majoritet där tre länder avstod (Belgien, Österrike och Italien) och ett land röstade emot (Spanien).
Rådet har inte haft en formell omröstning om överenskommelsen sedan dess, vilket inte endast beror på det växande motståndet från rörelsen för fria datorprogram, programvaruföretag, programmerare, forskare, små och medelstora företag och vissa nationella parlament, utan också på att Nederländernas parlament har uppmanat landets regering att dra tillbaka sitt stöd för förslaget till direktiv, d.v.s. rösta mot den politiska överenskommelse som ingåtts.
Mot bakgrund av den breda oppositionen mot konsekvenserna av detta förslag till direktiv som kommer att skapa hinder mot uppfinningar och teknisk utveckling, undrar jag varför kommissionen inte drar tillbaka förslaget?
MUNTLIG FRÅGA MED DEBATT O-0001/05
i enlighet med artikel 108 i arbetsordningen
från
Graham Watson
för ALDE -gruppen
till rådet
Angående: Hälsovårdare som sitter häktade i Libyen
Fem bulgariska sjuksköterskor och en palestinsk läkare dömdes i maj 2004 till döden av en libysk domstol och sedan dess har de väntat på att deras ärenden skall prövas på nytt i högsta domstolen.
Dessa hälsovårdare har suttit häktade sedan 1999 och anklagas för att avsiktligt ha smittat 400 barn med HIV vid Al Fateh-sjukhuset i Benghazi.
Under den rättsliga processen har det förekommit förfarandemässiga brister och framförts anklagelser om tortyr, och internationella experter har fastställt att sjukhusinfektion är den troligaste smittorsaken.
Vad har EU gjort för att bidra till att finna en tillfredsställande lösning i detta ärende?
MUNTLIG FRÅGA MED DEBATT O-0002/05
i enlighet med artikel 108 i arbetsordningen
från Baroness
Sarah Ludford
och
Alexander Alvaro
för ALDE -gruppen
till kommissionen
Angående: Överföring av uppgifter om passagerare
2003 och 2004 bestred parlamentet vid flera tillfällen, även inför domstolen, de amerikanska myndigheternas systematiska tillgång av säkerhetsskäl till vissa PNR-uppgifter om luftfartspassagerare.
Därefter, i samband med antagandet av 2005 års budget, antog parlamentet ett ändringsförslag till budgetpost 06 02 04 02 (passagerarnas rättigheter) för att föra en del av anslagen till reserven i väntan på att ett system för överföring av vissa personuppgifter inrättas.
Kan kommissionen, med hänsyn till de befogenheter den har i enlighet med fördragen och till de ”åtaganden” som gjorts redogöra för följande:
I vilket skede befinner sig varje enskild punkt i ”åtagandena”?
Hur kan kommissionen och de nationella myndigheter som ansvarar för skyddet av personuppgifter (Grupp 29) kontrollera hur ”åtagandena” fungerar i verkligheten?
Hur stora mängder uppgifter har de amerikanska myndigheterna fått tillgång till, förekommer det effektiv filtrering av känsliga uppgifter (punkt 10 i ”åtagandena”) och framför allt om flygningar inom gemenskapen utesluts?
Hur många misstänkta terrorister eller personer som gjort sig skyldiga till allvarliga brott har kunnat upptäckas sedan överenskommelsen trädde ikraft?
Har de europeiska passagerarna informerats på ett korrekt sätt och har det inkommit protester mot insamlingen och tillrättaläggandet av dessa uppgifter?
Har personuppgifter om passagerare från EU överförts från Förenta staterna till tredje land, och i så fall i vilken omfattning?
Har nya förhandlingar inletts med Förenta staterna om det projekt som skall ersätta CAPPS II?
Varför har Europaparlamentet aldrig informerats om de förhandlingar som förs i denna fråga inom Internationella civila luftfartsorganisationen (ICAO)?
Vad anser kommissionens ordförande om de frågor som rör de grundläggande rättigheterna?
MUNTLIG FRÅGA MED DEBATT O-0057/05
i enlighet med artikel 108 i arbetsordningen
från
Glyn Ford
,
Caroline Lucas
,
Vittorio Agnoletto
,
Harlem Désir
,
Daniel Cohn-Bendit
,
Monica Frassoni
,
Luisa Morgantini
,
Pierre Jonckheer
,
Frithjof Schmidt
,
Claude Turmes
,
Joost Lagendijk
,
Hiltrud Breyer
,
Rebecca Harms
,
Marie-Hélène Aubert
,
Evelin Lichtenberger
,
Sepp Kusstatscher
,
Raül Romeva i Rueda
,
Roberto Musacchio
,
Kyriacos Triantaphyllides
,
Giusto Catania
,
Jacky Henin
,
Tobias Pflüger
,
Daniel Stroz
,
Erik Meijer
,
André Brie
,
Gabriele Zimmer
,
Umberto Guidoni
,
Helmuth Markov
,
Bairbre de Brún
,
Sylvia-Yvonne Kaufmann
,
Vladimír Remek
,
Mary McDonald
,
Helga Trüpel
,
David Hammerstein Mintz
,
Carl Schlyter
,
Johannes Voggenhuber
,
Alain Lipietz
,
Angelika Beer
,
Jean Lambert
och
Elisabeth Schroedter
till rådet
Angående: Rådets ståndpunkt till en skatt på valutatransaktioner (Tobinskatt)
Lagstiftning om en skatt på valutatransaktioner (Tobinskatt) har antagits i Frankrike och Belgien och övervägs för närvarande i Italien.
Mot bakgrund av den växande enigheten i parlament, regeringar och det civila samhället om de potentiella fördelarna med internationella skatter som Tobinskatten, kan rådet redogöra för sina synpunkter i frågan?
Kan rådet särskilt ge svar på de förslag om internationell beskattning som president Chirac gav i sitt tal till Världsekonomiskt forum i Davos tidigare i år?
Har rådet för avsikt att stödja lagstiftningsinitiativen i Frankrike och Belgien att införa en Tobinskatt när en sådan skatt har införts i samtliga medlemsstater genom att uppmana samtliga medlemsstater att anta liknande nationella lagar?
Anser rådet att en sådan skatt kan bidra till att skapa intäkter för samhällsnyttiga investeringar i miljö, utbildning och utveckling över hela världen, och som ett viktigt bidrag till att millenniemålen uppnås?
Anser rådet att en sådan skatt kan bidra till att minska valutaspekulationer och stabilisera finansiella marknader?
Kommer rådet att vidta konkreta åtgärder i detta hänseende?
MUNTLIG FRÅGA MED DEBATT O-0127/06
i enlighet med artikel 108 i arbetsordningen
från
Simon Busuttil
,
Milan Cabrnoch
,
Petr Duchoň
,
Hynek Fajmon
,
Miroslav Ouzký
,
Nina Škottová
,
Ivo Strejček
,
Oldřich Vlasák
,
Jan Zahradil
,
Jaroslav Zvěřina
,
Valdis Dombrovskis
,
Aldis Kušķis
,
Rihards Pīks
,
Laima Liucija Andrikienė
,
Vytautas Landsbergis
,
Konstantinos Hatzidakis
,
Etelka Barsi-Pataky
,
Zsolt László Becsey
,
Antonio De Blasio
,
Kinga Gál
,
Béla Glattfelder
,
András Gyürk
,
Lívia Járóka
,
Péter Olajos
,
Csaba Őry
,
Pál Schmitt
,
György Schöpflin
,
László Surján
,
József Szájer
,
Edit Bauer
,
Árpád Duka-Zólyomi
,
Milan Gaľa
,
Ján Hudacký
,
Miroslav Mikolášik
,
Zita Pleštinská
,
Anna Záborská
,
Tunne Kelam
,
David Casa
,
Jerzy Buzek
,
Zdzisław Kazimierz Chmielewski
,
Małgorzata Handzlik
,
Stanisław Jałowiecki
,
Filip Kaczmarek
,
Barbara Kudrycka
,
Jan Olbrycht
,
Jacek Protasiewicz
,
Jacek Emil Saryusz-Wolski
,
Czesław Adam Siekierski
,
Bogusław Sonik
,
Zbigniew Zaleski
,
Tadeusz Zwiefka
,
Panayiotis Demetriou
,
Ioannis Kasoulides
,
Yiannakis Matsis
och
Peter Šťastný
till kommissionen
Angående: Förenta staternas viseringskrav för EU-medborgare från 10 medlemsstater
Förenta staterna kräver fortfarande inresevisum av medborgarna i nio av de tio nya medlemsstaterna (Cypern, Tjeckien, Estland, Ungern, Lettland, Litauen, Malta, Polen och Slovakien) samt Grekland.
Detta är en situation av icke-ömsesidighet, vilket innebär att dessa länder ger Förenta staternas medborgare rätt att resa utan visum medan Förenta staterna inte erbjuder samma möjlighet.
Av större betydelse är det faktum att denna situation är diskriminerande genom att viseringskravet tillämpas på tio av tjugofem EU-länder, vilket leder till en omotiverad åtskillnad mellan EU-medborgare som kommer från olika EU-länder.
Medborgarna i de berörda EU-länderna förväntar sig med rätta att de skall behandlas jämlikt med medborgarna i de femton andra länderna.
Trots kommissionens ansträngningar har det enligt den senaste rapporten om vissa tredjeländers avvikelser från ömsesidighetsprincipen när det gäller undantag från viseringskravet - KOM(2006)0568 - inte skett några framsteg.
Kommissionen ombeds mot denna bakgrund besvara följande frågor:
Vilka åtgärder är kommissionen beredd att vidta i syfte att rätta till denna situation?
När väntar sig kommissionen att Förenta staternas viseringskrav för de tio berörda länderna upphävs?
MUNTLIG FRÅGA MED DEBATT O-0049/07
i enlighet med artikel 108 i arbetsordningen
från
Miroslav Ouzký
för utskottet för miljö, folkhälsa och livsmedelssäkerhet
till rådet
Angående: Mål inför konferensen i Madrid för parterna i konventionen för bekämpning av ökenspridning den 3-14 september 2007
Kan rådet redogöra för Europeiska unionens mål inför den förestående åttonde konferensen för parterna i FN:s konvention för bekämpning av ökenspridning (COP 8) som kommer att äga rum i Madrid, Spanien den 3–14 september 2007?
MUNTLIG FRÅGA MED DEBATT O-0056/07
i enlighet med artikel 108 i arbetsordningen
från
Erika Mann
,
Carlos Carnero González
,
Javier Moreno Sánchez
och
Emilio Menéndez del Valle
för PSE -gruppen,
Daniel Varela Suanzes-Carpegna
och
Małgorzata Handzlik
för PPE-DE -gruppen,
Ignasi Guardans Cambó
och
Gianluca Susta
för ALDE -gruppen,
Cristiana Muscardini
och
Eugenijus Maldeikis
för UEN -gruppen,
Caroline Lucas
för Verts/ALE -gruppen,
Jens Holm
och
Helmuth Markov
för GUE/NGL -gruppen
till kommissionen
Angående: Förhandlingar om ett interregionalt associeringsavtal med Mercosur och det nya bilaterala strategiska partnerskapet med Brasilien
Under toppmötet mellan EU och Brasilien den 4 juli 2007 påminde EU och Brasilien om att de fäste stor vikt vid att förbindelserna mellan EU och Mercosur stärks och förpliktade sig att ingå ett associeringsavtal mellan EU och Mercosur.
I sin resolution INI/2006/2035 om EU:s ekonomiska och kommersiella förbindelser med Mercosur underströk Europaparlamentet att ett associeringsavtal mellan EU och Mercosur bör betraktas som ett prioriterat strategiskt mål för EU:s yttre förbindelser.
Icke desto mindre har kommissionen offentliggjort sitt meddelande av den 30 maj 2007 om ett bilateralt strategiskt partnerskap med Brasilien vilket skickar signaler som strider mot de regionala prioriteringar som fastställts ovan.
Mot bakgrund av ovanstående:
Skulle kommissionen kunna redogöra för den senaste utvecklingen i Mercosurförhandlingarna?
Skulle kommissionen kunna förklara hur det bilaterala strategiska partnerskapet med Brasilien som presenterades i meddelandet av den 30 maj 2007 skall kunna genomföras utan att det underminerar det bilaterala tillvägagångssätt som bör vara hörnstenen i våra förbindelser med Latinamerika i allmänhet och med Mercosur i synnerhet?
Skulle kommissionen kunna fastslå att detta nya partnerskap inte kommer att skada den regionala balansen och inte kommer att vara till skada för EU:s handel och ekonomiska förbindelser med andra Latinamerikanska partner?
MUNTLIG FRÅGA MED DEBATT O-0067/07
i enlighet med artikel 108 i arbetsordningen
från
Luis Manuel Capoulas Santos
för PSE -gruppen
till kommissionen
Angående: Konsumentskydd och prishöjningar
De senaste konsumentprishöjningarna till följd av de ökade kostnaderna för jordbruksråvaror har tvingat kommissionen att vidta vissa åtgärder, som att slopa kravet på träda för spannmål, och att börja överväga nödlösningar för andra branscher, exempelvis mjölkindustrin, som drabbats av de stigande foderpriserna.
Förutom att slå mot de europeiska produktionssektorerna får denna situation även kraftiga och direkta följder för konsumenterna och de europeiska hushållens ekonomi.
Europaparlamentet välkomnar åtgärder som det slopade kravet på träda och kommissionsledamotens tillkännagivande i plenum i Strasbourg att denna åtgärd om nödvändigt ska förlängas med ett regleringsår, men uttrycker samtidigt sin oro över den nuvarande situationen med stigande priser som kräver nya nödlösningar och som EU-institutionerna borde gå på djupet med, inte bara i form av en ”hälsokontroll”.
Kan kommissionen ange vilka åtgärder den tänker vidta tillsammans med de berörda sektorerna för att få bukt med denna situation?
Tänker sig kommissionen några konkreta åtgärder för att skydda konsumenterna och trygga hushållens ekonomi?
Anser inte kommissionen att de olika formerna av prishöjningar förtjänar ett helhetsgrepp som går längre än konkreta åtgärder för varje enskilt fall (spannmål, mjölk osv.)?
MUNTLIG FRÅGA MED DEBATT O-0118/08
i enlighet med artikel 108 i arbetsordningen
från
Elly de Groen-Kouwenhoven
och
Monica Frassoni
för Verts/ALE -gruppen,
Jan Marinus Wiersma
för PSE -gruppen,
Viktória Mohácsi
,
Renate Weber
och
Baroness Sarah Ludford
för ALDE -gruppen,
Vittorio Agnoletto
,
Giusto Catania
och
Lívia Járóka
till rådet
Angående: Krav på en EU-strategi för romer
I oktober 2007 sände parlamentsledamöter ett förslag till EU:s ordförandeskap (Slovenien) om ett nytt sätt att behandla romska frågor på EU-nivå.
Där föreslog man bland annat att det årligen skulle anordnas en EU-konferens om romska frågor där man kunde diskutera olika idéer, underlätta utbyte om bästa praxis och information och samordna samarbetet på EU-nivå.
Majoriteten i Europaparlamentet stödde en resolution ( P6_TA(2008)0035 ) där man i januari 2008 krävde en EU-strategi för romer.
Förbinder sig det franska ordförandeskapet att kräva en EU-strategi vid nästa EU-toppmöte i december 2008?
MUNTLIG FRÅGA MED DEBATT O-0028/09
i enlighet med artikel 108 i arbetsordningen
från
Johannes Blokland
för utskottet för miljö, folkhälsa och livsmedelssäkerhet
till kommissionen
Angående: IMO-förhandlingar i maj 2009 om villkoren för att konventionen om trygg och miljöriktig fartygsåtervinning ska kunna träda i kraft
Vilka initiativ tar kommissionen för att det oacceptabla tillvägagångssättet med upphuggning av uttjänta fartyg direkt på stranden ska frångås, såsom det klart rekommenderats av 170 parter i Baselkonventionen?
Ämnar kommissionen verka för att den konvention, som gäller trygg och miljöriktig fartygsåtervinning och är avsedd att förhandlas fram vid en diplomatisk konferens i maj 2009 under överinseende av Internationella sjöfartsorganisationen (IMO), tidigt och verkningsfullt kommer att införlivas med gemenskapslagstiftningen?
Vilka initiativ ämnar kommissionen ta för att denna IMO-konvention inte kommer att sänka den nivå på skydd mot skadliga effekter av farligt avfall, vilken i dag erbjuds av förordning (EG) nr 1013/2006 om transport av avfall?
EUT L 190, 12.7.2006, s.
1.
MUNTLIG FRÅGA MED DEBATT O-0048/09
i enlighet med artikel 108 i arbetsordningen
från
Helmuth Markov
och
Erika Mann
för utskottet för internationell handel
till kommissionen
Angående: Inledande avtal om ekonomiskt partnerskap mellan Europeiska gemenskapen och dess medlemsstater, å ena sidan, och Elfenbenskusten, å andra sidan
Kan kommissionen uppdatera Europaparlamentet om när ett "fullständigt" avtal om ekonomiskt partnerskap med den västafrikanska regionen kan komma att ingås?
Väntar sig kommissionen att underteckna ett heltäckande avtal för att ytterligare främja ekonomisk tillväxt, utveckling och goda styrelseformer i Elfenbenskusten och i den västafrikanska regionen som helhet?
Har man i förhandlingarna tagit hänsyn till några specifika intressen när det gäller denna region och hur skulle detta "fullständiga" avtal om ekonomiskt partnerskap skilja sig från Cariforumavtalet?
Kommer kommissionen att lova att tillhandahålla adekvat administrativt och tekniskt bistånd till Elfenbenskusten, inbegripet till dess privata sektor, för att underlätta övergången för landets näringsliv efter att interimsavtalet om ekonomiskt partnerskap undertecknats?
Kommer kommissionen att som villkor för ett ingående av ett "fullständigt" avtal om ekonomiskt partnerskap kräva att det ska finnas en ansvarsskyldig och demokratiskt vald regering på plats i landet?
Kan kommissionen förklara hur man bedömer följande aspekter med avseende på avtalet om ekonomiskt partnerskap mellan EU och Elfenbenskusten:
i) Finns det ett behov av och/eller garantier för starkare regler för skydd av nyetablerade industrier?
ii) Kommer man vid förhandlingarna om immaterialrätten att se till att inte bara europeisk/internationell immaterialrätt skyddas utan också traditionell kunskap?
iii) Bör det utarbetas regler för offentlig upphandling utifrån Elfenbenskustens särskilda behov?
iv) Hur långt har man kommit med utarbetandet av villkor för ”arbetsvisum” för Elfenbenskustens medborgare?
Kommer de att täcka en period på 24 månader?
För vilka slags yrken kommer de att gälla?
Kan kommissionen stödja kravet att parlamentet ska höras innan beslut fattas om den provisoriska tillämpningen av internationella avtal, såsom avtalen om ekonomiskt partnerskap, när samtyckesförfarandet ska tillämpas för att nå politisk förståelse för detta förfarande?
Kan kommissionen förklara hur man kommer att bedöma den politiska situationen i Elfenbenskusten med avseende på antingen ett interimsavtal eller ett slutligt avtal om ekonomiskt partnerskap?
Den politiska situationen i Elfenbenskusten uppfyller inte demokratiska standarder.
Hur kommer denna bedömning att påverka de övriga 15 västafrikanska ländernas möjlighet att komma i åtnjutande av ett viktigt biregionalt handels- och utvecklingsavtal?
Kan kommissionen klargöra tidsramen för utvecklingsbistånd till Elfenbenskusten i samband med avtalet om ekonomiskt partnerskap?
MUNTLIG FRÅGA MED DEBATT O-0078/09
i enlighet med artikel 115 i arbetsordningen
från
Sonia Alfano
,
Jeanine Hennis-Plasschaert
,
Sophia in 't Veld
och Baroness
Sarah Ludford
för ALDE -gruppen
till kommissionen
Angående: Lagen om uppskov av brottmål i Italien
Den italienska lagen 124/08 (Lodo Alfano) om uppskov av brottmål mot höga statstjänstemän, som föreslagits av Berlusconis regering, godkändes den 22 juli 2008 av det italienska parlamentet och undertecknades av republikens president.
Enligt lagen ska brottmål mot republikens president, ordförandena för senaten och deputeradekammaren samt premiärministern skjutas upp under deras ämbetsperiod.
Uppskovet omfattar även brott som dessa personer begått utanför tjänsten, eller innan de tillsattes, till och med om de tagits på bar gärning.
Italien är det enda landet i EU som ger premiärministern tillfällig immunitet mot straffrättslig lagföring.
Mot bakgrund av detta bör nämnas att Berlusconi har ätit middag med två domare från konstitutionsdomstolen samt justitieministern, understatssekreteraren för ministeriernas presidium och ordföranden för senatens konstitutionsutskott.
Är kommissionen medveten om detta?
Anser kommissionen att den italienska lagen är förenlig med mänskliga rättigheter och grundläggande friheter, demokrati och rättsstatsprincipen, som garanteras i bland annat Europeiska stadgan om de grundläggande rättigheterna och artiklarna 6 och 7 i EU-fördraget, samt medborgarnas grundläggande rätt till likhet inför lagen?
Anser kommissionen att det är förenligt med europeiska och demokratiska principer att den verkställande makten offentligt och våldsamt ger sig på domarkåren och försöker påverka konstitutionsdomstolen bara några månader innan denna ska ta ställning i en sådan viktig fråga som berör premiärministerns direkta intressen?
Vilka konkreta åtgärder kommer kommissionen i detta hänseende att vidta för att se till att grundläggande rättigheter, demokrati och rättsstatsprincipen respekteras i enlighet med EU:s fördrag och den italienska konstitutionen?
MUNTLIG FRÅGA MED DEBATT O-0164/09
i enlighet med artikel 115 i arbetsordningen
från
Raül Romeva i Rueda
,
Heidi Hautala
,
Jean Lambert
,
Hélène Flautre
,
Franziska Keller
och
Jan Philipp Albrecht
för Verts/ALE -gruppen
till kommissionen
Angående: Dröjsmål i stängningen av Guantánamo
Den amerikanska regeringen har meddelat att Guantánamo-fängelset inte kommer att stängas den 22 januari 2010, trots att president Obama gav ett löfte om att så skulle ske när han tillträdde presidentämbetet exakt ett år tidigare.
Försöken att väcka åtal mot vissa av fångarna i Guantánamo och att finna en plats på amerikansk mark där de kan tas emot har hittills misslyckats, bland annat på grund av att kongressen motsatt sig att före detta fångar beträder amerikansk mark.
Cirka 245 personer hölls fångna i Guantánamo vid den tidpunkt då Barack Obama tillträdde presidentämbetet.
Sedan dess har endast cirka 30 män lämnat fängelset och 215 hålls fortsättningsvis fångna.
Enligt media är det möjligt att Barack Obama under de närmaste veckorna kungör en plan för stängning av Guantánamo, vilket skulle kunna medföra att upp till 90 misstänka terrorister förblir häktade ”i preventivt syfte” och på obestämd tid, eftersom bevisen mot dem erhållits genom tortyr eller på grund av att en offentlig rättegång eventuellt skulle kunna innebära att ett omfattande sekretessbelagt material blottställs.
Efter en förfrågan från den amerikanska regeringen har Bermuda och Palau, samt bland europeiska stater Frankrike, Portugal, Irland, Belgien, Förenade kungariket, Italien och Ungern, gått med på att ta emot före detta fångar.
Vilka åtgärder har kommissionen vidtagit för att hjälpa EU och dess medlemsstater att bidra till att Guantánamo stängs, även när det gäller att ta emot före detta fångar?
Vilka konkreta åtgärder har kommissionen vidtagit när det gäller att garantera rätt till gottgörelse och rättvis och skälig ersättning för personer som förts bort i samband med extraordinära överlämnanden och för personer som utsatts för tortyr?
När och på vilket sätt har kommissionen meddelat de amerikanska myndigheterna EU:s oro över att fångarna kan komma att förbli häktade på obestämd tid och ställda inför en militärdomstol och att dödsstraff kan komma att tillämpas?
MUNTLIG FRÅGA MED DEBATT O-0057/10
i enlighet med artikel 115 i arbetsordningen
från
Gabriele Albertini
för utskottet för utrikesfrågor ,
Vital Moreira
för utskottet för internationell handel
till kommissionen
Angående: Verkställandet av rådets förordning (EG) nr 1236/2005
Rådets förordning (EG) nr 1236/2005 av den 27 juni 2005 berör kontrollen av EU:s handel med vissa varor som kan användas till dödsstraff, tortyr eller annan grym, omänsklig eller förnedrande behandling eller bestraffning, och innehåller en förteckning över utrustning som bör förbjudas eller kontrolleras noggrant.
Förordningen trädde i kraft den 30 juni 2006 och var det första multilaterala instrumentet för handelskontroll i världen som förbjöd internationell handel med utrustning som i praktiken inte har något annat användningsområde än dödsstraff, tortyr eller annan grym behandling.
Tyvärr finns det allvarliga farhågor för att verkställandet av förordningen inte har skett allt igenom exemplariskt.
Vilka åtgärder planerar kommissionen att vidta för att förbättra övervakningen av, rapporteringen om och verkställandet av förordningen?
Vilka åtgärder kan vidtas om så visar sig vara fallet?
EUT L 200, 30.7.2005, s.1.
MUNTLIG FRÅGA MED DEBATT O-0060/10
i enlighet med artikel 115 i arbetsordningen
från
Philippe Juvin
,
Damien Abad
,
Simon Busuttil
,
Ernst Strasser
och
Andreas Schwab
för PPE -gruppen
till kommissionen
Angående: Tillämpning av EU:s lagstiftning om personuppgiftsskydd och konkurrenslagstiftning gentemot Google och i frågor som gäller reklam på nätet
Kommissionen har för sin del nyligen meddelat att den utreder de inlämnade klagomålen utan att för tillfället inleda en officiell undersökning.
Tvivel råder om huruvida de sökresultat som sökmotorn föreslår är opartiska, och dess reklamhantering ifrågasätts.
Googles makt som sökmotor ger detta företag den unika fördelen av att ha tillgång till detaljerade uppgifter om sin publik och dess användning av Internet.
Google förfogar således över stora mängder känsliga och personliga uppgifter om Internetanvändarna, vilket oroar många människor i EU.
Även brittiska Information Commissioner's Office har sällat sig till den tyska uppgiftsskyddsmyndighetens kritik av Google Street View, när det gäller insamlingen av privata Wifi-nät och MAC-adresser.
Ett sådant tillvägagångssätt innebär verkliga risker såtillvida att Google utan medborgarnas vetskap skulle kunna samköra de införskaffade uppgifterna med de MAC-adresser som samlats in genom nättjänster, och på detta sätt fastställa Internetanvändarnas marknadsföringsprofil.
I detta sammanhang uppmanar Europaparlamentet kommissionen att besvara följande frågor:
1.
Anser inte kommissionen, med hänsyn till att ärendet hänskjutits till de nationella konkurrensmyndigheterna i tre medlemsstater, att man bör inleda en undersökning på EU-nivå för att utreda om Google eventuellt gjort sig skyldigt till missbruk av dominerande ställning när det gäller reklam på Internet?
2.
Hur ställer sig kommissionen till frågan om att erkänna Internetuppgifter som personuppgifter, inom ramen för strategin för att uppdatera direktiv 95/46/EG ?
3.
Anser kommissionen, med tanke på de territoriella problemen, att det är lämpligt och möjligt att lagstifta på EU-nivå i syfte att bemöta den osäkerhet som råder när det gäller skyddet av den personliga integriteten och ifråga om reklam på nätet?
EGT L 281, 23.11.1995, s.
31.
Fråga för muntligt besvarande O-0135/2010
till rådet
Artikel 115 i arbetsordningen
Herbert Reul
för utskottet för industrifrågor, forskning och energi Angående: Klimatkonferensen i Cancún (COP 16)
Vilka konkreta yttre åtgärder avser rådet att vidta för att återupprätta förtroendet för förhandlingarna före och under klimatkonferensen i Cancún (både vad gäller förhandlingarna om Kyotoprotokollets andra åtagandeperiod, dvs. 2013–2020, och om långsiktiga gemensamma åtgärder fram till 2050)?
Fråga för muntligt besvarande O-000001/2011
till kommissionen
Artikel 115 i arbetsordningen
Gaston Franco
,
José Manuel Fernandes
,
Véronique Mathieu
,
Theodoros Skylakakis
,
Danuta Maria Hübner
,
Sophie Auconie
,
Nuno Teixeira
,
Jolanta Emilia Hibner
,
Esther Herranz García
,
Giovanni La Via
,
Elisabeth Morin-Chartier
,
Veronica Lope Fontagné
,
Mariya Nedelcheva
,
Barbara Matera
,
Catherine Soullie
,
Cristina Gutiérrez-Cortines
,
Dominique Vlasto
,
Anne Delvaux
,
Jean-Pierre Audy
,
Michel Dantin
för PPE -gruppen Angående: Gemenskapsåtgärder för att förhindra skogsbränder
I EU förstörs i snitt 500 000 hektar skog varje år till följd av skogsbränder.
De medlemsstater som drabbas hårdast kan uppleva 50 000 bränder årligen.
Under de senaste tio åren har antalet bränder ökat och överskrider nu Medelhavsregionernas gränser, vilket innebär att det blir ett allmänt problem som berör hela Europa.
Skogsbränder uppkommer främst pga. mänsklig verksamhet: 90 procent av bränderna har människorelaterade orsaker.
Efter det att förordning (EEG) nr 2158/92 upphävdes finns det inte längre någon specifik skogspolitik för att förebygga brandrisker.
Kan kommissionen med beaktande av detta, och med beaktande av att grönboken ”Skogsskydd och skoglig information i EU: Att förbereda skogen för klimatförändring” offentliggjordes den 1 mars 2010, överväga åtgärder för att förhindra skogsbränder?
Vilka framsteg har gjorts i form av konkreta åtgärder?
Förbereder kommissionen ytterligare skyddsåtgärder på detta område?
Fråga för muntligt besvarande O-000013/2011
till kommissionen
Artikel 115 i arbetsordningen
Vital Moreira
,
Francesca Balzani
för utskottet för internationell handel Angående: Ingåendet av ett Genèveavtal om handel med bananer
Kan kommissionen tillförsäkra att den kommer att sända in en särskild rapport till Europaparlamentet, vid behov åtföljd av lämpliga förslag, för den händelse att de ekonomiska villkoren som påverkar utkomsten för EU:s bananproducenter, också producenterna i de yttersta randområdena och i AVS-länderna, skulle försämras?
Vad tänker kommissionen göra för att det vidtas speciella initiativ för att ge bananodlarna en starkare kommersiell ställning inom de olika leveranskedjorna?
Håller kommissionen med om att resurser från åtgärderna i samband med bananodling bör fördelas mellan olika länder utgående från vilket respektive bortfall av bananexport och bananproduktion som förväntas drabba dem, samt också utgående från ländernas utvecklingsnivå, viktade indikatorer samt handel med bananer med EU?
Kan kommissionen se till att den så snabbt som möjligt lägger fram en konsekvensbedömning av hur avtalen kommer att påverka bananproducerande utvecklingsländer samt EU:s yttersta randområden fram till 2020?
Vad tänker kommissionen göra för att anslagen med stöd såväl av åtgärderna i samband med bananodling som med stöd av Posei-ordningen är tillräckliga för att bananproducenterna inom AVS-länderna och EU ska kunna anpassa sig till förändringarna i EU:s importordning?
Kan kommissionen tillförsäkra att en bedömning av åtgärderna i samband med bananodling kommer att göras 18 månader innan dessa åtgärder upphör att gälla?
Vad tänker kommissionen göra för att samma tullsatser ska gälla för Ecuador som för dess huvudsakliga konkurrenter?
Fråga för muntligt besvarande O-000054/2011
till rådet
Artikel 115 i arbetsordningen
Manfred Weber
,
Simon Busuttil
,
Georgios Papanikolaou
för PPE -gruppen Angående: Inrättandet av ett gemensamt vidarebosättningsprogram för EU
Enligt UNHCR vidarebosätts varje år omkring 200 000 flyktingar i ett tredjeland.
Europaparlamentets utskott för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor (LIBE-utskottet) ställde sig vid sitt sammanträde den 23 februari 2010 bakom tanken om ett vidarebosättningsprogram för EU och lade fram två förslag till betänkanden: ett om kommissionens meddelande om vidarebosättningsprogrammet för EU och ett annat om de föreslagna förändringarna av Europeiska flyktingfonden.
Båda dessa betänkanden antogs med stor majoritet av Europaparlamentet i maj 2010 och det rådde verkligt samförstånd mellan kommissionen, rådet och parlamentet om det politiska innehållet i betänkandena.
Nästan ett år efter omröstningen i Europaparlamentet väntar parlamentet fortfarande på att rådet ska fullborda medbeslutandeförfarandet.
Avser rådet att prioritera att fullborda detta medbeslutandeförfarande?
Fråga för muntligt besvarande O-000094/2011
till kommissionen
Artikel 115 i arbetsordningen
Baroness
Sarah Ludford
,
Renate Weber
,
Stanimir Ilchev
,
Nadja Hirsch
,
Jan Mulder
,
Nathalie Griesbeck
,
Sonia Alfano
,
Cecilia Wikström
,
Louis Michel
,
Jens Rohde
,
Sophia in 't Veld
för ALDE -gruppen Angående: Medlemsstaternas svar på tillflödet av migranter och deras effekter på Schengensamarbetet
Förra veckan införde Frankrike gränskontroller nära den italienska staden Ventimiglia, sedan den italienska regeringen hade undertecknat ett dekret som gör det möjligt för myndigheterna att utfärda tillfälliga uppehållstillstånd till de 25 800 tunisiska flyktingar som har kommit till ön Lampedusa efter regimens fall.
Migrationskonflikten mellan Frankrike och Italien och den bristande solidariteten inom EU med de medlemsstater som har störst problem med migrationsflödena skadar Schengensystemet.
Frestelsen att stänga inre gränser eller ignorera situationen för de medlemsstater som direkt påverkas av migrationsflödena är bara en panikreaktion.
Det finns ingen enkel, långsiktig och heltäckande lösning.
I stället behövs en ansvarsfull, effektiv och samordnad bevakning av EU:s yttre gränser och ett samstämt asylsystem i EU där länderna erkänner att de är beroende av varandra.
Det som har skett är ett tydligt bevis på att det nu är dags att börja ta ansvar och visa solidaritet.
Detta innefattar en gemensam asylpolitik med gemensamma förfaranden för att ge internationellt skydd.
Vi skulle därför vilja ha svar på följande frågor:
– Kan kommissionen ange huruvida kontrollerna vid gränsen mellan Frankrike och Italien nära Ventimiglia är motiverade?
– Kan kommissionen ange huruvida de tillfälliga uppehållstillstånd som Italien har utfärdat är förenliga med Schengenreglerna och om de verkligen innebär att innehavaren får röra sig fritt inom Schengenområdet?
Fråga för muntligt besvarande O-000113/2011
till kommissionen
Artikel 115 i arbetsordningen
Isabella Lövin
för Verts/ALE -gruppen Angående: Kris i fiskeindustrin på grund av de stigande oljepriserna
Oljepriset stiger överallt, även för fiskefartygen.
Vissa delar av fiskeindustrin är mycket beroende av fossila bränslen, för vilka kostnaderna kan uppgå till över hälften av driftskostnaderna.
Andra delar av denna industri drabbas inte alls lika hårt eftersom de utnyttjar mycket mindre energikrävande fiskerimetoder.
Fiskeindustrin står för minst 4 procent av den totala oljeanvändningen i världen och för en motsvarande mängd koldioxidutsläpp.
Denna industri behöver helt klart befria sig från sitt beroende av fossila bränslen.
Fiskeindustrin får redan nu omfattande bränslesubventioner på grund av sin skattefria ställning och de nya reglerna för stöd av mindre betydelse.
Har kommissionen för avsikt att minska eller upphäva bränsleskattebefrielsen med målet att minska fiskeindustrins energiberoende?
Fråga för muntligt besvarande O-000121/2011
till rådet
Artikel 115 i arbetsordningen
Claude Moraes
,
Birgit Sippel
för S&D -gruppen Angående: Den europeiska arresteringsordern
Den europeiska arresteringsordern har visat sig vara ett effektivt instrument för att bekämpa gränsöverskridande brottslighet och terrorism.
Dess rykte har dock svärtats ned genom att den enligt uppgift ska ha använts för förhör och inte för lagföring eller verkställighet av domar samt för mindre allvarliga brott utan vederbörlig hänsyn till om utlämningen är proportionerlig, trots de mänskliga och ekonomiska kostnaderna (uppskattningsvis 25 000 euro per utlämningsförfarande).
Dessutom respekterar inte alltid medlemsstaten sitt beslut att inte utfärda en europeisk arresteringsorder, vilket innebär att personen grips på nytt när denne passerar gränsen.
Det finns inte heller något system för ett adekvat rättsligt bistånd för personer som är efterlysta enligt den europeiska arresteringsordern, varken i den utfärdande eller i den verkställande medlemsstaten.
Slutligen är förhållandena i fängelserna i många av EU:s medlemsstater dessvärre så dåliga att de allvarligt hotar förtroendet för en korrekt behandling av fångar, som utgör grundvalen för den europeiska arresteringsordern och det snart genomförda rambeslutet om överföring av dömda personer.
- Vad kommer rådet att göra för att se till att den oproportionerliga användningen av den europeiska arresteringsordern omedelbart upphör både i lag och i praktiken?
- Vad kommer rådet att göra för att garantera att personer som är efterlysta enligt den europeiska arresteringsordern har faktisk rätt att ifrågasätta den europeiska arresteringsordern både i den utfärdande och i den verkställande medlemsstaten och för att se till att ett beslut att inte verkställa en europeisk arresteringsorder leder till att Schengen-registreringen tas bort?
- Vad kommer rådet att göra för att se till att de straffrättsliga standarderna och förhållandena i fängelserna förbättras i EU innan domstolarna griper in och stoppar ytterligare överföringar på grund av att personens grundläggande rättigheter kan komma att kränkas?
Fråga för muntligt besvarande O-000149/2011
till kommissionen
Artikel 115 i arbetsordningen
Monica Luisa Macovei
,
Mariya Nedelcheva
,
Simon Busuttil
,
Manfred Weber
för PPE -gruppen Angående: Åtgärder för att minska klyftan mellan korruptionslagstiftningen och verkligheten
1.
Hur kommer kommissionen i sin rapporteringsmekanism att kontrollera, bedöma och angripa nyckelfrågan om en effektiv tillämpning av lagstiftningen mot korruption, tillsammans med avskräckande sanktioner, med tanke på att denna lagstiftning för närvarande inte tillämpas alls eller endast bristfälligt?
2.
3.
Hur kommer kommissionen att involvera Europaparlamentet i dessa ansträngningar?
Fråga för muntligt besvarande O-000250/2011
till rådet
Artikel 115 i arbetsordningen
Sonia Alfano
,
Alexander Alvaro
,
Gianni Vattimo
,
Jens Rohde
,
Sophia in 't Veld
, Baroness
Sarah Ludford
,
Louis Michel
,
Andrea Zanoni
,
Ramon Tremosa i Balcells
,
Giommaria Uggias
,
Cecilia Wikström
för ALDE -gruppen Angående: "Munkavlelagen" i Italien
Det italienska parlamentet håller på att behandla ett förslag från Berlusconis regering om att ändra avlyssningslagen (särskilt kriterierna och förfarandena i samband med tillstånd, de typer av brottslighet som omfattas, elektronisk övervakning, avlyssningstillståndens varaktighet, användning av avlyssnad information i samband med annan brottslighet, skyldighet att korrigera information i bloggar samt undantag för parlamentsledamöter, präster och ärkebiskopar) och att begränsa möjligheten att offentliggöra utskrifter av avlyssningar genom sträng bestraffning av medier – även nya medier – som återger information om rättsliga utredningar innan de förberedande förhören har hållits, dvs. under en period som i Italien kan sträcka sig från tre till sex och ibland upp till tio år.
Detta nya lagförslag har väckt stor oro i Italien: föredraganden har sagt upp sig i protest efter omröstningen i utskottet, och Wikipedia har stängt av sin italienska sajt i protest mot lagförslaget, som innebär att bloggar på begäran måste korrigera information inom 48 timmar, vilket annars kan leda till böter på upp till 12 000 euro (den s.k. bloggdödarartikeln) .
1.
Anser rådet att de planerade ändringarna av Italiens avlyssningslag är proportionerliga och överensstämmer med EU:s normer om informationsfrihet, mediefrihet och medborgarnas rätt till information, som garanteras genom artikel 11 i EU:s stadga om de grundläggande rättigheterna och artikel 10 i den europeiska konventionen om skydd för de mänskliga rättigheterna och därtill hörande rättspraxis?
2.
Anser rådet att de föreslagna ändringarna är förenliga med EU:s mål för bekämpning av brott och organiserad brottslighet i Europa?
3.
Anser rådet att de föreslagna ändringarna – som har som uttalat mål att förhindra överträdelser av rättegångssekretessen och skydda privatlivet – står i proportion till den effekt de kommer att få i praktiken, dvs. att allvarligt begränsa den nationella brottsbekämpande verksamheten, som ska garantera medborgarnas säkerhet genom att förebygga och bekämpa brott och organiserad brottslighet, och begränsa informationsfriheten?
4.
Vilka åtgärder kommer rådet att vidta för att se till att informationsfriheten, yttrandefriheten och tryckfriheten garanteras i Italien och i EU, och att bekämpningen av brott och organiserad brottslighet i Italien och EU är effektiv?
För några månader sedan uttryckte nationella domarförbundet farhågor för en försvagning av de verktyg som finns för att bekämpa brottslighet och skydda medborgarnas säkerhet.
Det italienska tidningsutgivarförbundet, det nationella pressförbundet och journalistförbundet påpekade att den nya lagen är en ”munkavlelag” och kritiserade särskilt de höga böter som föreslås.
Även amerikanska myndigheter, bland annat biträdande justitieministern Lanny Breuer, uttryckte oro över de planerade ändringarna.
Fråga för muntligt besvarande O-000272/2011
till rådet
Artikel 115 i arbetsordningen
Renate Weber
,
Marielle De Sarnez
,
Jan Mulder
,
Cecilia Wikström
,
Sonia Alfano
,
Nathalie Griesbeck
,
Ramon Tremosa i Balcells
,
Andrea Zanoni
, Baroness
Sarah Ludford
,
Nadja Hirsch
,
Louis Michel
för ALDE -gruppen Angående: Barns rättigheter i EU
Den 15 februari 2011 offentliggjorde kommissionen meddelandet ”En EU-agenda för barns rättigheter” där man beskriver vilka åtgärder som kommer att vidtas under de kommande åren för att stärka barns rättigheter.
Vad anser rådet om agendan och hur kommer det att se till
- att medlemsstaternas myndigheter utreder våld och övergrepp mot barn på ett mer effektivt och kraftfullt sätt och att immunitet mot rättslig lagföring aldrig beviljas,
- att frihetsberövande av barn förbjuds och att lämpliga alternativa åtgärder genomförs,
- att alla barn ges tillgång till utbildning, sociala tjänster, hälsovård och rättsväsendet,
- att särskilda kategorier av barn som befinner sig i mycket sårbara situationer får hjälp genom speciella stödsystem (romer, underåriga utan medföljande vuxen eller som separerats från vuxna, barn till invandrare, barn som växer upp i fattigdom osv.),
- att barns civilstånd i samband med reser inom EU erkänns i enlighet med principen om ömsesidigt erkännande, utan diskriminering på grundval av förälderns civilstånd eller typ av förhållande (äktenskap, civilt partnerskap etc.) eller sexuella läggning,
- att ett EU-omfattande alarmsystem för fall där barn har förts bort eller försvunnit införs och att journumret 116 000 genomförs samt att båda dessa mekanismer fungerar väl,
- att dialoger med barn uppmuntras, även inom familjen?
Fråga för muntligt besvarande O-000287/2011
till kommissionen
Artikel 115 i arbetsordningen
Judith Sargentini
,
Jan Philipp Albrecht
,
Rui Tavares
,
Tatjana Ždanoka
,
Raül Romeva i Rueda
för Verts/ALE -gruppen Angående: Förhållanden vid frihetsberövande inom EU
Grönboken lyfter fram kopplingarna mellan förhållanden vid frihetsberövande och olika EU-instrument, såsom den europeiska arresteringsordern och den europeiska övervakningsordern och beskriver hur EU skulle kunna göra satsningar inom områden som frihetsberövande före rättegång, barnens situation och fängelseförhållanden.
I grönboken ingår en bilaga som åskådliggör den mycket varierade och ofta bekymmersamma situationen i medlemsstaterna, framför allt i fråga om antalet intagna som är frihetsberövade före rättegång, beläggningsnivån, överfulla fängelser, antalet intagna på fängelser i förhållande till landets befolkning samt antalet intagna fångar som inte är medborgare i landet.
Europadomstolen har också upprepade gånger, bland annat på grundval av rapporter från Europeiska kommittén till förhindrande av tortyr och omänsklig eller förnedrande behandling eller bestraffning, fördömt EU:s medlemsstater vad gäller fängelseförhållanden, perioden för frihetsberövande före rättegång och domstolsförvaltningen.
Hur kommer kommissionen att agera på EU-nivå för att försäkra sig om att de intagnas grundläggande rättigheter respekteras och att fängelseförhållandena i medlemsstaterna förbättras?
Anser kommissionen att det finns ett samband mellan undermåliga fängelseförhållanden och verkställandet av en europeisk arresteringsorder, såsom underströks i de frågor som togs upp i fallet C-396/11, Radu?
Kan kommissionen lägga fram konkret statistik om hur lång tid personer som utlämnats under en europeisk arresteringsorder i genomsnitt var frihetsberövade före rättegång?
Är kommissionen villig att föreslå förfarandekrav för misstänkta som är frihetsberövade före rättegång, inklusive möjligheter till prövning och bestämmelser om maximitider innan de frisläpps?
Är kommissionen villig att lägga fram EU-lagstiftning som införlivar de europeiska fängelseregler som Europarådet utarbetat, särskilt vad gäller logi, tillgång till hälsovård och rättshjälp?
Fråga för muntligt besvarande O-000288/2011
till rådet
Artikel 115 i arbetsordningen
Lívia Járóka
,
Simon Busuttil
för PPE -gruppen Angående: Avskaffande av diskrimineringen av romer
Trots EU:s ram för nationella strategier för integrering av romer, som infördes av kommissionen och välkomnades av rådet, och de riktlinjer som kommissionen utfärdade till medlemsstaterna för utarbetandet av de nationella strategierna för integrering av romer, fortsätter diskrimineringen av romer i EU.
Med hänsyn till den utbredda fientligheten gentemot zigenare och det bristfälliga genomförandet av befintliga bestämmelser, återstår det mycket att göra när det gäller icke diskriminering.
Alla europeiska länder, både nuvarande och framtida medlemmar av Europeiska unionen, måste engagera sig i en gemensam insats för att komma till rätta med denna historiska och sociala utestängning av kontinentens största etniska minoritet och ansluta sig till EU:s strategi för integrering av romer.
Kan rådet förpliktiga sig till att vidta åtgärder i syfte att förhindra diskriminerande behandling och samtidigt garantera att EU:s strategi genomförs?
Fråga för muntligt besvarande O-000009/2012
till kommissionen
Artikel 115 i arbetsordningen
Cristian Silviu Buşoi
,
Jürgen Creutzmann
,
Sophia in 't Veld
,
Wolf Klinz
för ALDE -gruppen
Andreas Schwab
,
Hans-Peter Mayer
,
Anna Maria Corazza Bildt
,
Małgorzata Handzlik
,
Philippe Juvin
,
Evelyne Gebhardt
,
Heide Rühle
Angående: Ungerns särskilda krisskatt för detaljhandelssektorn
Den 18 oktober 2010 antog Ungerns regering en särskild krisskatt för detaljhandelssektorn som i och med sin struktur får negativa effekter för utländska företag och skulle kunna hota etableringsfriheten samt utgöra olagligt statligt stöd.
I och med skattens utformning är det de facto de utländska detaljhandlarna som får betala denna betydande finansiella börda, som inte läggs på deras ungerska konkurrenter som ingår i ett nätverk av franchiseföretag, utan att deras omsättning beräknas över hela nätverket.
Den högsta skattsatsen gäller följaktligen endast utländska företag, vilket strider mot EU-lagstiftningen och diskriminerar vissa företagsmodeller.
Denna selektiva skatt, som i särskilt hög grad har påverkat stora utländska företag och lett till ojämlika villkor för utländska och inhemska företag, skulle eventuellt kunna ses som en överträdelse mot bestämmelserna om statligt stöd.
Situationen för de utländska detaljhandlarna i Ungern, som betalar mycket för en diskriminerande skatt, är oförändrad mer än ett år efter att den särskilda krisskatten infördes.
Kommissionen bör, mot bakgrund av ovanstående och i egenskap av fördragens väktare, sätta stopp för sådana protektionistiska åtgärder vid en tidpunkt då respekten för inremarknadsreglerna är viktigare än någonsin, i enlighet med parlamentets begäran i resolutionen av den 5 juli 2011 om en effektivare och rättvisare detaljhandelsmarknad ( P7_TA(2011)0307 ).
1.
2.
Har kommissionen fått ytterligare information från de ungerska myndigheterna, vilket begärts för att bedöma om den särskilda detaljhandelsskatten är förenlig med EU-lagstiftningen?
3.
Kommer kommissionen att ytterligare undersöka skatten inom ramen för bestämmelserna om statligt stöd för att åtgärda den nuvarande betydande obalansen i konkurrenskraft?
4.
Vilka åtgärder avser kommissionen att vidta härnäst?
Kan kommission även ge en exakt tidsram för dessa undersökningar?
Föredragningslista
Strasbourg
Måndagen den 3 maj 2004 - onsdagen den 5 maj 2004
Måndagen den 3 maj 2004
18:00 - 19:00
Högtidligt öppnande av det utvidgade Europaparlamentets första sammanträde
Arbetsplan
Talartid ( artikel 120 i arbetsordningen)
Tisdagen den 4 maj 2004
10:00 - 11:00
Högtidlighållande av minnet av Jean Monnet samt av 20-årsdagen för förslaget till fördrag om upprättande av Europeiska unionen (1984 - Föredragande: Altiero Spinelli)
11:00 - 13:00
Allmän debatt
Det utvidgade EU:s framtid
Uttalanden av rådet och kommissionen
Mot en konstitution för Europa
13:00
Omröstning
15:00 - 20:00
Det utvidgade EU och dess grannskap
Uttalanden av kommissionen
Den europeiska ekonomiska och sociala modellen
EU-medborgarnas frihet och säkerhet
Talartid ( artikel 120 i arbetsordningen)
Onsdagen den 5 maj 2004
10:00 - 12:00
Kommissionens ordförande presenterar de nya ledamöterna av den utvidgade kommissionen
12:00 - 13:00
Omröstning
Talartid ( artikel 120 i arbetsordningen)
Tidsfrister
Artikel
40
Beredning av lagstiftningsdokument
1.
När ett förslag är upptaget i lagstiftningsprogrammet, kan ansvarigt utskott besluta att utse en föredragande som skall följa utarbetandet av förslaget.
När rådet eller kommissionen begär att parlamentet skall yttra sig, skall denna begäran vidarebefordras av talmannen till det utskott som ansvarar för beredningen av förslaget i fråga.
Bestämmelserna om första behandlingen i artiklarna 34-37, 49-56 och 66 skall tillämpas vid alla förslag till rättsakter, oavsett om de fordrar en, två eller tre behandlingar.
2.
Rådets gemensamma ståndpunkter skall hänvisas för beredning till det utskott som var ansvarigt vid första behandlingen.
Bestämmelserna om andra behandlingen i artiklarna 57-62 och 67 skall tillämpas vid gemensamma ståndpunkter.
3.
Under det förlikningsförfarande mellan parlamentet och rådet som följer på andra behandlingen får ingen återförvisning till utskott äga rum.
Bestämmelserna om tredje behandlingen i artiklarna 63-65 skall tillämpas vid förlikningsförfarandet.
4.
5.
Om en bestämmelse i arbetsordningen som rör andra och tredje behandlingen strider mot någon annan bestämmelse i arbetsordningen, skall de bestämmelser som rör andra och tredje behandlingen ha företräde.
Föredragningslista
Tisdagen den 14 september 2004
9:00 - 12:00 Omröstning om begäran om brådskande förfarande ( artikel 134 i arbetsordningen)
Begäran om brådskande förfarande
Internationella krigsförbrytartribunalen för f.d.
[ KOM(2004)0348 - C6-0041/2004 - 2004/0114(CNS)]
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Begäran om brådskande förfarande
Ekonomisk utveckling inom den turkcypriotiska befolkningsgruppen
Förslag till rådets förordning om införande av en stödordning för att stimulera den ekonomiska utvecklingen inom den turkcypriotiska befolkningsgruppen
[ KOM(2004)0465 - C6-0098/2004 - 2004/0145(CNS)]
Utskottet för utrikesfrågor
Tal av Europaparlamentets talman
Uttalande av kommissionen
Läget i Vitryssland
Lägesrapport om uppföljningen av kommissionens årliga politiska strategi för 2005
12:00 - 13:00 Omröstning
Bekräftelse av kalendern för Europaparlamentets sammanträdesperioder
2005
Begäran om samråd med Ekonomiska och sociala kommittén
Förslag till fördrag om en konstitution för Europa
Artikel 117 i arbetsordningen Begäran om samråd med Regionkommittén
Förslag till fördrag om en konstitution för Europa
Artikel 118 i arbetsordningen Betänkande Jan Mulder A6-0004/2004
Förslag till ändringsbudget nr 7/2004
om förslaget till Europeiska unionens ändringsbudget nr 7/2004 för budgetåret 2004
[11041/2004 - C6-0108/2004 - 2004/2039(BUD)]
Budgetutskottet
Betänkande Jan Mulder A6-0005/2004
Förslag till ändringsbudget nr 8/2004
om förslaget till Europeiska unionens ändringsbudget nr 8/2004 för budgetåret 2004
[11042/2004 – C6-0109/2004 – 2004/2066(BUD)]
Budgetutskottet
Förslag till beslut B6- /2004
Antalet ledamöter i de interparlamentariska delegationerna, delegationerna till de gemensamma parlamentariska kommittéerna och delegationerna till de parlamentariska samarbetskommittéerna
15:00 - 16:30 Rådets presentation av förslaget till allmän budget
Räkenskapsåret 2005
16:30 - 17:00 Meddelande från kommissionen
Mönsterskydd
17:00 - 18:30 Frågestund med frågor till kommissionen B6-0007/2004
18:30 - 19:30 Uttalanden av rådet och kommissionen
Humanitära situationen i Sudan
Talartid ( artikel 142 i arbetsordningen)
9:00 - 12:00 Tal av talmannen
De politiska gruppernas ordföranden:
PPE-DE: 4', PSE: 4', ALDE: 3', Verts/ALE: 2', GUE/NGL: 2', IND/DEM:2', UEN: 2', NI: 2'
Övriga punkter Kommissionen (inklusive repliker)
Ledamöter
PPE-DE
24
PSE
18
ALDE
9
Verts/ALE
5,5
GUE/NGL
5
IND/DEM
5
UEN
4
NI
4,5
15:00 - 16:30 Rådet (inklusive repliker)
Kommissionen (inklusive repliker)
Budgetutskottets ordförande
Föredragande (2 x 5')
De politiska gruppernas talesmän:
PPE-DE: 6', PSE: 6', ALDE: 5', Verts/ALE: 4', GUE/NGL: 4', IND/DEM:4', UEN: 4', NI: 4'
18:30 - 19:30 Rådet (inklusive repliker)
Kommissionen (inklusive repliker)
Ledamöter
PPE-DE
9
PSE
7
ALDE
3,5
Verts/ALE
2,5
GUE/NGL
2
IND/DEM
2
UEN
2
NI
2
Tidsfrister
Uttalande av kommissionen
Läget i Vitryssland
Resolutionsförslag
Måndagen den 13 september, 19:00
Ändringsförslag och gemensamma resolutionsförslag
Onsdagen den 15 september, 10:00
Betänkande Jan Mulder A6-0004/2004
Förslag till ändringsbudget nr 7/2004
Ändringsförslag till själva budgeten
har löpt ut
Återupptagande av ändringsförslag efter det att de förkastats i utskottet
har löpt ut
Förslag till fullständigt avslag
har löpt ut
Begäran om särskild omröstning, delad omröstning eller omröstning med namnupprop om ändringsförslagen till förslaget till budget
Måndagen den 13 september, 19:00
Betänkande Jan Mulder A6-0005/2004
Förslag till ändringsbudget nr 8/2004
Ändringsförslag till själva budgeten
har löpt ut
Återupptagande av ändringsförslag efter det att de förkastats i utskottet
har löpt ut
Förslag till fullständigt avslag
har löpt ut
Begäran om särskild omröstning, delad omröstning eller omröstning med namnupprop om ändringsförslagen till förslaget till budget
Måndagen den 13 september, 19:00
Förslag till beslut B6- /2004
Antalet ledamöter i de interparlamentariska delegationerna, delegationerna till de gemensamma parlamentariska kommittéerna och delegationerna till de parlamentariska samarbetskommittéerna
Ändringsförslag
Måndagen den 13 september, 19:00
Uttalanden av rådet och kommissionen
Humanitära situationen i Sudan
Resolutionsförslag
Tisdagen den 14 september, 10:00
Ändringsförslag och gemensamma resolutionsförslag
Onsdagen den 15 september, 10:00
Särskild omröstning - delad omröstning - omröstning med namnupprop Texter som kommer att gå till omröstning tisdag
Måndagen den 13 september, 19:00
Texter som kommer att gå till omröstning onsdag
Tisdagen den 14 september, 21:00
Texter som kommer att gå till omröstning torsdag
Onsdagen den 15 september, 21:00
Resolutionsförslag om debatter om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer ( artikel 115 i arbetsordningen)
Torsdagen den 16 september, 10:00
Föredragningslista
Strasbourg
Måndagen den 15 november 2004 - torsdag den 18 november 2004
Måndagen den 15 november 2004
17:00 - 18:00
Öppnande av sammanträdet samt arbetsplan
18:00 - 21:00
Utfrågningar av de nominerade kommissionsledamöterna
Tisdagen den 16 november 2004
9:00 - 12:00
Utfrågningar av de nominerade kommissionsledamöterna
15:00 - 18:00, 21:00 - 22:00
Gemensam debatt
Vapenhandel
Uttalande av rådet
Hävande av vapenembargot mot Kina
Betänkande Raül Romeva i Rueda A6-0022/2004
Vapenexport
Slut på den gemensamma debatten
Uttalanden av rådet och kommissionen
Operation Althea i Bosnien och Hercegovina
Gemensam debatt
Den turkcypriotiska befolkningsgruppen
Betänkande Anders Samuelsen A6-0031/2004
Europeiska byrån för återuppbyggnad
Betänkande Mechtild Rothe A6-0032/2004
Ekonomisk stödordning (Cypern)
Slut på den gemensamma debatten
Uttalanden av rådet och kommissionen
Klimatförändringar
22:00 - 24:00
Betänkande Dorette Corbey A6-0027/2004
Förpackningar och förpackningsavfall
Uttalande av kommissionen
Situationen i Kuba
Talartid ( artikel 142 i arbetsordningen)
Tidsfrister
Onsdagen den 17 november 2004
9:00 - 12:00
Rapport från Europeiska rådet och uttalande av kommissionen
Europeiska rådets möte (Bryssel den 4-5 november 2004)
12:00 - 12:30
Högtidligt möte
Sydafrika
12:00 - 13:00
Omröstning
15:00 - 18:30
Uttalande av Barroso, kommissionens ordförande
18:30 - 19:00
Frågestund med frågor till rådet B6-0132/2004
Talartid ( artikel 142 i arbetsordningen)
Tidsfrister
Torsdagen den 18 november 2004
10:00 - 11:00
Betänkande Proinsias De Rossa A6-0030/2004
Europeiska ombudsmannens verksamhet (2003)
11:00 - 13:00
Omröstning
15:00 - 16:00
Elfenbenskusten
Tibet (fallet Tenzin Deleg Rinpoche)
Mänskliga rättigheter i Eritrea
16:00 [eller efter de föregående debatterna]
Omröstning
Talartid ( artikel 142 i arbetsordningen)
Tidsfrister
-//EP//TEXT TA 20041216 ITEMS DOC XML V0//SV
Föredragningslista
Strasbourg
Måndagen den 7 mars 2005 - torsdag den 10 mars 2005
Måndagen den 7 mars 2005
17:00 - 21:00
Öppnande av sammanträdet samt arbetsplan
Betänkande Alain Lipietz A6-0032/2005
EIB:s verksamhetsberättelse (2003)
Andrabehandlingsrekommendation Esko Seppänen A6-0012/2005
Tillträde till naturgasöverföringsnät
Muntliga frågor
Alternativa energikällor
Betänkande Ingo Schmitt A6-0038/2005
Europeiskt flygledarcertifikat
Andrabehandlingsrekommendation Proinsias De Rossa A6-0003/2005
Sociala trygghetssystem
Talartid ( artikel 142 i arbetsordningen)
Tidsfrister
Tisdagen den 8 mars 2005
9:00 - 12:00, 21:00 - 24:00
Muntliga frågor
Uppföljningen av den fjärde världskvinnokonferensen om handlingsplanen från Peking (Beijing + 10)
Betänkande Ilda Figueiredo A6-0035/2005
Den sociala situationen i unionen
Betänkande Antolín Sánchez Presedo A6-0045/2005
Allmänna preferenssystemet
Betänkande Rainer Wieland A6-0040/2005
Överläggningar i utskottet för framställningar (2003-2004)
Betänkande John Bowis A6-0044/2005
Arbetet i den gemensamma parlamentariska församlingen AVS-EU (2004)
Gemensam debatt
Budgeten 2005 och 2006
Betänkande Valdis Dombrovskis A6-0043/2005
Budgetriktlinjer 2006
Eventuellt: Betänkande Salvador Garriga Polledo A6- /2005
Förslag till ändringsbudget 1/2005
Eventuellt: Betänkande Anne Elisabet Jensen A6- /2005
Beräknad budget inför det preliminära förslaget till ändringsbudget 2/2005
Slut på den gemensamma debatten
Uttalande av kommissionen
Handel med äggceller
12:00 - 13:00
Omröstning om färdigbehandlade texter (se omröstningsordningen sidan 2)
15:00 - 18:00
Uttalanden av rådet och kommissionen
Revidering av icke-spridningsavtalet - Kärnvapen i Nordkorea och Iran
Uttalanden av rådet och kommissionen
Situationen i Libanon
18:00 - 18:45
Meddelande från kommissionen
Tjänster på den inre marknaden / Patentbarhet av mjukvara
18:45 - 20:15
Frågestund med frågor till kommissionen B6-0019/2005
Talartid ( artikel 142 i arbetsordningen)
Tidsfrister
Onsdagen den 9 mars 2005
9:00 - 12:30
Uttalanden av rådet och kommissionen
Halvtidsöversyn av Lissabonstrategin
12:30 - 13:00
Omröstning om färdigbehandlade texter (se omröstningsordningen sidan 2)
15:00 - 17:30
Uttalanden av rådet och kommissionen
Förberedelser av Europeiska rådets möte (Bryssel, 22-23 mars 2005)
Uttalanden av rådet och kommissionen
Fängslad vårdpersonal i Libyen
17:30 - 19:00
Frågestund med frågor till rådet B6-0019/2005
21:00 - 24:00
Betänkande Pia Elda Locatelli A6-0046/2005
Politiska riktlinjer för forskningsstöd i Europeiska unionen
Gemensam debatt
Personuppgifter
Muntliga frågor
Överföring av passageraruppgifter
Muntliga frågor
Lagring och skydd av uppgifter
Slut på den gemensamma debatten
Eventuellt: Betänkande Margrete Auken A6- /2005
Finansiering av Natura 2000
Talartid ( artikel 142 i arbetsordningen)
Tidsfrister
Torsdagen den 10 mars 2005
10:00 - 12:00
Muntlig fråga
Den gemensamma organisationen av marknaden för socker
Betänkande Marie-Hélène Aubert A6-0039/2005
Ekologiska livsmedel och ekologiskt jordbruk
12:00 - 12:15
Parlamentet hedrar minnet av offren för terroristattentaten i Madrid den 11 mars 2004
12:15 - 13:00
Omröstning om färdigbehandlade texter (se omröstningsordningen sidan 2)
15:00 - 15:45
Uttalande av kommissionen
Situationen i Tibet
15:45 (eller efter avslutad debat) - 16:45
Vitryssland
Kambodja
Saudiarabien
16:45 [eller efter avslutad debatt]
Omröstning
Talartid ( artikel 142 i arbetsordningen)
Tidsfrister
-//EP//TEXT TA 20050526 ITEMS DOC XML V0//SV
Artikel
3
Valprövning
1.
Med utgångspunkt i ett betänkande från behörigt utskott skall parlamentet omgående granska de utfärdade bevisen och avgöra varje enskild ny ledamots mandat, samt eventuella tvister som uppkommer till följd av bestämmelserna i akten av den 20 september 1976 med undantag av invändningar som grundar sig på nationella vallagar.
2.
Behörigt utskotts betänkande skall grunda sig på de officiella kungörelserna från de enskilda medlemsstaterna om det samlade valresultatet, vilka innehåller namnen på de valda kandidaterna och deras ersättare samt en rangordning baserad på valresultatet.
Giltigheten av en ledamots mandat kan inte bekräftas förrän ledamoten har avgivit de skriftliga förklaringar som följer av artikel 7 i akten av den 20 september 1976 och bilaga I till arbetsordningen.
Parlamentet kan när som helst på grundval av ett betänkande från sitt behöriga utskott yttra sig om varje invändning mot ett mandats giltighet.
3.
4.
När behöriga myndigheter i medlemsstaterna inleder ett förfarande som kan leda till att en ledamot skiljs från sitt uppdrag, skall talmannen begära regelbunden information från dem om hur förfarandet framskrider.
Talmannen skall hänvisa ärendet till behörigt utskott, och parlamentet kan yttra sig på förslag av detta utskott.
5.
Varje ledamot, vars mandat inte har prövats eller för vilken det inte har fattats beslut i en tvist, får delta i parlamentets och dess organs sammanträden med oinskränkta rättigheter.
6.
I början av varje valperiod skall talmannen uppmana medlemsstaternas behöriga myndigheter att förse parlamentet med alla de upplysningar som krävs för att denna artikel skall kunna tillämpas.
Avtal om vinodling mellan Europeiska unionen och Amerikas förenta stater
Europaparlamentets resolution om vinavtalet mellan Europeiska unionen och Förenta staterna
Olja
Europaparlamentets resolution om oljeberoendet
Reform av Förenta nationerna och Millenieutvecklingsmålen
Europaparlamentets resolution om resultaten från Förenta nationernas världstoppmöte (14–16 september 2005)
Vitryssland
Europaparlamentets resolution om Vitryssland
Relationerna mellan EU och Indien
Europaparlamentets resolution om ett strategiskt partnerskap mellan EU och Indien (2004/2169(INI))
Andelen förnybar energi i EU
Europaparlamentets resolution om andelen förnybar energi i EU och förslag på konkreta åtgärder (2004/2153(INI))
Minska antalet dödsoffer i trafiken i EU
Europaparlamentets resolution om det Europeiska åtgärdsprogrammet för trafiksäkerhet: Att halvera antalet dödsoffer i trafiken i Europeiska unionen till år 2010: ett gemensamt ansvar (2004/2162(INI))
Nepal
Europaparlamentets resolution om Nepal
Tunisien
Europaparlamentets resolution om Tunisien
Vojvodina
Europaparlamentets resolution om skydd av den etniska mångfalden i Vojvodina
TECKENFÖRKLARING
*
Samrådsförfarandet
** I
** II
***
Samtyckesförfarandet
***I
Medbeslutandeförfarandet (första behandlingen)
***II
Medbeslutandeförfarandet (andra behandlingen)
***III
UPPLYSNINGAR ANGÅENDE OMRÖSTNINGAR
Om inget annat anges har föredraganden till talmannen skriftligen tillkännagivit sin inställning till ändringsförslagen.
FÖRKORTNINGAR FÖR UTSKOTTENS NAMN
AFET:
DEVE:
Utskottet för utveckling
INTA:
Utskottet för internationell handel
BUDG:
Budgetutskottet
CONT:
Budgetkontrollutskottet
ECON:
Utskottet för ekonomi och valutafrågor
EMPL:
Utskottet för sysselsättning och sociala frågor
ENVI:
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
ITRE:
Utskottet för industrifrågor, forskning och energi
IMCO:
Utskottet för den inre marknaden och konsumentskydd
TRAN:
Utskottet för transport och turism
REGI:
Utskottet för regional utveckling
AGRI:
PECH:
Fiskeriutskottet
CULT:
Utskottet för kultur och utbildning
JURI:
Utskottet för rättsliga frågor
LIBE:
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
AFCO:
Utskottet för konstitutionella frågor
FEMM:
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
PETI:
Utskottet för framställningar
FÖRKORTNINGAR FÖR DE POLITISKA GRUPPERNA
PPE-DE:
Gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater
PSE:
Europeiska socialdemokratiska partiets grupp
ALDE:
Gruppen Alliansen liberaler och demokrater för Europa
Verts/ALE:
Gruppen De gröna/Europeiska fria alliansen
GUE/NGL:
Gruppen Europeiska enade vänstern/Nordisk grön vänster
IND/DEM:
Gruppen Självständighet/Demokrati
UEN:
Gruppen Unionen för nationernas Europa
NI:
Grupplösa
Öppnande av sammanträdet
Det österrikiska ordförandeskapets program (debatt)
Parlamentets sammansättning
Omröstning
Budgetplan (omröstning)
Tillsättning av en undersökningskommitté beträffande bolaget Equitable Life Assurance Societys sammanbrott (omröstning)
Tillsättning av ett tillfälligt utskott för CIA:s påstådda användning av europeiska länder för transport och illegal internering av fångar (omröstning)
Restriktiva åtgärder mot vissa personer som misstänks för inblandning i mordet på Libanons före detta premiärminister Rafiq Hariri * (artikel 131 i arbetsordningen) (omröstning)
Hantering av avfall från utvinningsindustrin ***III (omröstning)
Kvalitet på badvatten ***III (omröstning)
Hur Århuskonventionen skall tillämpas på EG:s institutioner och organ ***II (omröstning)
Tillträde till marknaden för hamntjänster ***I (omröstning)
Afghanistan (omröstning)
Homofobin i Europa (omröstning)
Klimatförändring (omröstning)
Miljöaspekter på hållbar utveckling (omröstning)
Röstförklaringar
Rättelser till avgivna röster
Justering av protokollet från föregående sammanträde
Period av eftertanke (struktur, teman och ramar för en utvärdering av debatten om Europeiska unionen) (debatt)
Välkomsthälsning
Situationen i Tjetjenien efter valet och det civila samhället i Ryssland (debatt)
Frågestund (frågor till rådet)
Europeiska grannskapspolitiken (debatt)
Genomförande av Europeiska stadgan för småföretag (debatt)
Ordningsregler för Europaparlamentets ledamöter (ändring av arbetsordningen) (debatt)
Föredragningslista för nästa sammanträde
Avslutande av sammanträdet
NÄRVAROLISTA
PROTOKOLL
ORDFÖRANDESKAP: Josep BORRELL FONTELLES Talman
1 Öppnande av sammanträdet
Sammanträdet öppnades kl. 09.05.
2
Det österrikiska ordförandeskapets program (debatt)
Uttalande av rådet:
Det österrikiska ordförandeskapets program
Wolfgang Schüssel (rådets tjänstgörande ordförande) gjorde ett uttalande.
Talare:
José Manuel Barroso (kommissionens ordförande)
Talare:
Hans-Gert Poettering för PPE-DE-gruppen,
Martin Schulz för PSE-gruppen,
Graham Watson för ALDE-gruppen,
Daniel Marc Cohn-Bendit för Verts/ALE-gruppen,
Francis Wurtz för GUE/NGL-gruppen,
Roger Knapman för IND/DEM-gruppen,
Cristiana Muscardini för UEN-gruppen,
Hans-Peter Martin , grupplös,
Othmar Karas ,
Hannes Swoboda ,
Karin Resetarits ,
Johannes Voggenhuber ,
Kartika Tamara Liotard ,
Mario Borghezio ,
Konrad Szymański ,
Andreas Mölzer ,
Timothy Kirkhope ,
Poul Nyrup Rasmussen och
Silvana Koch-Mehrin .
ORDFÖRANDESKAP: Jacek Emil SARYUSZ-WOLSKI Vice talman
Talare:
Sepp Kusstatscher ,
Tobias Pflüger ,
Georgios Karatzaferis ,
Guntars Krasts ,
Sergej Kozlík ,
Jaime Mayor Oreja ,
Maria Berger ,
Patrick Louis ,
Jana Bobošíková ,
Antonio Tajani ,
Ralf Walter ,
Lena Ek ,
Françoise Grossetête ,
Csaba Sándor Tabajdi ,
Andrew Duff ,
João de Deus Pinheiro och
Nicola Zingaretti .
ORDFÖRANDESKAP: Josep BORRELL FONTELLES Talman
Talare:
Annemie Neyts-Uyttebroeck ,
Etelka Barsi-Pataky ,
Bernard Poignant ,
Bronisław Geremek ,
Gunnar Hökmark ,
Monika Beňová ,
Ria Oomen-Ruijten ,
Josef Zieleniec ,
Marianne Thyssen ,
Jacek Emil Saryusz-Wolski ,
Ursula Stenzel ,
Wolfgang Schüssel och
José Manuel Barroso .
Talmannen förklarade debatten avslutad.
ORDFÖRANDESKAP: Mario MAURO Vice talman
Talare:
Richard Howitt beklagade det faktum att en presskonferens som skulle äga rum samma eftermiddag, arrangerad av ledamöter från IND/DEM-gruppen, hade titeln ”Parlamentarisk autism” och begärde att denna titel skulle bytas ut.
Eija-Riitta Korhola opponerade sig mot titeln på resolutionsförslagen om homofobi.
3 Parlamentets sammansättning
4 Omröstning
4.1
Budgetplan (omröstning)
Resolutionsförslag som lagts fram av budgetutskottet i enlighet med artikel 54 i arbetsordningen
om Europeiska rådets gemensamma ståndpunkt avseende budgetplanen och förnyelsen av det interinstitutionella avtalet för 2007–2013 ( B6-0049/2006 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 1)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2006)0010
)
4.2
Tillsättning av en undersökningskommitté beträffande bolaget Equitable Life Assurance Societys sammanbrott (omröstning)
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 2)
FÖRSLAG TILL BESLUT
Antogs
(
P6_TA(2006)0011
)
Inlägg om omröstningen:
-
Heide Rühle för Verts/ALE-gruppen lade fram ett muntligt ändringsförslag till ändringsförslag 1, vilket beaktades.
4.3
Tillsättning av ett tillfälligt utskott för CIA:s påstådda användning av europeiska länder för transport och illegal internering av fångar (omröstning)
Förslag till beslut som lagts fram av talmanskonferensen i enlighet med artikel 176 i arbetsordningen
om tillsättning av ett tillfälligt utskott för CIA:s påstådda användning av europeiska länder för transport och illegal internering av fångar ( B6-0051/2006 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 3)
FÖRSLAG TILL BESLUT
Antogs
(
P6_TA(2006)0012
)
Inlägg om omröstningen:
-
-
4.4
Restriktiva åtgärder mot vissa personer som misstänks för inblandning i mordet på Libanons före detta premiärminister Rafiq Hariri * (artikel 131 i arbetsordningen) (omröstning)
Betänkande om rådets förslag till förordning om särskilda restriktiva åtgärder mot vissa personer som misstänks för inblandning i mordet på Libanons före detta premiärminister Rafiq Hariri [ KOM(2005)0614 - 15098/2005 - C6-0434/2005 - 2005/0234(CNS) ] - Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor.
Föredragande: Jean-Marie Cavada ( A6-0003/2006 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 4)
KOMMISSIONENS FÖRSLAG, ÄNDRINGSFÖRSLAG och FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs
(
P6_TA(2006)0013
)
4.5
Hantering av avfall från utvinningsindustrin ***III (omröstning)
Betänkande från Europaparlamentets delegation till förlikningskommittén
om förlikningskommitténs gemensamma utkast till Europaparlamentets och rådets direktiv om hantering av avfall från utvinningsindustrin och om ändring av direktiv 2004/35/EG [PE-CONS 3665/2005 - C6-0405/2005 - 2003/0107(COD) ] Föredragande: Jonas Sjöstedt ( A6-0001/2006 )
(Enkel majoritet erfordrades för godkännande)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 5)
GEMENSAMT UTKAST
Antogs (
P6_TA(2006)0014
)
4.6
Kvalitet på badvatten ***III (omröstning)
Betänkande från Europaparlamentets delegation till förlikningskommittén
om förlikningskommitténs gemensamma utkast till Europaparlamentets och rådets direktiv om förvaltning av badvattenkvaliteten och om upphävande av direktiv 76/160/EEG [PE-CONS 3659/2005 - C6 0373/2005 - 2002/0254(COD) ] Föredragande: Jules Maaten ( A6-0415/2005 )
(Enkel majoritet erfordrades för godkännande)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 6)
GEMENSAMT UTKAST
Antogs (
P6_TA(2006)0015
)
4.7
Hur Århuskonventionen skall tillämpas på EG:s institutioner och organ ***II (omröstning)
Andrabehandlingsrekommendation om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets förordning om tillämpning av bestämmelserna i Århuskonventionen om tillgång till information, allmänhetens deltagande i beslutsprocesser och tillgång till rättslig prövning i miljöfrågor på gemenskapens institutioner och organ [06273/2/2005 - C6-0297/2005 - 2003/0242(COD) ] - Utskottet för miljö, folkhälsa och livsmedelssäkerhet.
Föredragande: Eija-Riitta Korhola ( A6-0381/2005 )
(Kvalificerad majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 7)
RÅDETS GEMENSAMMA STÅNDPUNKT
Förklarades godkänt såsom ändrat av parlamentet
(
P6_TA(2006)0016
)
Inlägg om omröstningen:
-
Graham Booth yttrade sig om omröstningen om ändringsförslag 30.
4.8
Tillträde till marknaden för hamntjänster ***I (omröstning)
Betänkande om förslaget till Europaparlamentets och rådets direktiv om tillträde till marknaden för hamntjänster [ KOM(2004)0654 - C6-0147/2004 - 2004/0240(COD) ] - Utskottet för transport och turism.
Föredragande: Georg Jarzembowski ( A6-0410/2005 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 8)
KOMMISSIONENS FÖRSLAG
Talare:
Talare:
Martin Schulz för PSE-gruppen, och
Jens-Peter Bonde för IND/DEM-gruppen yttrade sig om denna begäran.
Parlamentet förkastade denna begäran genom omröstning med namnupprop (132 ja-röster, 523 nej-röster, 19 nedlagda röster).
Talare:
Willi Piecyk yttrade sig om omröstningsförfarandet.
Som en följd av att ändringsförslagen om förkastande antogs, förkastades kommissionens förslag.
Talare:
Jacques Barrot (kommissionens vice ordförande) yttrade sig om förkastandet av kommissionens förslag.
4.9
Afghanistan (omröstning)
Debatten hölls den 26.10.2005 (
punkt 11 i protokollet av den 26.10.2005 ).
-
Pasqualina Napoletano och
Emilio Menéndez del Valle för PSE-gruppen ,
om Afghanistan ( B6-0026/2006 ) ,
-
Emma Bonino för ALDE-gruppen ,
om Afghanistan ( B6-0030/2006 ) ,
-
José Ignacio Salafranca Sánchez-Neyra ,
João de Deus Pinheiro och
Jürgen Schröder för PPE-DE-gruppen ,
om Afghanistan ( B6-0042/2006 ) ,
-
Angelika Beer ,
Joost Lagendijk ,
Raül Romeva i Rueda och
Cem Özdemir för Verts/ALE-gruppen ,
om Afghanistan ( B6-0047/2006 ) ,
-
Cristiana Muscardini ,
Roberta Angelilli och
Inese Vaidere för UEN-gruppen ,
om Afghanistan ( B6-0048/2006 ) ,
-
André Brie och
Luisa Morgantini för GUE/NGL-gruppen ,
om Afghanistan ( B6-0054/2006 ) .
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 9)
RESOLUTIONSFÖRSLAG
RC-B6-0026/2006
(ersätter
B6-0026/2006 ,
B6-0030/2006 ,
B6-0042/2006 och
B6-0048/2006 ):
inlämnat av följande ledamöter:
José Ignacio Salafranca Sánchez-Neyra för PPE-DE-gruppen ,
Pasqualina Napoletano och
Emilio Menéndez del Valle för PSE-gruppen ,
Emma Bonino för ALDE-gruppen ,
Cristiana Muscardini ,
Roberta Angelilli ,
Inese Vaidere och
Konrad Szymański för UEN-gruppen
Antogs
(
P6_TA(2006)0017
)
Inlägg om omröstningen:
-
Emilio Menéndez del Valle för PSE-gruppen lade fram ett muntligt ändringsförslag till punkt 16, vilket beaktades.
(Resolutionsförslagen
B6-0047/2006 och
4.10
Homofobin i Europa (omröstning)
Resolutionsförslag
B6-0025/2006 ,
B6-0034/2006 ,
B6-0039/2006 ,
B6-0040/2006 och
B6-0043/2006
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 10)
RESOLUTIONSFÖRSLAG
RC-B6-0025/2006
(ersätter
B6-0025/2006 ,
B6-0039/2006 ,
B6-0040/2006 och
B6-0043/2006 ):
inlämnat av följande ledamöter:
Alexander Stubb för PPE-DE-gruppen ,
Martine Roure och
Michael Cashman för PSE-gruppen ,
Sophia in 't Veld för ALDE-gruppen ,
Kathalijne Maria Buitenweg ,
Jean Lambert ,
Monica Frassoni ,
Elisabeth Schroedter och
Raül Romeva i Rueda för Verts/ALE-gruppen ,
Giusto Catania ,
Jonas Sjöstedt ,
Vittorio Agnoletto ,
Roberto Musacchio och
Willy Meyer Pleite för GUE/NGL-gruppen .
Antogs
(
P6_TA(2006)0018
)
B6-0034/2006 bortföll.)
4.11
Klimatförändring (omröstning)
Resolutionsförslag
B6-0027/2006
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 11)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2006)0019
)
4.12
Miljöaspekter på hållbar utveckling (omröstning)
Betänkande om miljöaspekter på hållbar utveckling [ 2005/2051(INI) ] - Utskottet för miljö, folkhälsa och livsmedelssäkerhet.
Föredragande: Anne Ferreira ( A6-0383/2005 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 12)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2006)0020
)
Skriftliga röstförklaringar:
Muntliga röstförklaringar:
Betänkande Jules Maaten - A6-0415/2005
-
Andreas Mölzer
Betänkande Eija-Riitta Korhola - A6-0381/2005
-
Eija-Riitta Korhola
Betänkande Georg Jarzembowski - A6-0410/2005
-
Frank Vanhecke ,
Dirk Sterckx och
Christopher Heaton-Harris
Afghanistan (
RC-B6-0026/2006 )
-
Karin Scheele
Homofobin i Europa (
RC-B6-0025/2006 )
-
Eija-Riitta Korhola ,
Romano Maria La Russa och
Francesco Enrico Speroni
Klimatförändringar (
B6-0027/2006 )
-
Eija-Riitta Korhola
6 Rättelser till avgivna röster
Den elektroniska versionen på Europarl uppdateras regelbundet under högst två veckor efter den aktuella omröstningsdagen.
Därefter slutförs förteckningen över rättelserna till de avgivna rösterna för att översättas och offentliggöras i Europeiska unionens officiella tidning.
ORDFÖRANDESKAP: Josep BORRELL FONTELLES Talman
Martine Roure hade låtit meddela att hon hade varit närvarande men att hennes namn inte förekom på närvarolistan.
Protokollet från föregående sammanträde justerades.
8
Period av eftertanke (struktur, teman och ramar för en utvärdering av debatten om Europeiska unionen) (debatt)
Betänkande om perioden av eftertanke: struktur, teman och ramar för en utvärdering av debatten om Europeiska unionen [ 2005/2146(INI) ] - Utskottet för konstitutionella frågor. medföredragande: Johannes Voggenhuber och Andrew Duff ( A6-0414/2005 )
Andrew Duff och
Johannes Voggenhuber (medföredragande) redogjorde för betänkandet.
Talare:
Hans Winkler (rådets tjänstgörande ordförande) och
Margot Wallström (kommissionens vice ordförande) .
Talare:
Elmar Brok (föredragande av yttrande från utskottet AFET),
Hannes Swoboda (föredragande av yttrande från utskottet ITRE),
Paolo Costa (föredragande av yttrande från utskottet TRAN),
Vladimír Železný (föredragande av yttrande från utskottet REGI),
Willem Schuth (föredragande av yttrande från utskottet AGRI),
Maria Berger (föredragande av yttrande från utskottet JURI),
Jean-Marie Cavada (föredragande av yttrande från utskottet LIBE),
Edit Bauer (föredragande av yttrande från utskottet FEMM),
Alexander Stubb för PPE-DE-gruppen,
Richard Corbett för PSE-gruppen,
Bronisław Geremek för ALDE-gruppen,
Monica Frassoni för Verts/ALE-gruppen,
Francis Wurtz för GUE/NGL-gruppen, och
Jens-Peter Bonde för IND/DEM-gruppen .
ORDFÖRANDESKAP: Manuel António dos SANTOS Vice talman
Talare:
Brian Crowley för UEN-gruppen,
James Hugh Allister , grupplös,
Jean-Luc Dehaene ,
Carlos Carnero González ,
Ignasi Guardans Cambó ,
Sylvia-Yvonne Kaufmann ,
Bastiaan Belder ,
Irena Belohorská ,
Íñigo Méndez de Vigo ,
Jo Leinen ,
Jules Maaten ,
Roger Knapman ,
Jan Tadeusz Masiel ,
József Szájer ,
Pierre Moscovici ,
Nils Lundgren ,
Daniel Hannan ,
Genowefa Grabowska ,
Maria da Assunção Esteves ,
Pasqualina Napoletano ,
Panayiotis Demetriou ,
Stavros Lambrinidis ,
Reinhard Rack ,
Hans Winkler och
Margot Wallström .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 8.9 i protokollet av den 19.01.2006
.
10
Situationen i Tjetjenien efter valet och det civila samhället i Ryssland (debatt)
Uttalanden av rådet och kommissionen:
Situationen i Tjetjenien efter valet och det civila samhället i Ryssland
Hans Winkler (rådets tjänstgörande ordförande) och
Benita Ferrero-Waldner (ledamot av kommissionen) gjorde uttalanden.
Talare:
Charles Tannock för PPE-DE-gruppen,
Reino Paasilinna för PSE-gruppen,
Cecilia Malmström för ALDE-gruppen,
Bart Staes för Verts/ALE-gruppen,
Jonas Sjöstedt för GUE/NGL-gruppen,
Michał Tomasz Kamiński för UEN-gruppen,
Luca Romagnoli , grupplös,
Tunne Kelam ,
Richard Howitt ,
Milan Horáček ,
Aloyzas Sakalas ,
Józef Pinior ,
Hans Winkler och
Benita Ferrero-Waldner .
-
Michał Tomasz Kamiński och
Ģirts Valdis Kristovskis för UEN-gruppen ,
om situationen i Tjetjenien efter valen och det civila samhället i Ryssland ( B6-0028/2006 ) ;
-
Jan Marinus Wiersma ,
Reino Paasilinna ,
Richard Howitt och
Csaba Sándor Tabajdi för PSE-gruppen ,
om Tjetjenien efter valet och det civila samhället i Ryssland ( B6-0029/2006 ) ,
-
Cecilia Malmström för ALDE-gruppen ,
om Tjetjenien efter valet och det civila samhället i Ryssland ( B6-0032/2006 ) ,
-
Daniel Marc Cohn-Bendit ,
Milan Horáček ,
Tatjana Ždanoka ,
Marie Anne Isler Béguin ,
Hélène Flautre och
Bart Staes för Verts/ALE-gruppen ,
om Tjetjenien efter valet och det civila samhället i Ryssland ( B6-0037/2006 ) ,
-
Charles Tannock ,
Bogdan Klich och
Ari Vatanen för PPE-DE-gruppen ,
om Tjetjenien efter valet och det civila samhället i Ryssland ( B6-0041/2006 ) ,
-
Francis Wurtz för GUE/NGL-gruppen ,
om Tjetjenien efter valet och det civila samhället i Ryssland ( B6-0044/2006 ) .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 8.8 i protokollet av den 19.01.2006
.
ORDFÖRANDESKAP: Sylvia-Yvonne KAUFMANN Vice talman
11
Frågestund (frågor till rådet)
Parlamentet behandlade en rad frågor till rådet (
B6-0676/2005 ).
Talare:
Hans Winkler (rådets tjänstgörande ordförande) redogjorde närmare för vissa aspekter i det nya förfarandet.
Första delen
Fråga 1 (Liam Aylward): Klimatförändringar
H-1119/05 .
Liam Aylward ,
Paul Rübig och
Richard Seeber .
Fråga 2 hade dragits tillbaka.
Fråga 3 (Ursula Stenzel): Samordning mellan olika organ (EU, Europarådet, OSSE) och tillvaratagande av mänskliga rättigheter i samband med terroristbekämpning
H-1165/05 .
Ursula Stenzel ,
David Martin och
Reinhard Rack .
Fråga 4 (Diamanto Manolakou): Olaglig kidnappning och häktning av pakistanier som lever i Grekland
H-1178/05 .
Athanasios Pafilis (ersättare för frågeställaren) och
Dimitrios Papadimoulis .
Andra delen
Fråga 5 (Manuel Medina Ortega): Europa-Medelhavskonferensen i Barcelona
H-1110/05 .
Manuel Medina Ortega och
David Martin .
Fråga 6 (Bernd Posselt): Kosovos status
H-1126/05 .
H-1152/05 .
H-1177/05 .
Hans Winkler svarade på frågorna samt följdfrågor från
Bernd Posselt ,
Dimitrios Papadimoulis och
Othmar Karas .
Fråga 9 (John Bowis): Förföljelse och trakasserier av kristna
H-1149/05 .
John Bowis ,
Paul Rübig ,
James Hugh Allister och
Bernd Posselt .
Fråga 11 (Inger Segelström): Colombia
H-1159/05 .
Inger Segelström och
Paul Rübig .
H-1175/05 .
Athanasios Pafilis och
Paul Rübig .
De frågor som på grund av tidsbrist inte hade besvarats skulle erhålla skriftliga svar
(se bilagan till det fullständiga förhandlingsreferatet) .
Talmannen förklarade frågestunden med frågor till rådet avslutad.
ORDFÖRANDESKAP: Antonios TRAKATELLIS Vice talman
12
Europeiska grannskapspolitiken (debatt)
Betänkande om den Europeiska grannskapspolitiken [ 2004/2166(INI) ] - Utskottet för utrikesfrågor.
Föredragande: Charles Tannock ( A6-0399/2005 )
Charles Tannock redogjorde för sitt betänkande.
Talare:
Benita Ferrero-Waldner (ledamot av kommissionen) .
Talare:
Elmar Brok för PPE-DE-gruppen,
Pasqualina Napoletano för PSE-gruppen,
Paavo Väyrynen för ALDE-gruppen,
Marie Anne Isler Béguin för Verts/ALE-gruppen,
Erik Meijer för GUE/NGL-gruppen,
Bastiaan Belder för IND/DEM-gruppen,
Konrad Szymański för UEN-gruppen,
Ryszard Czarnecki , grupplös,
Paweł Bartłomiej Piskorski ,
Pierre Schapira ,
Diana Wallis , ordförande för delegationen för förbindelserna med Schweiz, Island och Norge samt till det Europeiska ekonomiska områdets (EEA) gemensamma parlamentarikerkommitté,
Cem Özdemir ,
Esko Seppänen ,
Gerard Batten ,
Ģirts Valdis Kristovskis ,
Frank Vanhecke ,
Francisco José Millán Mon ,
Panagiotis Beglitis ,
Cecilia Malmström ,
Hélène Flautre ,
Irena Belohorská ,
Anna Ibrisagic ,
Ana Maria Gomes ,
Jana Bobošíková ,
Alojz Peterle ,
Marianne Mikko ,
Christopher Beazley ,
Ioannis Varvitsiotis ,
Józef Pinior ,
Libor Rouček ,
Jana Hybášková ,
Bernd Posselt ,
Bogusław Sonik ,
Simon Busuttil ,
Benita Ferrero-Waldner och
Christopher Beazley som ställde en fråga vilken
Benita Ferrero-Waldner besvarade.
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 8.10 i protokollet av den 19.01.2006
.
13
Genomförande av Europeiska stadgan för småföretag (debatt)
Betänkande om genomförandet av Europeiska stadgan för småföretag [ 2005/2123(INI) ] - Utskottet för industrifrågor, forskning och energi.
Föredragande: Dominique Vlasto ( A6-0405/2005 )
Dominique Vlasto redogjorde för sitt betänkande.
Talare:
Günter Verheugen (kommissionens vice ordförande)
Talare:
Katerina Batzeli (föredragande av yttrande från utskottet ECON),
Philip Bushill-Matthews (föredragande av yttrande från utskottet EMPL),
Paul Rübig för PPE-DE-gruppen,
Pia Elda Locatelli för PSE-gruppen,
Jorgo Chatzimarkakis för ALDE-gruppen,
Ilda Figueiredo för GUE/NGL-gruppen,
Gerard Batten för IND/DEM-gruppen,
Guntars Krasts för UEN-gruppen,
Pilar del Castillo Vera ,
Reino Paasilinna ,
Jean Marie Beaupuy ,
Thomas Mann ,
Brigitte Douay ,
Šarūnas Birutis och
Edit Herczog .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 8.4 i protokollet av den 19.01.2006
.
ORDFÖRANDESKAP: Josep BORRELL FONTELLES Talman
14
Ordningsregler för Europaparlamentets ledamöter (ändring av arbetsordningen) (debatt)
Betänkande om ändring av Europaparlamentets arbetsordning gällande ordningsreglerna för Europaparlamentets ledamöter [ 2005/2075(REG) ] - Utskottet för konstitutionella frågor.
Föredragande: Gérard Onesta ( A6-0413/2005 )
Gérard Onesta redogjorde för sitt betänkande.
Talare:
Ingo Friedrich för PPE-DE-gruppen,
Richard Corbett för PSE-gruppen,
Ignasi Guardans Cambó för ALDE-gruppen,
Erik Meijer för GUE/NGL-gruppen,
Gerard Batten för IND/DEM-gruppen,
Íñigo Méndez de Vigo och
Rainer Wieland .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 8.3 i protokollet av den 19.01.2006
.
15 Föredragningslista för nästa sammanträde
Föredragningslistan för nästa sammanträde fastställdes ("Föredragningslista" PE 368.209/OJJE).
16 Avslutande av sammanträdet
Sammanträdet avslutades kl. 24.00.
Julian Priestley
Alejo Vidal-Quadras
Generalsekreterare
Vice talman
NÄRVAROLISTA
Följande skrev på:
Adamou
Agnoletto
Albertini
Allister
Alvaro
Andersson
Andrejevs
Andria
Andrikienė
Antoniozzi
Arif
Arnaoutakis
Ashworth
Assis
Atkins
Aubert
Audy
Auken
Ayala Sender
Aylward
Ayuso González
Bachelot-Narquin
Baco
Badia I Cutchet
Barón Crespo
Barsi-Pataky
Batten
Battilocchio
Batzeli
Bauer
Beaupuy
Beazley
Becsey
Beer
Beglitis
Belder
Belet
Belohorská
Bennahmias
Beňová
Berend
Berès
van den Berg
Berger
Berlato
Berman
Bersani
Bertinotti
Bielan
Birutis
Blokland
Bobošíková
Böge
Bösch
Bonde
Bonino
Bono
Booth
Borghezio
Borrell Fontelles
Bourlanges
Bourzai
Bowis
Bowles
Bozkurt
Bradbourn
Braghetto
Brejc
Brepoels
Breyer
Březina
Brie
Brok
Brunetta
Budreikaitė
van Buitenen
Buitenweg
Bullmann
van den Burg
Bushill-Matthews
Busk
Busquin
Busuttil
Buzek
Cabrnoch
Calabuig Rull
Callanan
Camre
Capoulas Santos
Carlotti
Carlshamre
Carnero González
Casa
Casaca
Cashman
Caspary
Castex
Castiglione
del Castillo Vera
Catania
Cavada
Cederschiöld
Cercas
Chatzimarkakis
Chichester
Chiesa
Chmielewski
Christensen
Chruszcz
Claeys
Clark
Cocilovo
Coelho
Cohn-Bendit
Corbett
Corbey
Cornillet
Costa
Cottigny
Coûteaux
Coveney
Cramer
Crowley
Marek Aleksander Czarnecki
Ryszard Czarnecki
D'Alema
Daul
Davies
de Brún
Degutis
Dehaene
Demetriou
Deprez
De Rossa
De Sarnez
Descamps
Désir
Deß
Deva
De Veyrac
De Vits
Díaz de Mera García Consuegra
Dičkutė
Didžiokas
Díez González
Dillen
Dimitrakopoulos
Dionisi
Di Pietro
Dobolyi
Dombrovskis
Doorn
Douay
Dover
Doyle
Drčar Murko
Duchoň
Dührkop Dührkop
Duff
Duka-Zólyomi
Duquesne
Ebner
Ehler
Ek
El Khadraoui
Elles
Esteves
Estrela
Ettl
Eurlings
Jill Evans
Robert Evans
Fajmon
Falbr
Farage
Fatuzzo
Fava
Fazakas
Ferber
Fernandes
Fernández Martín
Anne Ferreira
Elisa Ferreira
Figueiredo
Fjellner
Flasarová
Flautre
Florenz
Foglietta
Foltyn-Kubicka
Fontaine
Ford
Fourtou
Fraga Estévez
Frassoni
Freitas
Friedrich
Fruteau
Gahler
Gál
Gaľa
Galeote
García-Margallo y Marfil
García Pérez
Gargani
Garriga Polledo
Gaubert
Gauzès
Gawronski
Gebhardt
Gentvilas
Geremek
Geringer de Oedenberg
Gewalt
Gibault
Gierek
Giertych
Gill
Gklavakis
Glante
Glattfelder
Goebbels
Goepel
Golik
Gollnisch
Gomolka
Goudin
Grabowska
Grabowski
Graça Moura
Graefe zu Baringdorf
Gräßle
de Grandes Pascual
Grech
Griesbeck
Gröner
de Groen-Kouwenhoven
Groote
Grosch
Grossetête
Gruber
Guardans Cambó
Guellec
Guerreiro
Guidoni
Gurmai
Gutiérrez-Cortines
Guy-Quint
Gyürk
Hänsch
Hall
Hammerstein Mintz
Hamon
Hannan
Harangozó
Harkin
Harms
Hasse Ferreira
Hassi
Hatzidakis
Haug
Hazan
Heaton-Harris
Hedh
Hedkvist Petersen
Hegyi
Helmer
Henin
Hennicot-Schoepges
Hennis-Plasschaert
Herczog
Herranz García
Herrero-Tejedor
Hieronymi
Higgins
Hökmark
Honeyball
Hoppenstedt
Horáček
Hudacký
Hudghton
Hughes
Hutchinson
Hybášková
Ibrisagic
Ilves
in 't Veld
Isler Béguin
Itälä
Iturgaiz Angulo
Jackson
Jäätteenmäki
Jałowiecki
Janowski
Járóka
Jarzembowski
Jeggle
Jensen
Joan i Marí
Jöns
Jørgensen
Jonckheer
Juknevičienė
Kacin
Kaczmarek
Kallenbach
Kamall
Kamiński
Karas
Karatzaferis
Karim
Kasoulides
Kaufmann
Kauppi
Tunne Kelam
Kilroy-Silk
Kindermann
Kinnock
Kirkhope
Klamt
Klaß
Klinz
Knapman
Koch
Koch-Mehrin
Kohlíček
Konrad
Korhola
Kósáné Kovács
Koterec
Kozlík
Krahmer
Krasts
Kratsa-Tsagaropoulou
Krehl
Kreissl-Dörfler
Kristensen
Kristovskis
Krupa
Kuc
Kudrycka
Kuhne
Kułakowski
Kušķis
Kusstatscher
Kuźmiuk
Lagendijk
Laignel
Lamassoure
Lambert
Lambrinidis
Landsbergis
Lang
Langen
Langendries
Laperrouze
La Russa
Lauk
Lavarra
Lax
Lechner
Le Foll
Lehideux
Lehne
Lehtinen
Leichtfried
Leinen
Marine Le Pen
Le Rachinel
Letta
Lévai
Lewandowski
Liberadzki
Libicki
Lichtenberger
Lienemann
Liese
Liotard
Lipietz
Locatelli
Louis
Lucas
Ludford
Lulling
Lundgren
Lynne
Maat
Maaten
McAvan
McCarthy
McGuinness
McMillan-Scott
Madeira
Malmström
Manders
Maňka
Erika Mann
Thomas Mann
Manolakou
Markov
Marques
Martens
David Martin
Hans-Peter Martin
Martinez
Martínez Martínez
Masiel
Masip Hidalgo
Maštálka
Mastenbroek
Mato Adrover
Matsakis
Matsis
Matsouka
Mauro
Mavrommatis
Mayer
Mayor Oreja
Medina Ortega
Meijer
Méndez de Vigo
Menéndez del Valle
Meyer Pleite
Miguélez Ramos
Mikko
Mikolášik
Millán Mon
Mölzer
Montoro Romero
Moraes
Moreno Sánchez
Morgan
Morillon
Moscovici
Mote
Mulder
Musacchio
Muscardini
Muscat
Musotto
Musumeci
Myller
Napoletano
Nassauer
Nattrass
Navarro
Newton Dunn
Annemie Neyts-Uyttebroeck
Nicholson
Nicholson of Winterbourne
Niebler
van Nistelrooij
Novak
Obiols i Germà
Öger
Özdemir
Olajos
Olbrycht
Ó Neachtain
Onesta
Onyszkiewicz
Oomen-Ruijten
Ortuondo Larrea
Őry
Oviir
Paasilinna
Pack
Pafilis
Pahor
Paleckis
Panayotopoulos-Cassiotou
Pannella
Panzeri
Papadimoulis
Papastamkos
Parish
Patrie
Pavilionis
Pęk
Alojz Peterle
Pflüger
Piecyk
Pieper
Pīks
Pinheiro
Pinior
Piotrowski
Pirilli
Piskorski
Pistelli
Pittella
Pleguezuelos Aguilar
Pleštinská
Podkański
Poettering
Poignant
Polfer
Poli Bortone
Pomés Ruiz
Portas
Posdorf
Posselt
Prets
Procacci
Prodi
Protasiewicz
Purvis
Queiró
Quisthoudt-Rowohl
Rack
Radwan
Ransdorf
Rapkay
Rasmussen
Remek
Resetarits
Reul
Reynaud
Ribeiro e Castro
Riera Madurell
Ries
Riis-Jørgensen
Rivera
Rocard
Rogalski
Roithová
Romagnoli
Romeva i Rueda
Rosati
Roszkowski
Roth-Behrendt
Rothe
Rouček
Roure
Rudi Ubeda
Rübig
Rühle
Rutowicz
Ryan
Sacconi
Saïfi
Sakalas
Salafranca Sánchez-Neyra
Salinas García
Salvini
Samaras
Samuelsen
Sánchez Presedo
dos Santos
Sartori
Saryusz-Wolski
Savary
Savi
Sbarbati
Schapira
Scheele
Schenardi
Schierhuber
Schlyter
Schmidt
Schmitt
Schnellhardt
Schöpflin
Schröder
Schroedter
Schulz
Schuth
Schwab
Seeber
Seeberg
Segelström
Seppänen
Siekierski
Sifunakis
Silva Peneda
Sinnott
Sjöstedt
Skinner
Škottová
Smith
Sommer
Sonik
Sornosa Martínez
Spautz
Speroni
Staes
Staniszewska
Starkevičiūtė
Šťastný
Stenzel
Sterckx
Stevenson
Stockmann
Strejček
Strož
Stubb
Sturdy
Sudre
Surján
Swoboda
Szájer
Szejna
Szent-Iványi
Szymański
Tabajdi
Tajani
Takkula
Tannock
Tarabella
Tarand
Tatarella
Thomsen
Thyssen
Titford
Titley
Toia
Tomczak
Toubon
Toussas
Trakatellis
Trautmann
Triantaphyllides
Trüpel
Turmes
Tzampazi
Uca
Ulmer
Väyrynen
Vaidere
Vakalis
Valenciano Martínez-Orozco
Vanhecke
Van Hecke
Van Lancker
Van Orden
Varela Suanzes-Carpegna
Varvitsiotis
Vaugrenard
Ventre
Verges
Vergnaud
Vernola
Vidal-Quadras
de Villiers
Vincenzi
Virrankoski
Vlasák
Vlasto
Voggenhuber
Wagenknecht
Wallis
Walter
Watson
Henri Weber
Manfred Weber
Weiler
Weisgerber
Wieland
Wiersma
Wijkman
Wise
von Wogau
Wohlin
Bernard Piotr Wojciechowski
Janusz Wojciechowski
Wortmann-Kool
Wurtz
Wynn
Xenogiannakopoulou
Yañez-Barnuevo García
Záborská
Zahradil
Zaleski
Zani
Zapałowski
Zappalà
Zatloukal
Ždanoka
Železný
Zieleniec
Zīle
Zimmer
Zingaretti
Zvěřina
Zwiefka
Observatörer
Abadjiev Dimitar
Athanasiu Alexandru
Bărbuleţiu Tiberiu
Becşenescu Dumitru
Bliznashki Georgi
Buruiană Aprodu Daniela
Cappone Maria
Cioroianu Adrian Mihai
Corlăţean Titus
Coşea Dumitru Gheorghe Mircea
Creţu Corina
Creţu Gabriela
Dimitrov Martin
Dîncu Vasile
Duca Viorel
Dumitrescu Cristian
Ganţ Ovidiu Victor
Hogea Vlad Gabriel
Husmenova Filiz
Ilchev Stanimir
Ivanova Iglika
Kazak Tchetin
Kirilov Evgeni
Marinescu Marian-Jean
Mihăescu Eugen
Morţun Alexandru Ioan
Nicolae Şerban
Paparizov Atanas Atanassov
Parvanova Antonyia
Paşcu Ioan Mircea
Petre Maria
Podgorean Radu
Popa Nicolae Vlad
Popeangă Petre
Sârbu Daciana Octavia
Severin Adrian
Sofianski Stefan
Stoyanov Dimitar
Szabó Károly Ferenc
Tîrle Radu
Vigenin Kristian
Zgonea Valeriu Ştefan
EU vill öka arbetstagares rörlighet
Socialpolitik
2006-02-20 - 15:31
Dra nytta av EU:s inre marknad och arbeta utomlands.
Arbetstagares rörlighet är en vanlig förklaring till att den amerikanska ekonomin flyter bättre än den europeiska.
Det är troligt att en amerikan flyttar över kontinenten för ett jobb, medan endast 1,5 % av européerna lever och arbetar i ett annat land än deras eget.
På EU:s arbetsmarknad, som kännetecknas av hög arbetslöshet inom vissa regioner och sektorer och brist på färdigheter och arbetskraft inom andra, ses större rörlighet ofta som ett sätt att skapa bättre och fler jobb.
Större arbetskraftsrörlighet, både mellan och jobb och länder leder till högre sysselsättning.
Därför måste vi koncentrera oss på såväl jobb- som geografisk rörlighet".
EU statistik visar att under 2003 hade 8,2 % av EU:s totala arbetskraft bytt jobb efter ett år.
Det finns stora skillnader mellan länder.
I Storbritannien och Danmark är den årliga jobbrörligheten ungefär 13 %, jämfört med 5 % i Grekland och Sverige.
Anställda med erfarenhet av jobbrörlighet tenderar att vara bättre rustade att klara förändringar och att anpassa sig till nya miljöer.
"Globaliseringen förändrar arbetsmiljön och sätter press på arbetarna att bli flexiblare och bättre på att anpassa sig till förändringar.
Att det i nuläget saknas en verklig "mobilitetskultur" är därför en riktig barriär".
Med 1,5 % är antalet personer som arbetar i ett annat land ungefär på samma nivå som för 30 år sedan.
Trots gemensamma gränser och en ökning de senaste åren är gränsöverskridande pendling endast 0,2 %.
Europeiska året för arbetstagares rörlighet kommer att sammanfalla med en rad andra initiativ bland andra övergångsåtgärder för människors fria rörlighet i ett utvidgat EU och lanseringen av en ny webbportal med lediga tjänster från hela Europa.
I tillägg, förväntas framsteg att förbättra flytt av pensionsrättigheter och det gemensamma europeiska sjukförsäkringskortet, som redan används av 50 miljoner medborgare, kommer att bli tillängligt i alla 25 medlemsstaterna.
Webbportalen kommer att lanseras officiellt på måndag (20 februari) under en högnivåkonferens som kommer att inviga det europeiska året för arbetstagares rörlighet.
Jan Andersson, kommissionens ordförande José Manuel Barroso och kommissionär Spidla.
Jan Kulakowski, liberal Europaparlamentetsledamot och Jean Lambert, vice ordförande för Gruppen De Gröna kommer också att delta .
*Källa: Center för Europeiska politiska studier.
20060220STO05371 Webbplats Europeiska året för arbetstagares rörlighet: EURES webbplats: EP Utskott för sysselsättning och sociala frågor (EMPL):
SV
1
PHOTO
20060220PHT05368.jpg
SV
2
LINK
http://ec.europa.eu/employment_social/workersmobility2006/index_sv.htm
SV
3
LINK
http://europa.eu.int/eures/home.jsp?lang=en
SV
4
LINK
/activities/expert/committees/presentation.do?committee=1238&language=EN
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Internationella kvinnodagen: Avspark för kampanj mot tvångsprostitution
Kvinnors rättigheter/Lika möjligheter
2006-03-09 - 16:29
Kampen mot tvångsprostitution diskuteras i Europaparlamentet.
EU måste visa rött kort för påtvingad prostitution och bekämpa människohandel för sexuella ändamål.
Det sade deltagare i ett seminarium organiserat av Europaparlamentets utskott för kvinnors rättigheter på den internationella kvinnodagen 8 mars.
Med anledning av varningar om att stora evenemang, som sommarens fotbolls-VM i Tyskland, innebär en skarp ökning av tvångsprostitution ville utskottet utbyta åsikter och diskutera strategier och åtgärder för att bekämpa tvångsprostitution.
Utskottets ordförande Anna Záborská, slovakisk kristdemokrat, sade att "detta är inte slutet på debatten, debatten kommer att fortsätta tills tvångsprostitution upphör".
Modern form av slaveri
Margot Wallström, kommissionens vice ordförande, uttryckte djup oro och chock över denna moderna form av slaveri, då en människas kropp kanske kan säljas för ett pris lägre än en entrébiljett till fotbollsarenan.
Hennes kollega, vice ordförande Franco Frattini, gav vissa förslag på hur man kan tackla problemet, bland annat genom att införa temporära visum för en kort period under fotbolls-VM för medborgare från länder som kan vara ursprungsländer för människohandel.
Han kunde inte ge en exakt lista, men nämnde Latinamerika, länder söder om Sahara, Asien och Östeuropa.
Han föreslog dessutom en studie över hur lagstiftning för prostitution påverkar människohandelns omfattning, vidare sade han att det är viktigt att studera såväl efterfrågan som utbud.
Per Ravn Omdal, talade för den europeiska fotbollsorganisationen UEFA, han sade att "UEFA stöder EU:s arbete att bekämpa alla former av människohandel och utnyttjande".
Men han liksom FIFA:s ordförande Joseph Blatter konstaterade att fotbollsorganisationer inte kan kontrollera det som sker utanför fotbollsstadion.
NGO:s arbete
"Varje kvinna är viktig.
Detta är en lukrativ business som vi måste stoppa.
Visste du att en människohandlare kan tjäna upp till 67 000 dollar per år på bara en enda kvinna?" sade Brunhilde Raiser (Nationella rådet för Tysklands kvinnoorganisationer).
Frivillig prostitution?
"Man kan inte skilja på frivillig och påtvingad prostitution.
Den svenska lagstiftningen (kriminalisera sexköp) fungerar", sade Maria Carlshamre (ALDE, SE).
"I Tyskland, Österrike och Nederländerna orsakar prostitution problem", alla tre är länder där prostitution är legaliserat.
Tyska Hiltrud Breyer från Gruppen De gröna, bakom initiativet att lyfta upp frågan om tvångsprostitution, vädjade om "rent spel" under VM i fråga om påtvingad prostitution och uppmanade kommission att lägga fram ett direktiv om våld mot kvinnor.
"Detta är inte emot fotboll som sådant", sammanfattade Christa Prets (PSE, AT) - som är ansvarig för ett betänkande om människohandel som parlamentet antog i januari.
Hon tyckte att "det är oförståeligt att vissa trafikförseelser straffas hårdare än trafficking med människor".
När Europaparlamentet samlas 13-16 mars för plenarsammanträde i Strasbourg, kommer ledamöterna att använda en muntlig fråga till Europeiska kommissionen som en möjlighet att debattera möjliga åtgärder i kampen mot påtvingad prostitution under internationella idrottsevenemang.
20060309STO06004 Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män - Uttalande Europaparlamentets talman Borrell med anledning av Internationella kvinnodagen: Sessionsöversikt 13-16 mars 2006:
SV
1
PHOTO
20060309PHT06000.jpg
SV
2
LINK
/comparl/femm/womensday/2006/default_en.htm
SV
3
LINK
/president/Presidents_old/president_borrell/press_releases/en/files/cp0130.htm
-//EP//TEXT IM-PRESS 20060216BRI05330 FULL-TEXT NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Friare rörlighet i EU men begränsningar återstår
Sysselsättningspolitik
2006-06-01 - 11:16
Hantverkare från nya EU-länder kan dra nytta av nya arbetsmöjligheter.
"Gamla" och "nya" Europa tog ett steg närmare varandra den 1 maj.
Då öppnade Spanien, Portugal, Finland och Grekland sina arbetsmarknader för arbetstagare från de åtta central- och östeuropeiska länderna som anslöt till EU 2004.
På så sätt förenar de sig med Storbritannien, Irland och Sverige som öppnade sina arbetsmarknader vid utvidgningen.
2006 är det europeiska året för arbetstagares rörlighet, och nyheten mottogs med försiktig optimism från ledamöter som arbetar med frågan.
Jan Andersson, svensk socialdemokrat, och ordförande i Europaparlamentets utskott för sysselsättning och sociala frågor välkomnade öppnandet och sade att "det finns ett regelverk i EU för hur övergångsordningen ska hanteras och medlemsstaterna har att leva upp till detta.
Samtidigt anser jag att de EU-länder som ännu inte har avskaffat övergångsbestämmelserna för arbetstagare från de nya medlemsländerna, bör göra det så snart som möjligt."
Detta upprepades av Csaba Őry, ungersk ledamot från Gruppen för europeiska folkpartiet (kristdemokrater) och Europademokrater.
I april antog parlamentet Őrys betänkande om arbetstagares rörlighet.
Enligt betänkandet har bristande möjligheter för arbetstagare från de nya medlemsstaterna lett till att illegala arbeten, den svarta ekonomin och exploateringen av arbetstagare har ökat.
Att avveckla begränsningsåtgärder skulle, enligt betänkandet, skicka "en tydlig signal om solidaritet mellan medborgarna i västra och östra Europa".
2011 tidsfrist för de sista begränsningarna
Ekonomisk migration av arbetstagare är ett känsligt ämne, vilket förklarar varför, efter EU:s senaste utvidgning 2004, alla förutom tre av de femton gamla medlemsstaterna behöll "övergångperioder" för tillträdet till deras arbetsmarknader.
Den maximala tillåtna perioden för detta är sju år - men en "2+3+2"-årsformel gör det möjligt att gradvis införa rörlighet.
2011 är tidsfristen för att avlägsna alla begränsningar.
Frankrike, Italien och Luxembourg har anmält att de avser upphäva restriktionerna för svårrekryterade arbeten.
Nederländernas parlament ska ta ställning i frågan innan årets slut.
Tyskland och Österrike behåller begränsningarna till 2009.
Trots att Tyskland redan har beviljat 500 000 arbetstillstånd till migrerande arbetstagare från de nya EU-medlemmarna.
Från Warszawa till London, Dublin, Stockholm...
Frågan blir extra känslig eftersom "fri rörlighet av personer" är en av EU:s grundläggande rättigheter.
Arbetstagares rörlighet säkerställs i 1957 års Romfördrag.
Fördragets artikel 39 fastställer rätten att söka jobb, fritt ta anställning och vistas i en annan medlemsstat och rätt till lika behandling och tillgång till anställning.
De som planerar att arbeta utomlands hoppas på att alla EU-medlemsstater så snart som möjligt öppnar sina arbetsmarknader.
20060510STO08007 Europaparlamentets utskott för sysselsättning och sociala frågor: Csaba Őrys betänkande om övergångsbestämmelser på arbetsmarknaden (5 april 2006): Debatt om Őry-betänkandet (4 april 2006): Arbetstagares fria rörlighet - Fakta 2006 Europeiska året för arbetstagares rörlighet: Arbeta utomlands?
SV
1
PHOTO
20050818PHT00030.jpg
SV
2
LINK
/activities/expert/committees/presentation.do?committee=1238&language=SV
SV
5
LINK
http://ec.europa.eu/employment_social/free_movement/index_en.htm
SV
6
LINK
http://ec.europa.eu/employment_social/workersmobility_2006/index.cfm?language=SV
SV
7
LINK
http://ec.europa.eu/eures/
-//EP//TEXT TA P6-TA-2006-0129 0 NOT XML V0//SV
-//EP//TEXT CRE 20060404 ITEM-007 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Perioden av eftertanke - nästa steg
Europas framtid/Europeisk integration
2006-06-14 - 14:04
Beslut måste fattas om konstitutionen före slutet av 2007 så att överenskommelse om konstitutionen ska ligga färdig tills Europavalen 2009.
Europaparlamentet står i konstitutionsutskottets resolution fast vid sitt mål att en överenskommelse om konstitutionen ska ligga färdig när unionsmedborgarna röstar i valet till Europaparlamentet år 2009.
I dagsläget har sexton länder ratificerat det konstitutionella fördraget, medan två länder har röstat nej i nationella folkomröstningar.
Parlamentet upprepar sitt stöd för fördraget om upprättande av en konstitution för Europa och tror att försök att riva upp den övergripande kompromissen allvarligt skulle hota det europeiska politiska projektet.
Målet ska vara att man under andra halvan av 2007 fattar ett entydigt beslut om det konstitutionella fördragets öde.
De medlemsstater som ännu inte avslutat ratificeringsförfarandet måste ta fram trovärdiga alternativ för hur de har för avsikt att föra utvecklingen framåt.
En dialog bör också föras med representanterna för de länder i vilka folkomröstningen om det konstitutionella fördraget fick ett negativt resultat att utreda om och under vilka omständigheter det vore möjligt för dem att återuppta ratificeringsförfarandet.
Kommissionen uppmanas att stödja denna strategi och lägga fram en färdplan.
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
Föredragningslista
Torsdagen den 6 juli 2006
10:00 - 11:50, 15:00 - 16:00 Betänkande Marie-Arlette Carlotti A6-0210/2006
Utveckling och migration
om utveckling och migration
[ 2005/2244(INI) ]
Utskottet för utveckling
Betänkande Frithjof Schmidt A6-0207/2006
Rättvis handel och utveckling
om rättvis handel och utveckling
[ 2005/2245(INI) ]
Utskottet för utveckling
Muntlig fråga
Resultaten från WTO:s möte i Genève i slutet av april samt framtidsperspektiv
O-0036/2006 Enrique Barón Crespo B6-0314/2006 kommissionen Resultaten från WTO:s möte i Genève i slutet av april samt framtidsperspektiv
Utskottet för internationell handel
Muntlig fråga
Angivande av ursprungsland för vissa produkter som importeras från tredjeländer ("ursprungsmärkning")
O-0065/2006 Enrique Barón Crespo B6-0316/2006 kommissionen Angivande av ursprungsland för vissa produkter som importeras från tredjeländer ("ursprungsmärkning")
Utskottet för internationell handel
12:00 - 13:00 Omröstning
I enlighet med artikel 131 i arbetsordningen:
Betänkande Christoph Konrad A6-0209/2006
Uppbörden av mervärdesskatt och kampen mot skattefusk och skatteundandragande
om förslaget till rådets direktiv om ändring av direktiv 77/388/EEG när det gäller vissa åtgärder för att förenkla uppbörden av mervärdesskatt och för att förhindra skattefusk eller skatteundandragande samt om upphävande av vissa beslut om tillstånd till avvikelser
[ KOM(2005)0089 - C6-0100/2005 - 2005/0019(CNS) ]
Utskottet för ekonomi och valutafrågor
Artikel 131 i arbetsordningen
Betänkande Gabriele Zimmer A6-0211/2006
Ett partnerskap för tillväxt, stabilitet och utveckling mellan EU och Västindien
om ett partnerskap för tillväxt, stabilitet och utveckling mellan EU och Västindien
[ 2006/2123(INI) ]
Utskottet för utveckling
Artikel 131 i arbetsordningen
Betänkande 2 Stephen Hughes A6-0218/2006
Skydd för anställda inom hälsovårdssektorn i Europa mot infektioner som överförs via blodet till följd av skador orsakade av sprutor
om skydd för anställda inom hälsovårdssektorn i Europa mot infektioner som överförs via blodet till följd av skador orsakade av sprutor
[ 2006/2015(INI) ]
Utskottet för sysselsättning och sociala frågor
Artiklarna 39 och 131 i arbetsordningen
Betänkande Konrad Szymański A6-0164/2006
Europeiskt grannskaps- och partnerskapsinstrument
om förslaget till Europaparlamentets och rådets förordning om fastställande av de allmänna principerna för upprättandet av ett europeiskt grannskaps- och partnerskapsinstrument
[ KOM(2004)0628 - C6-0129/2004 - 2004/0219(COD) ]
Utskottet för utrikesfrågor
Debatt: 17 maj 2006
Betänkande Angelika Beer A6-0157/2006
Stabilitetsinstrument
om förslaget till Europaparlamentets och rådets förordning om upprättande av ett stabilitetsinstrument
[ KOM(2004)0630 - C6-0251/2004 - 2004/0223(COD) ]
Utskottet för utrikesfrågor
Debatt: 17 maj 2006
Betänkande István Szent-Iványi A6-0155/2006
Instrument för stöd inför anslutningen
om förslaget till rådets förordning om upprättande av ett instrument för stöd inför anslutningen
[ KOM(2004)0627 - C6-0047/2005 - 2004/0222(CNS) ]
Utskottet för utrikesfrågor
Debatt: 17 maj 2006
Betänkande Ingeborg Gräßle A6-0057/2006
Budgetförordning för Europeiska gemenskapernas allmänna budget
om förslaget till rådets förordning om ändring av rådets förordning (EG, Euratom) nr 1605/2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
[ KOM(2005)0181 - C6-0234/2005 - 2005/0090(CNS) ]
Budgetutskottet
Slutomröstning
Resolutionsförslag B6-0275/2006 /rev
Ändring av protokollet om privilegier och immunitet
Debatt: 26 april 2006
Somalia
Mauretanien
Yttrandefrihet på Internet
17:00 [eller efter att föregående debatter har avslutats] - 18:00 Omröstning
Talartid ( artikel 142 i arbetsordningen)
10:00 - 11:50, 15:00 - 16:00 Föredragande (2 x 5')
Föredragande av yttrande (5 x 1')
Frågeställare (2 x 5')
Kommissionen (inklusive repliker)
Ledamöter
PPE-DE
29
PSE
22
ALDE
11
Verts/ALE
6
GUE/NGL
6
UEN
5
IND/DEM
5
NI
6
16:00 [eller efter föregående debatt] - 17:00 Författare till varje resolutionsförslag
Kommissionen
Ledamöter
PPE-DE
7
PSE
6
ALDE
4
Verts/ALE
3
GUE/NGL
3
UEN
2
IND/DEM
2
NI
3
Tidsfrister
Betänkande Marie-Arlette Carlotti A6-0210/2006
Utveckling och migration
Ändringsförslag
har löpt ut
Betänkande Frithjof Schmidt A6-0207/2006
Rättvis handel och utveckling
Ändringsförslag
har löpt ut
Muntlig fråga
Angivande av ursprungsland för vissa produkter som importeras från tredjeländer ("ursprungsmärkning")
O-0065/2006 Enrique Barón Crespo B6-0316/2006 kommissionen Angivande av ursprungsland för vissa produkter som importeras från tredjeländer ("ursprungsmärkning")
Utskottet för internationell handel
Resolutionsförslag
Måndagen den 3 juli, 19:00
Ändringsförslag och gemensamma resolutionsförslag
Onsdagen den 5 juli, 10:00
Betänkande Konrad Szymański A6-0164/2006
Europeiskt grannskaps- och partnerskapsinstrument
Ändringsförslag
har löpt ut
Betänkande Angelika Beer A6-0157/2006
Stabilitetsinstrument
Ändringsförslag
har löpt ut
Betänkande István Szent-Iványi A6-0155/2006
Instrument för stöd inför anslutningen
Ändringsförslag
har löpt ut
Resolutionsförslag B6-0275/2006 /rev
Ändring av protokollet om privilegier och immunitet
Ändringsförslag
Måndagen den 3 juli, 19:00
Somalia
Resolutionsförslag ( artikel 115 i arbetsordningen)
Måndagen den 3 juli, 20:00
Ändringsförslag och gemensamma resolutionsförslag ( artikel 115 i arbetsordningen)
Onsdagen den 5 juli, 13:00
Mauretanien
Resolutionsförslag ( artikel 115 i arbetsordningen)
Måndagen den 3 juli, 20:00
Ändringsförslag och gemensamma resolutionsförslag ( artikel 115 i arbetsordningen)
Onsdagen den 5 juli, 13:00
Yttrandefrihet på Internet
Resolutionsförslag ( artikel 115 i arbetsordningen)
Måndagen den 3 juli, 20:00
Ändringsförslag och gemensamma resolutionsförslag ( artikel 115 i arbetsordningen)
Onsdagen den 5 juli, 13:00
Särskild omröstning - delad omröstning - omröstning med namnupprop Texter som kommer att gå till omröstning tisdag
Måndagen den 3 juli, 19:00
Texter som kommer att gå till omröstning onsdag
Tisdagen den 4 juli, 21:00
Texter som kommer att gå till omröstning torsdag
Onsdagen den 5 juli, 21:00
Resolutionsförslag om debatter om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer ( artikel 115 i arbetsordningen)
Torsdagen den 6 juli, 10:00
Pakistans president Musharraf besöker Europaparlamentet
Yttre förbindelser
2006-09-15 - 17:44
President Musharraf på Europaparlamentet.
Pakistans president, General Pervez Musharraf, avslutade ett tvådagarsbesök på Europaparlamentet med att träffa de politiska gruppernas ordförande och Europaparlamentets talman Josep Borrell.
Musharrafs huvudbudskap var en uppmaning till västvärlden att se Pakistan som en viktig bundsförvant i kriget mot terrorism och att EP-ledamöterna kan bidra till att främja handelsförbindelserna mellan EU och Pakistan.
Han tackade dessutom EU för dess humanitära stöd efter jordbävningen 2005.
Efter mötet i onsdags (13 september) uppmärksammade Borrell president Musharrafs ansträngningar att "bygga upp förtroendet" med Indien över det omtvistade Kashmir och lyfte även fram den pakistanska arméns kamp mot terrorister och talibanrörelsen.
Han sade att frågor om mänskliga rättigheter och kärnvapenspridning också tagits upp av de politiska gruppernas ordförande under mötet.
Musharraf efterlyser stärkt samarbete mellan EU-Pakistan
I tisdags (12 september) mötte Musharraf Europaparlamentets utskott för utrikesfrågor.
Under mötet redogjorde han för de utmaningar Pakistan står inför, och han fick också svara på en del tuffa frågor från ledamöterna om sitt styre (läs pressmeddelande om mötet genom att klicka på länken nedan).
Hans framförande handlade framförallt om Pakistans behov av hjälp från EU för att överkomma de svårigheter som landet står inför.
Pakistans demokratiska och ekonomiska utveckling är i behov av betydande stöd.
Och Musharraf ville gärna se en förbättrad marknadstillgång för pakistanska varor till EU.
På hemmaplan har Pakistans armé tagit upp kampen mot al-Qaida och talibanrörelsens medlemmar.
Musharraf lovade att fortsätta kampen mot "talibaniseringen" av vissa delar av Pakistan.
Han bad om EU:s hjälp att lösa den pågående tvisten om Kashmir som under nästan 60 år har lett till spända relationer med Indien.
Musharraf underströk sitt lands "måttliga, religiösa och toleranta" natur och sade att det endast har kärnvapen för att bemöta det indiska kärnvapenhotet.
Ledamöterna ifrågasatte Pakistans "demokratiska underskott" (inga demokratiska val, ingen separation mellan militär och politik) och bristen på religionstolerans.
De yrkade även på att dödsstraffets upphörande.
Ordföranden för utskottet för utrikesfrågor, tyske kristdemokraten Elmar Brok, framhöll att Pakistan går igenom en avgörande tid i sin historia, samtidigt som det spelar en viktig roll med sin "enorma omfattning av olika ansvar."
Neena Gill, brittisk socialist, och ordförande för parlamentets delegation för förbindelserna med länderna i Sydasien sade att Pakistan "är en viktig allierad för Europa i kampen mot internationell terrorism."
Men, hon uppmanade presidenten att vidta åtgärder för att "få ett slut på könsdiskriminering i alla dess former" i Pakistan liksom förekomsten av hedersmord på kvinnor (som exempelvis kan anklagas för otrohet).
Neena Gill sade att presidenten måste "se till att mänskliga rättigheter respekteras i hela Pakistan."
På frågor om hans egen framtid som general svarade Musharraf att han kommer att "fatta beslut 2007 i enlighet med Pakistans konstitution."
20060914STO10661 Pakistans president hoppas på mer handel med EU:
SV
1
PHOTO
20060913PHT10651.jpg
-//EP//TEXT IM-PRESS 20060908IPR10492 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Europaparlamentet och kampen mot bröstcancer
Folkhälsa
2006-10-03 - 14:45
Varannan minut får en kvinna i EU diagnosen bröstcancer, var sjätte minut dör en kvinna av sjukdomen.
Ett seminarium om yrkesutbildning för bröstsjukvårdspersonal anordnas i oktober, och plenum debatterar några dagar senare den senaste utvecklingen i kampen mot bröstcancer.
Cancer är den vanligaste dödsorsaken i EU.
35 % av de 275 000 kvinnor som varje år får diagnosen bröstcancer är under 55 år.
Internationella bröstcancermånaden
Internationella bröstcancermånaden, som äger rum årligen i oktober, syftar till att öka medvetenheten och kunskapen om sjukdomen och samla in pengar till forskning och till stöd för verksamhet för bröstcancerbehandlade.
I år (17 oktober) anordnas ett seminarium i Europaparlamentet i samarbete med "European Cancer Network".
Meningen är att identifiera grundläggande moment i bröstsjukvårdspersonals yrkesutbildning för framtida EU-riktlinjer.
Karin Jöns (tysk ledamot från socialdemokratiska gruppen) som utarbetade Europaparlamentets resolution om bröstcancer i EU från 2003 förklarar att enligt Världshälsoorganisationen (WHO) kan screening genom mammografiundersökningar minska antalet bröstcancerdödsfall med 35 %.
Det finns motsvarande EU-riktlinjer sedan 1992.
Men fortfarande erbjuder inte 14 av 25 medlemsstater landsomfattande screening.
Under oktober månads plenarsammanträde (23-26 oktober) röstar Europaparlamentet om en ny resolution om bröstcancer.
Förra året i oktober, för att uppmärksamma bröstcancermånaden, lyste Europaparlamentets byggnad i Bryssel rosa, den internationella färgen för kampen mot bröstcancer, för att öka kunskapen om sjukdomen även inom EU:s institutioner.
20061003STO11311 The European Parliamentary Group on Breast Cancer (EPGBC): EP:s resolution om bröstcancer: Bröstcancer: Screeningprogram kan halvera dödlighet (engelska och franska):
SV
1
PHOTO
20061003PHT11309.jpg
SV
2
LINK
http://www.epgbc.org/
-//EP//TEXT TA P5-TA-2003-0270 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20051017BKG01551 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Toomas Hendrik Ilves: Från ledamot till president
Institutioner
2006-10-10 - 11:39
Toomas Hendrik Ilves
Tidigare Europaparlamentsledamoten Toomas Hendrik Ilves är Estlands nya president.
Ilves konstaterar att de nya medlemsländernas synpunkter nu väger tyngre i Europaparlamentet än inledningsvis.
Att göra de nya medlemsstaternas röster hörda var enligt Ilves den största framgången.
"I början togs vi inte på allvar, men nu är jag övertygad om våra synpunkter fullt ut beaktas."
De nya medlemsstaternas svaga samarbete, exempelvis i fråga om tjänstedirektivet som inte är tillräckligt fördelaktigt för länderna, beskriver han som det största misslyckandet.
I fråga om medbeslutandeförfarandet förklarar Ilves att parlamentet nu har ett starkare utgångsläge.
"Men det finns alltid plats för mer.
Europaparlamentet är den första institutionen som representerar Europas medborgare", sade han.
Intresse för utrikesfrågor
Ilves, som är känd för att hellre bära fluga än slips, har arbetat mycket i utskottet för utrikesfrågor och bland annat med frågor som rör Östersjösamarbetet.
Några viktiga oavslutade frågor fick Ilves lämna bakom sig, exempelvis parlamentets yttrande om Rysslands visumregler och återtagandeavtalet.
De estniska rötterna är starka trots många år utomlands.
53-åriga Ilves är född i Sverige, dit hans föräldrar flydde från Estland under andra världskriget.
Skol- och studieåren tillbringade han i USA.
Ilves har en bakgrund som journalist för "Radio Free Europe", och har även varit Estlands USA-ambassadör och utrikesminister under två perioder.
Ilves är inte den första Europaparlamentsledamoten som blir president.
Ytterligare exempel är Frankrikes president Jacques Chirac och Italiens president Giorgio Napolitano.
20061010STO11505 Thomas Hendrik Ilves: Estlands president:
SV
1
PHOTO
20060914PHT10696.jpg
SV
2
LINK
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
115-miljardersfrågan: EU:s budgetprocess
Budget
2006-12-18 - 16:57
Europaparlamentet godkände den 14 december hur EU:s årsbudget för 2007 på 115 miljarder euro kommer att se ut.
Med talmannen Josep Borrells underskrift avslutas den första delen av budgetcykeln.
Men hur bestäms budgeten?
Hur finansieras den och vilka utgifter täcker den?
Läs mer om budgetprocessen i vår uppdaterade budgetfokus.
Den nya långtidsbudgeten för perioden 2007-2013 gäller för ett EU med 27 medlemsstater och dess finansieringsramar omfattar cirka 864,3 miljarder euro.
Inom ramen för den sjuåriga budgetplanen fastställs EU:s budget för varje enskilt år i den årliga budgetprocessen.
Budgeten 2007 uppgår till 115 miljarder euro.
Siffrorna kan tyckas höga men EU:s budget motsvarar endast ungefär 1 procent av EU-ländernas samlade BNI (bruttonationalinkomst).
Den två största utgiftsposten är jordbruksstöd (49 miljarder euro 2005) och strukturfonderna som finansierar EU:s regionalstöd till eftersatta regioner (32 miljarder euro 2005).
Övriga utgiftskategorier är: Inre politik, externa åtgärder, administration, reserver och föranslutningsstöd.
En hög procent av EU:s budget är investeringar snarare än konsumtionsutgifter.
Och till skillnad från statsbudgetar kan inte EU:s budget ha underutskott.
Alla utgifter måste finansieras med unionens inkomster.
20061106FCS12347
En årlig budget inom ramen för en flerårig budgetplan
Men för att effektivisera processen och undvika budgetkriser (som under 1980-talet) enas de båda institutionerna om en långtidsbudget som fastställer utgiftstak.
I december 2005 nådde EU :s medlemsstater en överenskommelse om den nya budgetplanen för 2007-2013.
Den var emellertid inte i linje med kommissionens ursprungliga förslag eller vad parlamentet ansåg nödvändigt för att möta de utmaningar som EU står inför.
En halvtidsöversyn äger rum 2009.
Tillväxt och sysselsättning (382 miljarder euro)
Frihet, säkerhet, rättvisa och medborgarskap (10,77 miljarder euro)
EU som global partner (49,5 miljarder euro)
Hur fattas beslut om budgeten?
Talmannen undertecknar budgetplanen 2007-2013 Europaparlamentet och ministerrådet, som utgör EU:s budgetansvariga myndighet, fattar gemensamt beslut om budgetens utformning och innehåll.
För 2007 års budget ansvarar James Elles (brittisk konservativ ledamot) för att utarbeta förslag till parlamentets position.
I april/maj presenterar kommissionen ett preliminärt budgetförslag.
Första behandlingen
Kommissionens preliminära budgetförslag överlämnas till ministerrådet (EU:s finansministrar) som gör sin första genomgång och antar sin första behandling av budgetförslaget i juli.
Trepartssamtal (parlamentet, kommissionen och rådet) hålls inför varje budgetförhandling för att underlätta en överenskommelse.
Därefter går parlamentet igenom rådets förslag.
I början av oktober har budgetutskottets ledamöter meterhöga staplar med ändringsförslagsdokument att ta ställning till.
Budgetutskottet lägger fram sitt förslag till betänkande för behandling i plenum där hela parlamentet röstar igenom ändringar.
Parlamentet antog sin första behandling av EU:s allmänna budget 2007 den 26 oktober i Strasbourg.
Andra behandlingen
Främst handlar det om utgifter på jordbruksområdet och kostnaderna för vissa avtal med tredje land.
På andra områden, så kallade icke-obligatoriska utgifter har däremot parlamentet sista ordet.
Rådet sänder därefter tillbaka den ändrade budgeten till parlamentet som antar sin andra behandling i december, vilket avslutar den årliga budgetprocessen.
Under 1980-talet, innan överenskommelserna om fleråriga budgetramar infördes, utnyttjade parlamentet vid tre tillfällen sin rätt att avvisa budgetutkastet och begära ett nytt utkast.
2007 års budget
Parlamentet vill öka EU:s budget för 2007.
2007 års budget är den första för EU 27 med och Bulgarien och Rumänien som nya medlemsstater.
Förslaget är mer än 7,4 miljarder euro under den nivå som den fleråriga budgetplanen 2007-2013 tillåter.
I parlamentets första behandling (som antogs den 26 oktober 2006) uppgick betalningarna till 122 miljarder.
Föredraganden Elles sade efter omröstningen: - Parlamentet har antagit en förnuftig, koherent och framåtblickande budget.
Samtidigt har vi låtit oss styras av principen om att man ska få valuta för pengarna.
Europaparlamentet sätter press på kommissionen
Europaparlamentet använde budgetförhandlingarna för att framhäva ett antal viktiga politiska frågor.
Parlamentet begärde exempelvis en gedigen genomgång eller utvärdering av kommissionens faktiska personalbehov.
Vilket kommissionen lovade att göra senast slutet av april 2007.
Vad gäller den gemensamma utrikes- och säkerhetspolitiken (GUSP) uttryckte parlamentet i första behandlingen oro över utökningen av verksamheter inom området "inte har åtföljts av ökad demokratisk ansvars- och redovisningsskyldighet samt granskning från parlamentets sida."
Genom föreslagna budgetändringar strävar parlamentet efter att främja en högre grad av insyn och samarbete i detta hänseende.
Frågan löstes i slutet av november genom en brevväxling mellan rådets ordförandeskap och Europaparlamentet enligt vilket parlamentet ska få information i rätt tid om planerade åtgärder.
Överenskommelse mellan EU-institutionerna
Redan vid det första mötet (21.11.06) kunde parterna nå en överenskommelse och den 14 december (i Strasbourg) kunde Europaparlamentet anta EU:s budget för 2007.
Samma dag undertecknade Europaparlamentets talman Josep Borrell och representanter för rådet och kommissionen budgeten.
EU:s budget 2007 fördelning per rubrik:
1.
Hållbar tillväxt: 44,86 miljarder euro (strukturfonder, forskning och utbildning) 2.
Administration: 6,94 miljarder euro
Den totala budgeten för 2007 är 115,15 miljarder euro i utgifter.
EU:s budget består av utgifter och åtaganden (som har ett större belopp).
Åtagandebemyndiganden är kommissionens utgiftsåtaganden - och motsvarar det belopp som kommissionen kan förbinda sig, utan att nödvändigtvis vara tvungen att betala hela summan under budgetåret.
2007 års budgets åtagandebemyndiganden uppgår till 126,55 miljarder euro.
Vem betalar?
EU:s egna medel 2005 uppgick till 105,684 miljarder euro.
EU-budgetens inkomster är främst det som kallas EU:s egna medel.
Dessa betalas in av medlemsländerna varje år och består av följande kategorier.
Direkta bidrag från medlemsstaterna baserade på bruttonationalinkomst
Jordbrukstullar och avgifter
Andra tullar (handel med tredje land)
Mervärdesskattebaserad avgift
Systemet med egna medel är en överenskommelse mellan medlemsstaterna och har ratificerats av alla nationella parlament.
Det är ett komplicerat system och att nå samsyn mellan medlemsstaterna om EU:s finansiering är sällan en lätt uppgift.
Parlamentet är därför övertygad om att det krävs ett nytt, öppet och mer rättvist system.
Parlamentet har efterlyst en konferens med nationella parlamentet för att se över och ersätta det nuvarande systemet.
Helst senast 2009.
Nettobetalarna
Stor del av importen till EU passerar Antwerpens hamn.
Ofta diskuteras vilka länder som "tjänar" eller "förlorar" på EU-budgeten.
I debatten talas det ofta om "nettobetalare".
Det vill säga om ett land betalar mer till EU än det får tillbaka i form av stöd.
Tyskland, Frankrike, Nederländerna, Storbritannien och Sverige är alla nettobetalare.
Men det är svårt att avgöra hur stora nettobetalningarna faktiskt är.
Exempelvis kan EU bidra med stöd till ett projekt i Frankrike som ett svenskt företag utför.
Ytterligare et exempel är tullavgifter.
Vad händer efter att budgeten godkänts?
EP efterlyser större ansvar på nationell nivå för användningen av EU-medel.
Kommissionen kan också föreslå ändringsbudgetar.
Parlamentet är den EU-institution som kan bevilja ansvarsfrihet för budgetens genomförande.
Beslutet om ansvarsfrihet fattas utifrån rekommendation från rådet och Europeiska revisionsrättens årsrapport.
SV
1
PHOTO
20061109PHT12446.jpg
SV
3
LINK
http://eur-lex.europa.eu/LexUriServ/site/sv/oj/2006/c_139/c_13920060614sv00010017.pdf
SV
6
LINK
http://ec.europa.eu/financial_perspective/index_en.htm
SV
7
PHOTO
20061109PHT12448.jpg
SV
9
LINK
/parliament/public/staticDisplay.do;jsessionid=DAF2A65B704676500366BDE967CC7028.node2?id=46&pageRank=7&language=SV
SV
10
LINK
/activities/expert/committees/presentation.do?committee=1235&language=SV
SV
13
LINK
SV
14
PHOTO
20061109PHT12450.jpg
SV
17
LINK
/comparl/budg/budg2007/2007_en.htm
SV
18
LINK
http://ec.europa.eu/budget/publications/budget_in_fig_en.htm
SV
19
PHOTO
20061109PHT12452.jpg
SV
22
PHOTO
20061109PHT12454.jpg
SV
23
PHOTO
20061109PHT12456.jpg
SV
25
LINK
http://ec.europa.eu/budget/publications/fin_reports_en.htm
-//EP//TEXT IM-PRESS 20060517STO08359 0 NOT XML V0//SV
-//EP//TEXT TA P6-TA-2006-0210 0 NOT XML V0//SV
-//EP//TEXT TA P6-TA-2005-0224 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061020IPR11896 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061020IPR11896 0 NOT XML V0//SV
-//EP//TEXT REPORT A6-2006-0223 0 NOT XML V0//SV
-//EP//TEXT TA P6-TA-2005-0224 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061011STO11555 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 FCS DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 FCS DOC XML V0//EN
Tjänstedirektivets sista tappning återspeglar parlamentets ståndpunkt
Fri rörlighet för tjänster
2006-11-15 - 14:03
Den slutgiltiga texten återspeglar nästan fullständigt parlamentets krav från första behandlingen och innebär en balans mellan konkurrens och sociala hänsyn.
Medlemsstaterna har tre år på sig att genomföra direktivet.
Endast tre ändringsförslag som rörde en teknisk anpassning antogs.
Två förslag om att helt förkasta den gemensamma ståndpunkten som lagts fram av grupperna De Gröna och GUE/NGL föll.
På presskonferensen efter omröstningen framhöll Europaparlamentets talman Josep BORRELL omröstningsresultatet som "en stor framgång för parlamentet som lagstiftare".
Borrell betonade vikten av det beslut parlamentet fattat som bidragit till att man "fått till stånd en välavvägd lagstiftningstext med brett stöd".
Tjänstesektorn generar nästan 70 % av BNP och sysselsättningen i EU.
Efter två års arbete antog Europaparlamentet i februari 2006 med bred majoritet den kompromiss som rådets ståndpunkt i allt väsentligt grundar sig på.
Kompromissen gällde bl.a. den övergripande målsättningen med direktivet (artikel 1), direktivets räckvidd (artikel 2) och bestämmelser för fritt tillhandahållande av tjänster (artikel 16, där kommissionen först mycket kontroversiellt föreslog att reglerna i ursprungslandet skulle gälla).
Rådet bedöms att till 90 procent ha respekterat parlamentets krav från första behandlingen.
Direktivets syfte (artikel 1)
Direktivet inrättar en rättslig ram för att avskaffa hindren för tjänstetillhandahållares fria etablering och fri rörlighet för tjänster mellan medlemsstaterna.
Det föreskriver administrativ förenkling, i synnerhet inrättande av gemensamma kontaktpunkter där tillhandahållarna av tjänsterna kan fullgöra de administrativa förfaranden som rör verksamheten och krav på att detta ska kunna göras på elektronisk väg, samt förenklat tillståndssystem för tjänsteverksamhet.
Samtidigt ska tjänsternas höga kvalitetsnivå garanteras.
Direktivet behandlar inte liberaliseringen av tjänster av allmänt ekonomiskt intresse som är förbehållna offentliga eller privata enheter, och inte heller privatiseringen av offentliga enheter som tillhandahåller tjänster.
Genom direktivet avskaffas inte heller monopol för tillhandahållande av tjänster eller statligt stöd från medlemsstater vilket omfattas av gemenskapens konkurrensregler.
Medlemsstaterna får själva definiera vad de anser vara tjänster av allmänt ekonomiskt intresse, hur dessa tjänster bör organiseras och finansieras i enlighet med bestämmelser om statligt stöd.
De påverkar inte heller medlemsstaternas lagstiftning om social trygghet.
Rätten att förhandla om, ingå och tillämpa kollektivavtal samt att vidta stridsåtgärder i enlighet med nationell lagstiftning och praxis påverkas inte heller.
Det skulle även ha varit ursprungslandets ansvar att kontrollera att dess gällande bestämmelser efterlevdes där tjänsterna utfördes.
Många medlemsstater och ledamöter fann detta orealistiskt och den kontroversiella artikeln ändrades därför av parlamentet och rådet har helt gått på parlamentets linje i fråga om "Frihet att tillhandahålla tjänster " som principen nu betecknas.
Enligt den nuvarande skrivningen ska medlemsstaterna respektera tjänsteleverantörernas rätt att tillhandahålla tjänster i en annan medlemsstat än den där de är etablerade.
Eventuella krav på tillstånd för tillträde till eller utövande av en tjänsteverksamhet på ett lands territorium måste vara icke diskriminerande ifråga om nationalitet eller, för juridiska personer, etableringsmedlemsstat, nödvändiga, d.v.s. motiverade med skäl som avser allmän ordning, allmän säkerhet, folkhälsa eller miljöskydd och proportionerliga.
Möjlighet att tillämpa särskilda nationella bestämmelser finns då "tvingande hänsyn till allmänintresset" föreligger.
Parlamentet lade till detta med stöd i domstolens rättspraxis.
Tjänster som omfattas av direktivet är företagsrelaterade tjänster, såsom konsulttjänster inom ledarskap och förvaltning, certifiering och testning, viss typ av fastighetsservice ("facilities management"), inklusive kontorsunderhåll och annan kontorsservice, reklam, rekryteringstjänster samt handelsagenter.
Icke ekonomiska tjänster av allmänt intresse.
- Finansiella tjänster såsom banktjänster och tjänster som avser krediter, försäkringar och återförsäkringar, tjänstepensioner och individuellt pensionssparande, värdepapper, investeringsfonder, betalningar och investeringsrådgivning.
- Elektroniska kommunikationstjänster och kommunikationsnät.
- Transporttjänster, inklusive lokaltrafik, taxi och ambulanser samt hamntjänster.
- Tjänster som tillhandahålls av bemanningsföretag.
- Hälso- och sjukvårdstjänster, oavsett om de tillhandahålls via sjukvårdsinrättningar eller inte, och oavsett hur de är organiserade och finansierade på nationell nivå eller om de är offentliga eller privata.
- Audiovisuella tjänster.
- Spelverksamhet, t.ex. lotterier, kasinospel och vadslagningar.
- Verksamhet som har samband med utövandet av offentlig makt.
- Sociala tjänster som rör subventionerat boende, barnomsorg och stöd till permanent eller tillfälligt behövande familjer och enskilda som tillhandahålls av staten, tjänsteleverantörer på uppdrag av staten eller av staten erkända välgörenhetsorganisationer.
- Privata säkerhetstjänster.
- Tjänster som tillhandahålls av officiellt utnämnda notarier och utmätningsmän.
Direktivet ska inte heller tillämpas på skatteområdet.
För att underlätta tillhandahållandet av tjänster åläggs medlemsstaterna att granska de förfaranden och formaliteter som är tillämpliga på tillträde till och utövande av en tjänsteverksamhet i syfte att förenkla dem.
Medlemsstaterna har tre år på sig att sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa direktivet sedan dagen efter att det offentliggjorts i Europeiska unionens officiella tidning.
Kommissionen ska fem år efter det att direktivet trätt i kraft och därefter vart tredje år lägga fram en övergripande rapport om tillämpningen av direktivet.
Evelyne GEBHARDT (PSE, DE) inledde med att tacka för all den konstruktiva hjälp hon fått från kollegor och nämnde särskilt sin skuggföredragande Malcolm HARBOUR (EPP-ED, UK).
Den kontroversiella principen om ursprungsland är helt struken, liksom de tidigare artiklarna 24 och 25, så att inte utstationeringsdirektivet ifrågasätts av det nya direktivet.
Direktivet rör kommersiella tjänster, fortsatte hon och betonade att merparten sociala tjänster därför inte berörs.
Enligt Gebhardt kommer alla tjänsteföretagen gagnas betydligt av direktivet och rörligheten kommer definitivt att underlättas genom friheten att tillhandahålla tjänster och den fria etableringsrätten som nu förbättras genom förenklade administrativa förfaranden, en gemensam kontaktpunkt o.s.v.
Gebhardt avslutade med att säga att hon nu förväntade sig en rad förtydliganden från kommissionen om arbetsrätten, sociala rättigheter straffrätten och om kommissionen riktlinjer till medlemsstaterna när det gäller vissa nationella bestämmelser.
Charlie MCCREEVY, med ansvar för den inre marknaden, talade om en milstolpe i EU:s och Europaparlamentets historia.
- Direktivet är viktigt för såväl konsumenter, arbetstagare och näringsliv.
Det behövs för den europeiska ekonomin och här har parlamentet gjort ett mycket viktigt arbete, sade McCreevy.
Samtidigt har medlemsstaterna fortfarande rätt att ställa krav med hänsyn till tvingande intressen.
De måste dock garantera friheten att tillhandahålla tjänster och den fria etableringsrätten.
Det var värre i rådet att få alla med.
McCreevy betonade att det är en mycket bräcklig kompromiss och en ny debatt i rådet vore ytterst riskabelt.
Parlamentet bör avstå från ändringar, endast de tre tekniska ändringsförslagen om kommittéförfarandet kan godkännas.
McCreevy avslutade med att göra de efterfrågade klargörandena.
Han sade att när det gäller översynen av de nationella krav som medlemsstaterna uppställer och hur dessa eventuellt ska ändras ska kommissionen företa en granskning, en "screening".
Detta tillkomer EG-domstolen.
Inga ändringar kan heller göras i direktivet utan parlamentets och rådets deltagande.
Om ytterligare åtgärder krävs på sikt inom vissa områden, eller om harmonisering behövs kommer parlamentet att göras delaktigt.
När det gäller arbetsrätten påminde kommissionären om att både parlamentet och rådet ville undanta denna.
Tjänstedirektivet påverkar alltså inte arbetsrätten och inte de kollektiva rättigheter som förhandlas fram av arbetsmarknadens parter enligt nationell praxis, med respekt för bestämmelserna i fördragen och annan EU-lagstiftning.
Straffrätten påverkas inte som sådan, däremot berörs utländska tjänsteleverantörer liksom alla andra av gällande nationella bestämmelser.
Men straffrätten får inte missbrukas för att kringgå bestämmelserna i direktivet.
De berörs därför inte.
Rådet
Finlands handels- och industriminister, Mauri PEKKARINEN, hänvisade till parlamentets historiska kompromiss i våras utan vilken man inte befunnit sig där man står idag.
Han påminde att det rörde sig om nästan tre års arbete och att sex ordförandeskap varit inblandade.
Föredragandens reaktion
GEBHARDT ansåg att kommissionens gjort nödvändiga förtydliganden och uppmanade därför kammaren att godkänna den gemensamma ståndpunkten och endast göra de tekniska tillägg som de tre ändringsförslagen om kommittéförfarandet innebär.
Gebhardt tog sedan tillfället i akt för att kritisera rådet för att det flera gånger hotat med den bräckliga kompromissen.
Det kommer att skapas ett större tjänsteutbud, men med bibehållna konsumenträttigheter.
Harbour betonade att det rörde sig om ett väldigt detaljerat direktiv med ett 40-tal åtgärder för att undanröja onödiga hinder och mer än 60 bestämmelser för att förenkla administrativa förfaranden.
Han tackade Gebhardt för att hon drivits av en stark övertygelse om behovet av detta direktiv och han nämnde också det samarbete som funnits med liberalerna och med det brittiska förbundet för små och medelstora företag.
Han beklagade den protektionism och nationalism som verkar florera och sade att EU:s ledare måste förklara innebörden av den inre marknaden för medborgarna, göra den begriplig.
Jäätteenmäki beklagade att rumänska och bulgariska medborgarna nu drabbas av samma restriktioner som de tio andra nya länderna vid utvidgningen 2004.
Om tjänstedirektivet nu utgör ett steg framåt innebär dessa restriktioner tyvärr ett steg tillbaka för den inre marknaden och den fria rörligheten för arbetstagare.
Hon hänvisade till vad Harbour sagt om att sociala tjänster inte omfattas, men påpekade att dessa definieras mycket olika i olika länder.
Detta kommer att skapa problem.
Hon betonade också att kommissionens förklaringar endast är bindande för den sittande kommissionen.
Wurtz varnade för gråzoner i texten och menade ett det blir domstolen som kommer att få avgöra.
Tjänster av allmänt intresse utesluts, men tjänster av allmänt ekonomiskt intresse omfattas och detta är känsligt.
Direktivet måste vara tydligare!
Romfördraget är snart femtio år och vi måste visa att vi värnar om våra medborgare, sade han avslutningsvis.
Adam Jerzy BIELAN (UEN, PL) sade att 70 % av unionens BNP genereras av tjänstesektorn, men tusentals byråkratiska hinder hämmar marknaden.
Han sade att han välkomnar arbetstagare och tillhandahållare av tjänster i Danmark, men sade att de måste ges danska löner för att undvika social dumpning.
Marine LE PEN (NI, FR) sade att EU avreglerar tjänster på ett farligt sätt och att vissa sociala tjänster omfattas.
Junilistan är emot nationell protektionism, byråkrati och skråväsendets kvarlevor i Europa.
Sådana restriktioner hindrar konkurrens, utveckling och tillväxt inom tjänstesektorn.
Junilistan välkomnar att rådet i likhet med parlamentet valde att förkasta ursprungslandsprincipen.
Den hade förvisso möjliggjort ökad konkurrens inom några tjänstesektorer, men nackdelarna var orimligt stora.
Ursprungslandsprincipen skulle ha tvingat medlemsländerna att ge upp nationellt självbestämmande på några av de viktigaste områdena av samhällslivet.
Det är självklart att de lagar, regler och traditioner som gäller på ett lands territorium har tillkommit i demokratisk ordning och måste följas av alla som verkar på dess territorium.
Junilistan välkomnar således rådets gemensamma ståndpunkt om tjänstedirektivet.
Jan ANDERSSON (PSE, SE) koncentrerade sig på arbetsrätten.
Även om han föredrog skrivningen i Europaparlamentets första behandling var han fullt nöjd med det som kvarstår.
Innebörden stärks dessutom av det McCreevy sade under debatten.
Charlotte CEDERSCHIÖLD (EPP-ED, SE) sade att Europaparlamentet idag tog ett stort principiellt steg, men påminde om att hon ansåg att direktivets starkaste livräddare varit EPP-ED och ALDE.
- Den nya svenska regeringen verkar för att göra det mer lönsamt att arbeta och den kommer att få bättre möjligheter att lyckas genom direktivet.
Kommissionär Charlie MCCREEVY sade att man nu måste börja inrikta sig på tillämpningen.
Medlemsstaterna har tre år på sig att genomföra direktivet.
Rådet
Betänkande: A6-0375/2006
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
EU:s nya kemikalielagstiftning Reach nu i hamn
Miljö
2006-12-13 - 13:22
Parlamentets omröstning idag innebär att Reach kan börja tillämpas den 1 juni 2007.
Registreringsprocessen kommer att ta 11 år eftersom omkring 30 000 ämnen berörs.
Kompromisspaketet antogs med 529 röster för, 98 emot och 24 nedlagda.
Enligt Europaparlamentets talman Josep Borrell "innebär Reach en lagstiftning som är av avgörande betydelse för folkhälsan och miljön i EU.
- Att inrätta ett enhetligt registreringssystem som utformats för att lämna grundinformation om farorna och riskerna med nya och befintliga ämnen som tillverkas i eller importeras till EU i mer än 1 ton.
- Att införa skyldighet att lämna information om användning och tillhörande riskhanteringsåtgärder avseende ämnena.
- Att upprätthålla det befintliga begränsningssystemet och införa ett tillståndsförfarande för de farligaste ämnena som ett nytt instrument.
- Att upprätta en central enhet för att underlätta förvaltningen av Reach och se till att systemet tillämpas på ett harmoniserat sätt i hela EU.
- En kemikaliemyndighet inrättas också.
Ytterst är det Europeiska kommissionen som beviljar de tillstånd som krävs för särskilt farliga ämnen.
Parlamentet kämpade in i det sista för att de allra farligaste ämnena ska ersättas, för att företagen ska tillämpa försiktighetsprincipen och för att minimera antalet djurförsök.
Parlamentet har nu ställt sig bakom den kompromiss som träffades med rådet den 30 november.
Sex år gäller för de ämnen som överskrider 100 ton och elva år för dem som överskrider 1 ton.
Principen om att dela information utökades till alla tester, inte bara djurförsök.
Parlamentet uppnådde att tillstånd ska vara tidsbegränsade och att när det gäller de farligaste substanserna måste en substitutionsplan finnas om tillstånd ska beviljas.
Om inga bättre alternativ finns att tillgå måste en forsknings- och utvecklingsplan tas fram av tillverkaren för att försöka hitta en ersättning.
Alternativa testmetoder ska godkännas av kommissionen så snart dessa erkänts av Kemikaliemyndigheten eller av behöriga internationella organisationer.
Kommissionen åläggs också att försöka inrätta en EU-kvalitetsmärkning för kemiska produkter.
Kemikaliemyndigheten .
Europaparlamentet ska utse två av medlemmarna i kemikaliemyndighetens styrelse som således ska bestå av en representant från varje medlemsstat och högst sex representanter som utses av kommissionen och två representanter som utses av Europaparlamentet.
Direktören kommer att höras av Europaparlamentet innan utnämningen godkänns.
Skyddet av immaterialrätten har stärkts och skyddet av dataskyddet förlängs från 3 år till 6 år.
Kemikalieinspektionens styrelse bör inte kunna vara hemlig och ha hemliga finansiella intressen.
- Reach borde nu byta namn till Risk, registrering men icke-substitution av kemikalier.
Schlyter förordade en ny kompromiss med rådet och uppmanade föredraganden Sacconi att gå vidare.
Lena Ek (ALDE/ADLE, SE) sade att hon hade mycket blandade känslor.
Det är viktigt att klargöra.
Avslutningsvis sade hon att u-länderna måste ges möjlighet att använda den samlade informationen, så att det inte skapas handelshinder för dem.
Akut metallförgiftning, sade doktorn att det var.
Det finns ingen rättsligt bindande ansvarsprincip och storföretagen kan fortsätta att hemlighålla sina fakta om kemikalier när EPP-ED fått igenom sina krav på stärkt immaterialrätt.
Denna princip, som säger att farliga kemikalier ska ersättas när det finns mindre farliga alternativ, är nu så begränsad att det är endast ett ytterst fåtal kemikalier som kommer att fasas ut.
För att minimera djurförsöken kräver vi också satsningar på helt nya djurfria metoder med ”toxygenomics”.
De stora partigrupperna har dock valt att vika sig inför rådet genom att godta den usla kompromiss som ligger på bordet, sade hon.
Hon kände sig överraskad över att den socialistiska gruppen valde att stödja kompromissen.
Mer substitution, mer information och datasäkerhetsblad för lågvolymkemikalier och fler kemikalier som borde registreras.
Den är det bästa vi kan få och innebär mycket bättre regler än de kemikalieregler som finns i Sverige och EU idag.
- Vi svenska socialdemokrater kommer att ta vårt ansvar och rösta för kompromissen.
Betänkande: A6-0352/2006 och A6-0345/2006
20061213IPR01493
SV
1
PHOTO
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
Föredragningslista - senaste utgåva
Måndagen den 18 december 2006
11:00 - 13:00 Gemensam debatt
Europeiska rådet / det finländska ordförandeskapet
Rapport från Europeiska rådet och uttalande av kommissionen
Europeiska rådets möte den 14 och 15 december 2006
Uttalande av rådets tjänstgörande ordförande
Arbetet under det gångna halvåret under det finländska ordförandeskapet
Slut på den gemensamma debatten
EU-debatt med tyska ungdomar
Institutioner
2006-12-20 - 18:12
Har utvidgningen försvagat EU?
Är EU en motpol till USA?
Och varför prioriteras inte utbildning i budgeten?
"Vi har byggt Europa för er, för den unga generationen.
Vi vill höra era förväntningar på EU-integrationen", sade Europaparlamentets talman Josep Borrell i samband med forumets öppnande.
Norbert Lammert tyska förbundsdagens talman sade: "EU:s framtid påverkar oss alla, men den påverkar särskilt den unga generationen."
Ledamöternas svar begränsades till 1,5 minuter.
Hans-Gert Pöttering (Gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater) underströk att EU:s förhållande till USA bygger på "vänskap och partnerskap", men han betonade samtidigt att "vi också måste säga ifrån, om vi inte håller med i vissa frågor, exempelvis om Guantanamo."
Martin Schulz (Socialdemokratiska gruppen i Europaparlamentet) betonade behovet att "stärka multilateralismen".
Han sade att kriget i Irak har lett till en "katastrof".
Och att Europa har ett ansvar för Irak och särskilt för det irakiska folket.
En student undrade om det inte kommer att bli ännu svårare med en EU-armé?
Jens-Peter Bonde (Gruppen Självständighet/Demokrati) höll absolut inte med, och sade: "Vi ska föra krig mot fattigdom."
Sylvia-Yvonne Kaufmann (Gruppen Europeiska enade vänstern/Nordisk grön vänster) menade att Europa måste "titta närmare på orsakerna för konflikter och ta itu med dessa.
Det är alltför enkelt att bara sända militärstyrkor."
Utvidgningen
De unga deltagarna var också nyfikna på utvidgningen och om den senaste stora utvidgningsrundan inte övergick EU:s förmåga.
Alla ledamöter underströk fördelarna av ett enat Europa.
Irena Belohorska ledamot från Slovakien som anslöt 2004 betonade att hon helt enkelt är "glad att vi idag är en del av denna gemenskap.
Vi var tvungna att vänta så länge."
Andra frågor som togs upp var den sociala modellen och ett åldrande EU:s ekonomiska utmaningar.
Det kan bli en fråga för Tyskland som den 1 januari tar över EU:s roterande sexmånadersordförandeskap.
Ungdomsforumet organiserades av Europaparlamentets informationskontor i Berlin tillsammans med det tyska parlamentet.
20061220STO01665
SV
1
PHOTO
20061220PHT01681.jpg
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
HÖJDPUNKTER 2004-2006
Institutioner
Sverige
2007-01-12 - 14:23
En översikt över Europaparlamentets verksamhet efter halva lagstiftningsperioden
INTRODUKTION
I januari 2007 är första hälften av Europaparlamentets innevarande lagstiftningsperiod till ända.
En ny talman och nya vice talmän ska väljas för den andra hälften liksom nya utskottsordförande.
Från den 1 januari 2007 då Bulgarien och Rumänien ansluter sig till EU ökar antalet ledamöter tillfälligt till 785 eftersom 35 nya rumänska ledamöter och 18 nya bulgariska ledamöter tillträder.
Från den 1 januari 2007 tillkommer tre nya språk bulgariska, rumänska och iriska.
Europaparlamentets presstjänst vill i detta sammanhang framhålla en rad höjdpunkter under den första perioden.
Sammanställningarna består dels av fullständiga artiklar på engelska och franska, dels av ett urval redan publicerade pressmeddelanden på svenska med länkar till den fullständiga texten.
20061221BKG01704
Fri rörlighet för tjänster
Tjänstedirektivets sista tappning återspeglar parlamentets ståndpunkt
Den slutgiltiga texten återspeglar nästan fullständigt parlamentets krav från första behandlingen och innebär en balans mellan konkurrens och sociala hänsyn.
Medlemsstaterna har tre år på sig att genomföra direktivet.
Television - inget förbud mot barn- och alkoholreklam
Parlamentet stödde vid sin första behandling kommissionens föreslagna modernisering av EU-bestämmelser om sändningsverksamhet för television.
Det rör sig om en uppdatering av direktivet Television utan gränser från 1989.
Parlamentet röstade för att även nya digitala audiovisuella tjänster ska omfattas.
Reklam kommer att få visas var 30:e minut och produktplacering tillåts i hela EU på gemensamma villkor.
Europaparlamentet förkastar mjukvarupatentet
Ledamöterna röstade med 648 röster för, 14 röster emot och 18 nedlagda röster, för ett förkastande av rådets gemensamma ståndpunkt.
Parlamentets förkastande innebär att lagstiftningsförfarandet avslutades.
Rådande praxis vid Europeiska patentverket och nationella patentverket kommer därmed fortsatt att gälla
Miljö
EU:s nya kemikalielagstiftning Reach nu i hamn
Europaparlamentet antog den 13 december 2006 en andrabehandlingskompromiss om Reach (registrering, utvärdering, godkännande och begränsning av kemikalier).
I juni 2007 inleds därmed registreringen av alla kemiska ämnen som produceras eller importeras i mer än ett ton per företag och år i EU.
För farliga ämnen måste en substitutionsplan tas fram och för de ämnen för vilka det för närvarande inte finns några alternativ måste en utvecklingsplan presenteras i syfte att försöka ersätta ämnet.
Registreringsprocessen kommer att ta 11 år eftersom omkring 30 000 ämnen berörs.
Man räknar med att ha avslutat till 2018.
Tillståndsförfarandet rör endast de bortåt 3 000 ämnen som bedöms vara särskilt farliga.
EU började riskbedöma nya ämnen först 1981.
Sedan dess har cirka 3 000 nya ämnen tillkommit.
För ämnen vars tillverkning inleddes före 1981 behövdes ingen bedömning.
Totalt handlar det om mer än 100 000 olika ämnen på EU-marknaden.
För 99 % av dessa saknar industrin och samhället tillräckliga kunskaper om riskerna och effekterna på miljö och hälsa.
Mindre fluorerade växthusgaser i atmosfären
Grundvatten - skärpta normer
Ledamöterna lyckades uppnå strängare normer och regler för att förhindra att grundvattnet förorenas i syfte att bättre skydda denna värdefulla dricksvattenskälla.
Insamling av batterier och ackumulatorer systematiseras i EU från 2008
Efter två års förhandlingar godkände parlamentet ett direktiv som innebär att det till 2008 i hela EU ska finnas system för insamling av använda batterier och ackumulatorer.
Hittills har bara sex medlemsstater, däribland Sverige, infört sådana system.
Renare luft genom ambitiösare mål och större flexibilitet
Luftföroreningar utgör en allvarlig sjukdomsfaktor och leder till ett stort antal förtida dödsfall i EU.
Europaparlamentet kräver därför ambitiösare mål för renare luft i Europa.
Samtidigt förespråkas större flexibilitet och mer tid för medlemsstaterna att vidta nödvändiga åtgärder så att fastställda mål verkligen uppnås.
Rent badvatten i sikte
Idag riskerar 12 badare av 100 att drabbas av t.ex. magsjukdomar eller andningsproblem.
I ett direktiv från 1976 finns 19 parametrar för vattenanalys vilka nu minskats ner till endast två i det nya direktiv som parlamentet antagit.
Parlamentet och rådet har ansträngt sig för att nå en balans mellan hälsoaspekter och rimliga administrativa och ekonomiska bördor kring kontrollen av kvaliteten.
Allmänheten ska ha tillgång till aktuell information, både på badplatsen och på Internet.
Översvämningsrisker - ledamöterna kräver samordning i EU
Med tanke på att nästan 80 % av de europeiska floderna och kusterna löper längs eller genom flera länder, yrkar ledamöterna på att EU-länderna på ett bättre sätt samordnar hanteringen av översvämningar.
Genom det betänkande som antagits om Europaparlamentets och rådets direktiv om bedömning och hantering av översvämningar vill parlamentet inrikta arbetet på riskförebyggande åtgärder.
Transport
Parlamentet stärker funktionshindrade personers rättigheter i samband med flygresor
Funktionshindrades rättigheter i samband med flygresor stärks tack vare bestämmelser i en förordning som godkänts av Europaparlamentet.
Föredragande Robert Evans (PSE, GB) Medbeslutande 1:a behandlingen
Europaparlamentet har antagit rådets gemensamma ståndpunkt.
För närvarande finns 110 olika modeller för körkort i EU, som successivt kommer att ersättas.
Den slutgiltiga texten återspeglar på ett balanserat sätt de olika traditioner och erfarenheter som finns i EU.
Föredragande: Mathieu GROSCH (EPP-ED, BE) Medbeslutande - 2:a behandlingen Omröstning: 14.12.2006
154 miljoner euro för att bekämpa föroreningar till havs
Europaparlamentet stöder kommissionens förslag om en finansieringsram på 154 miljoner euro för 2007–2013 för Europeiska sjösäkerhetsbyråns åtgärder mot föroreningar från fartyg.
Anslagen kommer att göra det möjligt för sjösäkerhetsbyrån, som blir operativ från den 14 september, att tillhandahålla medlemsstaterna fartyg för sanering och ta fram satellitbilder för att identifiera och lokalisera utsläpp.
Parlamentet vill att alla former av föroreningar omfattas och inte bara olja.
Parlamentet förkastar förslaget till hamndirektiv
Flertalet ledamöter sade sig föredra bestämmelser om bättre insyn och rättvis konkurrens mellan hamnarna.
Att kontroversiella frågor från kommissionens första förslag till hamndirektiv - exempelvis egenhantering och lotstjänster - fanns kvar i det nya förslaget väckte kritik.
I november 2003 förkastade parlamentet ett tidigare förslag till hamndirektiv.
Parlamentet kräver en översyn av centrala frågor som insyn i fråga om statsstöd och annat stöd till hamnar och rättvis konkurrens mellan hamnar.
Parlamentet och berörda inom sektorn ska delta i översynen.
En gemensam svart lista över osäkra flygbolag
Europaparlamentet stöder att en europeisk svart lista över flygbolag som brister i säkerhetskrav införs och att flygbolag som inte möter säkerhetskraven förbjuds inom EU.
Dessutom vill Europaparlamentet att flygresenärernas rätt till information om flygbolagens identitet ska stärkas.
Passagerare ska också ha rätt till ersättning om ett flygbolag förs upp på listan efter biljettreservation.
Föredragande: Christine De Veyrac (EPP-ED, FR), Medbeslutande 1:a behandlingen Omröstning: 17.11.2005
Hälsa och konsumentpolitik
EP skärper reglerna för närings- och hälsopåståenden om livsmedel - reglerna skärps
Europaparlamentet har godkänt skärpta bestämmelser för närings- och hälsopåståenden om livsmedel.
Ledamöterna vill ha tydliga definitioner för begrepp som lågt energivärde, låg fetthalt eller fiberrik.
Gemensamma bestämmelser för tillsättning av vitaminer och mineraler har också godkänts för att förbättra konsumentinformationen samtidigt som man underlättar för varors rörlighet på den inre marknaden.
Förordningen omfattar näringspåståenden och hälsopåståenden som används på märkning, presentation och i reklam för livsmedel.
Den största stötestenen har varit livsmedlens "näringsprofiler".
Incitament för läkemedelsföretagen att utveckla mediciner för barn
Genom dagens omröstning stimuleras läkemedelsföretag genom en förordning att ta fram medicin för barn.
Barn ska inte längre bara ges mindre doser av läkemedel för vuxna eftersom de kan var olämpliga eller t.o.m. skadliga för barns ämnesomsättning och utveckling.
Läkemedelsföretag som utvecklar effektiva och säkra test för barnläkemedel kommer att belönas med ett 6-månaders tilläggsskydd för sitt patent.
Endast företag som uppfyller mycket strikta normer kommer att ges tillstånd att sälja läkemedel för barn.
Europaparlamentet stöder ett utvidgat förbud mot ftalater i leksaker och barnvårdsartiklar.
De nya bestämmelserna innebär att tre ftalater - DEHP, DBP och BBP*- förbjuds i alla leksaker och barnvårdsartiklar om koncentrationen är över 0,1 %.
Detta kan jämföras med situationen före 1999 då det inte var ovanligt att upp till 30 % ibland förekom i vissa artiklar.
Också en andra kategori - DINP, DIDP och DNOP* - förbjuds, i samma koncentration, i leksaker och barnavårdsartiklar som kan stoppas i munnen, även utan att vara avsedda för detta.
Finansiering av program
Budgetplanen för 2007-2013 formellt godkänd av parlamentet
Kommissionen inledde förberedelserna för den nya budgetplanen och det nya interinstitutionella avtalet genom att lägga fram ett första förslag i februari 2004.
Parlamentet tillsatte i september 2004 ett tillfälligt utskott för politiska utmaningar och budgetmedel i ett utvidgat EU 2007–2013 med uppgift att fastställa parlamentets prioriteringar, föreslå en struktur för presentationen av den kommande budgetplanen, samt försöka beräkna de nödvändiga resurserna under respektive utgiftskategori för perioden 2007-2013.
Denna förkastades av parlamentet eftersom den inte ansågs kunna ge EU de kvantitativa och kvalitativa medel som behövs för att möta framtida utmaningar.
Föredragande: Reimer BÖGE (EPP-ED, DE) Budget Omröstning: 17.5.2006
Sjunde ramprogrammet för forskning 2007-2013
Den övergripande budgeten för det sjunde ramprogrammet uppgår till 54,582 miljarder euro i löpande priser för perioden 2007-2013.
Av dessa anslås 50,751 miljarder för den Europeiska gemenskapens program och 2 751 miljoner för Euratom-programmet som löper mellan 2007-2011.
Detta utgör EU:s tredje största budgetpost efter den gemensamma jordbrukspolitiken och strukturfonderna.
Programmet träder i kraft den 1 januari 2007.
Flera av parlamentets prioriteringar fick gehör under ärendets gång och bl.a. har små och medelstora företags deltagande underlättats på flera sätt genom parlamentets ändringar.
Föredragande: Jerzy BUZEK (EPP-ED, PL) Medbeslutande - 2:a behandlingen Omröstning: 30.11.2006
Rådet och parlamentet har enats om budgeten och innehållet i programmen så ärendena kunde slutföras genom denna andra behandling av parlamentet.
Programmen kan därmed börja användas den 1 januari 2007.
Föredragande: Hannu TAKKULA (ALDE, FI), Ruth HIERONYMI (EPP-ED, DE), Lissy GRÖNER (PSE, DE) Vasco GRAÇA MOURA (EPP-ED, PT) Doris PACK (EPP-ED, DE) Medbeslutande - 2:a behandlingen Omröstning: 25.10.2006
Parlamentet stöder EU:s strukturpaket på 308 miljarder euro för 2007-2013
Genom att anta fem betänkanden har Europaparlamentet godkänt de rättsliga grunderna för EU:s kommande paket med strukturfonder för perioden 2007-2013.
Förordningarna utgör gemenskapens rättsliga ramverk för att genomföra sin sammanhållningspolitik under perioden 2007-2013.
Strukturfonderna syftar till att öka solidariteten mellan EU:s olika regioner.
Medborgerliga fri- och rättigheter
Har europeiska flygplaster använts för transit av fångar som förts till hemliga läger där de riskerar att utsättas för tortyr?
Detta är de två viktigaste frågorna för det nya tillfälliga utskott som Europaparlamentet har beslutat att inrätta.
De 46 ledamöterna från de olika politiska grupperna ska också undersöka om några europeiska regeringar varit inblandade i den påstådda hanteringen av fångar.
Tre svenska ledamöter ska delta i utredningen - Anders Wijkman (EPP-ED), Inger Segelström (ESP) och Cecilia Malmström (ALDE) - bland de totalt 46 ledamöterna .
En mer samordnad invandringspolitik efterlyses
Ledamöterna anser vidare att jourtid i de flesta fall ska gälla som arbetstid.
Utstationering av arbetstagare - förtydliganden och bättre tillämpning behövs
För närvarande krävs inga ändringar av själva direktivet.
Föredragande: Elisabeth SCHROEDTER (De gröna/EFA, DE) Initiativbetänkande Omröstning: 26.10.2006
Institutionella frågor och utvidgningen
Val av kommissionen
Den nye ordföranden José Manuel Barroso fick tillsammans med rådet göra vissa förändringar i sammansättningen innan ledamöterna slutligen i mitten på november kunde godkänna den nya kommissionen i dess helhet.
Europaparlamentets ledamotsstadga
Europaparlamentet har antagit ett betänkande om en gemensam stadga för Europaparlamentets ledamöter (röstsiffrorna: 403 för, 89 emot och 92 nedlagda röster).
Betänkandet stöder rådets kompromiss som bl.a. innebär att ledamöternas arvode ska uppgå till 38,5 procent av grundlönen för en domare vid EG-domstolen (dvs. ungefär 7 000 euro i månaden före skatt).
På så sätt upphör skillnaden mellan ledamöterna, idag får de ett grundarvode som motsvarar det som ledamöterna i de nationella parlamenten har.
Ett klart och motiverat ja till konstitutionen för Europa
Parlamentet hoppas på dess snara ratificering.
Betänkandet är tänkt som ett bidrag i informationskampanjen om fördraget och framhåller fördelarna jämfört med tidigare fördrag.
En konstitution behövs senast 2009
Europaparlamentet vill att en ny konstitution ska finnas till 2009 så att EU även fortsättningsvis ska kunna fungera demokratiskt och rationellt.
Ett annat viktigt budskap i det initiativbetänkande som antagits är att EU, efter Bulgariens och Rumäniens anslutningar, inte bör kunna utvidgas ytterligare utan en översyn av de konstitutionella aspekterna.
Nicefördraget måste alltså ersättas på ett eller annat sätt.
Frågan är hur.
Ja till Bulgariens och Rumäniens begäran om anslutning till EU
Parlamentet gav den 13 april 2005 sitt formella samtycke till Rumäniens och Bulgariens anslutning till EU.
Rumäniens begäran om anslutning till EU erhöll 497 röster för, 93 emot och 71 nedlagda, medan Bulgariens begäran fick 522 röster för, 70 emot och 69 nedlagda röster.
Turkiet - förhandlingar bör inledas men utan garantier om medlemskap
EU bör utan onödigt dröjsmål inleda förhandlingar med Turkiet.
Två dagar före stats- och regeringschefernas toppmöte den 17 december 2004, då det formella beslutet i frågan ska fattas, antog parlamentet en resolution som framhåller Turkiets imponerande framsteg när det gäller uppfyllandet av de politiska Köpenhamnskriterierna.
Framstegen bedöms tillräckliga för att man ska kunna inleda förhandlingar.
Europaparlamentets Sacharovpris är en utmärkelse för en anmärkningsvärd prestation inom områdena mänskliga rättigheter och grundläggande friheter.
Den kubanska oppositionsrörelsen Kvinnor i vitt, Hauwa Ibrahim, advokat för mänskliga rättigheter i Nigeria, och Reportrar utan gränser delade alla tre på utmärkelsen 2005 och 2004 tilldelades Vitryska journalistförbundet priset
Förbindelserna mellan EU och Ryssland efter mordet på Anna Politkovskaja
Europaparlamentet har antagit en gemensam resolution om förbindelserna mellan EU och Ryssland efter mordet på den ryska journalisten Anna Politkovskaja.
Gemensam resolution Omröstning: 25.10.2006
Parlamentet har antagit en gemensam resolution om toppmötet mellan EU och Ryssland i Helsingfors den 24 november 2006.
Parlamentet uppmanar USA att stänga fånglägret på Guantanamo Bay
Europaparlamentet har mot bakgrund av löpande rapporter om övergrepp, tortyr, och nu nyligen tre självmord på Guantanamo Bay antagit en gemensam resolution för att på nytt uppmana USA:s regering att stänga fånglägret på Guantanamo Bay.
Europaparlamentet uttrycker i en gemensam resolution om situationen i Gazaremsan sin djupa indignation över den militära operation Israel genomfört i Beit Hanun och i Gaza.
Båda sidor uppmanas att försöka få stopp på det våld som drabbar civilbefolkningen, medan USA:s förvaltning uppmanas att se över sin roll i kvartetten
EU bör fortsätta att stödja den palestinska demokratiprocessen
Europaparlamentet har antagit en resolution om framtiden för den nordliga dimensionen.
Resolutionen poängterar att den nordliga dimensionen bättre måste synliggöras för att dess mål ska kunna nås och att förbättrad samordning mellan de olika aktörer som är involverade är en av de viktigaste utmaningarna.
Den nordliga dimensionen bör enligt Europaparlamentet få samma uppmärksamhet som övriga modeller för regionalt samarbete.
Den nordliga dimensionen är ett initiativ från 1999 för att utveckla EU:s yttre relationer och det regionala samarbetet på EU:s nordliga närområden.
Föredragande: Alexander STUBB (EPP-ED, FI) Initiativbetänkande Omröstning: 16.11.2006
Kvinnors rättigheter och jämställdhet
Det nya europeiska jämställdhetsinstitutet kan starta sitt arbete
Merparten av de uppgifter som parlamentet efterlyste i sin första behandling återfinns, exempelvis att institutet ska fokusera mer på analys.
Tack vare överenskommelsen kan nu institutet snart börja sitt arbete och senast tolv månader efter att förordningen trätt i kraft.
De övergripande målen för institutet är att bekämpa könsdiskriminering och främja jämställdhet samt att öka medvetenheten om dessa frågor bland EU:s medborgare
Daphne III - för att bekämpa våld mot barn, ungdomar och kvinnor
Europaparlamentet har antagit ett betänkande om Daphneprogrammet mot våld för perioden 2007–2013 och kräver att budgeten ökas till 125 miljoner euro, vilket är nästan 10 miljoner mer än vad kommissionen föreslog.
Enligt ledamöterna ska bl.a. även åtgärder som riktar sig till kvinnor i befolkningsgrupper med kulturella särdrag eller i etniska minoritetsgrupper omfattas av programmet.
Internationella bröstcancermånaden
Muntliga frågor och resolution Omröstning: 25.10.2006
Strategier för att bekämpa handeln med kvinnor och barn
Handeln med kvinnor och barn, som riskerar att utnyttjas sexuellt, är ett växande internationellt problem som måste bekämpas på global, europeisk och nationell nivå.
Det nya europeiska jämställdhetsinstitutet kan starta sitt arbete Daphne III - för att bekämpa våld mot barn, ungdomar och kvinnor Internationella bröstcancermånaden Strategier för att bekämpa handeln med kvinnor och barn
Parlamentet vill skärpa reglerna för djurskydd
Parlamentet har med bred majoritet antagit ett betänkande som kräver förbättrade regler för djurs välbefinnande.
Ledamöterna vill också att hund- och tuppfäktning ska förbjudas, medan kravet på att även tjurfäktning ska stoppas föll under omröstningen i plenum.
Förbud mot sälprodukter i EU
Korruption skadar fattiga - parlamentet antar en resolution om utvecklingsstöd och korruptionsbekämpning
Ledamöterna kräver tuffare tag mot korruptionen och ett effektivare utnyttjande av EU:s bistånd.
Kommande höjdpunkter
Inledningen av den andra hälften av lagstiftningsperioden sammanfaller med en ny utvidgning och ankomsten av 35 rumänska och 18 bulgariska ledamöter.
Efter Europaparlamentsvalen i juni 2009 minskar antalet till 736 genom en allmän omfördelning då Sverige kommer att mista en av sina 19 platser.
Under de månader som inleder den återstående halvtidsperioden fram till valen i juni 2009 kan nämnas det tredje järnvägspaketet vid januarisammanträdet 2007 och omröstningen i februari om slutbetänkandet från det tillfälliga utskottet för utredning av CIA:s påstådda användning av europeiska länder för transport och illegal internering av fångar.
Ett flertal ärenden kommer att röra klimatförändringarna och energipolitiken, där flera lagstiftningsinitiativ kommer att behandlas, t.ex. systemet med utsläppsrätter och planerna på att inbegripa transporter.
Bilavgaser, luft-, vatten och markkvalitet och biobränslen är andra områden.
Den 23 mars firas femtioårsdagen av EG-fördraget och under våren kommer debatten om EU:s framtid att fortsätta, liksom diskussionen om en reform av EU:s finansieringssystem.
EU:s yttre relationer i synnerhet med Ryssland och med arabvärlden kommer också att stå i fokus.
När det gäller den inre marknaden hoppas man att till 2008 få tillstånd ett direktiv om den fria rörligheten för patienter och hälsovårdstjänster.
En översyn av direktivet om avtal på tidsdelningsbasis (time-sharing) för nyttjande av andelar i fast egendom ska också göras.
Redan under våren kommer parlamentet att behandla kommissionens förslag i fråga om roaming vid gränsöverskridande mobilsamtal.
Parlamentet kommer att göra sin andra behandling av direktivet om audiovisuella tjänster som fastställer nya regler för reklam och produktplacering.
Frågan om märkning av alkoholdrycker (vodkakonflikten) beräknas kunna behandlas i mars.
Säkerheten på EU:s flygplatser ligger i medborgarnas intresse och här inväntar Europaparlamentet rådets gemensamma ståndpunkt.
-//EP//TEXT IM-PRESS 20061113IPR12540 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061207IPR01149 0 NOT XML V0//SV
-//EP//TEXT PRESS TW-20050704-S 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061213IPR01493 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060405IPR07094 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061207IPR01146 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060628IPR09335 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060922IPR10875 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060628IPR09334 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060118IPR04463 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060608IPR08811 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20051206BKG03221 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061207IPR01154 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060901IPR10226 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060113IPR04276 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20051117IPR02436 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060512IPR08047 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060530IPR08575 0 NOT XML V0//SV
-//EP//TEXT PRESS DN-20050705-1 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060524IPR08482 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061129IPR00712 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061020IPR11882 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061020IPR11880 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060628IPR09333 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060113IPR04295 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060628IPR09342 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060922IPR10897 0 NOT XML V0//SV
-//EP//TEXT PRESS TW-20050512-S 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060330IPR06869 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061021IPR11912 0 NOT XML V0//SV
-//EP//TEXT PRESS TW-20041115-S 0 NOT XML V0//SV
-//EP//TEXT PRESS TW-20050622-B 0 NOT XML V0//SV
-//EP//TEXT PRESS TW-20050110-S 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060119STO04525 0 NOT XML V0//SV
-//EP//TEXT PRESS TW-20050411-S 0 NOT XML V0//SV
-//EP//TEXT PRESS TW-20041213-S 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060922IPR10896 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061207IPR01148 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20051017FCS01528 0 NOT XML V0//SV
-//EP//TEXT PRESS TW-20041213-S 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061207IPR01153 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060608IPR08814 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061113IPR12542 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060131IPR04891 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20051111IPR02258 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061113BRI12514 ITEM-011-SV NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061024BRI12109 ITEM-013-SV NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061208IPR01264 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060901IPR10236 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061020IPR11875 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060113IPR04274 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060608IPR08828 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20061010IPR11536 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060906IPR10386 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20060331IPR06930 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 AVU DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 AVU DOC XML V0//EN
Avtal EG/Malaysia om vissa luftfartsaspekter *
Europaparlamentets lagstiftningsresolution av den 24 april 2007 om förslaget till rådets beslut om ingående av avtalet mellan Europeiska gemenskapen och Malaysias regering om vissa luftfartsaspekter (KOM(2006)0619 – C6-0004/2007 – 2006/0202(CNS))
Grundlöner och tillägg för Europols personal *
Europaparlamentets lagstiftningsresolution av den 24 april 2007 om Republiken Finlands initiativ inför antagandet av rådets beslut om justering av grundlöner och tillägg för Europols personal (16333/2006 – C6-0047/2007 – 2007/0801(CNS))
Tullkvoter för import till Bulgarien och Rumänien av rårörsocker *
Europaparlamentets lagstiftningsresolution av den 24 april 2007 om förslaget till rådets förordning om öppnande av tullkvoter för import till Bulgarien och Rumänien av rårörsocker för raffinering under regleringsåren 2006/2007, 2007/2008 och 2008/2009 (KOM(2006)0798 – C6-0003/2007 – 2006/0261(CNS))
Upphävande av Vural Ögers parlamentariska immunitet
Europaparlamentets beslut av den 24 april 2007 om begäran om upphävande av Vural Ögers immunitet (2006/2198(IMM))
Ansvarsfrihet 2005: Avsnitt IV, domstolen
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt IV – domstolen (C6-0467/2006 – 2006/2073(DEC))
2.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt IV – domstolen (C6-0467/2006 – 2006/2073(DEC))
Ansvarsfrihet 2005: Avsnitt V, Revisionsrätten
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt V - revisionsrätten (C6-0468/2006 – 2006/2074(DEC))
2.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt V – revisionsrätten (C6-0468/2006 – 2006/2074(DEC))
Ansvarsfrihet 2005: Avsnitt VI, Europeiska ekonomiska och sociala kommittén
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 200, avsnitt VI - Europeiska ekonomiska och sociala kommittén (C6-0469/2006 – 2006/2075(DEC))
2.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt VI − Europeiska ekonomiska och sociala kommittén (C6-0469/2006 – 2006/2075(DEC))
Ansvarsfrihet 2005: Avsnitt VIIIA - Europeiska ombudsmannen
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt VIIIA -Europeiska ombudsmannen (C6-0471/2006 – 2006/2063(DEC))
2.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt VIIIA − Europeiska ombudsmannen (C6-0471/2006 – 2006/2063(DEC))
Ansvarsfrihet 2005: Avsnitt VIIIB, Europeiska datatillsynsmannen
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt VIIIB - Europeiska datatillsynsmannen (C6-0472/2006 – 2006/2170(DEC))
2.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt VIIIB – Europeiska datatillsynsmannen (C6-0472/2006 – 2006/2170(DEC))
Ansvarsfrihet 2005: sjätte, sjunde, åttonde och nionde europeiska utvecklingsfonden (EUF)
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för sjätte, sjunde, åttonde och nionde Europeiska utvecklingsfonden för budgetåret 2005 (KOM(2006)0429 – C6-0264/2006 – 2006/2169(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna avseende genomförandet av budgeten för sjätte, sjunde, åttonde och nionde Europeiska utvecklingsfonden för budgetåret 2005 (KOM(2006)0429 – C6-0264/2006 – 2006/2169(DEC))
Ansvarsfrihet 2005: Europeiskt centrum för utveckling av yrkesutbildning
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska centrumet för utveckling av yrkesutbildning (Cedefop) för budgetåret 2005 (C6-0386/2006 – 2006/2153(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiskt centrum för utveckling av yrkesutbildning för budgetåret 2005 (C6-0386/2006 – 2006/2153(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiskt centrum för utveckling av yrkesutbildning för budgetåret 2005 (C6-0386/2006 – 2006/2153(DEC))
Ansvarsfrihet: Europeiska fonden för förbättring av levnads- och arbetsvillkor
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska fonden för förbättring av levnads- och arbetsvillkor för budgetåret 2005 (C6-0387/2006 – 2006/2154(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiska fonden för förbättring av levnads- och arbetsvillkor för budgetåret 2005 (C6-0387/2006 – 2006/2154(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska fonden för förbättring av levnads- och arbetsvillkor för budgetåret 2005 (C6-0387/2006 – 2006/2154(DEC))
Ansvarsfrihet 2005: Europeiskt centrum för övervakning av rasism och främlingsfientlighet
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska centrumet för övervakning av rasism och främlingsfientlighet för budgetåret 2005 (C6-0389/2006 – 2006/2156(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiskt centrum för övervakning av rasism och främlingsfientlighet för budgetåret 2005 (C6-0389/2006 – 2006/2156(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiskt centrum för övervakning av rasism och främlingsfientlighet för budgetåret 2005 (C6-0389/2006 – 2006/2156(DEC))
Ansvarsfrihet 2005: Europeiska centrumet för kontroll av narkotika och narkotikamissbruk
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska centrumet för kontroll av narkotika och narkotikamissbruk för budgetåret 2005 (C6-0390/2006 – 2006/2157(DEC))
2.Europaparlamentets beslut av den 24 april 2007 avslutande av räkenskaperna för Europeiska centrumet för kontroll av narkotika och narkotikamissbruk för budgetåret 2005 (C6-0390/2006 – 2006/2157(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska centrumet för kontroll av narkotika och narkotikamissbruk för budgetåret 2005 (C6-0390/2006 – 2006/2157(DEC))
Ansvarsfrihet 2005: Europeiska miljöbyrån
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska miljöbyrån för budgetåret 2005 (C6-0391/2006 – 2006/2158(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiska miljöbyrån för budgetåret 2005 (C6-0391/2006 – 2006/2158(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska miljöbyrån för budgetåret 2005 (C6-0391/2006 – 2006/2158(DEC))
Ansvarsfrihet 2005: Europeiska arbetsmiljöbyrån
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska arbetsmiljöbyrån för budgetåret 2005 (C6-0392/2006 – 2006/2159(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiska arbetsmiljöbyrån för budgetåret 2005 (C6-0392/2006 – 2006/2159(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska arbetsmiljöbyrån för budgetåret 2005 (C6-0392/2006 – 2006/2159(DEC))
Ansvarsfrihet 2005: Översättningscentrum för Europeiska unionens organ
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Översättningscentrumet för Europeiska unionens organ för budgetåret 2005 (C6-0393/2006 – 2006/2160(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Översättningscentrum för Europeiska unionens organ för budgetåret 2005 (C6-0393/2006 – 2006/2160(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Översättningscentrum för Europeiska unionens organ för budgetåret 2005 (C6-0393/2006 – 2006/2160(DEC))
Ansvarsfrihet 2005: Europeiska läkemedelsmyndigheten
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska läkemedelsmyndigheten för budgetåret 2005 (C6-0394/2006 – 2006/2161(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiska läkemedelsmyndigheten för budgetåret 2005 (C6-0394/2006 – 2006/2161(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska läkemedelsmyndigheten för budgetåret 2005 (C6-0394/2006 – 2006/2161(DEC))
Ansvarsfrihet 2005: Eurojust
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Eurojust för budgetåret 2005 (C6-0395/2006 – 2006/2162(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Eurojust för budgetåret 2005 (C6-0395/2006 – 2006/2162(DEC))
Ansvarsfrihet 2005: Europeiska yrkesutbildningsstiftelsen
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska yrkesutbildningsstiftelsen för budgetåret 2005 (C6-0396/2006 – 2006/2163(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiska yrkesutbildningsstiftelsen för budgetåret 2005 (C6-0396/2006 – 2006/2163(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska yrkesutbildningsstiftelsen för budgetåret 2005 (C6-0396/2006 – 2006/2163(DEC))
Ansvarsfrihet 2005: Europeiska sjösäkerhetsbyrån
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska sjösäkerhetsbyrån för budgetåret 2005 (C6-0397/2006 – 2006/2164(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiska sjösäkerhetsbyrån för budgetåret 2005 (C6-0397/2006 – 2006/2164(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska sjösäkerhetsbyrån för budgetåret 2005 (C6-0397/2006 – 2006/2164(DEC))
Ansvarsfrihet 2005: Europeiska byrån för luftfartssäkerhet
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska byrån för luftfartssäkerhet för budgetåret 2005 (C6-0398/2006 – 2006/2165(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiska byrån för luftfartssäkerhet för budgetåret 2005 (C6-0398/2006 – 2006/2165(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska byrån för luftfartssäkerhet för budgetåret 2005 (C6-0398/2006 – 2006/2165(DEC))
Ansvarsfrihet 2005: Europeiska myndigheten för livsmedelssäkerhet
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska myndigheten för livsmedelssäkerhet för budgetåret 2005 (C6-0399/2006 – 2006/2166(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiska myndigheten för livsmedelssäkerhet för budgetåret 2005 (C6-0399/2006 – 2006/2166(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska myndigheten för livsmedelssäkerhet för budgetåret 2005 (C6-0399/2006 – 2006/2166(DEC))
Ansvarsfrihet 2005: Europeiskt centrum för förebyggande och kontroll av sjukdomar
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska centrumet för förebyggande och kontroll av sjukdomar för budgetåret 2005 (C6-0400/2006 – 2006/2167(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiskt centrum för förebyggande och kontroll av sjukdomar för budgetåret 2005 (C6-0400/2006 – 2006/2167(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiskt centrum för förebyggande och kontroll av sjukdomar för budgetåret 2005 (C6-0400/2006 – 2006/2167(DEC))
Ansvarsfrihet 2005: Europeiska byrån för nät- och informationssäkerhet
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska byrån för nät- och informationssäkerhet för budgetåret 2005 (C6-0401/2006 – 2006/2168(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiska byrån för nät- och informationssäkerhet för budgetåret 2005 (C6-0401/2006 – 2006/2168(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska byrån för nät- och informationssäkerhet för budgetåret 2005 (C6-0401/2006 – 2006/2168(DEC))
Betaltjänster på den inre marknaden ***I
Europaparlamentets lagstiftningsresolution av den 24 april 2007 om förslaget till Europaparlamentets och rådets direktiv om betaltjänster på den inre marknaden och om ändring av direktiven 97/7/EG, 2000/12/EG och 2002/65/EG (KOM(2005)0603 – C6-0411/2005 – 2005/0245(COD))
Europaparlamentets ståndpunkt fastställd vid första behandlingen den 24 april 2007 om betaltjänster på den inre marknaden och om ändring av direktiven 97/7/EG, 2002/65/EG, 2005/60/EG och 2006/48/EG samt upphävande av direktiv 97/5/EG
Kvotsystem avseende produktionen av potatisstärkelse *
Europaparlamentets lagstiftningsresolution av den 24 april 2007 om förslaget till rådets förordning om ändring av förordning (EG) nr 1868/94 om inrättandet av ett kvotsystem avseende produktionen av potatisstärkelse (KOM(2006)0827 – C6-0046/2007 – 2006/0268(CNS))
Framtida utvidgningars konsekvenser för sammanhållningspolitikens effektivitet
Europaparlamentets resolution av den 24 april 2007 om framtida utvidgningars konsekvenser för sammanhållningspolitikens effektivitet (2006/2107(INI))
Kommissionens årliga politiska strategi för 2008
Europaparlamentets resolution av den 24 april 2007 om kommissionens årliga politiska strategi för budgetförfarandet för 2008 (2007/2017(BUD))
BILAGA I
BILAGA II
Ansvarsfrihet 2006: avsnitt III, kommissionen
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt III - kommissionen (SEK(2006)0916 – C6-0263/2006 – 2006/2070(DEC)) (SEK(2006)0915 – C6-0262/2006 – 2006/2070(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna avseende genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt III – kommissionen (SEK(2006)0916 – C6-0263/2006 – 2006/2070(DEC)) (SEK(2006)0915 – C6-0262/2006 – 2006/2070(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt III – kommissionen (SEK(2006)0916 – C6-0263/2006 – 2006/2070(DEC)) (SEK(2006)0915 – C6-0262/2006 – 2006/2070(DEC))
Ansvarsfrihet 2005: Avsnitt I, Europaparlamentet
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt I - Europaparlamentet (C6-0465/2006 – 2006/2071(DEC))
2.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt I – Europaparlamentet (C6-0465/2006 – 2006/2071(DEC))
Ansvarsfrihet 2005: Avsnitt II, rådet
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt II – rådet (C6-0466/2006 – 2006/2072(DEC))
2.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt II – rådet (C6-0466/2006 – 2006/2072(DEC))
Ansvarsfrihet 2005: Avsnitt VII, Regionkommittén
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005 - avsnitt VII - Regionkommittén(C6-0470/2006 – 2006/2076(DEC))
2.Europaparlamentets resolution av den 24 april 2007med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2005, avsnitt VII − Regionkommittén (C6-0470/2006 – 2006/2076(DEC))
Ansvarsfrihet 2005: Europeiska byrån för återuppbyggnad
1.Europaparlamentets beslut av den 24 april 2007 om ansvarsfrihet för genomförandet av budgeten för Europeiska byrån för återuppbyggnad för budgetåret 2005 (C6-0388/2006 – 2006/2155(DEC))
2.Europaparlamentets beslut av den 24 april 2007 om avslutande av räkenskaperna för Europeiska byrån för återuppbyggnad för budgetåret 2005 (C6-0388/2006 – 2006/2155(DEC))
3.Europaparlamentets resolution av den 24 april 2007 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska byrån för återuppbyggnad för budgetåret 2005 (C6-0388/2006 – 2006/2155(DEC))
Bekämpning av hiv/aids i Europeiska unionen och angränsande länder 2006-2009
Europaparlamentets resolution av den 24 april 2007 om bekämpning av hiv/aids i Europeiska unionen och angränsande länder 2006–2009 (2006/2232(INI))
Förenkling av gemenskapslagstiftning (ändring av arbetsordningen)
Europaparlamentets beslut av den 10 maj 2007 om ändring av Europaparlamentets arbetsordning för att anpassa de interna förfarandena till kravet på en förenkling av gemenskapslagstiftningen (2005/2238(REG))
Kollektivtrafik på järnväg och väg ***II
Europaparlamentets lagstiftningsresolution av den 10 maj 2007 om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets förordning om kollektivtrafik på järnväg och väg och om upphävande av rådets förordningar (EEG) nr 1191/69 och (EEG) nr 1107/70 (13736/1/2006 – C6-0042/2007 – 2000/0212(COD))
Bestämmelser för färdigförpackade varors nominella mängder ***II
Europaparlamentets lagstiftningsresolution av den 10 maj 2007 om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets direktiv om fastställande av bestämmelser för färdigförpackade varors nominella mängder, om upphävande av rådets direktiv 75/106/EEG och 80/232/EEG samt om ändring av rådets direktiv 76/211/EEG (13484/1/2006 – C6-0039/2007 – 2004/0248(COD))
Godkännande av fordon och släpvagnar ***II
Europaparlamentets lagstiftningsresolution av den 10 maj 2007 om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets direktiv om fastställande av en ram för godkännande av motorfordon och släpvagnar till dessa fordon samt av system, komponenter och separata tekniska enheter som är avsedda för sådana fordon ("ramdirektiv") (9911/3/2006 – C6-0040/2007 – 2003/0153(COD))
Montering i efterhand av backspeglar på tunga lastbilar ***I
Europaparlamentets lagstiftningsresolution av den 10 maj 2007 om förslaget till Europaparlamentets och rådets direktiv om eftermontering av speglar på tunga fordon registrerade i gemenskapen (KOM(2006)0570 – C6-0332/2006 – 2006/0183(COD))
Europaparlamentets ståndpunkt fastställd vid första behandlingen den 10 maj 2007 inför antagandet av Europaparlamentets och rådets direktiv
2007/.../EG
om eftermontering av speglar på tunga fordon registrerade i gemenskapen
Toppmötet mellan EU och Ryssland
Europaparlamentets resolution av den 10 maj 2007 om toppmötet mellan EU och Ryssland i Samara den 18 maj 2007
Reformerna i arabvärlden: Vilken strategi bör EU följa?
Europaparlamentets resolution av den 10 maj 2007 om reformer i arabvärlden: vilken strategi bör EU följa? (2006/2172(INI))
Afrikas horn: EU:s regionala politiska partnerskap för fred, säkerhet och utveckling
Europaparlamentets resolution av den 10 maj 2007 om Afrikas horn: EU:s regionala politiska partnerskap för fred, säkerhet och utveckling (2006/2291(INI))
Utvärdering av Euratom
Europaparlamentets resolution av den 10 maj 2007 om utvärdering av Euratom – femtio år av gemensam kärnkraftspolitik (2006/2230(INI))
Skydd av miljön mot strålning till följd av en olycka med ett militärflygplan på Grönland
Europaparlamentets resolution av den 10 maj 2007 om konsekvenserna för folkhälsan av Thule-olyckan 1968 (framställning nr 720/2002) (2006/2012(INI))
Bostäder och regionalpolitik
Europaparlamentets resolution av den 10 maj 2007 om bostäder och regionalpolitik (2006/2108(INI))
Den framtida regionalpolitiken och innovation
Europaparlamentets resolution av den 10 maj 2007 om den framtida regionalpolitikens bidrag till Europeiska unionens innovativa kapacitet (2006/2104(INI))
Förstärkning av gemenskapsrätten beträffande information och samråd med arbetstagare
Europaparlamentets resolution av den 10 maj 2007 om förstärkning av gemenskapsrätten beträffande information och samråd med arbetstagare
Enade i mänsklig värdighet: EU:s talman möter religiösa ledare
Kultur
2007-05-15 - 17:54
Talman Hans-Gert Poettering, Angela Merkel och den tyske rabbin Chaim Soussan.
Ett Europa byggt på mänsklig värdighet var temat för ett möte mellan ledarna av de tre monoteistiska religionerna och ledarna av tre EU-institutioner i dag den 15 maj i kommissionen.
Talman Pöttering representerade Europaparlamentet under diskussionen, Barroso kommissionen samt Angela Merkel rådet.
Det var första gången som de tre europeiska institutionerna mötte de 20 ledande representanterna av den kristna, judiska och islamska tron i Europa.
Vilken roll kan religion och religiösa samhällen spela i Europa, baserat på mänsklig värdighet?
Värden som demokrati, lagen, tolerans, rättvisa, solidaritet, ömsesidig respekt och mänsklig värdighet är det som binder européer samman.
Representanterna för de olika religiösa inriktningarna och representanterna från EU-institutionerna kom överens om att genom dessa värden kommer de alla att arbeta mot samma mål, det gemensamma goda.
"Underbar upplevelse"
Talman Pöttering sa att det var en "underbar upplevelse att lyssna till kristna, judiska och muslimska röster.
Han lade till: "till trots för alla våra olikheter så finns där en gemensam punkt: mänsklig värdighet, och vi är överens om att den behöver försvaras och det borde vara basen för vårt politiska arbete".
Han sa att europeiska institutioner är ansvariga för att omsätta mänsklig värdighet i praktik.
Barroso reagerade på denna fråga genom att säga att kommissionen kommer att föreslå ett direktiv för flyktingars rättigheter i EU.
Pöttering sa att när detta förslag är skrivet kommer det att komma till Europaparlamentet för att ta ett beslut på lika villkor som rådet.
"Europaparlamentet kommer att se till att dessa principer av mänsklig värdighet är inkluderade".
Barroso betonade också temat med mänsklig värdighet "som en kärnfråga för de tre religionerna men också för EU-institutionerna: frihet, fred, rättvisa och solidaritet".
Han lade till: "Vi diskuterade behovet av att respektera religionsfrihet, i EU och i alla länder som vill bli del av EU.
Angela Merkel sa att "dialog mellan politiker och religioner är essentiell".
Hon berättade att de diskuterade Berlinförklaringen och 50-årsfirandet av Romfördraget.
När hon svarade på en fråga från en journalist om inkluderandet av "Gud" i det nya konstitutionella fördraget sa hon: "Personligen skulle jag vilja ha en sådan referens, men jag tror att det är liten chans att det blir inkluderat.
Det finns redan en referens till kyrkor i förslaget till det konstitutionella fördraget, vilket är viktigt.
Men tyvärr kan jag inte lova någonting annat".
Hon sa också: "Vi är alla överens om att mänsklig värdighet är okränkbart men det finns olika synsätt på de praktiska implikationerna av det".
Ledarna sa att ett liknande möte kommer att organiseras under det slovenska ordförandeskapet (januari-juni 2008).
20070514STO06592 Pressmeddelande från talman Pöttering
SV
1
PHOTO
20070515PHT06677.jpg
SV
2
LINK
/president/defaulten.htm
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//TEXT TA 20070522 ITEMS DOC XML V0//SV
TECKENFÖRKLARING
*
Samrådsförfarandet
** I
** II
***
Samtyckesförfarandet
***I
Medbeslutandeförfarandet (första behandlingen)
***II
Medbeslutandeförfarandet (andra behandlingen)
***III
UPPLYSNINGAR ANGÅENDE OMRÖSTNINGAR
Om inget annat anges har föredraganden till talmannen skriftligen tillkännagivit sin inställning till ändringsförslagen.
FÖRKORTNINGAR FÖR UTSKOTTENS NAMN
AFET:
DEVE:
Utskottet för utveckling
INTA:
Utskottet för internationell handel
BUDG:
Budgetutskottet
CONT:
Budgetkontrollutskottet
ECON:
Utskottet för ekonomi och valutafrågor
EMPL:
Utskottet för sysselsättning och sociala frågor
ENVI:
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
ITRE:
Utskottet för industrifrågor, forskning och energi
IMCO:
Utskottet för den inre marknaden och konsumentskydd
TRAN:
Utskottet för transport och turism
REGI:
Utskottet för regional utveckling
AGRI:
PECH:
Fiskeriutskottet
CULT:
Utskottet för kultur och utbildning
JURI:
Utskottet för rättsliga frågor
LIBE:
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
AFCO:
Utskottet för konstitutionella frågor
FEMM:
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
PETI:
Utskottet för framställningar
FÖRKORTNINGAR FÖR DE POLITISKA GRUPPERNA
PPE-DE:
Gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater
PSE:
Europeiska socialdemokratiska partiets grupp
ALDE:
Gruppen Alliansen liberaler och demokrater för Europa
UEN:
Gruppen Unionen för nationernas Europa
Verts/ALE
Gruppen De gröna/Europeiska fria alliansen
GUE/NGL:
Gruppen Europeiska enade vänstern/Nordisk grön vänster
IND/DEM:
Gruppen Självständighet/Demokrati
ITS
Gruppen Identitet, tradition och suveränitet
NI:
Grupplösa
Öppnande av sammanträdet
Inkomna dokument
Roaming i allmänna mobilnät ***I (debatt)
Anständigt arbete för alla (debatt)
Omröstning
Gemenskapens finansiella stöd på området transeuropeiska nät på transportområdet och energiområdet ***II (omröstning)
Roaming i allmänna mobilnät ***I (omröstning)
Avtalet om ekonomiskt partnerskap, politisk samordning och samarbete EG/Mexiko * (omröstning)
Tillnärmning av punktskattesatser på alkohol och alkoholdrycker * (omröstning)
Sammansättning av delegationen till EUROLAT (omröstning)
Effekterna och konsekvenserna av att undanta vårdtjänster från direktivet om tjänster på den inre marknaden (omröstning)
Strukturpolitikens effekter på sammanhållningen i EU (omröstning)
EU:s handelsrelaterade bistånd (omröstning)
Avtal om ekonomiskt partnerskap (omröstning)
Gemensam utrikes- och säkerhetspolitik 2005 (omröstning)
Anständigt arbete för alla (omröstning)
Röstförklaringar
Rättelser/avsiktsförklaringar till avgivna röster
Justering av protokollet från föregående sammanträde
Débat sur le futur de l'Europe (debatt)
Situationen i Nigeria (debatt)
Internationell handel med utrotningshotade arter av vilda djur och växter (CITES) (debatt)
Frågestund (frågor till rådet)
Valprövning av Beniamino Donnici (debatt)
Innovationsstrategi (debatt)
Bekämpande av organiserad brottslighet (debatt)
Gemensam organisation av jordbruksmarknaderna * (debatt)
Den gemensamma organisationen av marknaden för spannmål * (debatt)
Föredragningslista för nästa sammanträde
Avslutande av sammanträdet
NÄRVAROLISTA
PROTOKOLL
ORDFÖRANDESKAP: Alejo VIDAL-QUADRAS Vice talman
1 Öppnande av sammanträdet
Sammanträdet öppnades kl. 09.00.
2 Inkomna dokument
Följande dokument hade kommit in från utskottet JURI:
- Betänkande om valprövning av Beniamino Donnici ( 2007/2121(REG) ) - utskottet JURI - Föredragande: Giuseppe Gargani ( A6-0198/2007 )
3
Roaming i allmänna mobilnät ***I (debatt)
Betänkande om förslaget till Europaparlamentets och rådets förordning om roaming i allmänna mobilnät i gemenskapen och om ändring av direktiv 2002/21/EG om ett gemensamt regelverk för elektroniska kommunikationsnät och kommunikationstjänster [ KOM(2006)0382 - C6-0244/2006 - 2006/0133(COD) ] - Utskottet för industrifrågor, forskning och energi.
Föredragande: Paul Rübig ( A6-0155/2007 )
Talare:
Viviane Reding (ledamot av kommissionen) .
Paul Rübig redogjorde för sitt betänkande.
Talare:
Joachim Wuermeling (rådets tjänstgörande ordförande) .
Talare:
Andrea Losco (föredragande av yttrande från utskottet ECON),
Joseph Muscat (föredragande av yttrande från utskottet IMCO),
Manolis Mavrommatis (föredragande av yttrande från utskottet CULT),
Angelika Niebler för PPE-DE-gruppen,
Reino Paasilinna för PSE-gruppen,
Šarūnas Birutis för ALDE-gruppen,
Romano Maria La Russa för UEN-gruppen,
David Hammerstein för Verts/ALE-gruppen,
Umberto Guidoni för GUE/NGL-gruppen,
Nigel Farage för IND/DEM-gruppen,
Giles Chichester ,
Robert Goebbels ,
Toine Manders ,
Adam Bielan ,
Gisela Kallenbach ,
Miloslav Ransdorf och
Gunnar Hökmark .
ORDFÖRANDESKAP: Luigi COCILOVO Vice talman
Talare:
Hannes Swoboda ,
Lena Ek ,
Roberts Zīle ,
Claude Turmes ,
Vittorio Agnoletto ,
Pilar del Castillo Vera ,
Andres Tarand ,
Alexander Alvaro ,
Alyn Smith ,
Ivo Belet ,
Evelyne Gebhardt ,
Anneli Jäätteenmäki ,
Herbert Reul ,
Arlene McCarthy ,
Karin Riis-Jørgensen ,
Marianne Thyssen ,
Eluned Morgan ,
Nikolaos Vakalis ,
Katerina Batzeli ,
Zita Pleštinská ,
Béatrice Patrie ,
Françoise Grossetête ,
Silvia-Adriana Ţicău ,
Jerzy Buzek ,
Dorette Corbey ,
Zuzana Roithová ,
Dariusz Rosati ,
Lambert van Nistelrooij ,
Mia De Vits ,
Werner Langen ,
Edit Herczog och
Joachim Wuermeling .
ORDFÖRANDESKAP: Luisa MORGANTINI Vice talman
Omröstning:
punkt 5.2 i protokollet av den 23.05.2007
.
4
Anständigt arbete för alla (debatt)
Betänkande om anständigt arbete för alla [ 2006/2240(INI) ] - Utskottet för sysselsättning och sociala frågor.
Föredragande: Marie Panayotopoulos-Cassiotou ( A6-0068/2007 )
Marie Panayotopoulos-Cassiotou redogjorde för sitt betänkande.
Talare:
Vladimír Špidla (ledamot av kommissionen) .
Talare:
Feleknas Uca (föredragande av yttrande från utskottet DEVE),
Harlem Désir (föredragande av yttrande från utskottet INTA),
Philip Bushill-Matthews för PPE-DE-gruppen,
Stephen Hughes för PSE-gruppen,
Ona Juknevičienė för ALDE-gruppen,
Zdzisław Zbigniew Podkański för UEN-gruppen,
Sepp Kusstatscher för Verts/ALE-gruppen,
Kyriacos Triantaphyllides för GUE/NGL-gruppen,
Derek Roland Clark för IND/DEM-gruppen,
Cristian Stănescu för ITS-gruppen,
Alessandro Battilocchio , grupplös,
José Albino Silva Peneda ,
Anne Van Lancker ,
Marian Harkin ,
Ilda Figueiredo ,
Kathy Sinnott ,
Jean-Claude Martinez ,
Jan Andersson ,
Georgios Karatzaferis ,
Magda Kósáné Kovács ,
Ole Christensen och
Vladimír Špidla .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 5.11 i protokollet av den 23.05.2007
.
ORDFÖRANDESKAP: Edward McMILLAN-SCOTT Vice talman
5 Omröstning
Omröstningsresultaten (ändringsförslag, särskilda omröstningar, delade omröstningar etc.) återfinns i bilagan ”Omröstningsresultat” som bifogas protokollet.
5.1
Gemenskapens finansiella stöd på området transeuropeiska nät på transportområdet och energiområdet ***II (omröstning)
Andrabehandlingsrekommendation om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets förordning om allmänna regler för gemenskapens finansiella stöd på området för transeuropeiska nät på transportområdet och energiområdet [17032/2/2006 - C6-0101/2007 - 2004/0154(COD) ] - Budgetutskottet.
Föredragande: Mario Mauro ( A6-0169/2007 )
(Kvalificerad majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 1)
RÅDETS GEMENSAMMA STÅNDPUNKT
Förklarades godkänt såsom ändrat av parlamentet
(
P6_TA(2007)0198
)
5.2
Roaming i allmänna mobilnät ***I (omröstning)
Betänkande om förslaget till Europaparlamentets och rådets förordning om roaming i allmänna mobilnät i gemenskapen och om ändring av direktiv 2002/21/EG om ett gemensamt regelverk för elektroniska kommunikationsnät och kommunikationstjänster [ KOM(2006)0382 - C6-0244/2006 - 2006/0133(COD) ] - Utskottet för industrifrågor, forskning och energi.
Föredragande: Paul Rübig ( A6-0155/2007 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 2)
KOMMISSIONENS FÖRSLAG
Godkändes såsom ändrat av parlamentet
(
P6_TA(2007)0199
)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs
(
P6_TA(2007)0199
)
Inlägg om omröstningen:
-
Martin Callanan och
-
Richard Corbett om dessa inlägg.
-
Paul Rübig (föredragande) , efter omröstningen.
5.3
Avtalet om ekonomiskt partnerskap, politisk samordning och samarbete EG/Mexiko * (omröstning)
Betänkande om förslaget till rådets beslut om ingående av ett andra tilläggsprotokoll till avtalet om ekonomiskt partnerskap, politisk samordning och samarbete mellan Europeiska gemenskapen och dess medlemsstater, å ena sidan, och Mexikos förenta stater, å andra sidan, med anledning av Republiken Bulgariens och Rumäniens anslutning till Europeiska unionen [ KOM(2006)0777 - C6-0077/2007 - 2006/0259(CNS) ] - Utskottet för internationell handel.
Föredragande: Helmuth Markov ( A6-0138/2007 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 3)
KOMMISSIONENS FÖRSLAG
Godkändes såsom ändrat av parlamentet
(
P6_TA(2007)0200
)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs
(
P6_TA(2007)0200
)
5.4
Tillnärmning av punktskattesatser på alkohol och alkoholdrycker * (omröstning)
Betänkande om förslaget till rådets direktiv om ändring av direktiv 92/84/EEG om tillnärmning av punktskattesatser på alkohol och alkoholdrycker [ KOM(2006)0486 - C6-0319/2006 - 2006/0165(CNS) ] - Utskottet för ekonomi och valutafrågor.
Föredragande: Astrid Lulling ( A6-0148/2007 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 4)
KOMMISSIONENS FÖRSLAG
Förkastades
Inlägg om omröstningen:
-
Ieke van den Burg och
Astrid Lulling (föredragande)
.
5.5 Sammansättning av delegationen till EUROLAT (omröstning)
om tillsättning av delegationen till den parlamentariska församlingen EU-Latinamerika och antalet ledamöter i delegationen
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 5)
TALMANSKONFERENSENS FÖRSLAG
Antogs
Talmannen meddelade att PPE-DE-gruppen hade meddelat att den hade utsett
Antonio Tajani till ordinarie ledamot av delegationen.
5.6
Effekterna och konsekvenserna av att undanta vårdtjänster från direktivet om tjänster på den inre marknaden (omröstning)
Betänkande om effekterna och konsekvenserna av att undanta vårdtjänster från direktivet om tjänster på den inre marknaden [ 2006/2275(INI) ] - Utskottet för den inre marknaden och konsumentskydd.
Föredragande: Bernadette Vergnaud ( A6-0173/2007 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 6)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2007)0201
)
Inlägg om omröstningen:
-
Bernadette Vergnaud (föredragande) meddelade för omröstningen att det förelåg ett fel som rörde punkterna 47 och3 (talmannen meddelade att en korrekt version av texten hade delats ut).
5.7
Strukturpolitikens effekter på sammanhållningen i EU (omröstning)
Betänkande om strukturpolitikens effekter på sammanhållningen i EU [ 2006/2181(INI) ] - Utskottet för regional utveckling.
Föredragande: Francisca Pleguezuelos Aguilar ( A6-0150/2007 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 7)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2007)0202
)
5.8
EU:s handelsrelaterade bistånd (omröstning)
Betänkande om EU:s handelsrelaterade bistånd [ 2006/2236(INI) ] - Utskottet för internationell handel.
Föredragande: David Martin ( A6-0088/2007 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 8)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2007)0203
)
5.9
Avtal om ekonomiskt partnerskap (omröstning)
Betänkande om avtal om ekonomiskt partnerskap [ 2005/2246(INI) ] - Utskottet för internationell handel.
Föredragande: Robert Sturdy ( A6-0084/2007 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 9)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2007)0204
)
Inlägg om omröstningen:
-
Margrietus van den Berg lade fram ett muntligt ändringsförslag till ändringsförslag 23, vilket beaktades.
5.10
Gemensam utrikes- och säkerhetspolitik 2005 (omröstning)
Betänkande om rådets årliga rapport till Europaparlamentet om de viktigaste aspekterna och de grundläggande vägvalen när det gäller GUSP, inbegripet de finansiella konsekvenserna för Europeiska unionens allmänna budget 2005 [ 2006/2217(INI) ] - Utskottet för utrikesfrågor.
Föredragande: Elmar Brok ( A6-0130/2007 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 10)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2007)0205
)
Inlägg om omröstningen:
-
Vittorio Agnoletto meddelade att han hade blandat ihop punkt 10 och punkt 11 och därför röstat fel.
5.11
Anständigt arbete för alla (omröstning)
Betänkande om anständigt arbete för alla [ 2006/2240(INI) ] - Utskottet för sysselsättning och sociala frågor.
Föredragande: Marie Panayotopoulos-Cassiotou ( A6-0068/2007 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 11)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2007)0206
)
6 Röstförklaringar
Skriftliga röstförklaringar:
Muntliga röstförklaringar:
Betänkande Mario Mauro - A6-0169/2007 :
Hubert Pirker och
Andreas Mölzer
Betänkande Paul Rübig - A6-0155/2007 :
Gyula Hegyi och
Ivo Strejček
Betänkande Astrid Lulling - A6-0148/2007 :
Danutė Budreikaitė och
Andreas Mölzer
Betänkande Bernadette Vergnaud - A6-0173/2007 :
Miroslav Mikolášik
Betänkande Elmar Brok - A6-0130/2007 :
Hubert Pirker
Betänkande Marie Panayotopoulos-Cassiotou - A6-0068/2007 :
Hubert Pirker och
John Attard-Montalto .
7 Rättelser/avsiktsförklaringar till avgivna röster
Den elektroniska versionen på Europarl uppdateras regelbundet under högst två veckor efter den aktuella omröstningsdagen.
Därefter slutförs förteckningen över rättelserna till de avgivna rösterna för att översättas och offentliggöras i Europeiska unionens officiella tidning.
Följande ledamöter meddelade att de av tekniska skäl inte hade kunnat delta i följande omröstningar:
Betänkande Mario Mauro - A6-0169/2007 :
- ändringsförslag 2:
Mario Mauro
Betänkande Astrid Lulling - A6-0148/2007 :
- ändrat förslag:
Othmar Karas
Rapport Bernadette Vergnaud - A6-0173/2007 :
- punkt 4:
Guido Podestà
- ändringsförslag 20:
Bruno Gollnisch
- punkt 71:
Bernadette Vergnaud
Betänkande Francisca Pleguezuelos Aguilar - A6-0150/2007 :
- ändringsförslag 12:
Bernadette Vergnaud
- ändringsförslag 4:
Roberta Angelilli
Betänkande David Martin - A6-0088/2007 :
- slutomröstning:
Marie Anne Isler Béguin
ORDFÖRANDESKAP: Hans-Gert PÖTTERING Talman
Maria Petre hade låtit meddela att hon hade varit närvarande men att hennes namn inte förekom på närvarolistan.
Protokollet från föregående sammanträde justerades.
9 Débat sur le futur de l'Europe (debatt)
Talmannen gjorde ett kort inlägg som inledning på debatten.
Talare:
Jan Peter Balkenende , Nederländernas premiärminister.
Talare:
Joseph Daul för PPE-DE-gruppen,
Martin Schulz för PSE-gruppen,
Graham Watson för ALDE-gruppen,
Brian Crowley för UEN-gruppen,
Kathalijne Maria Buitenweg för Verts/ALE-gruppen,
Erik Meijer för GUE/NGL-gruppen,
Bastiaan Belder för IND/DEM-gruppen,
Philip Claeys för ITS-gruppen,
Jim Allister , grupplös,
Jan Peter Balkenende ,
Maria Martens ,
Margrietus van den Berg ,
Andrew Duff ,
Konrad Szymański ,
Johannes Voggenhuber ,
Sylvia-Yvonne Kaufmann ,
Jens-Peter Bonde ,
Andreas Mölzer ,
Timothy Kirkhope ,
Richard Corbett ,
Jules Maaten ,
Guntars Krasts ,
Vladimír Remek ,
Nils Lundgren ,
Jean-Luc Dehaene ,
Enrique Barón Crespo ,
Sophia in 't Veld ,
Hanna Foltyn-Kubicka ,
Adrian Severin och
Jan Peter Balkenende .
Talmannen förklarade debatten avslutad.
ORDFÖRANDESKAP: Mechtild ROTHE Vice talman
10
Situationen i Nigeria (debatt)
Uttalanden av rådet och kommissionen:
Situationen i Nigeria
Günter Gloser (rådets tjänstgörande ordförande) och
Benita Ferrero-Waldner (ledamot av kommissionen) gjorde uttalanden.
Talare:
Filip Kaczmarek för PPE-DE-gruppen,
Margrietus van den Berg för PSE-gruppen,
Johan Van Hecke för ALDE-gruppen,
Marie-Hélène Aubert för Verts/ALE-gruppen,
Vittorio Agnoletto för GUE/NGL-gruppen,
Bastiaan Belder för IND/DEM-gruppen,
Andreas Mölzer för ITS-gruppen,
Edward McMillan-Scott ,
Libor Rouček ,
Fiona Hall ,
Urszula Krupa ,
Bogusław Sonik ,
Pierre Schapira ,
Toomas Savi ,
Luís Queiró ,
Karin Scheele ,
András Gyürk ,
Ryszard Czarnecki ,
Günter Gloser och
Benita Ferrero-Waldner .
-
Filip Kaczmarek och
Edward McMillan-Scott för PPE-DE-gruppen ,
Margrietus van den Berg ,
John Attard-Montalto och
Libor Rouček för PSE-gruppen ,
Toomas Savi ,
Thierry Cornillet och
Johan Van Hecke för ALDE-gruppen ,
Ryszard Czarnecki ,
Eoin Ryan ,
Adam Bielan och
Michał Tomasz Kamiński för UEN-gruppen ,
Margrete Auken för Verts/ALE-gruppen, och
Vittorio Agnoletto för GUE/NGL-gruppen ,
om de nyligen hållna valen i Nigeria ( B6-0201/2007 ) .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 7.4 i protokollet av den 24.05.2007
.
11
Internationell handel med utrotningshotade arter av vilda djur och växter (CITES) (debatt)
Muntlig fråga (
O-0018/2007 ) från
Miroslav Ouzký , för utskottet ENVI, till rådet:
Huvudmålen för konferensen för parterna i konventionen om internationell handel med utrotningshotade arter av vilda djur och växter (CITES) i Haag den 3-15 juni 2007 ( B6-0020/2007 )
Muntlig fråga (
O-0019/2007 ) från
Miroslav Ouzký , för utskottet ENVI, till kommissionen:
Huvudmålen för konferensen för parterna i konventionen om internationell handel med utrotningshotade arter av vilda djur och växter (CITES) i Haag den 3-15 juni 2007 ( B6-0121/2007 )
Marie Anne Isler Béguin (ersättare för frågeställaren) utvecklade de muntliga frågorna.
ORDFÖRANDESKAP: Diana WALLIS Vice talman
Günter Gloser (rådets tjänstgörande ordförande) besvarade frågan (
B6-0020/2007 ).
Benita Ferrero-Waldner (ledamot av kommissionen) besvarade frågan (
B6-0121/2007 ).
Talare:
John Bowis för PPE-DE-gruppen,
Dorette Corbey för PSE-gruppen,
Mojca Drčar Murko för ALDE-gruppen,
Marie Anne Isler Béguin för Verts/ALE-gruppen,
Johannes Blokland för IND/DEM-gruppen,
Karin Scheele ,
Alfonso Andria och
Benita Ferrero-Waldner .
-
Miroslav Ouzký , för utskottet ENVI,
om EU:s strategiska mål för det fjortonde mötet i partskonferensen för konventionen om internationell handel med utrotningshotade arter av vilda djur och växter (CITES-konventionen), avsedd att hållas i Haag den 3-15 juni 2007 ( B6-0200/2007 ) .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 7.5 i protokollet av den 24.05.2007
.
12
Frågestund (frågor till rådet)
B6-0018/2007 ).
Fråga 1 (Rodi Kratsa-Tsagaropoulou): Politisk kris i Turkiet och utsikterna till medlemskap
H-0339/07 .
Rodi Kratsa-Tsagaropoulou ,
Reinhard Rack och
H-0278/07 .
Manuel Medina Ortega ,
Simon Busuttil och
H-0280/07 .
Marie Panayotopoulos-Cassiotou ,
Robert Evans ,
Justas Vincas Paleckis och
H-0285/07 .
Sarah Ludford .
H-0287/07 .
Bernd Posselt .
H-0291/07 .
Philip Bushill-Matthews .
H-0294/07 .
Marie Anne Isler Béguin och
Justas Vincas Paleckis .
(
) .
ORDFÖRANDESKAP: Edward McMILLAN-SCOTT Vice talman
Betänkande om valprövning av Beniamino Donnici - Utskottet för rättsliga frågor.
Föredragande: Giuseppe Gargani ( A6-0198/2007 )
Giuseppe Gargani redogjorde för sitt betänkande.
Talare:
Manuel Medina Ortega för PSE-gruppen,
Luigi Cocilovo för ALDE-gruppen,
Salvatore Tatarella för UEN-gruppen, och
Nicola Zingaretti .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 7.3 i protokollet av den 24.05.2007
.
14
Innovationsstrategi (debatt)
Betänkande om meddelandet "Kunskap i praktiken: en brett upplagd innovationsstrategi för EU" ( 2006/2274(INI) ) - Utskottet för industrifrågor, forskning och energi.
Föredragande: Adam Gierek ( A6-0159/2007 )
Adam Gierek redogjorde för sitt betänkande.
Talare:
Günter Verheugen (kommissionens vice ordförande) .
Talare:
Sharon Bowles (föredragande av yttrande från utskottet ECON),
Barbara Weiler (föredragande av yttrande från utskottet IMCO),
Christa Prets (föredragande av yttrande från utskottet REGI),
Jaroslav Zvěřina (föredragande av yttrande från utskottet JURI),
Ján Hudacký för PPE-DE-gruppen,
Silvia-Adriana Ţicău för PSE-gruppen,
Patrizia Toia för ALDE-gruppen,
Mieczysław Edmund Janowski för UEN-gruppen,
David Hammerstein för Verts/ALE-gruppen,
Lambert van Nistelrooij ,
Gábor Harangozó ,
Šarūnas Birutis och
Zbigniew Krzysztof Kuźmiuk .
ORDFÖRANDESKAP: Rodi KRATSA-TSAGAROPOULOU Vice talman
Talare:
Zita Pleštinská ,
Jorgo Chatzimarkakis och
Jerzy Buzek .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 9.1 i protokollet av den 24.05.2007
.
15
Bekämpande av organiserad brottslighet (debatt)
Betänkande om rekommendationen till rådet om utarbetande av ett strategiskt koncept för bekämpande av organiserad brottslighet [ 2006/2094(INI) ] - Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor.
Föredragande: Bill Newton Dunn ( A6-0152/2007 )
Bill Newton Dunn redogjorde för sitt betänkande.
Talare:
Franco Frattini (kommissionens vice ordförande) .
Talare:
Giuseppe Castiglione för PPE-DE-gruppen,
Magda Kósáné Kovács för PSE-gruppen,
Marios Matsakis för ALDE-gruppen,
Giusto Catania för GUE/NGL-gruppen,
Petre Popeangă för ITS-gruppen,
Jim Allister , grupplös,
Carlos Coelho och
Adina-Ioana Vălean .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 9.2 i protokollet av den 24.05.2007
.
16
Gemensam organisation av jordbruksmarknaderna * (debatt)
Betänkande om förslaget till rådets förordning om upprättande av en gemensam organisation av jordbruksmarknaderna och om särskilda bestämmelser för vissa jordbruksprodukter [ KOM(2006)0822 - C6-0045/2007 - 2006/0269(CNS) ] - Utskottet för jordbruk och landsbygdens utveckling.
Föredragande: Niels Busk ( A6-0171/2007 )
Talare:
Benita Ferrero-Waldner (ledamot av kommissionen) .
ORDFÖRANDESKAP: Luisa MORGANTINI Vice talman
Omröstning:
punkt 7.1 i protokollet av den 24.05.2007
.
17
Den gemensamma organisationen av marknaden för spannmål * (debatt)
Betänkande om förslaget till rådets förordning om ändring av förordning (EG) nr 1784/2003 om den gemensamma organisationen av marknaden för spannmål [ KOM(2006)0755 - C6-0044/2007 - 2006/0256(CNS) ] - Utskottet för jordbruk och landsbygdens utveckling.
Föredragande: Béla Glattfelder ( A6-0141/2007 )
Talare:
Benita Ferrero-Waldner (ledamot av kommissionen) .
Béla Glattfelder redogjorde för sitt betänkande.
Talare:
James Nicholson för PPE-DE-gruppen,
Bogdan Golik för PSE-gruppen,
Leopold Józef Rutowicz för UEN-gruppen,
Czesław Adam Siekierski ,
Monica Maria Iacob-Ridzi och
Benita Ferrero-Waldner .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 7.2 i protokollet av den 24.05.2007
.
18 Föredragningslista för nästa sammanträde
Föredragningslistan för nästa sammanträde fastställdes ("Föredragningslista" PE 389.455/OJJE).
19 Avslutande av sammanträdet
Sammanträdet avslutades kl. 24.00.
Harald R
ømer
Gérard Onesta
Generalsekreterare
Vice talman
NÄRVAROLISTA
Följande skrev på:
Adamou
Agnoletto
Aita
Albertini
Ali
Allister
Alvaro
Anastase
Andersson
Andrejevs
Andria
Andrikienė
Angelilli
Antoniozzi
Arif
Arnaoutakis
Ashworth
Assis
Athanasiu
Atkins
Attard-Montalto
Attwooll
Aubert
Audy
Auken
Ayuso
Baco
Badia i Cutchet
Bărbuleţiu
Barón Crespo
Batten
Battilocchio
Batzeli
Bauer
Beaupuy
Beazley
Becsey
Belder
Belet
Belohorská
Bennahmias
Beňová
Berend
Berès
van den Berg
Berlinguer
Berman
Bielan
Birutis
Bliznashki
Blokland
Bloom
Bobošíková
Böge
Bösch
Bonde
Bono
Bonsignore
Booth
Borghezio
Borrell Fontelles
Bourlanges
Bourzai
Bowis
Bowles
Bozkurt
Bradbourn
Braghetto
Brejc
Brepoels
Breyer
Březina
Brie
Brok
Budreikaitė
van Buitenen
Buitenweg
Bulfon
Bullmann
van den Burg
Buruiană-Aprodu
Bushill-Matthews
Busk
Buşoi
Busquin
Busuttil
Buzek
Calabuig Rull
Callanan
Camre
Capoulas Santos
Cappato
Carlotti
Carnero González
Casa
Casaca
Casini
Caspary
Castex
Castiglione
del Castillo Vera
Catania
Cavada
Cederschiöld
Cercas
Chatzimarkakis
Chervenyakov
Chichester
Chiesa
Chmielewski
Christensen
Christova
Chruszcz
Claeys
Clark
Cocilovo
Coelho
Cohn-Bendit
Corbett
Corbey
Correia
Coşea
Costa
Cottigny
Coûteaux
Cramer
Corina Creţu
Gabriela Creţu
Crowley
Marek Aleksander Czarnecki
Ryszard Czarnecki
Daul
Davies
De Blasio
Degutis
Dehaene
De Keyser
Deprez
Descamps
Désir
Deß
Deva
De Veyrac
De Vits
Díaz de Mera García Consuegra
Dičkutė
Didžiokas
Díez González
Dillen
Dimitrakopoulos
Konstantin Dimitrov
Martin Dimitrov
Philip Dimitrov Dimitrov
Dîncu
Dobolyi
Dombrovskis
Doorn
Douay
Dover
Doyle
Drčar Murko
Duchoň
Dührkop Dührkop
Duff
Duka-Zólyomi
Dumitrescu
Ebner
Ek
El Khadraoui
Elles
Esteves
Estrela
Ettl
Jill Evans
Jonathan Evans
Robert Evans
Färm
Fajmon
Farage
Fava
Ferber
Fernandes
Fernández Martín
Anne Ferreira
Elisa Ferreira
Figueiredo
Fjellner
Flasarová
Flautre
Florenz
Foltyn-Kubicka
Fontaine
Ford
Fourtou
Fraga Estévez
Frassoni
Freitas
Friedrich
Fruteau
Gahler
Gál
Gaľa
Galeote
Ganţ
Gargani
Gaubert
Gauzès
Gawronski
Gebhardt
Gentvilas
Geremek
Geringer de Oedenberg
Gewalt
Gibault
Gierek
Giertych
Gill
Gklavakis
Glante
Glattfelder
Goebbels
Goepel
Golik
Gomes
Gomolka
Gottardi
Goudin
Grabowska
Grabowski
Graça Moura
Graefe zu Baringdorf
Gräßle
de Grandes Pascual
Griesbeck
Gröner
de Groen-Kouwenhoven
Groote
Grosch
Grossetête
Gruber
Guardans Cambó
Guellec
Guerreiro
Guidoni
Gurmai
Gutiérrez-Cortines
Guy-Quint
Gyürk
Hänsch
Hall
Hammerstein
Hamon
Handzlik
Hannan
Harangozó
Harbour
Harkin
Harms
Hassi
Hatzidakis
Haug
Hazan
Hedh
Hegyi
Hellvig
Helmer
Henin
Hennicot-Schoepges
Hennis-Plasschaert
Herczog
Herranz García
Herrero-Tejedor
Hieronymi
Hökmark
Holm
Honeyball
Hoppenstedt
Horáček
Howitt
Hudacký
Hudghton
Hughes
Hutchinson
Iacob-Ridzi
Ibrisagic
in 't Veld
Isler Béguin
Itälä
Iturgaiz Angulo
Jackson
Jäätteenmäki
Jałowiecki
Janowski
Jarzembowski
Jeggle
Jensen
Jöns
Jørgensen
Jonckheer
Jordan Cizelj
Juknevičienė
Kacin
Kaczmarek
Kallenbach
Kamall
Kamiński
Karas
Karatzaferis
Karim
Kaufmann
Kauppi
Kazak
Tunne Kelam
Kelemen
Kilroy-Silk
Kindermann
Kinnock
Kirilov
Kirkhope
Klamt
Klaß
Klich
Knapman
Koch
Koch-Mehrin
Kohlíček
Konrad
Kónya-Hamar
Korhola
Kósáné Kovács
Koterec
Kozlík
Krahmer
Krasts
Kratsa-Tsagaropoulou
Krehl
Kreissl-Dörfler
Kristovskis
Krupa
Kuc
Kudrycka
Kuhne
Kułakowski
Kušķis
Kusstatscher
Kuźmiuk
Lagendijk
Laignel
Lamassoure
Lambert
Lambrinidis
Lambsdorff
Lang
De Lange
Langen
Langendries
La Russa
Lavarra
Lax
Lechner
Le Foll
Lehideux
Lehne
Lehtinen
Leichtfried
Leinen
Jean-Marie Le Pen
Marine Le Pen
Le Rachinel
Lévai
Lewandowski
Liberadzki
Libicki
Lichtenberger
Lienemann
Liese
Liotard
Locatelli
Lombardo
López-Istúriz White
Losco
Louis
Lucas
Ludford
Lulling
Lundgren
Lynne
Lyubcheva
Maaten
McAvan
McCarthy
McMillan-Scott
Madeira
Maldeikis
Manders
Maňka
Erika Mann
Thomas Mann
Manolakou
Mantovani
Marinescu
Markov
Marques
Martens
David Martin
Hans-Peter Martin
Martinez
Martínez Martínez
Masiel
Mastenbroek
Mathieu
Matsakis
Matsouka
Mauro
Mavrommatis
Mayer
Medina Ortega
Meijer
Méndez de Vigo
Menéndez del Valle
Miguélez Ramos
Mihăescu
Mihalache
Mikko
Mikolášik
Millán Mon
Mölzer
Mohácsi
Moisuc
Montoro Romero
Moraes
Moreno Sánchez
Morgan
Morgantini
Morillon
Morţun
Moscovici
Mote
Mulder
Musacchio
Muscardini
Muscat
Musotto
Musumeci
Napoletano
Nassauer
Nattrass
Navarro
Newton Dunn
Nicholson
Nicholson of Winterbourne
Niebler
van Nistelrooij
Novak
Obiols i Germà
Öger
Özdemir
Olajos
Olbrycht
Onesta
Onyszkiewicz
Oomen-Ruijten
Ortuondo Larrea
Őry
Ouzký
Oviir
Paasilinna
Pack
Paleckis
Pannella
Panzeri
Papadimoulis
Paparizov
Papastamkos
Parish
Parvanova
Paşcu
Patrie
Pęk
Alojz Peterle
Petre
Pflüger
Pieper
Pīks
Pinheiro
Piotrowski
Pirker
Piskorski
Pistelli
Pittella
Pleštinská
Podestà
Podgorean
Podkański
Pöttering
Pohjamo
Poignant
Polfer
Pomés Ruiz
Popeangă
Portas
Posdorf
Posselt
Post
Prets
Vittorio Prodi
Protasiewicz
Purvis
Queiró
Quisthoudt-Rowohl
Rack
Radwan
Ransdorf
Rapkay
Rasmussen
Remek
Resetarits
Reul
Ribeiro e Castro
Riera Madurell
Ries
Riis-Jørgensen
Rivera
Rizzo
Rocard
Rogalski
Roithová
Romeva i Rueda
Rosati
Roszkowski
Roth-Behrendt
Rothe
Rouček
Roure
Rudi Ubeda
Rübig
Rühle
Rutowicz
Sacconi
Saïfi
Sakalas
Saks
Samaras
Samuelsen
Sánchez Presedo
dos Santos
Sârbu
Saryusz-Wolski
Savary
Savi
Schaldemose
Schapira
Scheele
Schenardi
Schierhuber
Schlyter
Olle Schmidt
Frithjof Schmidt
Schmitt
Schnellhardt
Schöpflin
Jürgen Schröder
Schroedter
Schuth
Schwab
Seeber
Seeberg
Segelström
Seppänen
Şerbu
Severin
Siekierski
Silva Peneda
Simpson
Sinnott
Siwiec
Škottová
Smith
Sofianski
Sommer
Søndergaard
Sonik
Sornosa Martínez
Sousa Pinto
Spautz
Speroni
Staes
Stănescu
Staniszewska
Starkevičiūtė
Šťastný
Stauner
Sterckx
Stevenson
Stihler
Stockmann
Stoyanov
Strejček
Strož
Stubb
Sturdy
Sudre
Sumberg
Surján
Susta
Svensson
Szabó
Szájer
Szejna
Szent-Iványi
Szymański
Tabajdi
Tajani
Takkula
Tannock
Tarabella
Tarand
Tatarella
Thomsen
Thyssen
Ţicău
Ţîrle
Titford
Titley
Toia
Toma
Tomczak
Toubon
Toussas
Trakatellis
Trautmann
Triantaphyllides
Trüpel
Turmes
Tzampazi
Uca
Ulmer
Vaidere
Vakalis
Vălean
Van Hecke
Van Lancker
Varela Suanzes-Carpegna
Vatanen
Vaugrenard
Veneto
Ventre
Veraldi
Vergnaud
Vernola
Vidal-Quadras
de Villiers
Virrankoski
Vlasák
Vlasto
Voggenhuber
Wagenknecht
Wallis
Walter
Watson
Henri Weber
Manfred Weber
Weiler
Weisgerber
Westlund
Wieland
Wiersma
Wijkman
Willmott
Wise
von Wogau
Bernard Wojciechowski
Janusz Wojciechowski
Wortmann-Kool
Wurtz
Yañez-Barnuevo García
Záborská
Zahradil
Zaleski
Zani
Zapałowski
Zatloukal
Ždanoka
Železný
Zieleniec
Zīle
Zimmer
Zingaretti
Zvěřina
Zwiefka
Microsoftdom gynnar konsumenterna, säger EP-ledamöter
Konkurrens
2007-09-20 - 17:56
Microsoft förlorar EU-konkurrensmål
Europeiska kommissionens framgång i konkurrensmålet mot Microsoft gynnar konsumenterna.
Domen välkomnas av flera Europaparlamentsledamöter eftersom den leder till ett större utbud på mjukvarumarknaden.
EU:s förstainstansrätt gick på kommissionens linje och slog fast att Microsoft har missbrukat sin dominerande ställning - 90 procent av mjukvaruindustrin.
Kommissionen krävde i mars 2004 Microsoft på 497 miljoner euro på böter.
Datajätten anklagas för att inte dela med sig information, så att andra företags program kan användas i Microsofts operativsystem Windows.
EU:s förstainstansrätt dömde i måndags (17 september) Microsoft.
Microsoft har nu två månader på sig att överklaga domen till EG-domstolen.
Konsumenternas valfrihet garanteras
Internationella handelsutskottets ordförande Helmuth Markov (Gruppen Europeiska enade vänstern/Nordisk grön vänster, Tyskland) välkomnar "alla domslut som hindrar att oligopol skapas.
Konsumenterna ska ha möjlighet att välja mellan olika produkter från olika tillverkare."
Beslutet garanterar "konsumenternas valfrihet och en rättvis konkurrens på IT-marknaden", sa hon.
Alain Lipietz (Gruppen De gröna/Europeiska fria alliansen, Frankrike), som sitter i utskottet för rättsliga frågor, ansåg att domen "är en stor seger för upprätthållandet av konkurrensrätten."
Inremarknadsutskottets vice ordförande Graf Alexander Lambsdorff (Gruppen Alliansen liberaler och demokrater för Europa, Tyskland) påpekade att domen var "en viktig seger för Europas konsumenter.
Den stärker konkurrensen på mjukvarumarknaden och sänder en klar signal till andra företag att EU konsekvent tillämpar sin konkurrenslagstiftning."
Vissa amerikanska reaktioner är inte lika positiva.
Thomas Barnett, chef för amerikanska justitiedepartements konkurrensenhet, sa att domen "kan hämma innovation" och på så sätt missgynna konsumenterna.
Kommer vi i framtiden att se fler domar mot utnyttjande av marknadsposition?
Exempelvis har det påpekats från vissa håll att samma argument kan användas mot Apples "ipod" och "itunes".
Redan nu kan emellertid Europas medborgare glädja sig åt att hela bötessumman från Microsoft går till EU:s gemensamma kassa.
20070920STO10523 EU:s förstainstansrätts dom mot Microsoft (engelska) Europaparlamentets utskott Europeiska kommissionen: konkurrens Microsofts reaktion (engelska)
SV
1
PHOTO
20070920PHT10521.jpg
SV
2
LINK
http://www.curia.europa.eu/en/actu/communiques/cp07/aff/cp070063en.pdf
SV
3
LINK
/activities/expert/committees.do?language=SV
SV
4
LINK
http://www.microsoft.com/presspass/press/2007/sep07/09-17Statement.mspx
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
EP-veckan 22-25 oktober 2007, Strasbourg
2007-10-31 - 16:53
EP-veckan 22-25 oktober 2007
Europaparlamentet beslutade att Salih Mahmoud Osman ska motta 2007 års Sacharovspris och att Vid himlens utkant av Fatih Akin får filmpriset Lux.
Resultaten från toppmötet i Lissabon välkomnades och Turkiet och afghanskt opium behandlades också.
20071019BRI11923
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-001-SV DOC XML V0//SV
Miljö
En mer hållbar användning av bekämpnings­medel
2007-10-31 - 16:53
Flygbesprutning förbjuds och buffertzoner ska finnas runt vattendrag.
Bostadsområden och rekreationsområden ska i princip hållas fria från bekämpningsmedel.
Bekämpningsmedel ökar jordbrukets avkastning och jordbruksprodukternas kvalitet och minskar arbetsinsatsen.
De har dessutom många användningsområden utanför jordbrukssektorn, alltifrån skydd av trä och textilier till skydd av folkhälsan.
Den nya lagstiftningen ska förbättra hälso- och miljöskyddet, gagna jordbruket, minska djurförsöken och öka konkurrensen mellan tillverkarna.
Ledamöterna ställer sig bakom substitutionsprincipen som säger att produkter i princip inte ska godkännas om de innehåller ämnen som skulle kunna ersättas med alternativa ämnen som är avsevärt säkrare för miljön och för djurs och människors hälsa.
Ämnen som betraktas som lågriskämnen ska godkännas för 15 år, godkännandet ska kunna förlängas, en eller flera gånger, för en period på högst 10 år och inte utan tidsbegränsning som kommissionen föreslår.
För ämnen där det finns säkrare alternativ bör godkännandet endast gälla i fem år och inte sju som kommissionen föreslår.
"Folk vill inte ha gift på sina tallrikar"
Parlamentet stöder kommissionen när det gäller förbud av cancerogena, reproduktionstoxiska och mutagena ämnen och ämnen som kan förorsaka endokrina störningar eller har toxikologisk betydelse för människor.
Till de förbjudna kategorierna ska man enligt ledamöterna även föra ämnen med utvecklingsmässiga, neurotoxiska och immuntoxiska risker.
- Folk inte vill ha gift på sina tallrikar, sade föredraganden under debatten.
Då så är nödvändigt ska ett acceptabelt dagligt intag (ADI), en godtagbar användarexponering (AOEL) och en akut referensdos (ARfD) fastställas.
Möjliga kombinerade effekter samt sårbarheten hos specifika befolkningsgrupper i riskzonen ska också beaktas.
Det föreslagna direktivet kommer att innehålla regler om:
– nationella handlingsplaner för att fastställa mål för minskning av faror, risker och beroendet av kemisk bekämpning för växtskydd,
– system för utbildning och information till distributörer och yrkesmässiga användare av bekämpningsmedel samt bättre information till allmänheten,
– regelbunden inspektion av spridningsutrustning,
– förbud mot flygbesprutning med möjlighet till undantag,
– särskilda åtgärder för att skydda vattenmiljön från att förorenas av bekämpningsmedel,
– fastställande av områden med kraftigt minskad eller ingen användning av bekämpningsmedel (jfr ramdirektivet för vatten, fågeldirektivet, habitatdirektivet m.fl.) eller för att skydda känsliga grupper,
– hantering och lagring av bekämpningsmedel samt deras förpackningar och rester,
– utveckling av standarder på gemenskapsnivå för integrerat växtskydd.
Parlamentet stöder idén om nationella handlingsplaner och anger att för andra än biologiska bekämpningsmedel och ämnen med låg risk ska kvantitativa mål för minskad användning, anges i form av ett index för behandlingsfrekvens.
Indexet för behandlingsfrekvens ska anpassas till de specifika förhållandena i varje medlemsstat.
För verksamma ämnen som inger mycket stora betänkligheter ska minskningsmålet vara en reducering på minst 50 procent i förhållande till indexet för behandlingsfrekvens beräknat för år 2005 före utgången av 2013 och för beredningar av bekämpningsmedel som klassificeras som giftiga eller mycket giftiga ska målet vara en minskning på minst 50 procent.
Utskottets krav på en 25-procentig allmän minskning inom fem år och en 50-procentig inom tio år föll.
När det gäller information till allmänheten kan medlemsstaterna välja att införa ett krav på att berörda grannar ska informeras om planerad besprutning.
För att skydda vattendrag föreslår kommissionen att man inrättar buffertzoner där bekämpningsmedel inte får användas eller lagras.
- Jag håller naturligtvis med om att en informationsplikt på 48 timmar före besprutning är opraktiskt, men att därav dra slutsatsen att vi inte behöver någon informationsplikt alls är inte rimligt.
Han sade att en annan viktig fråga gäller de s.k. cut off criteria för särskilt känsliga substanser.
- Vi måste vara konsekventa i förhållande till vårt beslut om den nya kemikalielagstiftningen Reach, där en av utgångspunkterna består i att fasa ut ämnen där tröskelvärden är svåra att etablera.
Det gäller riskerna hos ämnen som anses särskilt oroväckande och dessa ska inte komma i kontakt med livsmedel.
Wijkman fann i princip kommissionens förslag att försöka dela in Europa i zoner som är relativt lika vad gäller vegetationsförhållanden, klimat osv intressant.
Många av de mest miljö- och hälsofarliga ämnena har förbjudits, och den totala förbrukningen räknat i mängd aktiv substans har minskat kraftigt.
Kemisk bekämpning är trots detta fortfarande den helt dominerande växtskyddsmetoden i Sverige.
De nya, mer koncentrerade medlen innebär att man med mindre mängder kan bekämpa en lika stor areal som tidigare.
Kemikalieinspektionen har också de senaste åren genomfört en omregistrering av jordbrukets bekämpningsmedel, som lett till att drygt 80 av de hälso- och miljöfarligaste ämnena förbjudits helt.
Här har Sverige varit ett föregångsland och antalet tillåtna ämnen är idag lägre än i de flesta jämförbara länder.
Utrensningen har möjliggjorts av den lagfästa substitutionsprincipen, som innebär att kemiska medel kan totalförbjudas om det finns ett mindre farligt med motsvarande effekt.
I samband med omregistreringen har också de rekommenderade doserna för många medel justerats ned.
Tidigare rekommendationer låg ofta högre än vad som krävdes för full bekämpningseffekt.
Kravet på harmonisering av vilka medel som är tillåtna inom EU hotar den svenska situationen eftersom andra länder i EU inte har lika restriktiva regler.
Beslutsförfarande: Medbeslutande - 1:a behandlingen (***I)
Omröstning: 23.10.2007 Antagna texter Antagna texter
-//EP//TEXT TA P6-TA-2007-0445 0 NOT XML V0//SV
-//EP//TEXT TA P6-TA-2007-0444 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-COVER-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-002-SV DOC XML V0//SV
Miljö
Parlamentet kräver en ambitiös strategi för en hållbar användning av bekämpnings­medel
2007-10-31 - 16:53
Parlamentet anser att ambitionsnivån ska höjas ytterligare.
Uppmuntra till minskad användning
Europaparlamentet inser behovet av en europeisk rättslig ram för användningen av bekämpningsmedel eftersom gällande lagstiftning inte har räckt till för att minimera de faror och risker som bekämpningsmedel medför för hälsa och miljö.
Felanvändning, överanvändning och förgiftningsolyckor måste förebyggas och parlamentet välkomnar därför inrättandet av ett system för utbildning av yrkesmässiga användare av bekämpningsmedel.
Den globala uppvärmningen kommer sannolikt att leda till en ökad population av skadegörare och parlamentet efterlyser en undersökning av hur klimatförändringen påverkar jordbruksproduktionen, men också miljöskyddet.
Medlemsstaterna uppmanas att främja både jordbruk med liten användning av bekämpningsmedel och ekologiskt jordbruk samt att se till att yrkesmässiga användare av bekämpningsmedel går över till en miljövänligare användning av tillgängliga växtskyddsmetoder, där icke-kemiska växtskydds- och odlingsmetoder, exempelvis växelbruk och ogräsrensning, ges företräde framför systematisk användning av bekämpningsmedel.
Starkare koppling till hälsofrågor
Bättre information om möjliga miljö- och hälsorisker måste finnas anser ledamöterna och all fortsatt användning av bekämpningsmedel bör ske endast om försiktighetsprincipen respekteras.
De beklagar för övrigt att hälsoaspekten bara berörs flyktigt i den temainriktade strategin, trots att bekämpningsmedel kan ha ett samband med skador på immunförsvaret, endokrina störningar, neurotoxiska skador och cancer.
Bin och former för frukt och grönt
Ledamöterna uppmanar kommissionen att genast utvidga den temainriktade strategins räckvidd till att även omfatta biocidprodukter, eftersom dessa också medför risker för människors hälsa och miljön.
Bortskaffande av gamla lager
Europaparlamentet kräver att befintliga gemenskapsmedel ska användas för säkert bortskaffande av gamla bekämpningsmedel, med tanke på att mer än 200 000 ton bekämpningsmedel i EU ännu lagras såväl under jord som utomhus.
Föredragande: Irena BELOHORSKÁ (NI, SK)
-//EP//TEXT TA P6-TA-2007-0467 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-001-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-003-SV DOC XML V0//SV
Miljö
Bindande tak för bilavgaser ska vara 125 g koldioxid/km till 2015
2007-10-31 - 16:53
Parlamentet yrkar i ett initiativbetänkande på att koldioxidutsläppen från personbilar ska hållas under 125 g koldioxid/km från 2015.
Ett bindande tak bör fastställas eftersom bilindustrin misslyckats med att uppfylla sina frivilliga åtaganden.
Nästan en femtedel av koldioxidutsläppen i EU kommer från personbilar och mindre transportbilar.
Om vi gör detta på rätt sätt kan båda miljön, konsumenterna och bilindustrins framtid gagnas.
Parlamentet rekommenderar därför att varje tillverkare eller importör ska ha rätt att undanta 500 identifierade fordon per år från de uppgifter som används för att fastställa de genomsnittliga utsläppen.
Koldioxidkrediter Slutligen föreslår parlamentet att en ny stängd marknadsmekanism i form av ett system för minskningar av utsläppskvoter för koldioxid (CARS) ska införas den 1 januari 2011, så att tillverkare och importörer får böta utifrån hur mycket varje såld bil överskrider gränsvärdena för utsläpp.
Jag tror att det är marknadsföringen som påverkar konsumenternas efterfrågan.
Studier visar att en stor andel av utgifterna för marknadsföringen går till att framhäva bilens styrka, storlek och hastighet.
Europaparlamentet rekommenderar att obligatoriska och enhetliga minimikrav ska fastställas för den information som ska visas om bränsleekonomi (l/100 km) och koldioxidutsläpp (g/km) för nya bilar i allt marknadsförings- och reklammaterial och i visningshallar.
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-002-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-004-SV DOC XML V0//SV
Miljö
Rökfria arbetsplatser i Europa
2007-10-31 - 16:53
Parlamentet förespråkar i ett initiativbetänkande en rad restriktioner när det gäller rökning på offentliga platser och regler som ska göra det svårare för minderåriga att skaffa sig tobak och cigaretter.
Det initiativbetänkande av Karl-Heinz FLORENZ (EPP-ED, DE) som parlamentet antagit är ledamöternas svar på kommissionens grönbok om grönboken ”Mot ett rökfritt Europa: policyalternativ på EU-nivå.
Minst 650 000 människor dör årligen i EU på grund av rökning och cirka 80 000 människor uppskattas dö till följd av passiv rökning.
Tobaksrök skadar bland annat luftvägarna och orsakar irriterade slemhinnor, hosta, heshet, andnöd, nedsatt lungfunktion, astma, lunginflammationer, bronkit och kronisk obstruktiv lungsjukdom.
Parlamentet välkomnar kommissionens grönbok som utgångspunkt för en ansvarsfull europeisk politik, men vill att man går längre.
Det upprepar sin uppmaning till kommissionen att snarast möjligt klassificera tobaksrök i miljön som en cancerogen ämnesblandning av klass 1 enligt direktivet om farliga ämnen från 1967.
Medlemsstaterna uppmanas att inom två år införa ett generellt rökförbud på alla slutna arbetsplatser, inbegripet arbetsplatser i serveringsbranschen, samt i alla slutna offentliga lokaler och kollektiva färdmedel i EU.
Parlamentet uppmanar kommissionen, om de nämnda målen inte uppnås av alla medlemsstater, att senast 2011 överlämna ett förslag till parlamentet och rådet med bestämmelser om skydd av icke rökare på området för arbetarskydd samt att i detta sammanhang erkänna medlemsstaternas gällande nationella bestämmelser.
E uropaparlamentet uppmanar kommissionen att undersöka vilka hälsorisker som är förknippade med användning av snus och vilken inverkan denna användning har på cigarettkonsumtionen.
Kommissionen uppmanas också att till 2008 lägga fram ett förslag om ändring av direktiv 2001/37/EG (”tobaksvarudirektivet”) så att detta omfattar ett omedelbart förbud mot alla beroendeförstärkande tillsatsämnen, samt mot alla de tillsatsämnen som man på grundval av befintliga toxikologiska uppgifter har identifierat som cancerframkallande, mutagena eller reproduktionstoxiska, samt en rad skyldigheter om uppgiftslämning och delade hälsokostnader för tillverkarna.
Beviljande av tillstånd att ställa upp cigarettautomater bör endast ges om dessa görs otillgängliga för ungdomar under 18 år.
Tobaksvaror ska inte kunna köpas genom självbetjäning i butiker och distansförsäljning (t.ex. via Internet) av tobaksvaror till ungdomar under 18 år bör förhindras.
Medlemsstaterna bör åta sig att till 2025 minska rökning bland ungdomar med minst 50 procent.
Ledamöterna föreslår också att en EU omfattande högsta minimiskattenivå för alla tobaksprodukter införs och att hårdare kontroller görs mot tobakssmuggling.
Kommissionen uppmanas också att till 2008 lägga fram ett förslag om ändring av direktiv 2001/37/EG (”tobaksvarudirektivet”) så att detta omfattar ett omedelbart förbud mot alla beroendeförstärkande tillsatsämnen, samt mot alla de tillsatsämnen som man på grundval av befintliga toxikologiska uppgifter har identifierat som cancerframkallande, mutagena eller reproduktionstoxiska, samt en rad skyldigheter om uppgiftslämning och delade hälsokostnader för tillverkarna.
– 650 000 personer dör av rökning varje år, och 80 000 avlider årligen av passiv rökning, endast i EU.
Bara dessa svarta siffror ger oss en klar bild av att vi måste göra allt vi kan för att motarbeta rökningen, sade Jens HOLM (GUE/NGL, SE).
Holm konstaterade att föredragande Florenz lagt fram en serie bra åtgärdsförslag, exempelvis skärpning av befintlig lagstiftning, avskräckande märkning på cigarettpaket, åtgärder för att förhindra att ungdomar börjar röka, åtgärder för att hjälpa rökare som vill bli kvitt sitt beroende, men påpekade att han samtidigt är motståndare till att flytta upp mer makt till EU på folkhälsoområdet.
- Minst tio EU-länder har redan idag någon form av förbud mot rökning på restauranger och krogar.
Det började med Irland 2004 och spred sig snabbt vidare till Sverige, Italien, Finland, Malta, Belgien osv. och många fler är på gång.
Ska vi nu stoppa denna process av goda exempel och vänta in central EU-lagstiftning?
Nej, det tycker jag inte, utan låt de goda exemplen fortsätta att sprida sig.
Holm lyfte också fram EU:s subventioner av tobaksodlingar.
– Finns det inte risk för att vi tar med den ena handen och att vi ger med den andra?
Å den ena sidan uppmanar vi människor att sluta röka, å den andra sidan fortsätter EU att subventionera tobaksodlingar på över en 1 miljard euro årligen.
Dessa subventioner måste förstås snarast avvecklas, sade Holm.
Även Carl SCHLYTER (De gröna/EFA, SE) berörde EU:s tobakssubventioner och sade att alla subventioner måste avvecklas.
– Vi måste se till att våra tobaksbolag inte förstör arbetet mot rökning genom en massiv marknadsföring i u-länderna, påpekade han.
Enligt Schlyter är det också viktigt att tillsatserna i cigaretter nämns i betänkandet.
Därför väntar vi nu på ett snabbt förslag från kommissionen för att bli av med dessa hemska tillsatser som gör cigaretter ännu värre.
Christofer FJELLNER (EPP-ED, SE) påpekade att han i grunden är skeptisk till idén att EU ska förbjuda rökning på allmän plats i hela unionen.
– Även den som är för denna typ av rökförbud måste se problemet med att vi gör det på EU-nivå.
Det finns dock saker som vi kan göra här i EU för att minska skadorna av tobaksrök i hela Europa, sade han.
– Vi kan t.ex. avskaffa EU:s obegripliga förbud mot svenskt snus.
Jag kommer återigen med en dåres envishet att ta tillfället i akt och påpeka den svenska erfarenheten.
Vi har den lägsta andelen rökare i hela Europa, vi har den minsta andelen av alla tobaksrelaterade sjukdomar i hela Europa och vet ni vad?
Vi har trots detta ungefär samma förbrukning av tobak som resten av Europa, men vi förbrukar snus istället för cigaretter.
Faktum är att om resten av Europa skulle ersätta cigaretter med snus i samma utsträckning som vi har gjort i Sverige så skulle 200 000 européer slippa lugncancer varje år.
Därför tycker jag att det är omoraliskt att fortsätta blunda, sade Fjellner avslutningsvis.
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-003-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-005-SV DOC XML V0//SV
Mänskliga rättigheter
Sacharovpriset 2007 till Salih Mahmoud Osman
2007-10-31 - 16:53
Den sudanesiske människorättsadvokaten Salih Mahmoud Osman får Europaparlaments Sacharovpris för tankefrihet.
Namnet på årets Sacharovpristagare tillkännagavs i Europaparlamentets kammare i Strasbourg torsdagen den 25 oktober, kl. 11.30 av Europaparlamentets talman Hans-Gert PÖTTERING som motiverade valet så här.
Europaparlamentet delar varje år sedan 1988 ut Sacharovpriset för tankefrihet till individer och organisationer som har gjort anmärkningsvärda insatser mot förtryck, intolerans och orättvisa.
Priset är ett sätt för Europaparlamentet att främja och uppmärksamma kampen för mänskliga rättigheter och demokrati i världen.
I år sker prisutdelningen den 11 december.
Salih Mahmoud Osman
Salih Mahmoud Osman är advokat och människorättsaktivist.
Han arbetar för en sudanesisk organisation mot tortyr - "Sudan Organisation Against Torture"- som erbjuder kostnadsfri rättshjälp för personer som drabbats av människorättsövergrepp och stridigheterna i Sudan.
Personer i hans familj har torterats och dödats till följd av hans engagemang.
Han har varit ledamot i Sudans parlament, men har fråntagits sitt mandat.
Förteckning över tidigare Sacharovpristagare
2006 - Alexander Milinkevitj
2005 - Kvinnor i vitt, Hauwa Ibrahim och Reportrar utan gränser
2004 - Zhanna Litvina, ordförande för vitryska journalistförbundet
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-004-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-006-SV DOC XML V0//SV
Budget
Parlamentets första behandling av EU:s budget för 2008 klar
2007-10-31 - 16:53
Rådet vill sänka beloppet till 0,95 %.
Anslagen för Galileo och för Europeiska tekniska institutet höjs avsevärt och de ursprungliga anslagen för satsningar inom Lissabonstrategin återinförs.
I EU:s budget för 2008 utgör jordbrukspolitiken för första gången mindre än hälften av utgifterna.
Europaparlamentet har behandlat kommissionens budget i ett betänkande av Kyösti VIRRANKOSKI (ALDE, FI) som antogs med 487 röster för, 73 emot och 15 nedlagda och ett betänkande av Ville ITÄLÄ (EPP-ED, FI) om övriga institutioner som antogs med 499 röster för, 24 emot och 42 nedlagda.
Ledamöterna var inte nöjda med budgetens storlek och vill se en total ökning av budgeten för nästa år.
Ökade medel föreslogs bland annat till Galileo, Europeiska tekniska institutet och för att finansiera vissa utrikespolitiska prioriteringar som Kosovo och Palestina.
Det totala beloppet bör enligt parlamentet uppgå till 124 201 365 130 euro i betalningsbemyndiganden och 129 693 891 505 euro i åtagandebemyndiganden.
När det gäller betalningsbemyndiganden anser Europaparlamentet att ett belopp motsvarande 0,95 procent av EU:s BNI är otillräckligt med tanke på de politiska utmaningar som EU står inför.
Parlamentet vill öka den totala betalningsnivån till ett belopp motsvarande 0,99 procent av EU:s BNI.
Parlamentets allmänna linje är att återställa utgiftstaken till den nivå som anges i det preliminära förslaget till budget och utnyttja de ramar som ges i det interinstitutionella avtalet för perioden 2007-2013.
Anslagsfördelning per rubrik
1.
1a.
Sammanhållning för tillväxt och sysselsättning - 42,447 miljarder euro i betalningsbemyndiganden
3a Frihet, säkerhet och rättvisa - 533 miljoner euro i betalningsbemyndiganden
EU som global partner - 8,132 miljarder i betalningsbemyndiganden
Reserver - 206, 6 miljoner
Varken ledamöterna eller kommissionen är nöjda med det belopp på 151 miljoner euro i åtagandebemyndiganden som rådet föreslagit i sin första behandling av budgeten.
Kommissionen lade fram en ny finansieringsplan för Galileo i september som bl.a. bygger på en omfördelning av outnyttjade medel inom jordbrukspolitiken.
Ledamöterna anser att man bör höja de åtagandebemyndiganden som föreslagits av rådet för Galileo och EIT från 739 miljoner euro till totalt 890 miljoner euro för 2008 (varav 400 miljoner i betalningsbemyndiganden).
Ledamöterna anser att detta är nödvändigt om projektet ska kunna fullföljas enligt utsatt tidsplan.
Parlamentet menar att projektet måste finansieras helt med gemenskapsmedel, eftersom risken är att hela projektet går om intet om erforderliga medel saknas.
För att finansiera EIT och Galileo yrkar ledamöterna på en översyn av den fleråriga budgetplanen för 2007-2013.
Om rådet inte kan övertygas, finns ett ändringsförslag som säger att anslagen för Galileo ska föras till det sjunde ramprogrammet för forskning.
Europaparlamentet motsätter sig de nedskärningar som rådet föreslagit i många budgetposter under denna budgetramsrubrik.
Parlamentet återinför det preliminära budgetförslaget på många ställen, men konstaterar att rådet kommer att ha sista ordet när det gäller dessa poster eftersom de avser obligatoriska utgifter enligt fördragen.
Parlamentet begär att flexibilitetsmekanismen används till ett belopp av 87 miljoner euro för andra prioriteringar, bland annat Kosovo och Palestina.
Således skulle det ursprungliga beloppet på 200 miljoner euro för GUSP kvarstå, eftersom de 40 miljoner euro som skulle kunna frigöras exakt motsvarar den sänkning med 20 % för GUSP som parlamentet förordar.
5.
Europaparlamentets fastställdes i omröstningen till 1 452 miljoner euro.
Debatt
-//EP//TEXT TA P6-TA-2007-0474 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-005-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-007-SV DOC XML V0//SV
Europeiska rådet
Ledamöterna nöjda med resultaten från Lissabon
2007-10-31 - 16:53
Europaparlamentet har den 23 oktober 2007 debatterat resultaten från det informella Europeiska rådet i Lissabon den 18-19 oktober med det portugisiska ordförandeskapet och kommissionen.
Stats- och regeringscheferna träffade en slutgiltig uppgörelse om det nya ändringsfördraget och om antalet platser i Europaparlamentets som fastställdes till 751.
Europaparlamentets talman Hans-Gert PÖTTERING välkomnade inledningsvis resultaten från toppmötet och överenskommelsen om det nya fördraget.
Han betonade att utan Europaparlamentet och dess stöd under hela processen hade EU inte nått ända fram.
Han berörde Ioannina-klausulen som utgjort en av de största stötestenarna.
Socrates preciserade att regeringskonferensen även antog en förklaring som förtydligar den befogenhetsuppdelning mellan union och medlemsstaterna som fastsälls i fördragen.
Socrates påminde om att det nya fördraget, Lissabonfördraget, kommer att undertecknas den 13 december i Lissabon och han gladde sig över att tidsplanen har kunnat respekteras.
- Vi har ett nytt fördrag som löser EU:s kris och banar väg för framtiden.
Europaparlamentets befogenheter och de nationella parlamentens inflytande stärks vilket ökar demokratin.
Rådets beslutsprocesser förbättras, främst på området rättvisa, säkerhet och frihet, sade han vidare och framhöll den rättsliga inramning som det europeiska medborgarskapet får genom stadgan för de grundläggande rättigheterna.
Socrates tackade ledamöterna, talmannen och de tre observatörerna vid regeringskonferensen för deras stöd och konstruktiva bidrag.
Han sade sedan att andra dagen av toppmötet ägnades den externa dimensionen av Lissabonstrategin.
Klimatförändringarna behandlades och han sade att stats- och regeringscheferna varit eniga om att EU har alla förutsättningar och därmed ett särskilt ansvar när det gäller kampen för att skydda miljön och motverka klimatförändringarna.
Kommissionen hade två oeftergivliga villkor - man kunde inte acceptera en mindre ambitiös text än Nicefördraget och kommissionens roll som motor fick inte ifrågasättas.
Barroso berörde sedan Lissabonstrategin och dess externa aspekter och EU:s ledande roll när det gäller en hållbar utveckling och en hållbar energipolitik.
Han berörde också det möte som hållits på EU-nivå samma dag som toppmötet mellan arbetsmarknadens parter där man enats om att acceptera begreppet "flexicurity".
Politiska grupper
Joseph DAUL (EPP-ED, FR) sade att han själv och gruppen var väldigt nöjda med Tysklands och Portugals ordförandeskap, trots att de egentligen skulle vilja ha haft en mer ambitiös text.
- Det väsentliga är innehållet, som är bra, trots den opraktiska förpackningen.
Medborgarnas förväntningar bemöts, nu måste vi förklara innehållet och dess fördelar och hur parlamentets befogenhet stärks, bl.a. i fråga om invandring och rättsliga och inrikes frågor.
En slags utrikesminister kommer också att finnas som ska samordna den gemensamma utrikes- och säkerhetspolitiken, gladde han sig.
EU måste agera konsekvent i internationella frågor även på handelsområdet, sade han.
Vi fick mindre än konstitutionen men mer än Nicefördraget och vi stöder fördragstexten.
Graham WATSON (ALDE, GB) gladde sig också över att fördraget undertecknats.
Det blir mindre vetorätt och flera andra förbättringar även om texten inte är lättläst.
EU kommer bättre att kunna bemöta globaliseringens utmaningar.
Ratificeringsprocessen blir ett tillfälle att bättre involvera medborgarna.
- De gröna kommer att uppriktigt förklara för- och nackdelar med fördraget för att upplysa medborgarna men vi hoppas att fördraget ratificeras som ett första steg på vägen mot något bättre på sikt.
Nigel FARAGE (IND/DEM, GB) sade det inte var första gången som kommissionen och rådet slår sig för bröstet i kammaren och betonar hur framgångsrikt EU är och hur bra ekonomin går och att full sysselsättning snart råder.
Låt oss hoppas att de kräver folkomröstningar.
Det är ett avskyvärt beteende, ansåg han, och hoppades på folkomröstning i Storbritannien.
- Är det en för viktig text för att man ska konsultera befolkningen?
Tvärtom är den just så viktig att den förtjänar att folket godkänner den först.
EU måste garantera grundläggande fri- och rättigheter om medborgarnas förtroende för EU ska bibehållas.
Elmar BROK (EPP-ED, DE) menade att det rörde sig om ett genombrott för demokratin.
Europaparlamentet blir medlagsstiftare i 95 % av lagstiftningen i EU.
Parlamentet kommer också att välja kommissionens ordförande inte längre bara godkänna honom eller henne.
Den tredje pelaren som rör inrikes och rättsliga frågor kommer att omfattas av medbeslutandeförfarandet.
Brok varnade avslutningsvis för att övergångarna mellan ett fördrag till ett annat inte får innebära möjligheter för rådet att rucka på den institutionella balansen.
Han betonade att talmannens rätt att rösta som en av de 751 folkvalda ledamöterna efter 2009 inte ifrågasätts.
Han berörde också tillsättningen av viktiga ämbeten och parlamentets roll vid val och utnämningar.
Alla principer har bibehållits i texten även om utformningen är mindre lyckad.
De vill inskränka EU:s befogenheter såväl vad gäller den gemensamma utrikes- och säkerhetspolitiken som samarbetet inom rättsliga och inrikes frågor.
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-006-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-008-SV DOC XML V0//SV
Kultur
Filmen Vid himlens utkant får Europa­parlamentets Luxpris
2007-10-31 - 16:53
Den tysk-turkiska filmen Vid himlens utkant av Fatih Akin tilldelas den 24 oktober 2007 Europaparlamentets nya filmpris Lux.
Den tyska skådespelerskan Hanna Schygulla, som innehar en av huvudrollerna i filmen, mottog priset i kammaren i närvaro och ledamöterna och representanter från de övriga nominerade filmerna.
Den tyska skådespelerskan Hanna Schygulla, som representerade den vinnande filmen, mottog priset i kammaren i närvaro av ledamöterna och representanter för de övriga filmer som konkurrerat om priset.
- Femtio år efter att Romfördraget undertecknades delar Europaparlamentet för första gången ut sitt nyinstiftade filmpris Lux.
Med vårt filmpris och valet av film vill vi varje år belysa utvecklingen i Europa och framhålla det europeiska skapandet, inledde talmannen ceremonin.
Prisstatyetten åkallar Babels torn och symboliserar språklig mångfald.
Men vi vill vända på den trend som uppstod i den bibliska berättelsen om byggandet av Babels torn och visa att språklig mångfald fungerar.
Vi vill med priset bidra till denna mångfald och gör dessutom filmen möjlig att ses för personer med nedsatt hörsel.
Hanns Schygulla mottog statyetten och sade:
- Det gläder mig mycket att man i Europaparlamentet talar om film idag.
Jag tackar å hela filmbranschens vägnar för att ni instiftat detta pris.
Hon tackade även å regissören Fatih Akins vägnar, som bad om ursäkt för att han inte kunde närvara.
Lux betyder ljus och utan ljus ingen film, fortsatte hon.
Ni har valt en film som ger hopp, men inte blint hopp.
Våld och konflikter skildras också, försoning och förståelse är dock möjligt.
De övriga två filmer som Europaparlamentets ledamöter sett och röstat om var
- 4 månader, 3 veckor och 2 dagar av Cristian Mungiu och
För att stödja europeisk film lanserar Europaparlamentet i år ett filmpris kallat Lux (ljus) som syftar till en bättre spridning av europeisk film över landsgränser och språkbarriärer.
Filmpriset Lux har som mål att främja européernas kunskap om Europa genom att förbättra deras möjligheter att se varandras filmer.
Europaparlamentet bidrar konkret genom att bryta språkbarriärer eftersom den film som utses till vinnare kommer att få textning på EU:s officiella 23 språk finansierad.
Dessutom förses originalversionen med en textning som är anpassad för döva och hörselskadade personer och med hjälpmedel för personer med nedsatt syn.
Europaparlamentets kulturutskott har utsett en jury på 17 personer verksamma inom filmbranschen.
Juryn fick i uppdrag att utnämna tre filmer, varav vinnaren sedan röstats fram av Europaparlamentet ledamöter:
Mellan den 1-18 oktober 2007 visades varje film nio gånger i Europaparlamentets lokaler i Bryssel.
Alla ledamöter som sett samtliga tre filmer i Europaparlamentet eller någon annanstans har kunnat rösta.
Film är ett universalt medium och en spegel av den värld vi lever i.
I EU är 70 procent av de filmer som ses amerikanska, 20 procent är nationella filmer och endast 10 kommer från andra europeiska länder.
I USA svarar europeisk film endast för 4,6 % av marknaden.
Nio av tio filmer som faktiskt distribueras i ett annat land i EU än ursprungslandet är beroende av stöd från EU-programmet Media.
Från den 24.10.2007
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-007-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-009-SV DOC XML V0//SV
Energi
EU fortfarande beroende av konventionella energikällor
2007-10-31 - 16:53
Ledamöterna efterlyser i ett initiativbetänkande om konventionell energi säkrare, effektivare och mer hållbara metoder för att producera energi inom EU.
Fossila energikällor kommer enligt alla prognoser att utgöra en central beståndsdel av EU:s energimix även 2020 och därefter, påminner ledamöterna i ett initiativbetänkande av Herbert REUL (EPP-ED, DE) som antogs med röstsiffrorna .
Ledamöterna betonar att man för att tillgodose grundbehoven inte kan avstå från kärnenergi i Europa på medellång sikt, eftersom kärnenergin är en viktig del av kraftförsörjningen i 15 av 27 medlemsstater, och därmed är viktig för hela EU där den tillhandahåller en tredjedel av elförsörjningen.
Kärnkraften utgör enligt ledamöterna den största koldioxidfattiga energikällan i Europa och de betonar dess potentiella roll i klimatskyddet.
Finland, Frankrike, Bulgarien, Rumänien, Slovakien, Litauen (i samarbete med Lettland och Estland), Förenade kungariket, Polen och Tjeckien håller enligt betänkandet på att bygga, planerar att bygga eller undersöker möjligheten att bygga nya kärnkraftverk.
För att nå de utsläppsmål som EU ställt upp för att motverka klimatförändringarna måste medlemsstaterna öka FoU-insatserna på energiområdet, framför allt i syfte att förbättra effektiviteten i energiproduktion och energiförsörjning, öka miljövänligheten, göra befintlig teknik säkrare, utveckla lagringstekniken i samband med förnybara energikällor och utveckla nya generationer av kärnreaktorer och ny energiteknik, inklusive kärnfusion, kräver ledamöterna.
Andris PIEBALGS, kommissionär för energifrågor, som talade i debatten före omröstningen, sade även han att det kommer att blir svårt för EU att uppnå sina utsläppsmål om man inte använder kärnenergin.
Tekniska, miljömässiga och rättsliga frågor om lagring av koldioxid är utmaningar som endast kan klargöras genom forskningsinsatser och politiska initiativ, anser ledamöterna.
Det är dock viktigt att CCS-anordningar så tidigt som det är praktiskt möjligt anpassas till kraftverk som drivs med fossila bränslen.
Piebalgs uppgav att kommissionen planerar att lägga fram ett lagstiftningsförslag om dessa tekniker.
- Målet är att det i EU till 2015 ska finnas flera storskaliga demonstrationsanläggningar och att tekniken ska kunna användas 2020.
Europaparlamentet framhåller i betänkandet den betydande potential för energi som framställts från biomassa.
Kommissionen uppmanas vidare att stödja syntetisk bränsleteknik med tanke på dess potential att öka energiförsörjningstryggheten och minska utsläppen från vägtransportsektorn i EU.
Ledamöterna varnar också för ett ensidigt beroende av vissa leverantörer eller leveranssätt när det gäller gas och betonar betydelsen av kondenserad naturgas för diversifiering av gasimporten.
Oljan stod för den största andelen (37,2 procent), åtföljd av gas (23,9 procent) och kol (17,9 procent).
-//EP//TEXT TA P6-TA-2007-0468 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-008-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-010-SV DOC XML V0//SV
Yttre förbindelser
Turkiet - den nya regeringens reformåtaganden välkomnas
2007-10-31 - 16:53
Europaparlamentet välkomnar i en resolution valresultaten och den nya regeringens starka engagemang för fortsatta reformer.
Det påminner dock om att det finns områden där mer framsteg behövs, i synnerhet när det gäller konstitutionella reformer och spänningarna vid gränsen mot norra Irak.
Turkiet debatterades också med rådet och kommissionen i plenum.
Parlamentet har antagit en resolution av Ria OOMEN-RUIJTEN (EPP-ED, NL) om förbindelserna mellan EU och Turkiet inför kommissionens kommande framstegsrapport som väntas den 7 november 2007.
Anslutningsförhandlingarna inleddes för ganska exakt två år sedan.
Ledamöterna välkomnar att fria och rättvisa val genomfördes och gläder sig över att Turkiets nya regering förbundit sig att påskynda reformprocessen så att man uppfyller åtagandena i partnerskapet för anslutning.
Regeringens planer på att anta en civil författning som bättre skyddar grundläggande mänskliga fri- och rättigheter ses också som mycket positivt.
Parlamentet välkomnar den turkiska regeringens ansträngningar att anpassa sig till EU:s energilagstiftning.
Det förespråkar ett stärkt energisamarbete mellan EU och Turkiet och uppmanar Turkiet att ansluta sig till den europeiska energigemenskapen.
Turkiet utgör en viktig länk när det gäller främst gasleveranser till EU.
Politiska reformer
Ledamöterna fördömer starkt mordet på Hrant Dink och Andrea Santoro och betonar att brådskande åtgärder måste vidtas för att bekämpa alla former av extremism och våldshandlingar med politiska förtecken.
För övrigt påminner parlamentet om att alla Köpenhamnskriterier måste vara helt uppfyllda för att man ska få ansluta sig till EU.
Varje anslutning är dessutom beroende av unionens integrationsförmåga, i enlighet med slutsatserna från Europeiska rådets möte i december 2006.
Ett ändringsförslag med en vädjan till Turkiet att erkänna folkmordet på armenierna, i överensstämmelse med parlamentets resolution från september 2005 om inledandet av förhandlingar med Turkiet förkastades.
Europaparlamentet fördömer starkt de våldshandlingar som PKK och andra terroristgrupper gjort sig skyldiga till på turkisk mark.
Parlamentet uttrycker sin solidaritet med Turkiet i dess kamp mot terrorismen och upprepar sin uppmaning till PKK om att utlysa ett omedelbart och ovillkorligt eldupphör och respektera det.
Parlamentet understryker behovet att gå vidare i kampen mot terrorismen på ett sätt som står i proportion till den aktuella hotbilden och som till fullo är förenligt med internationella rättsliga instrument och standarder.
Parlamentet understryker att det aldrig finns någon ursäkt för våld mot civila.
Europaparlamentet är djupt bekymrat över konsekvenserna av eventuella gränsöverskridande militära åtgärder från de turkiska styrkornas sida i norra Irak.
Turkiet och Irak uppmanas att utöka det militära och polisiära samarbetet för att effektivt förhindra terroristverksamhet från norra Irak och därmed minska spänningarna vid den turkisk-irakiska gränsen.
Parlamentet uppmanar rådet att verka för ett konkret samarbete mellan Turkiet och den kurdiska regionala regeringen i Irak, som måste påta sig sitt ansvar att förhindra terroristattacker från norra Irak.
Ledamöterna välkomnar dialogen mellan det civila samhället i EU och Turkiet och uppmanar kommissionen att informera om de insatser som gjorts i detta sammanhang.
Kommissionen uppmanas att vara mer närvarande i de olika regionerna i Turkiet och att ge riktat stöd till det civila samhället.
Parlamentet välkomnar att det inrättats ett instrument för ekonomiskt stöd för att uppmuntra den ekonomiska utvecklingen i det turkcypriotiska samhället.
Kommissionen uppmanas att lägga fram en särskild rapport om detta instruments effektivitet.
Kommissionen
Olli REHN, kommissionär för EU:s utvidgning, välkomnade valen i Turkiet.
Han konstaterade att Turkiet har genomlevt en svår period med en konstitutionell kris och politiska spänningar.
Rehn påpekade att Turkiet måste reformera paragraf 301 (om yttrandefriheten) i brottsbalken samt förbättra religionsfriheten i landet.
– Kvinnornas situation i landet, fackliga organisations situation och kampen mot korruption är andra områden som måste förbättras, sade Rehn.
Rehn kommenterade också den aktuella situationen och attackerna från PKK och konstaterade att landet oavbrutet ställs inför gränsöverskridande terrorattacker från PKK.
– Vi fördömer dessa terrorattacker, poängterade Rehn.
Föredragande
– Resolutionen tar upp de framsteg som uppnåtts men den beskriver också det som inte uppnåtts.
Vi har stora förväntningar på den nya turkiska regeringen, sade föredragande Ria OOMEN-RUIJTEN (EPP-ED, NL) i sitt inledningsanförande.
Hon lyfte fram den nya turkiska författningen och poängterade att den inte får bli en förevändning att undvika att med alla medel se till att få till stånd förändringar.
Framförallt måste Turkiet få till stånd en förändring av artikel 301 i brottsbalken och förbättra yttrandefriheten i landet, konstaterade Oomen-Ruijten.
Föredragande Oomen-Ruijten poängterade också att Turkiet måste erkänna sin förflutna historia i förhållande till Armenien.
Politiska grupper
Även Hannes SWOBODA (PSE, AT) poängterade att reformerna i Turkiet måste fortsätta, i synnerhet artikel 301 i den turkiska brottsbalken och andra reformer som garanterar yttrandefriheten.
Han lyfte även fram kurdernas situation och betonade att det nu är möjligt att lösa den politiskt och parlamentariskt och avstå från våld.
– Vi måste ge tydliga signaler att vi vill ha en fredlig lösning, sade han.
Han påpekade att det är viktigt att den turkiska regeringen utnyttjar sitt mandat för att driva på reformerna i landet.
– Regeringen måste se till att kvinnornas situation blir bättre och hedersmorden måste avskaffas.
Landsdorff påpekade också att 10-procentsspärren i det turkiska parlamentet är problematisk och att valrätten måste reformeras.
Regeringen måste ändra artikel 301 i brottsbalken och det finns fortfarande folkmord som inte har blivit erkända, poängterade han.
Joost LAGENDIJK (Verts/ALE, NL) fördömde den senaste tidens attacker från PKK.
– PKK:s attacker riktar sig mot den turkiska staten men de är också en attack på det kurdiska partiet, sade han.
– Turkiet måste erkänna cypriotiska institutioner.
Landet måste också öppna sina hamnar och flygplatser för cypriotiska fartyg och flyg.
Georgios GEORGIOU (IND/DEM, GR) kritiserade kommissionär Olli Rehn för att han betecknar alla som kämpar för frihet för terrorister.
– Jag undrar om vi inte förhastar oss när vi anser att Turkiet attackeras.
Låt oss inse att Turkiet har trupper utplacerade i ett annat EU-medlemsland och att Turkiet inte uppfyller EU:s krav, sade Georgiou.
Philip CLAEYS (ITS, BE) konstaterade att inga framsteg har gjorts sedan medlemskapsförhandlingarna inleddes.
– Vi är emot att Turkiet ansluter sig till Europa för det tillhör inte Europa, sade han.
Resolutionsförslag: B6- 0376/2007
-//EP//TEXT TA P6-TA-2007-0472 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-009-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-011-SV DOC XML V0//SV
Yttre förbindelser
Afghansk opiumproduktion för medicinska ändamål
2007-10-31 - 16:53
Europaparlamentet avger på uppmaning av utskottet för utrikesfrågor en rekommendation till rådet om opiumproduktion för medicinska ändamål i Afghanistan i syfte att skapa alternativ till den olagliga produktionen i landet som fortsätter att öka.
EU är den största biståndsgivaren när det gäller insatserna för att minska utbudet av opium genom projekt för att främja alternativa inkomstkällor som kan ersätta illegala odlingar.
År 2007 uppgick det sammanlagda priset för opiumskörden till 13 procent av Afghanistans lagliga BNP.
Enligt nya siffror från både Världsbanken och Internationella valutafonden beräknas nästan 40 procent av Afghanistans BNP vara kopplad till opiumhandeln och cirka 2,9 miljoner människor är verksamma inom vallmosektorn.
Afghanistan har i praktiken blivit den enda leverantören av världens farligaste drog, med 93 procent av världsmarknaden för opiater.
Parlamentet har med 368 röster för 49 emot och 25 nedlagda antagit ett initiativbetänkande av Marco CAPPATO (ALDE, IT) om en rekommendation från Europaparlamentet till rådet om opiumproduktion för medicinska ändamål i Afghanistan.
Parlamentet hänvisar till dokumenterade bevis om att upprorsmän, krigsherrar, talibaner och terroristgrupper har handeln med illegal narkotika som sin främsta finansieringskälla.
- att inom ramen för integrerade utvecklingsprogram motsätta sig användningen av desinfektion som ett sätt att utrota vallmoodlingar i Afghanistan,
- att utarbeta en omfattande plan och strategi, som syftar till att kontrollera produktionen av narkotika i Afghanistan genom att förbättra styrelseformerna och bekämpa korruptionen på hög nivå inom den afghanska statsförvaltningen, att läggas fram för den afghanska regeringen.
-//EP//TEXT TA P6-TA-2007-0485 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-010-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-012-SV DOC XML V0//SV
Utbildning
Yrkeskvalifikationer bör enkelt kunna jämföras i EU till 2012
2007-10-31 - 16:53
Yrkeskvalifikationer eller examensbevis som erhållits i ett EU-land bör lätt kunna jämföras mellan olika EU-länder senast 2012 tack vare en gemensam referensram som samtliga behöriga myndigheter bör referera till.
Däremot bör medlemsstaterna få ytterligare ett år på sig att koppla sina nationella kvalifikationssystem till den europeiska referensramen som dessutom bör kompletteras med system på yrkesutbildningens område, anser Europaparlamentet.
Europaparlamentet har inom medbeslutandeförfarandet antagit ett kompromisspaket av ändringar till ett betänkande av Mario MANTOVANI (EPP-ED, IT) om en rekommendation till medlemsstaterna om en europeisk referensram för kvalifikationer för livslångt lärande.
Sedan en kompromiss träffats med rådet kan ärendet avslutas genom en enda behandling.
Referensramen består av åtta vertikala nivåer, så kallade referensnivåer, som definieras genom tre horisontella nivåer – kunskap, färdigheter och förmåga – för att kunna klassificera de enskilda personerna på ett bättre sätt enligt resultatet av lärandet.
Parlamentet anser att medlemsstaterna behöver fram till 2010 (ett år mer än kommissionen föreslår) för att koppla sina nationella kvalifikationssystem till den europeiska referensramen för kvalifikationer, och på ett tydligt sätt göra hänvisningar från nationella kvalifikationsnivåer till de nivåer som ange referensramen.
Föreliggande rekommendation bygger på de riktlinjer som har tagits fram inom den så kallade Bologna-processen som inleddes 1999 och där totalt 45 europeiska stater deltar.
Betänkande: A6-0245/2007
Beslutsförfarande: Medbeslutande - 1:a behandlingen (***I)
Antagna texter
-//EP//TEXT TA P6-TA-2007-0463 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-011-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-013-SV DOC XML V0//SV
Konsumenter
Stigande livsmedelspriser
2007-10-31 - 16:53
Europaparlamentet har antagit en gemensam resolution om de stigande livsmedelspriserna och yrkar på ökade kvoter för spannmål och mjölk.
Världsmarknadspriserna på spannmål har ökat dramatiskt de senaste månaderna, och spannmålslagren har sjunkit till den lägsta nivån på 40 år.
Spannmålsskörden i EU–27 ser dessutom ut att bli ca 8 miljoner ton lägre än förra året.
Enligt jordbrukskommissionär Fischer Boels kan priserna på kött och köttprodukter komma att öka med upp till 30 procent under 2008 p.g.a. ökande foderkostnader.
Europaparlamentet välkomnar i sin resolution EU:s jordbruksministrars beslut nyligen att skjuta upp kraven på arealuttag för 2008.
Ledamöterna beklagar att rådet inte antog parlamentets ändringsförslag med syftet att skjuta upp kraven på arealuttag även för 2009, och förväntar sig att denna fråga tas upp vid den nära förestående översynen av den gemensamma jordbrukspolitiken.
Ledamöterna uppmanar även kommissionen att utan dröjsmål tillfälligt öka mjölkkvoterna för att stabilisera priserna på den inre marknaden.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att analysera skillnaderna mellan producentpriserna och de priser som tas ut av stormarknadskedjorna.
Effekterna av koncentrationen inom detaljhandelssektorn, som främst är till nackdel för små producenter, små företag och konsumenterna, bör analyseras och kommissionen bör utnyttja erforderliga lagliga åtgärder om man skulle konstatera att det förekommer missbruk av dominerade ställning på marknaden.
Biobränslen
Endast en mycket liten del av EU:s spannmålsproduktion utnyttjas för närvarande för framställning av biobränsle och endast 15 procent av odlingsarealen i EU skulle behöva tas i anspråk för att uppfylla EU:s biobränslemål 2020.
Kommissionen och medlemsstaterna uppmanas ändå att göra mera för att främja användning och framställning av andra generationens bioenergi, som bl.a. utvinns ur gödsel och avfallsprodukter från jordbruket i stället för ur primära jordbruksprodukter.
Import och export
Rådet har för avsikt att utarbeta ett förslag om att ta bort importavgifterna på spannmål 2008, som en åtgärd för att möta den svåra situationen i boskapssektorn, särskilt inom svinuppfödningen.
Europaparlamentet förkastar vidare varje försök att införa exportkvoter och avgifter för EU:s jordbruksprodukter.
Minskade livsmedelslager globalt får allvarliga följder särskilt för utvecklingsländer med låga inkomster och livsmedelunderskott.
Kommissionen bör föreslå instrument och åtgärder som kan förhindra störningar i livsmedelsförsörjningen och inflationseffekter av ytterligare prisökningar.
Slutligen uppmanar Europaparlamentet kommissionen att göra en fördjupad analys av trenderna på världsmarknaderna, inklusive den ökande efterfrågan på livsmedel i utvecklingsländerna, för att inom ramen för översynen av den gemensamma jordbrukspolitiken överväga inrättandet av en permanent mekanism för att i framtiden garantera adekvat utbud på marknaderna.
Gemensamt resolutionsförslag: B6-0400/2007/RC
-//EP//TEXT TA P6-TA-2007-0480 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-ITEM DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 FULL-TEXT DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-012-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-COVER-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-001-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-002-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-003-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-004-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-005-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-006-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-007-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-008-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-009-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-010-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-011-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-012-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-013-SV DOC XML V0//SV
-//EP//DTD IM-PRESS 20050901 PBR-FULL DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 PBR-FULL DOC XML V0//EN
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-COVER-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-001-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-002-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-003-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-004-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-005-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-006-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-007-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-008-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-009-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-010-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-011-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-012-SV DOC XML V0//SV
-//EP//TEXT IM-PRESS 20071019BRI11923 ITEM-013-SV DOC XML V0//SV
Föredragningslista - senaste utgåva
Tisdagen den 23 oktober 2007
9:00 - 10:00 Betänkande Sahra Wagenknecht A6-0391/2007
Skattepolitikens och tullpolitikens bidrag till Lissabonstrategin
om skattepolitikens och tullpolitikens bidrag till Lissabonstrategin
[ 2007/2097(INI) ]
Utskottet för ekonomi och valutafrågor
Omröstningen kommer att äga rum onsdag
10:00 - 12:20 Uttalanden av rådet och kommissionen
Resultat från det informella toppmötet mellan stats- och regeringschefer (Lissabon, 18-19 oktober 2007)
12:30 - 13:30 Omröstning
Rekommendation Helmuth Markov A6-0361/2007
Ingående av protokollet till avtalet om associering EG/Chile med anledning av Bulgariens och Rumäniens anslutning till EU
om förslaget till rådets beslut om ingående av ett andra tilläggsprotokoll till avtalet om upprättandet av en associering mellan Europeiska gemenskapen och dess medlemsstater, å ena sidan, och Republiken Chile, å andra sidan, för att ta hänsyn till Republiken Bulgariens och Rumäniens anslutning till Europeiska unionen
[12550/2007 - C6-0325/2007 - 2007/0083(AVC) ]
Utskottet för internationell handel
Betänkande Angelika Niebler A6-0377/2007
Avtal om vetenskapligt och tekniskt samarbete mellan EG och Schweiz
om förslaget till rådets och kommissionens beslut om ingående på Europeiska gemenskapens och Europeiska atomenergigemenskapens vägnar av avtalet om vetenskapligt och tekniskt samarbete mellan Europeiska gemenskaperna, å ena sidan, och Schweiziska edsförbundet, å andra sidan
[ KOM(2007)0305 - C6-0227/2007 - 2007/0106(CNS) ]
Utskottet för industrifrågor, forskning och energi
Betänkande Neil Parish A6-0373/2007
Gemenskapens växtförädlarrätt
om förslaget till rådets förordning om ändring av förordning (EG) nr 2100/94 med avseende på rätten att ansöka om gemenskapens växtförädlarrätt
[ KOM(2007)0445 - C6-0274/2007 - 2007/0161(CNS) ]
Utskottet för jordbruk och landsbygdens utveckling
Rekommendation Giuseppe Gargani A6-0369/2007
Sloveniens ratificering av protokollet av den 12 februari 2004 om ändring av Pariskonventionen av den 29 juli 1960 om skadeståndsansvar på atomenergins område
om förslaget till rådets beslut om bemyndigande för Republiken Slovenien att i Europeiska gemenskapens intresse ratificera protokollet av den 12 februari 2004 om ändring av Pariskonventionen av den 29 juli 1960 om skadeståndsansvar på atomenergins område
[9453/2007 - C6-0180/2007 - 2006/0260(AVC) ]
Utskottet för rättsliga frågor
Artikel 131 i arbetsordningen
Betänkande Miroslav Ouzký A6-0395/2007
Godkännande av den första och andra ändringen av UNECE:s Esbokonvention
om förslaget till rådets beslut om godkännande, på Europeiska gemenskapens vägnar, av den första och andra ändringen av UNECE:s Esbokonvention om miljökonsekvensbeskrivningar i ett gränsöverskridande sammanhang
[ KOM(2007)0470 - C6-0291/2007 - 2007/0169(CNS) ]
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Artikel 131 i arbetsordningen
Betänkande Jean-Marie Cavada A6-0360/2007
Bulgariens och Rumäniens anslutning till konventionen av den 26 juli 1995 om skydd av Europeiska gemenskapernas finansiella intressen och till diverse protokoll till denna konvention
om rekommendationen till rådets beslut om Bulgariens och Rumäniens anslutning till konventionen av den 26 juli 1995, som utarbetats på grundval av artikel K 3 i fördraget om Europeiska unionen, om skydd av Europeiska gemenskapernas finansiella intressen, anslutning till dess protokoll av den 27 september 1996, som utarbetats på grundval av artikel K 3 i fördraget om Europeiska unionen, till konventionen om skydd av Europeiska gemenskapernas finansiella intressen, anslutning till protokollet av den 29 november 1996, som utarbetats på grundval av artikel K 3 i fördraget om Europeiska unionen, anslutning till protokollet om förhandsavgörande av Europeiska gemenskapernas domstol angående tolkningen av konventionen om skydd av Europeiska gemenskapernas finansiella intressen, samt anslutning till det andra protokollet, som utarbetats på grundval av artikel K 3 i fördraget om Europeiska unionen, till konventionen om skydd av Europeiska gemenskapernas finansiella intressen
[ KOM(2007)0277 - C6-0238/2007 - 2007/0100(CNS) ]
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Artikel 131 i arbetsordningen
Betänkande Carlos Coelho A6-0357/2007
Kommunikationsinfrastruktur för Schengens informationssystem (SIS) (beslut)
om förslaget till rådets beslut om installation, drift och ledning av en kommunikationsinfrastruktur för SIS-sammanhang (Schengens informationssystem)
[ KOM(2007)0306 - C6-0215/2007 - 2007/0104(CNS) ]
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Artikel 131 i arbetsordningen
Betänkande Reimer Böge A6-0378/2007
Utnyttjande av Europeiska fonden för justering för globaliseringseffekter
om förslaget till Europaparlamentets och rådets beslut om utnyttjandet av Europeiska fonden för justering för globaliseringseffekter med tillämpning av punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
[ 2007/2168(ACI) ]
Budgetutskottet
Betänkande Christa Klaß A6-0347/2007
Ramdirektiv om hållbar användning av bekämpningsmedel
om förslaget till Europaparlamentets och rådets direktiv om upprättande av en ram för gemenskapens åtgärder för att uppnå en hållbar användning av bekämpningsmedel
[ KOM(2006)0373 - C6-0246/2006 - 2006/0132(COD) ]
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Betänkande Hiltrud Breyer A6-0359/2007
Utsläppande av växtskyddsmedel på marknaden
om förslaget till Europaparlamentets och rådets förordning om utsläppande av växtskyddsmedel på marknaden
[ KOM(2006)0388 - C6-0245/2006 - 2006/0136(COD) ]
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Betänkande Sharon Bowles A6-0327/2007
Rådgivande organet för styrning av den europeiska statistiken
om förslaget till Europaparlamentets och rådets beslut om inrättande av det rådgivande organet för styrning av den europeiska statistiken
[ KOM(2006)0599 - C6-0348/2006 - 2006/0199(COD) ]
Utskottet för ekonomi och valutafrågor
Betänkande Ieke van den Burg A6-0328/2007
Europeisk rådgivande kommitté för gemenskapens politik inom statistisk information
om förslaget till Europaparlamentets och rådets beslut om att inrätta en europeisk rådgivande kommitté för gemenskapens politik inom statistisk information
[ KOM(2006)0653 - C6-0379/2006 - 2006/0217(COD) ]
Utskottet för ekonomi och valutafrågor
Betänkande Carlos Coelho A6-0358/2007
Kommunikationsinfrastruktur för Schengens informationssystem (SIS) (förordning)
om förslaget till rådets förordning om installation, drift och ledning av en kommunikationsinfrastruktur för SIS sammanhang (Schengens informationssystem)
[ KOM(2007)0311 - C6-0216/2007 - 2007/0108(CNS) ]
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Betänkande Irena Belohorská A6-0291/2007
Temainriktad strategi för hållbar användning av bekämpningsmedel
om en temainriktad strategi för hållbar användning av bekämpningsmedel
[ 2007/2006(INI) ]
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Betänkande Herbert Reul A6-0348/2007
Konventionella energikällor och energiteknik
om konventionella energikällor och energiteknik
[ 2007/2091(INI) ]
Utskottet för industrifrågor, forskning och energi
15:00 - 18:00 Gemensam debatt
Budgetförfarande 2008
Betänkande Kyösti Virrankoski A6-0397/2007
Förslag till allmän budget 2008 (avsnitt III)
Budgetutskottet
Omröstningen kommer att äga rum torsdag
Betänkande Ville Itälä A6-0394/2007
Förslag till allmän budget 2008 (avsnitt I, II, IV, V, VI, VII, VIII, IX)
om förslaget till Europeiska unionens allmänna budget för budgetåret 2008
Avsnitt I, Europaparlamentet
Avsnitt II, Rådet
Avsnitt IV, Domstolen
Avsnitt V, Revisionsrätten
Avsnitt VI, Europeiska ekonomiska och sociala kommittén
Avsnitt VII, Regionkommittén
Avsnitt VIII, Ombudsmannen
Avsnitt IX, Europeiska datatillsynsmannen
[ C6-0288/2007 – 2007/2019B(BUD) ]
Budgetutskottet
Omröstningen kommer att äga rum torsdag
Slut på den gemensamma debatten
18:00 - 19:30 [eller efter avslutad debatt] Frågestund med frågor till kommissionen B6-0318/2007
21:00 - 24:00 Muntliga frågor
Stigande livsmedelspriser, konsumentskydd
O-0065/2007 Joseph Daul Lutz Goepel Neil Parish B6-0321/2007 kommissionen De stigande livsmedelspriserna
Gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater
O-0067/2007 Luis Manuel Capoulas Santos B6-0377/2007 kommissionen Konsumentskydd och prishöjningar
Socialdemokratiska gruppen i Europaparlamentet
O-0069/2007 Sergio Berlato Janusz Wojciechowski Gintaras Didžiokas Liam Aylward B6-0378/2007 kommissionen Avsevärt högre livsmedelspriser och konsumentskydd
Gruppen Unionen för nationernas Europa
Betänkande Karl-Heinz Florenz A6-0336/2007
Grönbok: Mot ett rökfritt Europa: policyalternativ på EU-nivå
om grönboken "Mot ett rökfritt Europa: policyalternativ på EU-nivå"
[ 2007/2105(INI) ]
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Rekommendation Gianluca Susta A6- /2007
Protokoll om ändring av avtalet om handelsrelaterade aspekter av immaterialrätter (TRIPS)
om förslaget till rådets beslut om godkännande på Europeiska gemenskapens vägnar av protokollet om ändring av TRIPS-avtalet, undertecknat i Genève den 6 december 2005
[8934/2006 - C6-0359/2006 - 2006/0060(AVC) ]
Utskottet för internationell handel
Betänkande Mario Mantovani A6-0245/2007
Europeisk referensram för kvalifikationer för livslångt lärande
om förslaget till Europaparlamentets och rådets rekommendation om en europeisk referensram för kvalifikationer för livslångt lärande
[ KOM(2006)0479 - C6-0294/2006 - 2006/0163(COD) ]
Utskottet för sysselsättning och sociala frågor
Föredragande av yttrande:
Milan Gaľa, utskottet för kultur och utbildning
Artikel 47 i arbetsordningen
Sacharovpriset 2007 till Salih Mahmoud Osman
Mänskliga rättigheter
2007-10-25 - 12:24
Sakharovpriset till Saleh Mahmud Osman © BELGA
Den sudanesiske människorättsadvokaten Salih Mahmoud Osman får Europaparlaments Sacharovpris för tankefrihet.
Årets Sacharovpristagare tillkännagavs i Europaparlamentets kammare i Strasbourg torsdagen den 25 oktober, kl. 11.30 av Europaparlamentets talman Hans-Gert PÖTTERING som motiverade valet så här.
- Salih Mahmoud Osman är en stark förkämpe för mänskliga rättigheter som arbetar sedan mer än tjugo år för att hjälpa och försvara personer som fördrivits, torterats eller hotas av dödsstraff.
Salih Mahmoud Osman kommer att får ta emot priset tisdagen den 11 december i samband med en officiell ceremoni i Europaparlamentets kammare i Strasbourg.
Europaparlamentet delar varje år sedan 1988 ut Sacharovpriset för tankefrihet till individer och organisationer som har gjort anmärkningsvärda insatser mot förtryck, intolerans och orättvisa.
Utmärkelsen är uppkallad efter den ryske fysikern och dissidenten Andrej Sacharov (1921-1989), som tilldelades Nobels fredspris 1975.
Priset är ett sätt för Europaparlamentet att främja och uppmärksamma kampen för mänskliga rättigheter och demokrati i världen.
I anslutning till årsdagen av undertecknandet den 10 december 1948 av FN:s deklaration om mänskliga rättigheter, delas priset ut vid en högtidlig ceremoni i Europaparlamentets plenisal i Strasbourg.
I år sker prisutdelningen den 11 december.
Pristagaren får ett certifikat och en check med prissumman 50 000 euro.
Europaparlamentets politiska grupper och en grupp individuella ledamöter (minst 40 stycken) utser varje år till att börja med fem kandidaterna till Sacharovpriset som tillkännages vid ett särskilt möte mellan utrikesutskottet, utvecklingsutskottet och underutskottet för mänskliga rättigheter.
Alla utnämningar måste åtföljas av en motivering.
Beslutet om vem som får ta emot utmärkelsen i år fattades idag den 25 oktober av talmanskonferensen (Europaparlamentets talman och ledarna för de politiska grupperna).
Salih Mahmoud Osman
Personer i hans familj har torterats och dödats till följd av hans engagemang.
Han har varit ledamot i Sudans parlament, men har fråntagits sitt mandat.
2006 - Alexander Milinkevitj
2005 - Kvinnor i vitt, Hauwa Ibrahim och Reportrar utan gränser
2004 - Zhanna Litvina, ordförande för vitryska journalistförbundet
2003 - FN:s personal och generalsekreterare Kofi Annan
2002 - Oswaldo José Payá Sardiñas
2001 - Izzat Ghazzawi, Nurit Peled-Elhanan och Dom Zacarias Kamwenho
2000 - ¡ Basta Ya!
1999 - Xanana Gusmão
1998 - Ibrahim Rugova
1997 - Salima Ghezali
1996 - Wei Jingsheng
1995 - Leyla Zana
1994 - Taslima Nasrin
1993 - Tidningen Oslobodjenje
1992 - Mödrarna från Plaza de Mayo
1991 - Adem Demaçi
1990 - Aung Sang Suu Kyi
1989 - Alexander Dubcek
SV
1
PHOTO
SV
4
MULTIMEDIA
20071025MLT12485.wmv
SV
5
MULTIMEDIA
20071025MLT12501.asf
SV
6
MULTIMEDIA
20071025MLT12503.asf
SV
7
MULTIMEDIA
20071025MLT12507.mp3
-//EP//TEXT IM-PRESS 20070702IPR08709 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
Nicolas Sarkozy i Europaparlamentets kammare
Institutioner
2007-11-13 - 16:42
Nicolas Sarkozy och Hans-Gert Pöttering i Europaparlamentet
Frankrikes president Nicolas Sarkozy upprepade inför Europaparlamentets ledamöter sitt engagemang för Europa och Frankrikes strävan efter att stå i centrum av den europeiska integrationen.
Han talade i kammaren inom ramen för ett högtidligt möte.
Europaparlamentets talman Hans-Gert PÖTTERING inledde på franska då han välkomnade Frankrikes president Nicolas Sarkozy.
Pöttering omnämnde sedan den franske författaren Victor Hugo som redan 1849 sade att Europas stater borde enas och ett antal andra fransmän vars betydelse varit avgörande för EU:s utveckling.
Ändå var det i Frankrike, påpekade han, som medborgarna förkastade konstitutionen.
- Det franska nejet var inte ett förkastade av EU, försäkrade presidenten, utan snarare ett uttryck för att EU måste leva upp mot andra krav och erbjuda något mer.
Sarkozy påminde om EU:s uppkomst efter de två världskrigen och det mod som unionens grundare uppvisade då de lyckades få ledarna i Europa och befolkningarna med sig mot en gemensam framtid.
- EU är ett uttryck för en gemensam vilja, en union grundade på gemensamma värden och en gemensam civilisation.
Misstro och besvikelse inför EU har uppstått och nu måste vi visa att vi förtjänar EU-medborgarnas förtroende.
De har intrycket av att EU inte innebär det skydd de behöver och att EU är likgiltigt inför deras dagliga problem.
Sarkozy betonade dock att EU uppnått mycket sedan kol- och stålgemenskapen.
"Utan att glömma - ty det vore att häda - har vi beslutat att ge oss in på ett stort äventyr som, om företaget lyckas, ska göra det möjligt för oss att bevara det vackraste och mest värdefulla som vi har gemensamt."
- Nu har detta äventyr pågått under mer än ett halvt sekel och olika parlamentariska församlingar har följt efter varandra.
EU fick lämna konstitutionstexten bakom sig och ta fram ett nytt fördrag för att komma ur den institutionella krisen.
- Att anta det förenklade fördraget innebar det politiska Europas seger över sig självt.
All EU-politik inom alla områden bör bli föremål för en demokratisk debatt.
Sarkozy nämnde sitt förslag om at inrätta ett "de vises råd" som ska diskutera olika utvecklingsmöjligheter för EU
- Det var ett genidrag av unionens fäder att börja med ekonomin och handeln med kol och stål, men sedan gick tiden och politiken släpade efter för att inte tala om kulturaspekten.
Men vi måste också vara kapabla att skydda vår medborgare mot ekonomiska faktorer.
- Illojal konkurrens och dumpning är inte acceptabelt.
Många länder har en stark industripolitik, en jordbrukspolitik som gagnar det egna landet, och en positiv särbehandling av nationella små och medelstora företag.
Vi vill inte ha någon protektionism, men vi måste kräva ömsesidighet.
Vi vill trygga vår energiförsörjning och vår livsmedelsförsörjning och vi vill gå i täten i klimatfrågan, men vi kan inte acceptera illojal konkurrens från länder som inte vidtar några åtgärder alls i kampen mot klimatförändringarna.
EU är mycket fäst vid fri konkurrens, men detta får inte göras till en religion.
Solidaritet bör råda när det gäller säkerheten och om man är med i Schengensamarbetet ska man inte ensidigt kunna fatta beslut om att göra ett stort antal f.d. olagliga invandrare till lagliga invandrare eftersom detta berör hela EU genom den fria rörligheten.
I slutet av sitt tal upprepade Nicolas Sarkozy sitt åtagande som president att se till att Frankrike ska stå i centrum för den europeiska integrationen och han hänvisade till en rad konkreta steg han tagit för att förbättra relationerna med de europeiska institutionerna och för att få alla ombord.
Barcelonaprocessen har inte nått ända fram och det behövs mer dynamik och nya idéer för att regionen ska utvecklas och förbindelserna mellan EU och Afrika ska stärkas, ansåg han.
Allra sist sade han:
Vi har ingen tid att förlora.
20071109IPR12787 Audio, 04:25 Audio, 31:27
SV
1
PHOTO
20071113PHT12924.jpg
SV
2
MULTIMEDIA
20071113MLT12961.asf
SV
3
MULTIMEDIA
20071113MLT12965.asf
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//TEXT TA P6-TA-2007-0507 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0508 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0509 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0510 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0511 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0512 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0513 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0514 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0515 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0516 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0517 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0518 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0519 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0520 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0521 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0522 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0523 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0524 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0525 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0526 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0527 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0528 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0529 0 DOC XML V0//SV
Kommissionens lagstiftnings- och arbetsprogram för 2008
Institutioner
2007-12-12 - 19:11
Vissa brister påpekas dock också.
Satsningar på tillväxt och sysselsättning, hållbar utveckling, klimatförändringar, energi och migration samt betoningen av bättre lagstiftning, korrekt genomförande och stärkande av Europas roll som världspartner under 2008 får oförbehållt parlamentets stöd, men kommissionen uppmanas att vara mer ambitiös i sina initiativ som syftar till att garantera grundläggande rättigheter, frihet, rättvisa och social integration.
Kommissionens åtagande att stödja ratificeringen av ändringsfördraget välkomnas.
Fördraget kommer att stärka demokratin i EU och minska avståndet mellan EU och medborgarna.
Lissabonstrategin
Tjänstedirektivet måste genomföras på ett konsekvent sätt och effektiva gemensamma kontaktpunkter inrättas för att främja tillträdet till den inre marknaden.
Parlamentet påminner om de allvarliga konsekvenserna av krisen med subprime-lånen i USA för de europeiska finansmarknaderna.
Europaparlamentet välkomnar kommissionens beslutsamma avsikt att uppnå målet med att minska de administrativa bördorna för företagen som uppstår i EU och medlemsstaterna med 25 procent senast 2012.
Översynen av telekommunikationspaketet framhålls av ledamöterna som en nyckelprioritering under det kommande året.
Ett hållbart Europa och en Östersjöstrategi
Kommissionens åtagande att inrätta en inre energimarknad och avreglera den välkomnas liksom kommissionens ambitiösa förslag om klimatförändringar.
Europaparlamentet efterlyser en omfattande och övergripande lagstiftningsram för främjande och användning av förnybar energi i EU, med bindande mål.
De två prioriterade initiativen om sjöfart och luftfart välkomnas i detta sammanhang.
Parlamentet uppmanar kommissionen att välja en tydlig och konstruktiv strategi i dialogen med Ryssland.
Europaparlamentet betonar behovet av en Östersjöstrategi för EU och uppmanar kommissionen att lägga fram en omfattande EU-strategi för Östersjöregionen under 2008.
En integrerad syn på invandring
Arbetsprogrammet nämner inte EU:s framtida system för passageraruppgifter, men ledamöterna efterlyser ökat operativt samarbete på europeisk nivå för att bekämpa terrorism.
Externa relationer
Kommissionen bör även i fortsättningen göra medborgarna uppmärksamma på vikten av kulturell mångfald och interkulturell dialog.
Debatt och omröstning: 12.12.2007
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//TEXT TA P6-TA-2007-0578 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0579 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0580 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0581 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0582 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0583 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0584 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0585 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0586 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0587 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0588 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0589 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0590 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0591 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0592 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0593 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0594 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0595 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0596 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0597 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0598 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2007-0599 0 DOC XML V0//SV
ENVI
Presentation och befogenheter
Utskottet är behörigt i frågor som rör följande områden:
2.
20071217CDE15712
Föredragningslista - dagens
Tisdagen den 15 januari 2008
LAGSTIFTNINGSDEBATT:
9:00-11:20 och 15:00-17:30
9:00 - 11:20 [LAGSTIFTNINGSDEBATT] Betänkande Glenis Willmott A6-0518/2007
Gemenskapens arbetsmiljöstrategi 2007–2012
om gemenskapens arbetsmiljöstrategi 2007–2012
[ 2007/2146(INI) ]
Utskottet för sysselsättning och sociala frågor
Betänkande Csaba Őry A6-0515/2007
Tillämpningen av systemen för social trygghet när anställda, egenföretagare eller deras familjemedlemmar flyttar inom gemenskapen
om förslaget till Europaparlamentets och rådets förordning om ändring av rådets förordning (EEG) nr 1408/71 om tillämpningen av systemen för social trygghet när anställda, egenföretagare eller deras familjemedlemmar flyttar inom gemenskapen
[ KOM(2007)0159 - C6-0104/2007 - 2007/0054(COD) ]
Utskottet för sysselsättning och sociala frågor
Andrabehandlingsrekommendation Kurt Lechner A6-0504/2007
Konsumentkrediter
om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets direktiv om konsumentkreditavtal och upphävande av rådets direktiv 87/102/EEG
[9948/2/2007 - C6-0315/2007 - 2002/0222(COD) ]
Utskottet för den inre marknaden och konsumentskydd
Omröstningen kommer att äga rum onsdag
11:30 - 12:00 Omröstning
Betänkande Jacek Saryusz-Wolski A6-0517/2007
Partnerskap inom ramen för stabiliserings- och associeringsprocessen
om förslaget till rådets förordning om ändring av förordning (EG) nr 533/2004 om upprättande av partnerskap inom ramen för stabiliserings- och associeringsprocessen
[ KOM(2007)0662 - C6-0471/2007 - 2007/0239(CNS) ]
Utskottet för utrikesfrågor
Betänkande Bogusław Liberadzki A6-0506/2007
Vägtransporter av farligt gods (kommissionens genomförandebefogenheter)
om förslaget till Europaparlamentets och rådets direktiv om ändring av direktiv 95/50/EG när det gäller kommissionens genomförandebefogenheter
[ KOM(2007)0509 - C6-0278/2007 - 2007/0184(COD) ]
Utskottet för transport och turism
Artikel 131 i arbetsordningen
Betänkande Paolo Costa A6-0513/2007
Avskaffande av diskriminering såvitt avser fraktsatser och befordringsvillkor
[ KOM(2007)0090 - C6-0086/2007 - 2007/0037(COD) ]
Utskottet för transport och turism
Betänkande Ulrich Stockmann A6-0497/2007
Flygplatsavgifter
om förslaget till Europaparlamentets och rådets direktiv om flygplatsavgifter
[ KOM(2006)0820 - C6-0056/2007 - 2007/0013(COD) ]
Utskottet för transport och turism
Betänkande Johannes Blokland A6-0406/2007
Export och import av farliga kemiska produkter
om förslaget till Europaparlamentets och rådets förordning om export och import av farliga kemikalier
[ KOM(2006)0745 - C6-0439/2006 - 2006/0246(COD) ]
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Betänkande Csaba Őry A6-0515/2007
Tillämpningen av systemen för social trygghet när anställda, egenföretagare eller deras familjemedlemmar flyttar inom gemenskapen
om förslaget till Europaparlamentets och rådets förordning om ändring av rådets förordning (EEG) nr 1408/71 om tillämpningen av systemen för social trygghet när anställda, egenföretagare eller deras familjemedlemmar flyttar inom gemenskapen
[ KOM(2007)0159 - C6-0104/2007 - 2007/0054(COD) ]
Utskottet för sysselsättning och sociala frågor
Betänkande Jorgo Chatzimarkakis A6-0494/2007
CARS 21: Ett konkurrenskraftigt motorfordonsregelverk
om CARS 21: Ett konkurrenskraftigt motorfordonsregelverk
[ 2007/2120(INI) ]
Utskottet för industrifrågor, forskning och energi
Betänkande Piia-Noora Kauppi A6-0481/2007
Skattemässig behandling av förluster i gränsöverskridande situationer
om skattemässig behandling av förluster i gränsöverskridande situationer
[ 2007/2144(INI) ]
Utskottet för ekonomi och valutafrågor
Betänkande Glenis Willmott A6-0518/2007
Gemenskapens arbetsmiljöstrategi 2007–2012
om gemenskapens arbetsmiljöstrategi 2007–2012
[ 2007/2146(INI) ]
Utskottet för sysselsättning och sociala frågor
12:00 - 12:30 Högtidligt möte
Syriens stormufti
12:30 - 13:00 Fortsättning på omröstningen
15:00 - 17:30 [LAGSTIFTNINGSDEBATT]
Betänkande Michael Cashman A6-0514/2007
Flerårigt ramprogram för Europeiska unionens byrå för grundläggande rättigheter för 2007–2012
om förslaget till rådets beslut om genomförande av förordning (EG) nr 168/2007 vad beträffar antagandet av ett flerårigt ramprogram för Europeiska unionens byrå för grundläggande rättigheter för 2007–2012
[ KOM(2007)0515 - C6-0322/2007 - 2007/0189(CNS) ]
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Omröstningen kommer att äga rum torsdag
Betänkande Roberta Angelilli A6-0520/2007
Mot en EU-strategi för barnets rättigheter
om en EU-strategi för barnets rättigheter
[ 2007/2093(INI) ]
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Associerat utskott: utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
Föredragande av yttrande: Marie Panayotopoulos-Cassiotou
Artikel 47 i arbetsordningen
17:30 - 19:00 Frågestund med frågor till kommissionen B6-0001/2008
21:00 - 24:00 Uttalande av kommissionen
Alarmerande avfallssituation i regionen Kampanien
Betänkande Doris Pack A6-0502/2007
Vuxenutbildning: Det är aldrig för sent att lära
om vuxenutbildning: Det är aldrig för sent att lära
[ 2007/2114(INI) ]
Utskottet för kultur och utbildning
Associerat utskott: utskottet för sysselsättning och sociala frågor
Föredragande av yttrande: Jan Andersson
Artikel 47 i arbetsordningen
Betänkande Friedrich-Wilhelm Graefe zu Baringdorf A6-0508/2007
Åtgärder att vidta genom fjärranalystillämpningar som inrättats inom ramen för den gemensamma jordbrukspolitiken
om förslaget till rådets förordning om de åtgärder som kommissionen avseende perioden 2008–2013 skall vidta med hjälp av det system för fjärranalys som inrättats inom ramen för den gemensamma jordbrukspolitiken
[ KOM(2007)0383 - C6-0273/2007 - 2007/0132(CNS) ]
Utskottet för jordbruk och landsbygdens utveckling
Muntlig fråga
Den rättsliga ställningen för en ledamot av Europaparlamentet som valts i Polen
O-0082/2007 Giuseppe Gargani B6-0002/2008 kommissionen Den rättsliga ställningen för en ledamot av Europaparlamentet som valts i Polen
Utskottet för rättsliga frågor
TECKENFÖRKLARING
*
Samrådsförfarandet
** I
** II
***
Samtyckesförfarandet
***I
Medbeslutandeförfarandet (första behandlingen)
***II
Medbeslutandeförfarandet (andra behandlingen)
***III
UPPLYSNINGAR ANGÅENDE OMRÖSTNINGAR
Om inget annat anges har föredraganden till talmannen skriftligen tillkännagivit sin inställning till ändringsförslagen.
FÖRKORTNINGAR FÖR UTSKOTTENS NAMN
AFET:
DEVE:
Utskottet för utveckling
INTA:
Utskottet för internationell handel
BUDG:
Budgetutskottet
CONT:
Budgetkontrollutskottet
ECON:
Utskottet för ekonomi och valutafrågor
EMPL:
Utskottet för sysselsättning och sociala frågor
ENVI:
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
ITRE:
Utskottet för industrifrågor, forskning och energi
IMCO:
Utskottet för den inre marknaden och konsumentskydd
TRAN:
Utskottet för transport och turism
REGI:
Utskottet för regional utveckling
AGRI:
PECH:
Fiskeriutskottet
CULT:
Utskottet för kultur och utbildning
JURI:
Utskottet för rättsliga frågor
LIBE:
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
AFCO:
Utskottet för konstitutionella frågor
FEMM:
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
PETI:
Utskottet för framställningar
FÖRKORTNINGAR FÖR DE POLITISKA GRUPPERNA
PPE-DE:
Gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater
PSE:
Europeiska socialdemokratiska partiets grupp
ALDE:
Gruppen Alliansen liberaler och demokrater för Europa
UEN:
Gruppen Unionen för nationernas Europa
Verts/ALE
Gruppen De gröna/Europeiska fria alliansen
GUE/NGL:
Gruppen Europeiska enade vänstern/Nordisk grön vänster
IND/DEM:
Gruppen Självständighet/Demokrati
NI:
Grupplösa
Återupptagande av sessionen
Uttalande av talmannen
Justering av protokollet från föregående sammanträde
Invändning mot giltigheten av mandatet för en ledamot av Europaparlamentet
Begäran om fastställelse av parlamentarisk immunitet
Utskottens och delegationernas sammansättning
Tillfälliga utskottet för klimatförändringar (förlängning av mandat)
Rättelser
Undertecknande av rättsakter som antagits genom medbeslutandeförfarandet
Maktmissbruk som stormarknader med verksamhet i Europeiska unionens utövar (skriftlig förklaring)
Avtalstexter översända av rådet
Bortfallna skriftliga förklaringar
Inkomna dokument
Muntliga frågor och skriftliga förklaringar (ingivande)
Framställningar
Anslagsöverföringar
Kommissionens åtgärder till följd av parlamentets resolutioner
Arbetsplan
Anföranden på en minut om frågor av politisk vikt
Begäran om fastställelse av Witold Tomczaks immunitet (debatt)
Insyn i finansiella frågor (debatt)
Skydd av gemenskapernas ekonomiska intressen - Bedrägeribekämpning - Årsrapporter 2005 -2006 (debatt)
Ömsesidigt bistånd och samarbete mellan medlemsstaternas administrativa myndigheter och kommissionen vid tillämpningen av tull- och jordbrukslagstiftningen ***I (debatt)
Gemenskapens tullkodex ***II (debatt)
Faktorer som bidrar till ökat stöd för terrorism och en ökad rekrytering av terrorister (debatt)
EU:s strategi för bättre marknadstillträde för europeiska företag (debatt)
Reform av instrumenten för skydd av handeln (debatt)
Föredragningslista för nästa sammanträde
Avslutande av sammanträdet
NÄRVAROLISTA
EUROPAPARLAMENTET
STRASBOURG
PROTOKOLL
ORDFÖRANDESKAP: Hans-Gert PÖTTERING Talman
1 Återupptagande av sessionen
Sammanträdet öppnades kl. 17.00.
2 Uttalande av talmannen
Talmannen uttalade sig till följd av att parlamentet i Kosovo förklarat landet självständigt dagen innan den 17 februari 2008.
Han uppmuntrade framför allt de styrande i Kosovo att ta sitt politiska ansvar och välkomnade rådets beslut att sända Eulex (EU:s polis- och rättinsats) till Kosovo för att övervaka och skapa en ram för den nyvunna självständigheten.
3 Justering av protokollet från föregående sammanträde
Protokollet från föregående sammanträde justerades.
4 Invändning mot giltigheten av mandatet för en ledamot av Europaparlamentet
Giulietto Chiesa s nominering till ledamot av Europaparlamentet som lagts fram av
Beniamino Donnici .
Motiveringen till detta beslut framgår av skrivelsen av den 16 januari 2008 som ordföranden i utskottet JURI sänt till parlamentets talman.
Talmannen konstaterade att det inte finns något som talar emot utskottet JURIs beslut och beslutet godkändes därför.
5 Begäran om fastställelse av parlamentarisk immunitet
Talmannen meddelade att han hade tagit emot en begäran från
Tatjana Ždanoka om skydd av hennes privilegier och immunitet till följd av en händelse som hon råkat ut för på en resa i Estland.
6 Utskottens och delegationernas sammansättning
Grupperna PPE-DE och PSE hade begärt att följande utnämningar skulle godkännas:
utskottet IMCO:
Syed Kamall i stället för
Daniel Hannan
utskottet AGRI:
James Nicholson
utskottet PECH:
Daniel Hannan i stället för
James Nicholson
delegationen till den parlamentariska församlingen EU-Latinamerika:
Charles Tannock i stället för
Daniel Hannan ,
Iuliu Winkler i stället för
Georgios Papastamkos
delegationen till den gemensamma parlamentarikerkommittén EU-Chile:
Nicolae Vlad Popa
Mihaela Popa
delegationen för förbindelserna med Maghrebländerna och Arabiska Maghrebunionen:
Rareş-Lucian Niculescu
delegationen för förbindelserna med Mercosur:
Richard James Ashworth i stället för
Daniel Hannan
delegationen för förbindelserna med Japan:
John Attard-Montalto
delegationen för förbindelserna med Folkrepubliken Kina:
Marian Zlotea
delegationen för förbindelserna med Afghanistan:
Daniel Hannan
Dessa utnämningar skulle betraktas som godkända om det inte framställdes några invändningar mot detta före justeringen av detta protokoll.
7 Tillfälliga utskottet för klimatförändringar (förlängning av mandat)
På begäran av tillfälliga utskottet för klimatförändringar föreslog talmanskonferensen vid sitt sammanträde den 14 februari 2008 att detta tillfälliga utskotts mandat skulle förlängas med 9 månader från och med den 10 maj 2008.
Det har för övrigt lagts fram ett förslag om att en interimsrapport, som enbart skulle behandla de vetenskapliga uppgifterna rörande klimatförändringen, skulle kunna läggas fram före sammanträdesperioden i maj.
Den slutgiltiga rapporten kommer att läggas fram för parlamentet efter att det nya mandatet gått ut.
Talmannen konstaterade att det inte fanns några invändningar mot förslaget.
8 Rättelser
IMCO-utskottet hade lämnat följande rättelse:
Europaparlamentets och rådets direktiv 2005/36/EG av den 7 september 2005 om erkännande av yrkeskvalifikationer Dokument 12470/2007 - 2002/0061 (COD) - LEX 637
° ° ° °
ECON-utskottet hade lämnat följande rättelser till de texter som Europaparlamentet antagit:
- Rättelse
Europaparlamentets och rådets direktiv 2008/.../EG om ändring av direktiv 2006/48/EG om rätten att starta och driva verksamhet i kreditinstitut vad gäller kommissionens genomförandebefogenheter
P6_TA-PROV(2007)0513 - ( KOM(2006)0902 – C6-0023/2007 – 2006/0284(COD) )
- Rättelse
P6_TA-PROV(2007)0517 - ( KOM(2006)0910 – C6-0018/2007 – 2006/0305(COD) )
Talmannen meddelade att han tillsammans med rådets ordförande under tisdagen skulle underteckna följande rättsakter som antagits genom medbeslutandeförfarandet, i enlighet med artikel 68 i parlamentets arbetsordning:
- Europaparlamentets och rådets förordning om fastställande av gemensamma bestämmelser på det civila luftfartsområdet och inrättande av en europeisk byrå för luftfartssäkerhet, och om upphävande av rådets direktiv 91/670/EEG, förordning (EG) nr 1592/2002 och direktiv 2004/36/EG (03697/2007/LEX - C6-0072/2008 - 2005/0228(COD) )
- Europaparlamentets och rådets direktiv om ändring av direktiv 97/67/EG beträffande fullständigt genomförande av gemenskapens inre marknad för posttjänster (03605/2008/LEX - C6-0071/2008 - 2006/0196(COD) )
- Europaparlamentets och rådets förordning om inrättande av en gemensam ram för företagsregister för statistiska ändamål och om upphävande av rådets förordning (EEG) nr 2186/93 (03665/2007/LEX - C6-0070/2008 - 2005/0032(COD) )
- Europaparlamentets och rådets förordning om ändring av förordning (EG) nr 1059/2003 om inrättande av en gemensam nomenklatur för statistiska territoriella enheter (Nuts) med anledning av Bulgariens och Rumäniens anslutning till Europeiska unionen (03645/2007/LEX - C6-0069/2008 - 2007/0038(COD) )
10 Maktmissbruk som stormarknader med verksamhet i Europeiska unionens utövar (skriftlig förklaring)
Rådet hade översänt vidimerade kopior av följande dokument:
-
-
12 Bortfallna skriftliga förklaringar
13 Inkomna dokument
Talmannen hade mottagit följande dokument:
1) från parlamentets utskott
1.1) betänkanden:
- Betänkande om EU:s strategi för att få till stånd marknadstillträde för europeiska företag ( KOM(2007)0183 - 2007/2185(INI) ) - utskottet INTA - Föredragande: Ignasi Guardans Cambó ( A6-0002/2008 )
- Betänkande om begäran om fastställelse av Claudio Favas immunitet och privilegier ( 2007/2155(IMM) ) - utskottet JURI - Föredragande: Klaus-Heiner Lehne ( A6-0007/2008 )
- Betänkande om begäran om fastställelse av Witold Tomczaks immunitet och privilegier ( 2007/2130(IMM) ) - utskottet JURI - Föredragande: Aloyzas Sakalas ( A6-0008/2008 )
- Betänkande om skydd av gemenskapernas ekonomiska intressen samt bedrägeribekämpning – årsrapporterna 2005 och 2006 ( KOM(2006)0378 - 2006/2268(INI) ) - utskottet CONT - Föredragande: Francesco Musotto ( A6-0009/2008 )
- Betänkande om öppenhet i ekonomiska frågor ( 2007/2141(INI) ) - utskottet CONT - Föredragande: José Javier Pomés Ruiz ( A6-0010/2008 )
- Betänkande om Lissabonfördraget ( 2007/2286(INI) ) - utskottet AFCO ( A6-0013/2008 )
- Betänkande om en hållbar europeisk transportpolitik, med beaktande av EU:s energi- och miljöpolitik ( 2007/2147(INI) ) - utskottet TRAN - Föredragande: Gabriele Albertini ( A6-0014/2008 )
- Betänkande med ett förslag till Europaparlamentets rekommendation till rådet om de faktorer som bidrar till ett ökat stöd för terrorism och en ökad rekrytering av terrorister ( B6-0677/2005 - 2006/2092(INI) ) - utskottet LIBE - Föredragande: Gérard Deprez ( A6-0015/2008 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets direktiv om föreskrivna skyltar och märkningar samt deras placering och fastsättningssätt på motorfordon och släpvagnar till dessa fordon (kodifierad version) ( KOM(2007)0344 - C6-0193/2007 - 2007/0119(COD) ) - utskottet JURI - Föredragande: Hans-Peter Mayer ( A6-0016/2008 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets direktiv om bakre skyltlyktor för motorfordon och släpvagnar till dessa fordon (kodifierad version) ( KOM(2007)0451 - C6-0252/2007 - 2007/0162(COD) ) - utskottet JURI - Föredragande: Hans-Peter Mayer ( A6-0017/2008 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets direktiv om dämpning av radiostörningar (elektromagnetisk kompatibilitet) som orsakas av jordbruks- eller skogsbrukstraktorer (kodifierad version) ( KOM(2007)0462 - C6-0256/2007 - 2007/0166(COD) ) - utskottet JURI - Föredragande: Francesco Enrico Speroni ( A6-0018/2008 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets direktiv om bullernivån på förarplatsen i hjulburna jordbruks- eller skogstraktorer (kodifierad version) ( KOM(2007)0588 - C6-0344/2007 - 2007/0205(COD) ) - utskottet JURI - Föredragande: Francesco Enrico Speroni ( A6-0019/2008 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets förordning om inrättande av Europeiska miljöbyrån och Europeiska nätverket för miljöinformation och miljöövervakning (kodifierad version) ( KOM(2007)0667 - C6-0397/2007 - 2007/0235(COD) ) - utskottet JURI - Föredragande: Francesco Enrico Speroni ( A6-0020/2008 )
- * Betänkande om förslaget till rådets direktiv om strukturen och skattesatserna för punktskatten på tobaksvaror (kodifierad version) ( KOM(2007)0587 - C6-0392/2007 - 2007/0206(CNS) ) - utskottet JURI - Föredragande: Francesco Enrico Speroni ( A6-0021/2008 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets direktiv om installationen av belysnings- och ljussignalanordningar på jordbruks- och skogsbrukstraktorer med hjul (kodifierad version) ( KOM(2007)0192 - C6-0108/2007 - 2007/0066(COD) ) - utskottet JURI - Föredragande: Hans-Peter Mayer ( A6-0022/2008 )
- Betänkande om fjärde rapporten om ekonomisk och social sammanhållning ( KOM(2007)0273 - 2007/2148(INI) ) - utskottet REGI - Föredragande: Ambroise Guellec ( A6-0023/2008 )
- Betänkande om Europas demografiska framtid ( KOM(2006)0571 - 2007/2156(INI) ) - utskottet EMPL - Föredragande: Françoise Castex ( A6-0024/2008 )
- *** Rekommendation om förslaget till rådets beslut om ingående av protokollet till Europa-Medelhavsavtalet om upprättande av en associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Staten Israel, å andra sidan, för att ta hänsyn till Republiken Bulgariens och Rumäniens anslutning till Europeiska unionen (15061/2007 - C6-0445/2007 - 2007/0165(AVC) ) - utskottet AFET - Föredragande: Jacek Saryusz-Wolski ( A6-0025/2008 )
- *** Rekommendation om förslaget till rådets beslut om ingående av ett protokoll till Europa-Medelhavsavtalet om upprättande av en associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Arabrepubliken Egypten, å andra sidan, för att ta hänsyn till Republiken Bulgariens och Rumäniens anslutning till Europeiska unionen (13199/2007 - C6-0438/2007 - 2007/0180(AVC) ) - utskottet AFET - Föredragande: Jacek Saryusz-Wolski ( A6-0026/2008 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets beslut om gemenskapens deltagande i ett forsknings- och utvecklingsprogram som syftar till att öka livskvaliteten för äldre människor genom användning av informations- och kommunikationsteknik (IKT) och som inletts av flera medlemsstater ( KOM(2007)0329 - C6-0178/2007 - 2007/0116(COD) ) - utskottet ITRE - Föredragande: Neena Gill ( A6-0027/2008 )
- Betänkande om en uppföljning av EU:s territoriella agenda och Leipzigstadgan – ett europeiskt handlingsprogram för fysisk planering och territoriell sammanhållning ( 2007/2190(INI) ) - utskottet REGI - Föredragande: Gisela Kallenbach ( A6-0028/2008 )
- Betänkande om de integrerade riktlinjerna för tillväxt och sysselsättning (del: allmänna riktlinjer för medlemsstaternas och gemenskapens ekonomiska politik): start för den nya treårsperioden (2008–2010) ( 2007/2275(INI) ) - utskottet ECON - Föredragande: Margarita Starkevičiūtė ( A6-0029/2008 )
- Betänkande om kvinnornas situation i EU:s landsbygdsområden ( 2007/2117(INI) ) - utskottet FEMM - Föredragande: Christa Klaß ( A6-0031/2008 )
- Betänkande om en EU-strategi för Centralasien ( 2007/2102(INI) ) - utskottet AFET - Föredragande: Cem Özdemir ( A6-0503/2007 )
1.2) andrabehandlingsrekommendationer:
- ***II Andrabehandlingsrekommendation om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets förordning om fastställande av en tullkodex för gemenskapen (Moderniserad tullkodex) (11272/6/2007 - C6-0354/2007 - 2005/0246(COD) ) - utskottet IMCO - Föredragande: Janelly Fourtou ( A6-0011/2008 )
2) från ledamöterna
2.1) muntliga frågor inför frågestunden (artikel 109 i arbetsordningen) ( B6-0010/2008 )
till rådet:
till kommissionen: - Jensen Anne E., Leichtfried Jörg, Gutiérrez-Cortines Cristina, Panayotopoulos-Cassiotou Marie, Posselt Bernd, Ó Neachtain Seán, Kirilov Evgeni, Moraes Claude, Higgins Jim, Crowley Brian, Martin David, Papadimoulis Dimitrios, Kuźmiuk Zbigniew Krzysztof, Geringer de Oedenberg Lidia Joanna, Ebner Michl, Angelakas Emmanouil, Papastamkos Georgios, Corda Giovanna, Mitchell Gay, Burke Colm, McGuinness Mairead, Arnaoutakis Stavros, Hieronymi Ruth, Badia i Cutchet Maria, van Nistelrooij Lambert, Chatzimarkakis Jorgo, Medina Ortega Manuel, Doyle Avril, Hutchinson Alain, Ludford Sarah, McAvan Linda, Vălean Adina-Ioana, Dillen Koenraad, Farage Nigel, Öger Vural, Ryan Eoin, Aylward Liam, Claeys Philip, Mavrommatis Manolis, Schlyter Carl, Toussas Georgios, Nicholson James, Harkin Marian, Filip Petru, Irujo Amezaga Mikel, Sonik Bogusław, Newton Dunn Bill, Van Hecke Johan, Vanhecke Frank, Paleckis Justas Vincas, Pleštinská Zita, Ayala Sender Inés, Rack Reinhard, Georgiou Georgios, Salinas García María Isabel, Podimata Anni, Bushill-Matthews Philip, Czarnecki Marek Aleksander, Budreikaitė Danutė, Czarnecki Ryszard, Botopoulos Costas, de Brún Bairbre, Evans Robert, Andrikienė Laima Liucija, Pafilis Athanasios, Manolakou Diamanto, Schmidt Olle, Martin Hans-Peter, Batzeli Katerina, Ţicău Silvia-Adriana
hänvisat till
ansvarigt utskott :
ENVI
hänvisat till
ansvarigt utskott :
LIBE
hänvisat till
ansvarigt utskott :
LIBE
hänvisat till
ansvarigt utskott :
IMCO
rådgivande utskott :
INTA, REGI
14 Muntliga frågor och skriftliga förklaringar (ingivande)
Talmannen hade mottagit följande dokument från ledamöterna::
1) muntliga frågor (artikel 108 i arbetsordningen):
-
( O-0009/2008 ) från
Arlene McCarthy , för utskottet IMCO, till kommissionen:
Säkerhetsmärkning av konsumentprodukter ( B6-0009/2008 )
2) skriftliga förklaringar införda i registret (artikel 116 i arbetsordningen):
-
Filiz Hakaeva Hyusmenova ,
Metin Kazak ,
Vladko Todorov Panayotov ,
Bilyana Ilieva Raeva och
Iliana Malinova Iotova ,
om en gemensam europeisk politik för uppfostran och omsorg av missgynnade barn
(0014/2008) ;
-
Marian Zlotea och
Sebastian Valentin Bodu ,
om full återbetalning av registreringsavgiften för fordon som registreras för första gången till dem som i strid med gemenskapslagstiftningen fått betala denna avgift
(0015/2008) .
15 Framställningar
Den 28.01.2008
från Takis Onisiforou (Sintonistiki Epitropi Agona Ton Idioktiton Temachion Gia Tis Archaiotites Sti Periochi Amathountas) (2 underskrifter) (nr 1374/2007);
från Dimitrios Hatzinas (nr 1375/2007);
från Eleni Kalamboka (nr 1376/2007);
från Aleksander Bicanic Plut (nr 1377/2007);
från Georgiou Apostoliki (nr 1378/2007);
från Georgios Giorgopoulos (Panellinio Somatio Ethnikon diethnon Epivatikon Mataforon o Dromeas) (2 underskrifter) (nr 1379/2007);
från Javier Gomez Gonzalez (nr 1380/2007);
från Antero Oliveiro Resende (Partido Ecologista "Os Verdes") (nr 1381/2007);
från Ioan Dascaliuc (nr 1382/2007);
från Stefania Anna Sulkowska (nr 1383/2007);
från Malina Ioncova Ivanova (nr 1384/2007);
från Antonio Cuevas Benitez (nr 1385/2007);
från Alfonso Santos Roman (Esquerda Unida - Izquierda Unida) (nr 1386/2007);
från Pedro Dominguez Gento (nr 1387/2007);
från Valeriu Melinte (nr 1388/2007);
från William Lanzoni (4 underskrifter) (nr 1389/2007);
från Thomas Pankauke (5 underskrifter) (nr 1390/2007);
från Miguel Angel Ortiz López (Plataforma para la difensa del Rio Castril) (690 underskrifter) (nr 1391/2007);
från Iago Patino (Izquierda unida del ayuntamiento de Ames) (nr 1392/2007);
från Silvia Leal Acevedo (nr 1393/2007);
från Miguel Angel Gea Rifá (Izquierda Unida Los Verdes-Convocatoria por Andalucía) (nr 1394/2007);
från Zoltan Baghy (nr 1395/2007);
från Csaba Vetésy (nr 1396/2007);
från Mircea Nicusor Purcareata (Mostenitori Fam.
Rata) (nr 1397/2007);
från Nicolae Dragulanescu (Romanian Foundation for Quality Promotion) (nr 1398/2007);
från Gyula Implom (nr 1399/2007);
från Maria Donciu Ivanov (nr 1400/2007);
från Frédérique Carnaroli (nr 1401/2007);
från Amerigo Rutigliano (nr 1402/2007);
från Dobrinka Pavlova (nr 1403/2007);
från Ivan Shumkov (Инициативен комитет за борба с терора на преминаващите тирове през град Габрово (Initiative committee against the passing trucks through the town)) (nr 1404/2007);
från Ivaylo Krastev Assenov (ЗАЩИТА ЗДРАВЕТО И ЖИВОТА НА НАСЕЛЕНИЕТО И ОКОЛНАТА СРЕДА (Protection of the health and life of the population and environment)) (1061 underskrifter) (nr 1405/2007);
från Carlos Santos (nr 1406/2007);
från (konfidentiellt namn) (nr 1407/2007);
från Vicente Felipe Sanchez Pedrosa (nr 1408/2007);
från Willi Waxweiler (nr 1409/2007);
från Dominique Couprie (nr 1410/2007);
från Bernd Fritz (nr 1411/2007);
från Angelo Romano (nr 1412/2007);
från (konfidentiellt namn) (nr 1413/2007);
från Elad Shetreet (nr 1414/2007);
från (konfidentiellt namn) (nr 1415/2007);
från Roland Blomeyer (nr 1416/2007);
från Konstantinos Skoufis (372 underskrifter) (nr 1418/2007);
från Christos Nikoloutsopoulos (3 underskrifter) (nr 1419/2007);
från Rolf Hecht (nr 1420/2007);
från (konfidentiellt namn) (nr 1421/2007);
från Inge Rosenberger (nr 1422/2007);
från Stephanie Bleck (nr 1423/2007);
från Wayne Pendle (nr 1424/2007);
från (konfidentiellt namn) (nr 1425/2007);
från (konfidentiellt namn) (nr 1426/2007);
från (konfidentiellt namn) (nr 1427/2007);
från Erich Klein (nr 1428/2007);
från Gabriela Dana Olaneanu (S.C. Prestige Trading Srl) (nr 1429/2007);
från Rita Fahle (nr 1430/2007);
från Rumiana Ivanova (nr 1431/2007);
från Maria Domenica Cerfeda (2 underskrifter) (nr 1432/2007);
från Michael Scheeder (2 underskrifter) (nr 1433/2007);
från Klaus Dieter Grothe (nr 1434/2007);
från Robert Cautain (2 underskrifter) (nr 1435/2007);
från Ioan Berfela (nr 1436/2007);
från Terry McHugh (nr 1437/2007);
från Christos Savvas (nr 1438/2007);
från Timothy Guy Neville (nr 1439/2007);
från Josep Vicent Requena Diez (Agrupament Progressiste de Manises (APM)) (10 underskrifter) (nr 1440/2007);
från Grigorios Mentis (4 underskrifter) (nr 1441/2007);
från Radu Miron Costin (Parohia Unita cu Roma Greco Catolica) (2 underskrifter) (nr 1442/2007);
från Carlos Enrique Gozalo Ara (nr 1443/2007);
från Werner Gottstein (nr 1444/2007);
från Bodo Prüfer (nr 1445/2007);
från Markus Huber (2 underskrifter) (nr 1446/2007);
från Edith Mézière (nr 1447/2007);
från Henryk Demps (nr 1448/2007);
från Chan Tsz Wai (nr 1449/2007);
från Peter Penchev (Association for the freedom of speech "Anna Politkovskaia" (Асоциация на свободното слово “Анна Политковская”)) (nr 1452/2007);
från Milan Jaros (nr 1454/2007);
från Stamatis Pantelidis (nr 1455/2007);
Den 06.02.2008
från Manuel Joaquim Monteiro de Barros (Union Pan-Européenne de la Propriété Immobilière) (nr 1456/2007);
från Andreas Radicke (Humanitas - Human Aid (Dachverband Berlin)) (2 underskrifter) (nr 1457/2007);
från Luis de la Rasilla Sánchez-Arjona (Proyector INTER/SUR para la Ecociudadanía y la Democracia Ecociudadana) (nr 1458/2007);
från Roberto Giurastante (Greenaction Transnational) (nr 1459/2007);
från René Merite (nr 1460/2007);
från Ion Falcuta (nr 1461/2007);
från Antonio Rodriguez Perez (Federación Ben Magec-Ecologistas en Acción) (nr 1462/2007);
från Frédéric Brozdziak (FFMC (Fédération Française des Motards en Colère)) (nr 1463/2007);
från Ramiro Pinto Cañón (Asociación Renta Ciudadana (Arenci)) (nr 1464/2007);
från Luis de la Rasilla Sánchez-Arjona (Proyector INTER/SUR para la Ecociudadanía y la Democracia Ecociudadana) (nr 1465/2007);
från Jan Naumów (nr 1466/2007);
från Odysseas Nikou (nr 1467/2007);
från Fotini Dermitzaki (34 underskrifter) (nr 1468/2007);
från Ioannis Kartsidimas (nr 1469/2007);
från Kiriakos Daraktsis (Συλλογοσ αλιεων κεραμωτησ) (nr 1470/2007);
från Theodoros Pitikaris (nr 1471/2007);
från Peter Reitbauer (nr 1472/2007);
från Lucia Bogdan (nr 1473/2007);
från Manuela Neugeschwandtner (nr 1474/2007);
från Christo Sofianidi (Panpontiakos Sillogos "Argo" ) (nr 1475/2007);
från (konfidentiellt namn) (nr 1476/2007);
från (konfidentiellt namn) (nr 1477/2007);
från Penny Konitsioti (nr 1478/2007);
från Franz Rehbein (nr 1479/2007);
från Gabriele Menzel (Tierfreunde ohne Grenzen e.V.) (2 underskrifter) (nr 1480/2007);
The Metropolitan Pavlos of Kyrenia (-) (nr 1481/2007);
från Justice Livingstone (African-Migrants Victims Support Organisation) (nr 1482/2007);
från Gina Diaconu (nr 1483/2007);
från Constantin Predescu (nr 1484/2007);
från Teofil Perneac Gheorghe (nr 1485/2007);
från Nella Manofu (nr 1486/2007);
från Sylvain Sieauvy (nr 1487/2007);
från Jurij Rudanovai (nr 1488/2007);
från Stefanos Modeas (nr 1491/2007);
från Helmut Bruns (nr 1492/2007);
från António Araújo Jacome (nr 1493/2007);
från Plamena Naydenova (nr 1494/2007);
från Franco Quinti (nr 1495/2007);
från Aimo Lahdelma (nr 1496/2007);
från Naveed Iqbal Hashmi (12 underskrifter) (nr 1497/2007);
från Yosheba Sainz de la Higuera y Gartzia (nr 1498/2007);
från Yosheba Sainz de la Higuera y Gartzia (nr 1499/2007);
från Apostolos Ziakas (nr 1500/2007);
från Helmut Musiala (nr 1501/2007);
från Theodoros Papoulakos (nr 1502/2007);
från Asztrik Várszegi (Bishop, archabbot of Pannonhalma, archabbot of Hungarian Benedectine Congregation) (nr 1504/2007);
från Sindicato dos Profissionais dos Transportes, Turismo e Outros Serviços de Angra do Heroísmo (nr 1505/2007);
från Aikaterini Tsamadia (Sillogos Alilleggiis ip Mesologgiou) (2 underskrifter) (nr 1506/2007);
Den 11.02.2008
från David Bacchetta (nr 0001/2008);
från Marc Sasiek (2 underskrifter) (nr 0002/2008);
från (konfidentiellt namn) (nr 0003/2008);
från (konfidentiellt namn) (nr 0004/2008);
från Heiner Holzapfel (nr 0005/2008);
från Massimo Poggi (nr 0006/2008);
från Christopher Celegrat (Mavero Recruitment) (nr 0007/2008);
från Jennifer Harvey (nr 0008/2008);
från Corinne Jaussaud (nr 0009/2008);
från Marie-France Legas (nr 0010/2008);
från Monica Kinsella (nr 0011/2008);
från Francesco Miglino (Partito Internettiano) (nr 0012/2008);
från John McElligott (Kilcolgan Residents Association) (nr 0013/2008);
från Svitlana Hluvko (nr 0014/2008);
från Mario Carassale (nr 0015/2008);
från (konfidentiellt namn) (nr 0016/2008);
från Alexandra Bougé (nr 0017/2008);
från Constanta Dumitrascu (nr 0018/2008);
från (konfidentiellt namn) (nr 0019/2008);
från Sebastian Ochieng Onyango (Kenyans for Democracy) (nr 0020/2008);
från (konfidentiellt namn) (nr 0021/2008);
från Hartmut Schmidt (nr 0022/2008);
från Felipe Xosé Larino Noia (nr 0023/2008);
från Daniela Hepe (nr 0024/2008);
från (konfidentiellt namn) (nr 0025/2008);
från Manuel Francisco Oliveira Gonçalves (Rancho Folclórico de Canidelo) (nr 0026/2008);
från (konfidentiellt namn) (nr 0027/2008);
från Juan Carlos Anguita Raigon (nr 0028/2008);
från Mihai Anisoara (nr 0029/2008);
från Robert Walczak (nr 0030/2008);
från Ilie Carzon (nr 0031/2008);
från Pietro Borsellino (nr 0032/2008);
från Michael Kramer (nr 0033/2008);
från (konfidentiellt namn) (nr 0034/2008);
från (konfidentiellt namn) (nr 0035/2008);
från (konfidentiellt namn) (nr 0036/2008);
från Wolfgang Kottwitz (3 underskrifter) (nr 0038/2008);
från (konfidentiellt namn) (nr 0039/2008);
från Fergal Mee (nr 0040/2008);
Den 12.02.2008
från Giovanni Ceravola (nr 0041/2008);
från Mihaela-Ioana Matei (nr 0043/2008);
från (konfidentiellt namn) (nr 0044/2008);
från Andy Vermaut (De Missie) (nr 0045/2008);
från (konfidentiellt namn) (nr 0046/2008);
från Victor Ciustea (SC "Trans-Service" Srl.) (nr 0047/2008);
från Karl Windisch (nr 0048/2008);
från Jeanine Wallace (nr 0049/2008);
från Michel Abate (nr 0050/2008);
från (konfidentiellt namn) (nr 0051/2008);
från Nadine Schmissek (nr 0052/2008);
från Gabriel Kevers (nr 0053/2008);
från Niko Linsa (nr 0054/2008);
från Gennaro Ciancio (nr 0055/2008);
från Rainer Kunze (nr 0056/2008);
från (konfidentiellt namn) (nr 0057/2008);
från Genaro Pens Souto (nr 0058/2008);
från Georg Krulik (nr 0059/2008);
från Alfred Weiss (nr 0060/2008);
från Royston Goodwin (nr 0061/2008);
från Dietmar Gehrmann (nr 0062/2008);
från Judith Hejda (nr 0063/2008);
från Sotiris Balagiannis (nr 0064/2008);
från Jozef Blazejczyk (nr 0065/2008);
från Wolfgang Lange (2 underskrifter) (nr 0066/2008);
från Thomas Koenig (nr 0067/2008);
från Maria Gzabanowska (nr 0068/2008);
från Lahoucine Hindi (nr 0069/2008);
från European Citizens' Initiative (1 000 000 underskrifter) (nr 0070/2008);
från Karl Berger (93 underskrifter) (nr 0071/2008);
från Theodoros Papoulakos (nr 0072/2008);
från (konfidentiellt namn) (nr 0073/2008);
från (konfidentiellt namn) (nr 0074/2008);
från (konfidentiellt namn) (nr 0075/2008);
från Bernadette Faherty (Óstán Inís Meáin (Inishmaan Hotel)) (nr 0076/2008);
16 Anslagsöverföringar
Budgetutskottet hade behandlat kommissionens förslag till anslagsöverföring DEC 01/2008 (
C6-0032/2008 - SEC(2008)0014 final ).
Kommissionens meddelande om de åtgärder som kommissionen vidtagit till följd av resolutioner som parlamentet antagit under sammanträdesperioden oktober I och II 2007 finns nu tillgängligt.
18 Arbetsplan
Nästa punkt på föredragningslistan var fastställandet av arbetsplanen.
Det slutgiltiga förslaget till föredragningslista för sammanträdesperioderna i februari I (PE 401.169/PDOJ) hade delats ut.
Följande ändringar hade föreslagits i enlighet med artikel 132 i arbetsordningen:
Sammanträdena den 18.02.2008
− 21.02.2008
måndagen
- inga ändringar
tisdagen
- inga ändringar
onsdagen
- begäran från gruppen IND/DEM om att skjuta fram omröstningen om betänkandet av
Richard Corbett och Íñigo Méndez de Vigo
om Lissabonfördraget (
A6-0013/2008 )
(punkt 29 i PDOJ)
Talare:
Jens-Peter Bonde för IND/DEM-gruppen , som motiverade begäran,
Richard Corbett (föredragande),
Hannes Swoboda för PSE-gruppen, och
Jens-Peter Bonde om dessa två inlägg.
Genom omröstning med namnupprop (IND/DEM) (24 för, 220 emot, 11 nedlagda röster), parlamentet förkastade begäran.
Talmannen,
Piia-Noora Kauppi och
Brigitte Fouré meddelade att de hade velat rösta mot begäran.
Omröstningen kommer således att äga rum på onsdagen kl. 12.00.
torsdagen
- inga ändringar
Arbetsplanen var därmed fastställd.
19 Anföranden på en minut om frågor av politisk vikt
Följande ledamöter höll, i enlighet med artikel 144 i arbetsordningen, ett anförande på en minut för att uppmärksamma parlamentet på frågor av politisk vikt:
Georgios Papastamkos ,
Ioan Mircea Paşcu ,
Ignasi Guardans Cambó ,
Jan Tadeusz Masiel ,
Claude Turmes ,
Daniel Strož ,
Slavi Binev ,
Nicolae Vlad Popa ,
Csaba Sándor Tabajdi ,
Tunne Kelam ,
Neena Gill ,
Viktória Mohácsi ,
Hanna Foltyn-Kubicka ,
Urszula Gacek ,
Jörg Leichtfried ,
Toomas Savi ,
Bogusław Rogalski ,
Milan Horáček ,
Zsolt László Becsey ,
Proinsias De Rossa ,
Csaba Sógor ,
Marusya Ivanova Lyubcheva ,
Marie Panayotopoulos-Cassiotou ,
Magor Imre Csibi ,
Jaromír Kohlíček ,
László Tőkés ,
Anna Záborská ,
Ioannis Gklavakis och
Silvia-Adriana Ţicău .
ORDFÖRANDESKAP: Manuel António dos SANTOS Vice talman
Talare:
Péter Olajos ,
Iuliu Winkler ,
Milan Gaľa ,
Colm Burke ,
Jean-Claude Martinez ,
Ján Hudacký och
Avril Doyle .
20
Begäran om fastställelse av Witold Tomczaks immunitet (debatt)
Betänkande om begäran om fastställelse av Witold Tomczaks immunitet och privilegier [ 2007/2130(IMM) ] - Utskottet för rättsliga frågor.
Föredragande: Aloyzas Sakalas ( A6-0008/2008 )
Aloyzas Sakalas presenterade sitt betänkande.
Talare:
Lidia Joanna Geringer de Oedenberg för PSE-gruppen,
Marek Aleksander Czarnecki för UEN-gruppen,
Jens-Peter Bonde och
Aloyzas Sakalas .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 6.13 i protokollet av den 19.02.2008
.
21
Insyn i finansiella frågor (debatt)
Betänkande om insyn i finansiella frågor [ 2007/2141(INI) ] - Budgetkontrollutskottet.
Föredragande: José Javier Pomés Ruiz ( A6-0010/2008 )
José Javier Pomés Ruiz redogjorde för sitt betänkande.
Talare:
Siim Kallas (kommissionens vice ordförande).
Talare:
Ingeborg Gräßle för PPE-DE-gruppen,
Dan Jørgensen för PSE-gruppen ,
Janusz Wojciechowski för UEN-gruppen ,
Bart Staes för Verts/ALE-gruppen,
Esko Seppänen för GUE/NGL-gruppen,
Nils Lundgren för IND/DEM-gruppen,
Esther De Lange ,
Paulo Casaca ,
Wiesław Stefan Kuc ,
Alexander Stubb ,
Inés Ayala Sender och
Ville Itälä .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Paul Rübig ,
Jens-Peter Bonde ,
Czesław Adam Siekierski ,
Zbigniew Zaleski och
Alexander Stubb .
Talare:
Siim Kallas och
José Javier Pomés Ruiz .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 6.16 i protokollet av den 19.02.2008
.
22
Skydd av gemenskapernas ekonomiska intressen - Bedrägeribekämpning - Årsrapporter 2005 -2006 (debatt)
Betänkande om skydd av gemenskapernas ekonomiska intressen - Bedrägeribekämpning - Årsrapporter 2005-2006 [ 2006/2268(INI) ] - Budgetkontrollutskottet.
Föredragande: Francesco Musotto ( A6-0009/2008 )
Francesco Musotto redogjorde för sitt betänkande.
ORDFÖRANDESKAP: Mario MAURO Vice talman
Talare:
Siim Kallas (kommissionens vice ordförande).
Talare:
Jan Březina (föredragande av yttrande från utskottet REGI),
Kyösti Virrankoski (föredragande av yttrande från utskottet AGRI) ,
Ingeborg Gräßle för PPE-DE-gruppen ,
Szabolcs Fazakas för PSE-gruppen,
Zbigniew Krzysztof Kuźmiuk för UEN-gruppen,
Bart Staes för Verts/ALE-gruppen,
Derek Roland Clark för IND/DEM-gruppen,
Andreas Mölzer , grupplös,
Ville Itälä ,
Herbert Bösch och
Mairead McGuinness .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Bart Staes ,
Dumitru Oprea och
Ingeborg Gräßle .
Talare:
Siim Kallas och
Francesco Musotto .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 6.17 i protokollet av den 19.02.2008
.
23
Ömsesidigt bistånd och samarbete mellan medlemsstaternas administrativa myndigheter och kommissionen vid tillämpningen av tull- och jordbrukslagstiftningen ***I (debatt)
Betänkande om förslaget till Europaparlamentets och rådets förordning om ändring av rådets förordning (EG) nr 515/97 om ömsesidigt bistånd mellan medlemsstaternas administrativa myndigheter och om samarbete mellan dessa och kommissionen för att säkerställa en korrekt tillämpning av tull- och jordbrukslagstiftningen [ KOM(2006)0866 – C6-0033/2007 – 2006/0290(COD) ] - Utskottet för den inre marknaden och konsumentskydd.
Föredragande: Bill Newton Dunn ( A6-0488/2007 )
Talare:
Siim Kallas (kommissionens vice ordförande).
Bill Newton Dunn redogjorde för sitt betänkande.
Talare:
Véronique Mathieu (föredragande av yttrande från utskottet CONT),
Christopher Heaton-Harris för PPE-DE-gruppen, och
Catherine Neris för PSE-gruppen .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Mairead McGuinness .
Talare:
Siim Kallas och
Bill Newton Dunn .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 6.15 i protokollet av den 19.02.2008
.
24
Gemenskapens tullkodex ***II (debatt)
Andrabehandlingsrekommendation om den gemensamma ståndpunkten antagen av rådet inför antagandet av Europaparlamentets och rådets förordning om fastställande av en tullkodex för gemenskapen (Moderniserad tullkodex) [11272/6/2007 - C6-0354/2007 - 2005/0246(COD) ] - Utskottet för den inre marknaden och konsumentskydd.
Föredragande: Janelly Fourtou ( A6-0011/2008 )
Janelly Fourtou redogjorde för andrabehandlingsrekommendationen.
Talare:
László Kovács (ledamot av kommissionen) .
Talare:
Christopher Heaton-Harris för PPE-DE-gruppen,
Manuel Medina Ortega för PSE-gruppen,
Othmar Karas och
Andreas Schwab .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Zuzana Roithová ,
Bill Newton Dunn och
Mairead McGuinness .
Talare:
László Kovács och
Janelly Fourtou .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 6.14 i protokollet av den 19.02.2008
.
25
Faktorer som bidrar till ökat stöd för terrorism och en ökad rekrytering av terrorister (debatt)
Betänkande innehållande ett förslag till Europaparlamentets rekommendation till rådet om faktorer som bidrar till ett ökat stöd för terrorism och en ökad rekrytering av terrorister [ 2006/2092(INI) ] - Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor.
Föredragande: Gérard Deprez ( A6-0015/2008 )
Gérard Deprez redogjorde för sitt betänkande.
Talare:
Franco Frattini (kommissionens vice ordförande) .
Talare:
Manfred Weber för PPE-DE-gruppen,
Claudio Fava för PSE-gruppen,
Ignasi Guardans Cambó för ALDE-gruppen,
Ryszard Czarnecki för UEN-gruppen,
Georgios Georgiou för IND/DEM-gruppen,
Jim Allister , grupplös,
Carlos Coelho ,
Inger Segelström och
Alexander Alvaro .
ORDFÖRANDESKAP: Adam BIELAN Vice talman
Talare:
Bárbara Dührkop Dührkop ,
Sarah Ludford ,
Jan Marinus Wiersma och
Olle Schmidt .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Hubert Pirker ,
Manfred Weber ,
Alexander Alvaro ,
Ignasi Guardans Cambó och
Sarah Ludford .
Talare:
Franco Frattini och
Gérard Deprez .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 6.18 i protokollet av den 19.02.2008
.
26
EU:s strategi för bättre marknadstillträde för europeiska företag (debatt)
Betänkande om EU:s strategi för bättre marknadstillträde för europeiska företag [ 2007/2185(INI) ] - Utskottet för internationell handel.
Föredragande: Ignasi Guardans Cambó ( A6-0002/2008 )
Ignasi Guardans Cambó redogjorde för sitt betänkande.
Talare:
Peter Mandelson (ledamot av kommissionen) .
Talare:
Silvia-Adriana Ţicău (föredragande av yttrande från utskottet ITRE),
Corien Wortmann-Kool för PPE-DE-gruppen,
Carlos Carnero González för PSE-gruppen,
Cristiana Muscardini för UEN-gruppen,
Carl Schlyter för Verts/ALE-gruppen,
Christofer Fjellner ,
Leopold Józef Rutowicz och
Georgios Papastamkos .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Zuzana Roithová ,
Mairead McGuinness ,
Zbigniew Krzysztof Kuźmiuk och
Czesław Adam Siekierski .
Talare:
Peter Mandelson och
Ignasi Guardans Cambó
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 6.19 i protokollet av den 19.02.2008
.
27
Reform av instrumenten för skydd av handeln (debatt)
Uttalande av kommissionen:
Reform av instrumenten för skydd av handeln
Peter Mandelson (ledamot av kommissionen) gjorde ett uttalande.
Talare:
Christofer Fjellner för PPE-DE-gruppen,
Jan Marinus Wiersma för PSE-gruppen,
Carl Schlyter för Verts/ALE-gruppen,
Helmuth Markov för GUE/NGL-gruppen,
Daniel Caspary ,
Erika Mann ,
Tokia Saïfi ,
Kader Arif och
Elisa Ferreira .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Mairead McGuinness ,
Zbigniew Zaleski ,
Czesław Adam Siekierski ,
Corien Wortmann-Kool ,
Kader Arif och
Elisa Ferreira .
Talare:
Peter Mandelson .
Talmannen förklarade debatten avslutad.
28 Föredragningslista för nästa sammanträde
Föredragningslistan för nästa sammanträde fastställdes ("Föredragningslista" PE 401.169/OJMA).
29 Avslutande av sammanträdet
Sammanträdet avslutades kl. 23.10.
Harald R
ømer
Hans-Gert Pöttering
Generalsekreterare
Talman
NÄRVAROLISTA
Följande skrev på:
Adamou
Agnoletto
Aita
Albertini
Allister
Alvaro
Anastase
Andersson
Andrejevs
Andrikienė
Angelakas
Angelilli
Antoniozzi
Arif
Ashworth
Atkins
Attwooll
Aubert
Audy
Auken
Ayala Sender
Aylward
Ayuso
Baco
Badia i Cutchet
Baeva
Barón Crespo
Batten
Battilocchio
Batzeli
Bauer
Beaupuy
Beazley
Becsey
Belder
Belohorská
Beňová
Berend
Berès
Berlato
Berlinguer
Bielan
Binev
Blokland
Bloom
Bobošíková
Bodu
Bösch
Bonde
Booth
Borrell Fontelles
Boştinaru
Bourzai
Bowis
Bowles
Bradbourn
Braghetto
Brejc
Brepoels
Breyer
Březina
Brie
Brok
Brunetta
Budreikaitė
van Buitenen
Buitenweg
Bulfon
Bullmann
Bulzesc
van den Burg
Burke
Bushill-Matthews
Busk
Buşoi
Buzek
Cabrnoch
Calabuig Rull
Callanan
Camre
Capoulas Santos
Cappato
Carlotti
Carnero González
Carollo
Casaca
Cashman
Caspary
Castex
del Castillo Vera
Cederschiöld
Cercas
Chichester
Chmielewski
Christensen
Chruszcz
Claeys
Clark
Cocilovo
Coelho
Cohn-Bendit
Corbett
Corbey
Corda
Cornillet
Paolo Costa
Cottigny
Coûteaux
Cramer
Corina Creţu
Gabriela Creţu
Crowley
Csibi
Marek Aleksander Czarnecki
Ryszard Czarnecki
Dăianu
Daul
David
Davies
De Blasio
de Brún
Degutis
De Keyser
Deprez
De Rossa
De Sarnez
Descamps
Désir
Deß
Deva
De Veyrac
De Vits
Dičkutė
Didžiokas
Dillen
Dimitrakopoulos
Dombrovskis
Doorn
Dover
Doyle
Drčar Murko
Duchoň
Dührkop Dührkop
Duff
Duka-Zólyomi
Dumitriu
Ehler
Ek
Elles
Estrela
Ettl
Jill Evans
Jonathan Evans
Färm
Falbr
Farage
Fava
Fazakas
Ferber
Fernandes
Fernández Martín
Ferrari
Anne Ferreira
Elisa Ferreira
Figueiredo
Flautre
Florenz
Foglietta
Foltyn-Kubicka
Fontaine
Ford
Fouré
Fourtou
Fraga Estévez
França
Frassoni
Friedrich
Frunzăverde
Gacek
Gál
Gaľa
Galeote
Garcés Ramón
García Pérez
Garriga Polledo
Gaubert
Gauzès
Gawronski
Gebhardt
Gentvilas
Georgiou
Geremek
Geringer de Oedenberg
Gewalt
Gierek
Giertych
Gill
Gklavakis
Glante
Glattfelder
Goebbels
Goepel
Golik
Gollnisch
Gomolka
Gottardi
Goudin
Grabowska
Graça Moura
Graefe zu Baringdorf
Gräßle
Grech
Griesbeck
de Groen-Kouwenhoven
Groote
Grosch
Grossetête
Guardans Cambó
Guellec
Guerreiro
Guidoni
Gurmai
Gutiérrez-Cortines
Guy-Quint
Gyürk
Hall
Hammerstein
Hamon
Handzlik
Hannan
Harbour
Harkin
Hassi
Haug
Heaton-Harris
Hedh
Helmer
Hennicot-Schoepges
Hennis-Plasschaert
Herczog
Herranz García
Hieronymi
Higgins
Hökmark
Honeyball
Hoppenstedt
Horáček
Howitt
Hudacký
Hudghton
Hughes
Hutchinson
Hyusmenova
Iacob-Ridzi
in 't Veld
Irujo Amezaga
Itälä
Iturgaiz Angulo
Jackson
Jacobs
Jäätteenmäki
Jałowiecki
Janowski
Járóka
Jeggle
Jeleva
Jensen
Jöns
Jørgensen
Jordan Cizelj
Jouye de Grandmaison
Kacin
Kaczmarek
Kallenbach
Kamall
Karas
Kaufmann
Kauppi
Kazak
Tunne Kelam
Kindermann
Kinnock
Kirilov
Klamt
Klaß
Knapman
Koch
Kohlíček
Konrad
Koterec
Kozlík
Krahmer
Krasts
Kratsa-Tsagaropoulou
Krehl
Kreissl-Dörfler
Kristovskis
Krupa
Kuc
Kuhne
Kušķis
Kusstatscher
Kuźmiuk
Laignel
Lamassoure
Lambert
Lambrinidis
Lambsdorff
Lang
De Lange
Langen
Langendries
Laperrouze
La Russa
Lavarra
Lax
Lebech
Le Foll
Lefrançois
Lehideux
Lehne
Lehtinen
Leichtfried
Jean-Marie Le Pen
Le Rachinel
Lewandowski
Liberadzki
Libicki
Lienemann
Lipietz
Locatelli
López-Istúriz White
Louis
Ludford
Lulling
Lundgren
Lynne
Lyubcheva
Maaten
McAvan
McCarthy
McGuinness
McMillan-Scott
Madeira
Maldeikis
Manders
Maňka
Erika Mann
Thomas Mann
Marinescu
Markov
Marques
David Martin
Hans-Peter Martin
Martinez
Martínez Martínez
Masiel
Masip Hidalgo
Maštálka
Mathieu
Mato Adrover
Matsakis
Mauro
Mavrommatis
Mayer
Mayor Oreja
Medina Ortega
Meijer
Méndez de Vigo
Menéndez del Valle
Miguélez Ramos
Mikolášik
Millán Mon
Mitchell
Mölzer
Mohácsi
Moreno Sánchez
Morgan
Morgantini
Morillon
Morin
Mote
Mulder
Musacchio
Muscardini
Musotto
Mussolini
Musumeci
Napoletano
Nassauer
Nattrass
Navarro
Nechifor
Neris
Newton Dunn
Neyts-Uyttebroeck
Nicholson
Niculescu
Niebler
van Nistelrooij
Novak
Olajos
Olbrycht
Ó Neachtain
Onesta
Onyszkiewicz
Oomen-Ruijten
Oprea
Őry
Ouzký
Oviir
Paasilinna
Pack
Pahor
Paleckis
Panayotopoulos-Cassiotou
Panayotov
Pannella
Panzeri
Papadimoulis
Paparizov
Papastamkos
Parish
Paşcu
Patriciello
Patrie
Peillon
Alojz Peterle
Petre
Pflüger
Piecyk
Pieper
Pīks
Pinheiro
Pinior
Piotrowski
Pirker
Pittella
Pleguezuelos Aguilar
Pleštinská
Plumb
Podimata
Podkański
Pöttering
Pohjamo
Pomés Ruiz
Mihaela Popa
Nicolae Vlad Popa
Posselt
Prets
Vittorio Prodi
Protasiewicz
Purvis
Queiró
Quisthoudt-Rowohl
Rack
Radwan
Raeva
Ransdorf
Rapkay
Rasmussen
Remek
Resetarits
Reul
Ribeiro e Castro
Riera Madurell
Ries
Riis-Jørgensen
Rivera
Rizzo
Rogalski
Roithová
Romeva i Rueda
Rosati
Roszkowski
Roth-Behrendt
Rothe
Rouček
Roure
Rovsing
Rudi Ubeda
Rübig
Rühle
Rutowicz
Ryan
Sacconi
Saïfi
Sakalas
Saks
Salafranca Sánchez-Neyra
Sánchez Presedo
dos Santos
Sartori
Saryusz-Wolski
Savi
Sbarbati
Schaldemose
Scheele
Schenardi
Schierhuber
Schinas
Schlyter
Frithjof Schmidt
Olle Schmidt
Schnellhardt
Schöpflin
Jürgen Schröder
Schroedter
Schulz
Schuth
Schwab
Seeber
Segelström
Seppänen
Severin
Siekierski
Silva Peneda
Simpson
Sinnott
Siwiec
Skinner
Škottová
Smith
Sógor
Sommer
Søndergaard
Sonik
Speroni
Staes
Staniszewska
Starkevičiūtė
Šťastný
Stavreva
Sterckx
Stevenson
Stihler
Stockmann
Stolojan
Strejček
Strož
Stubb
Sturdy
Sudre
Sumberg
Surján
Svensson
Szájer
Szejna
Szent-Iványi
Szymański
Tabajdi
Tajani
Takkula
Tannock
Tarand
Tatarella
Thomsen
Thyssen
Ţicău
Titford
Titley
Toia
Tőkés
Tomaszewska
Trakatellis
Trautmann
Triantaphyllides
Trüpel
Turmes
Ulmer
Vakalis
Vălean
Vanhecke
Van Orden
Varela Suanzes-Carpegna
Varvitsiotis
Vatanen
Vaugrenard
Ventre
Veraldi
Vergnaud
Vernola
Vidal-Quadras
Vigenin
de Villiers
Virrankoski
Visser
Vlasto
Voggenhuber
Wallis
Walter
Watson
Henri Weber
Manfred Weber
Renate Weber
Weisgerber
Westlund
Whittaker
Wiersma
Willmott
Iuliu Winkler
Wise
von Wogau
Wohlin
Bernard Wojciechowski
Janusz Wojciechowski
Wortmann-Kool
Wurtz
Yañez-Barnuevo García
Záborská
Zaleski
Zapałowski
Zappalà
Ždanoka
Zdravkova
Železný
Zieleniec
Zingaretti
Zlotea
Zvěřina
Zwiefka
Lissabonfördraget
Europaparlamentets resolution av den 20 februari 2008 om Lissabonfördraget (2007/2286(INI))
Folk- och bostadsräkningar
Europaparlamentets ståndpunkt fastställd vid första behandlingen den 20 februari 2008 inför antagandet av Europaparlamentets och rådets förordning (EG) nr .../2008 om folk- och bostadsräkningar
Lissabonstrategin
Europaparlamentets resolution av den 20 februari 2008 om bidraget till diskussionerna om Lissabonstrategin vid Europeiska rådets vårmöte 2008
Riktlinjerna för den allmänna ekonomiska politiken 2008–2010
Europaparlamentets resolution av den 20 februari 2008 om de integrerade riktlinjerna för tillväxt och sysselsättning (del: allmänna riktlinjer för medlemsstaternas och gemenskapens ekonomiska politik): start för den nya treårsperioden (2008–2010) (KOM(2007)0803 – 2007/2275(INI))
En EU-strategi för Centralasien
Europaparlamentets resolution av den 20 februari 2008 om en EU-strategi för Centralasien (2007/2102(INI))
TECKENFÖRKLARING
*
Samrådsförfarandet
** I
** II
***
Samtyckesförfarandet
***I
Medbeslutandeförfarandet (första behandlingen)
***II
Medbeslutandeförfarandet (andra behandlingen)
***III
UPPLYSNINGAR ANGÅENDE OMRÖSTNINGAR
Om inget annat anges har föredraganden till talmannen skriftligen tillkännagivit sin inställning till ändringsförslagen.
FÖRKORTNINGAR FÖR UTSKOTTENS NAMN
AFET:
DEVE:
Utskottet för utveckling
INTA:
Utskottet för internationell handel
BUDG:
Budgetutskottet
CONT:
Budgetkontrollutskottet
ECON:
Utskottet för ekonomi och valutafrågor
EMPL:
Utskottet för sysselsättning och sociala frågor
ENVI:
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
ITRE:
Utskottet för industrifrågor, forskning och energi
IMCO:
Utskottet för den inre marknaden och konsumentskydd
TRAN:
Utskottet för transport och turism
REGI:
Utskottet för regional utveckling
AGRI:
PECH:
Fiskeriutskottet
CULT:
Utskottet för kultur och utbildning
JURI:
Utskottet för rättsliga frågor
LIBE:
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
AFCO:
Utskottet för konstitutionella frågor
FEMM:
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
PETI:
Utskottet för framställningar
FÖRKORTNINGAR FÖR DE POLITISKA GRUPPERNA
PPE-DE:
Gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater
PSE:
Europeiska socialdemokratiska partiets grupp
ALDE:
Gruppen Alliansen liberaler och demokrater för Europa
UEN:
Gruppen Unionen för nationernas Europa
Verts/ALE
Gruppen De gröna/Europeiska fria alliansen
GUE/NGL:
Gruppen Europeiska enade vänstern/Nordisk grön vänster
IND/DEM:
Gruppen Självständighet/Demokrati
NI:
Grupplösa
Öppnande av den årliga sessionen
Öppnande av sammanträdet
Uttalande av talmannen
Kommissionens åtgärder till följd av parlamentets resolutioner
Inkomna dokument
Debatt om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer (tillkännagivande av ingivna resolutionsförslag)
Årlig politisk strategi 2009 (debatt)
Europeiska institutet för innovation och teknik ***II (debatt)
Valprövning
Omröstning
Förvaltningen av tillgångarna i EKSG och Kol- och stålforskningsfonden * (artikel 131 i arbetsordningen) (omröstning)
Avtal mellan EG och Förenade Arabemiraten om vissa luftfartsaspekter * (artikel 131 i arbetsordningen) (omröstning)
Gemensam organisation av jordbruksmarknaderna (ändring av enda förordningen om de gemensamma organisationerna av marknaden) * (artikel 131 i arbetsordningen) (omröstning)
Gemensam organisation av jordbruksmarknaderna (enda förordningen om de gemensamma organisationerna av marknaden) * (artikel 131 i arbetsordningen) (omröstning)
Statistisk näringsgrensindelning i EG (kodifierad version) ***I (artikel 131 i arbetsordningen) (omröstning)
Identifikation och registrering av svin (kodifierad version) * (artikel 131 i arbetsordningen) (omröstning)
Saluförande av plantmaterial av grönsaker (kodifierad version) * (artikel 131 i arbetsordningen) (omröstning)
Gemensamma skyddsregler för den civila luftfarten ***III (omröstning)
Europeiska institutet för innovation och teknik ***II (omröstning)
Utnyttjande av EU:s solidaritetsfond (omröstning)
Ändringsbudget nr 1/2008 - Solidaritetsfonden (omröstning)
Partnerskapsavtal om fiske mellan EG och Guinea-Bissau * (omröstning)
Partnerskapsavtal om fiske mellan EG och Elfenbenskusten * (omröstning)
En hållbar europeisk transportpolitik (omröstning)
Högtidligt möte - Estland
Röstförklaringar
Rättelser/avsiktsförklaringar till avgivna röster
Föredragningslista
Justering av protokollet från föregående sammanträde
Gemensam organisation av jordbruksmarknaderna och särskilda bestämmelser för de nationella kvoterna för mjölk * (debatt)
"Hälsokontroll" av den gemensamma jordbrukspolitiken (debatt)
Uppföljning efter översynen av Lamfalussyprocessen (debatt)
Frågestund (frågor till kommissionen)
Kvinnornas situation i EU:s landsbygdsområden (debatt)
Hållbart jordbruk och biogas: behov av översyn av EU-lagstiftningen (debatt)
Energistatistik ***I (debatt)
Statistik om växtskyddsmedel ***I (debatt)
Föredragningslista för nästa sammanträde
Avslutande av sammanträdet
NÄRVAROLISTA
EUROPAPARLAMENTET
STRASBOURG
PROTOKOLL
ORDFÖRANDESKAP: Hans-Gert PÖTTERING Talman
2 Öppnande av sammanträdet
Sammanträdet öppnades kl. 09.00.
3 Uttalande av talmannen
Talmannen fördömde ännu en gång alla terrordåd och uttryckte på parlamentets vägnar sin medkänsla med offrens familjer.
Parlamentet höll en tyst minut för att hedra minnet av alla dem som fallit offer för terrorismen.
5 Inkomna dokument
Talmannen hade mottagit följande dokument:
1) från rådet och kommissionen
- Förslag till Europaparlamentets och rådets direktiv om leksakers säkerhet ( KOM(2008)0009 - C6-0039/2008 - 2008/0018(COD) )
hänvisat till
ansvarigt utskott :
IMCO
rådgivande utskott :
ENVI, ITRE
- Förslag till Europaparlamentets och rådets direktiv om skyddsbågar på jordbruks- eller skogsbrukstraktorer med hjul (statisk provning) (kodifierad version) ( KOM(2008)0025 - C6-0044/2008 - 2008/0008(COD) )
hänvisat till
ansvarigt utskott :
JURI
- Förslag till Europaparlamentets och rådets förordning om livsmedelsinformation till konsumenterna ( KOM(2008)0040 - C6-0052/2008 - 2008/0028(COD) )
hänvisat till
ansvarigt utskott :
ENVI
rådgivande utskott :
IMCO
- Förslag till Europaparlamentets och rådets beslut om ändring av rådets direktiv 76/769/EEG med avseende på begränsningar för utsläppande på marknaden och användning av vissa farliga ämnen och preparat (diklormetan) (Ändring av rådets direktiv 76/769/EEG) ( KOM(2008)0080 - C6-0068/2008 - 2008/0033(COD) )
hänvisat till
ansvarigt utskott :
ENVI
rådgivande utskott :
IMCO
- Förslag till anslagsöverföring DEC 03/2008 - Avsnitt III - Kommissionen ( SEK(2008)0016 - C6-0077/2008 - 2008/2042(GBD))
hänvisat till
ansvarigt utskott :
BUDG
hänvisat till
ansvarigt utskott :
CONT
rådgivande utskott :
DEVE, BUDG
hänvisat till
ansvarigt utskott :
CONT
rådgivande utskott :
DEVE, BUDG
hänvisat till
ansvarigt utskott :
CONT
rådgivande utskott :
DEVE, BUDG
hänvisat till
ansvarigt utskott :
CONT
rådgivande utskott :
DEVE, BUDG
- Rådets rekommendation om beviljande av ansvarsfrihet för kommissionen för genomförandet av budgeten för budgetåret 2006 (05842/2008 - C6-0082/2008 - 2007/2037(DEC) )
hänvisat till
ansvarigt utskott :
CONT
rådgivande utskott :
PETI, FEMM, AFCO, DEVE, CULT, AFET, PECH, AGRI, ENVI, EMPL, BUDG, ITRE, JURI, ECON, LIBE, INTA, IMCO, TRAN, REGI
- Rådets rekommendation om beviljande av ansvarsfrihet för genomförandeorganen för genomförandet av budgeten för budgetåret 2006 (05855/2008 - C6-0083/2008 - 2007/2037(DEC) )
hänvisat till
ansvarigt utskott :
CONT
rådgivande utskott :
PETI, FEMM, AFCO, DEVE, CULT, AFET, PECH, AGRI, ENVI, EMPL, BUDG, ITRE, JURI, ECON, LIBE, INTA, IMCO, TRAN, REGI
- Ansvarsfrihet för Europeiska gemenskapernas organ för genomförandet av budgeten för budgetåret 2006 (05843/2008 - C6-0084/2008 - 2007/2046(DEC) )
hänvisat till
ansvarigt utskott :
CONT
rådgivande utskott :
EMPL
- Förslag till Europaparlamentets och rådets beslut om att utnyttja Europeiska fonden för justering för globaliseringseffekter ( KOM(2008)0094 - C6-0085/2008 - 2008/2043(ACI) )
hänvisat till
ansvarigt utskott :
BUDG
rådgivande utskott :
EMPL
- Förslag till Europaparlamentets och rådets förordning om ändring av förordning (EG) nr 562/2006 när det gäller användningen av informationssystemet för viseringar (VIS) enligt kodexen om Schengengränserna ( KOM(2008)0101 - C6-0086/2008 - 2008/0041(COD) )
hänvisat till
ansvarigt utskott :
LIBE
rådgivande utskott :
DEVE, AFET
- Anpassning till det föreskrivande förfarandet med kontroll - Förslag till Europaparlamentets och rådets förordning om ändring av rådets förordning (EG) nr 338/97 om skyddet av arter av vilda djur och växter genom kontroll av handeln med dem när det gäller kommissionens genomförandebefogenheter ( KOM(2008)0104 - C6-0087/2008 - 2008/0042(COD) )
hänvisat till
ansvarigt utskott :
ENVI
rådgivande utskott :
JURI
- Anpassning till det föreskrivande förfarandet med kontroll - Förslag till Europaparlamentets och rådets direktiv om ändring av kommissionens genomförandebefogenheter enligt rådets direktiv 79/409/EEG om bevarande av vilda fåglar ( KOM(2008)0105 - C6-0088/2008 - 2008/0038(COD) )
hänvisat till
ansvarigt utskott :
ENVI
rådgivande utskott :
JURI
- Förslaget till rådets och kommissionens beslut om ingående av protokollet till stabiliserings- och associeringsavtalet mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och f.d. jugoslaviska republiken Makedonien, å andra sidan, med anledning av Republiken Bulgariens och Rumäniens anslutning till Europeiska unionen (16731/2007 - C6-0093/2008 - 2007/0218(AVC) )
hänvisat till
ansvarigt utskott :
AFET
rådgivande utskott :
INTA
- Förslag till Europaparlamentets och rådets direktiv om provning av motorfordons och tillhörande släpfordons trafiksäkerhet (omarbetad version) ( KOM(2008)0100 - C6-0094/2008 - 2008/0044(COD) )
hänvisat till
ansvarigt utskott :
JURI
rådgivande utskott :
TRAN
- Förslag till rådets direktiv om allmänna regler för punktskatt ( KOM(2008)0078 - C6-0099/2008 - 2008/0051(CNS) )
hänvisat till
ansvarigt utskott :
ECON
rådgivande utskott :
AGRI, ITRE, CONT, IMCO, REGI
- Förslag till ändringsbudget nr 1 för budgetåret 2008 - Avsnitt III – Kommissionen (07259/2008 - C6-0124/2008 - 2008/2017(BUD) )
hänvisat till
ansvarigt utskott :
BUDG
hänvisat till
ansvarigt utskott :
JURI
2) från parlamentets utskott
2.1) betänkanden:
- Betänkande om begäran om upphävande av Hans-Peter Martins immunitet ( 2007/2215(IMM) ) - utskottet JURI - Föredragande: Diana Wallis ( A6-0071/2008 )
6 Debatt om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer (tillkännagivande av ingivna resolutionsförslag)
Nedanstående ledamöter eller politiska grupper hade, i enlighet med artikel 115 i arbetsordningen, begärt en debatt om följande resolutionsförslag:
I.
Armenien
-
Marie Anne Isler Béguin för Verts/ALE-gruppen
, om Armenien (
B6-0110/2008
),
-
Pasqualina Napoletano ,
Jan Marinus Wiersma ,
Hannes Swoboda och
Alexandra Dobolyi för PSE-gruppen
, om situationen i Armenien (
B6-0113/2008
),
-
Árpád Duka-Zólyomi ,
Urszula Gacek ,
Bernd Posselt och
Eija-Riitta Korhola för PPE-DE-gruppen
, om Armenien (
B6-0114/2008
),
-
Jaromír Kohlíček för GUE/NGL-gruppen
, om Armenien (
B6-0119/2008
),
-
Marios Matsakis ,
Annemie Neyts-Uyttebroeck och
Marco Cappato för ALDE-gruppen
, om situationen i Armenien (
B6-0120/2008
),
-
Ryszard Czarnecki ,
Adam Bielan och
Ewa Tomaszewska för UEN-gruppen , om Armenien (
B6-0121/2008 ).
II.
Gripande av demonstranter efter presidentvalet i Ryssland
-
Bernd Posselt ,
Jana Hybášková ,
Christopher Beazley ,
Tunne Kelam och
Thomas Mann för PPE-DE-gruppen , om gripandet av demonstranter efter presidentvalet i Ryssland (
B6-0124/2008 ),
-
Janusz Onyszkiewicz och
Annemie Neyts-Uyttebroeck för ALDE-gruppen
, om gripandet av demonstranter efter presidentvalet i Ryssland (
B6-0127/2008
),
-
Bart Staes och
Milan Horáček för Verts/ALE-gruppen
, om gripandet av demonstranter efter presidentvalet i Ryssland (
B6-0128/2008
),
-
Jan Marinus Wiersma och
Hannes Swoboda för PSE-gruppen
, om demonstrationerna i Ryssland efter presidentvalet (
B6-0129/2008
),
-
Ryszard Czarnecki ,
Adam Bielan ,
Hanna Foltyn-Kubicka ,
Ģirts Valdis Kristovskis ,
Ewa Tomaszewska ,
Konrad Szymański ,
Marcin Libicki ,
Roberts Zīle och
Mieczysław Edmund Janowski för UEN-gruppen , om gripandet av demonstranter efter presidentvalet i Ryssland (
B6-0130/2008 ).
III.
Fallet med journalisten Perwez Kambakhsh - Fallet med den iranske medborgaren Seyed Mehdi Kazemi
Perwez Kambakhsh
-
Angelika Beer ,
Joost Lagendijk och
Hélène Flautre för Verts/ALE-gruppen , om Afghanistan (
B6-0112/2008 ),
-
Thomas Mann ,
Guido Podestà ,
Eija-Riitta Korhola och
Nicole Fontaine för PPE-DE-gruppen
, om den afghanske medborgare som dömts av islamiska domstolar (
B6-0115/2008
),
-
Adam Bielan ,
Ryszard Czarnecki och
Ewa Tomaszewska för UEN-gruppen , om fallet med journalisten Perwez Kambakhsh (
B6-0116/2008 ),
-
Pasqualina Napoletano ,
Ana Maria Gomes ,
Robert Evans ,
Elena Valenciano Martínez-Orozco och
Emilio Menéndez del Valle för PSE-gruppen , om fallet med journalisten Perwez Kambakhsh (
B6-0118/2008 );
-
Francis Wurtz och
André Brie för GUE/NGL-gruppen
, om Afghanistan: fallet med journalisten Perwez Kambakhsh (
B6-0123/2008
),
-
Jules Maaten ,
Marios Matsakis och
Marco Cappato för ALDE-gruppen , om Afghanistan (
B6-0125/2008 ).
Seyed Mehdi Kazemi
-
Jean Lambert och
Raül Romeva i Rueda för Verts/ALE-gruppen , om fallet Mehdi Kazemi (
B6-0111/2008 ),
-
Pasqualina Napoletano och
Michael Cashman för PSE-gruppen , om fallet Mehdi Kazemi (
B6-0117/2008 ),
-
Vittorio Agnoletto för GUE/NGL-gruppen , om fallet Mehdi Kazemi (
B6-0122/2008 ),
-
Marco Cappato ,
Marco Pannella ,
Sophia in 't Veld ,
Jeanine Hennis-Plasschaert ,
Sarah Ludford och
Marios Matsakis för ALDE-gruppen , om fallet Mehdi Kazemi (
B6-0126/2008 ).
Talartiden fördelas i enlighet med artikel 142 i arbetsordningen.
7
Årlig politisk strategi 2009 (debatt)
Uttalande av kommissionen:
Årlig politisk strategi 2009
José Manuel Barroso (kommissionens ordförande) gjorde ett uttalande.
Talare:
Hartmut Nassauer för PPE-DE-gruppen,
Hannes Swoboda för PSE-gruppen,
Diana Wallis för ALDE-gruppen,
Brian Crowley för UEN-gruppen,
Eva Lichtenberger för Verts/ALE-gruppen,
Helmuth Markov för GUE/NGL-gruppen,
Godfrey Bloom för IND/DEM-gruppen,
Frank Vanhecke , grupplös,
José Ignacio Salafranca Sánchez-Neyra ,
Catherine Guy-Quint ,
Adina-Ioana Vălean ,
Jan Tadeusz Masiel ,
Jens-Peter Bonde ,
Luca Romagnoli ,
László Surján ,
Véronique De Keyser ,
Ingeborg Gräßle ,
Alain Hutchinson ,
Lambert van Nistelrooij ,
Göran Färm ,
Lutz Goepel ,
Carmen Fraga Estévez ,
John Bowis ,
Maria Martens ,
Jacek Saryusz-Wolski och
Othmar Karas .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Mairead McGuinness ,
Luís Queiró ,
Katalin Lévai ,
Zuzana Roithová och
Danutė Budreikaitė .
Talare:
Margot Wallström (kommissionens vice ordförande) .
Då de resolutionsförslag som lagts fram ännu inte fanns tillgängliga, skulle de tillkännages vid en senare tidpunkt.
Talmannen förklarade debatten avslutad.
Omröstning:
8
Europeiska institutet för innovation och teknik ***II (debatt)
Andrabehandlingsrekommendation om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets förordning om inrättande av Europeiska institutet för innovation och teknik [15647/1/2007 - C6-0035/2008 - 2006/0197(COD) ] - Utskottet för industrifrågor, forskning och energi.
Föredragande: Reino Paasilinna ( A6-0041/2008 )
Reino Paasilinna redogjorde för andrabehandlingsrekommendationen.
Talare:
Ján Figeľ (ledamot av kommissionen) .
ORDFÖRANDESKAP: Luigi COCILOVO Vice talman
Talare:
Romana Jordan Cizelj för PPE-DE-gruppen,
Hannes Swoboda för PSE-gruppen,
Jorgo Chatzimarkakis för ALDE-gruppen,
Konrad Szymański för UEN-gruppen,
Miloslav Ransdorf för GUE/NGL-gruppen,
Jana Bobošíková , grupplös,
Angelika Niebler ,
Gyula Hegyi ,
Lena Ek ,
Ryszard Czarnecki ,
Zdzisław Kazimierz Chmielewski ,
Teresa Riera Madurell ,
Grażyna Staniszewska och
Pierre Pribetich .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Lambert van Nistelrooij ,
Lidia Joanna Geringer de Oedenberg ,
Jacek Protasiewicz ,
Erna Hennicot-Schoepges ,
Marusya Ivanova Lyubcheva ,
Sylwester Chruszcz ,
Miroslav Mikolášik ,
Nina Škottová och
Czesław Adam Siekierski .
Talare:
Ján Figeľ och
Reino Paasilinna .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 10.9 i protokollet av den 11.03.2008
.
11.15
, i avvaktan på omröstningen, och återupptogs kl.
11.30
.)
ORDFÖRANDESKAP: Edward McMILLAN-SCOTT Vice talman
9 Valprövning
Giuseppe Gargani , ordförande för utskottet JURI, redogjorde muntligen för utskottets förslag beträffande valprövning av följande ledamöter:
Roberta Alma Anastase ,
Sebastian Valentin Bodu ,
Victor Boştinaru ,
Nicodim Bulzesc ,
Cristian Silviu Buşoi ,
Titus Corlăţean ,
Corina Creţu ,
Gabriela Creţu ,
Magor Imre Csibi ,
Daniel Dăianu ,
Dragoş Florin David ,
Constantin Dumitriu ,
Petru Filip ,
Sorin Frunzăverde ,
Monica Maria Iacob-Ridzi ,
Ramona Nicole Mănescu ,
Marian-Jean Marinescu ,
Cătălin-Ioan Nechifor ,
Rareş-Lucian Niculescu ,
Dumitru Oprea ,
Ioan Mircea Paşcu ,
Maria Petre ,
Rovana Plumb ,
Mihaela Popa ,
Nicolae Vlad Popa ,
Daciana Octavia Sârbu ,
Adrian Severin ,
Csaba Sógor ,
Theodor Dumitru Stolojan ,
Silvia-Adriana Ţicău ,
László Tőkés ,
Adina-Ioana Vălean ,
Renate Weber ,
Iuliu Winkler och
Urszula Gacek och
Parlamentet beslutade att godkänna mandaten för dessa ledamöter.
10 Omröstning
Omröstningsresultaten (ändringsförslag, särskilda omröstningar, delade omröstningar etc.) återfinns i bilagan ”Omröstningsresultat” som bifogas protokollet.
Bilagan med resultaten av omröstningarna med namnupprop finns endast i elektronisk form på Europarl.
10.1
Förvaltningen av tillgångarna i EKSG och Kol- och stålforskningsfonden * (artikel 131 i arbetsordningen) (omröstning)
Betänkande om förslaget till rådets beslut om ändring av rådets beslut 2003/77/EG om fastställande av fleråriga ekonomiska riktlinjer för förvaltningen av tillgångarna i EKSG under avveckling och, efter slutförd avveckling, av Kol- och stålforskningsfondens tillgångar [ KOM(2007)0435 - C6-0276/2007 - 2007/0150(CNS) ] - Budgetutskottet.
Föredragande: Reimer Böge ( A6-0062/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 1)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs genom en enda omröstning
(
P6_TA(2008)0073
)
10.2
Avtal mellan EG och Förenade Arabemiraten om vissa luftfartsaspekter * (artikel 131 i arbetsordningen) (omröstning)
Betänkande om förslaget till rådets beslut om ingående av ett avtal mellan Europeiska gemenskapen och Förenade Arabemiraten om vissa luftfartsaspekter [ KOM(2007)0134 - C6-0472/2007 - 2007/0052(CNS) ] - Utskottet för transport och turism.
Föredragande: Paolo Costa ( A6-0043/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 2)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs genom en enda omröstning
(
P6_TA(2008)0074
)
10.3
Gemensam organisation av jordbruksmarknaderna (ändring av enda förordningen om de gemensamma organisationerna av marknaden) * (artikel 131 i arbetsordningen) (omröstning)
Betänkande om förslaget till rådets förordning om ändring av förordning (EG) nr 1234/2007 om upprättande av en gemensam organisation av jordbruksmarknaderna och om särskilda bestämmelser för vissa jordbruksprodukter (”enda förordningen om de gemensamma organisationerna av marknaden”) [ KOM(2007)0854 - C6-0033/2008 - 2007/0290(CNS) ] - Utskottet för jordbruk och landsbygdens utveckling.
Föredragande: Neil Parish ( A6-0044/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 3)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs genom en enda omröstning
(
P6_TA(2008)0075
)
10.4
Gemensam organisation av jordbruksmarknaderna (enda förordningen om de gemensamma organisationerna av marknaden) * (artikel 131 i arbetsordningen) (omröstning)
Betänkande om förslaget till rådets förordning om ändring av förordning (EG) nr 1234/2007 om upprättande av en gemensam organisation av jordbruksmarknaderna och om särskilda bestämmelser för vissa jordbruksprodukter (enda förordningen om de gemensamma organisationerna av marknaden) [ KOM(2008)0027 - C6-0061/2008 - 2008/0011(CNS) ] - Utskottet för jordbruk och landsbygdens utveckling.
Föredragande: Neil Parish ( A6-0045/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 4)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs genom en enda omröstning
(
P6_TA(2008)0076
)
10.5
Statistisk näringsgrensindelning i EG (kodifierad version) ***I (artikel 131 i arbetsordningen) (omröstning)
Betänkande om förslaget till Europaparlamentets och rådets förordning om statistisk näringsgrensindelning i Europeiska gemenskapen (kodifierad version) [ KOM(2007)0755 - C6-0437/2007 - 2007/0256(COD) ] - Utskottet för rättsliga frågor.
Föredragande: Lidia Joanna Geringer de Oedenberg ( A6-0055/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 5)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs genom en enda omröstning
(
P6_TA(2008)0077
)
10.6
Identifikation och registrering av svin (kodifierad version) * (artikel 131 i arbetsordningen) (omröstning)
Betänkande om förslaget till rådets direktiv om identifikation och registrering av svin (kodifierad version) [ KOM(2007)0829 - C6-0037/2008 - 2007/0294(CNS) ] - Utskottet för rättsliga frågor.
Föredragande: Lidia Joanna Geringer de Oedenberg ( A6-0057/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 6)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs genom en enda omröstning
(
P6_TA(2008)0078
)
10.7
Saluförande av plantmaterial av grönsaker (kodifierad version) * (artikel 131 i arbetsordningen) (omröstning)
Betänkande om förslaget till rådets direktiv om saluförande av annat föröknings- och plantmaterial av grönsaker än utsäde (kodifierad version) [ KOM(2007)0852 - C6-0038/2008 - 2007/0296(CNS) ] - Utskottet för rättsliga frågor.
Föredragande: Lidia Joanna Geringer de Oedenberg ( A6-0056/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 7)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs genom en enda omröstning
(
P6_TA(2008)0079
)
10.8
Gemensamma skyddsregler för den civila luftfarten ***III (omröstning)
Betänkande om förlikningskommitténs gemensamma utkast till Europaparlamentets och rådets förordning om gemensamma skyddsregler för den civila luftfarten och om upphävande av förordning (EG) nr 2320/2002 [PE-CONS 3601/2008 – C6 0029/2008 – 2005/0191(COD) ] - Europaparlamentets delegation till förlikningskommittén - Föredragande:
Paolo Costa (
A6-0049/2008 )
(Enkel majoritet erfordrades för godkännande)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 8)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs (
P6_TA(2008)0080
)
10.9
Europeiska institutet för innovation och teknik ***II (omröstning)
Andrabehandlingsrekommendation om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets förordning om inrättande av Europeiska institutet för innovation och teknik [15647/1/2007 - C6-0035/2008 - 2006/0197(COD) ] - Utskottet för industrifrågor, forskning och energi.
Föredragande: Reino Paasilinna ( A6-0041/2008 )
(Kvalificerad majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 9)
RÅDETS GEMENSAMMA STÅNDPUNKT
Förklarades godkänt
(
P6_TA(2008)0081
)
10.10
Utnyttjande av EU:s solidaritetsfond (omröstning)
Betänkande om förslaget till Europaparlamentets och rådets beslut om utnyttjande av EU:s solidaritetsfond, med tillämpning av punkt 26 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning [ KOM(2008)0014 – C6 0036/2008 – 2008/2019(ACI) ] - Budgetutskottet.
Föredragande: Reimer Böge ( A6-0065/2008 )
(Kvalificerad majoritet och tre femtedelar av de avgivna rösterna erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 10)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2008)0082
)
10.11
Ändringsbudget nr 1/2008 - Solidaritetsfonden (omröstning)
Betänkande om ändringsbudget nr 1/2008 - Solidaritetsfonden Avsnitt III - Kommissionen [ 2008/2017(BUD) ] - Budgetutskottet.
Föredragande: Kyösti Virrankoski ( A6-0058/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 11)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2008)0083
)
10.12
Partnerskapsavtal om fiske mellan EG och Guinea-Bissau * (omröstning)
Betänkande om förslaget till rådets förordning om ingående av ett partnerskapsavtal om fiske mellan Europeiska gemenskapen och Republiken Guinea-Bissau [ KOM(2007)0580 - C6-0391/2007 - 2007/0209(CNS) ] - Fiskeriutskottet.
Föredragande: Luis Manuel Capoulas Santos ( A6-0053/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 12)
KOMMISSIONENS FÖRSLAG
Godkändes såsom ändrat av parlamentet
(
P6_TA(2008)0084
)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs
(
P6_TA(2008)0084
)
10.13
Partnerskapsavtal om fiske mellan EG och Elfenbenskusten * (omröstning)
Betänkande om förslaget till rådets förordning om ingående av ett partnerskapsavtal om fiske mellan Europeiska gemenskapen, å ena sidan, och Elfenbenskusten, å andra sidan [ KOM(2007)0648 - C6-0429/2007 - 2007/0226(CNS) ] - Fiskeriutskottet.
Föredragande: Daniel Varela Suanzes-Carpegna ( A6-0054/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 13)
KOMMISSIONENS FÖRSLAG
Godkändes såsom ändrat av parlamentet
(
P6_TA(2008)0085
)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs
(
P6_TA(2008)0085
)
10.14
En hållbar europeisk transportpolitik (omröstning)
Betänkande om en hållbar europeisk transportpolitik, med beaktande av EU:s energi- och miljöpolitik [ 2007/2147(INI) ] - Utskottet för transport och turism.
Föredragande: Gabriele Albertini ( A6-0014/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 14)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2008)0086
)
ORDFÖRANDESKAP: Hans-Gert PÖTTERING Talman
11 Högtidligt möte - Estland
ORDFÖRANDESKAP: Edward McMILLAN-SCOTT Vice talman
12 Röstförklaringar
Skriftliga röstförklaringar:
Muntliga röstförklaringar:
Betänkande Paolo Costa - A6-0049/2008 :
Hubert Pirker ,
Bernard Wojciechowski och
Jan Březina
Betänkande Reino Paasilinna - A6-0041/2008 :
Hubert Pirker ,
Zuzana Roithová ,
Tomáš Zatloukal ,
Hannu Takkula ,
Syed Kamall och
Christopher Heaton-Harris
Betänkande Reimer Böge - A6-0065/2008 :
Zuzana Roithová och
Glyn Ford
Betänkande Kyösti Virrankoski - A6-0058/2008 :
Zuzana Roithová ,
Bernard Wojciechowski och
Christopher Heaton-Harris
Betänkande Luis Manuel Capoulas Santos - A6-0053/2008 och
Betänkande Daniel Varela Suanzes-Carpegna - A6-0054/2008 :
Christopher Heaton-Harris
Betänkande Gabriele Albertini - A6-0014/2008 :
Christopher Heaton-Harris ,
Richard Seeber och
Zuzana Roithová
13 Rättelser/avsiktsförklaringar till avgivna röster
Den elektroniska versionen på Europarl uppdateras regelbundet under högst två veckor efter den aktuella omröstningsdagen.
Därefter slutförs förteckningen över rättelserna till de avgivna rösterna för att översättas och offentliggöras i Europeiska unionens officiella tidning.
° ° ° °
Victor Boştinaru hade låtit meddela att hans omröstningsapparat inte hade fungerat under hela omröstningen.
ORDFÖRANDESKAP: Miguel Angel MARTÍNEZ MARTÍNEZ Vice talman
14 Föredragningslista
Diana Wallis om begäran om upphävande av Hans-Peter Martins immunitet (
15 Justering av protokollet från föregående sammanträde
Protokollet från föregående sammanträde justerades.
16
Gemensam organisation av jordbruksmarknaderna och särskilda bestämmelser för de nationella kvoterna för mjölk * (debatt)
Betänkande om förslaget till rådets förordning om ändring av förordning (EG) nr 1234/2007 om upprättande av en gemensam organisation av jordbruksmarknaderna och om särskilda bestämmelser för vissa jordbruksprodukter ("enda förordningen om de gemensamma organisationerna av marknaden") vad gäller de nationella kvoterna för mjölk [ KOM(2007)0802 - C6-0015/2008 - 2007/0281(CNS) ] - Utskottet för jordbruk och landsbygdens utveckling.
Föredragande: Elisabeth Jeggle ( A6-0046/2008 )
Elisabeth Jeggle redogjorde för sitt betänkande.
Talare:
Czesław Adam Siekierski för PPE-DE-gruppen,
Rosa Miguélez Ramos för PSE-gruppen,
Niels Busk för ALDE-gruppen,
Alyn Smith för Verts/ALE-gruppen,
Dimitar Stoyanov , grupplös,
James Nicholson ,
Csaba Sándor Tabajdi ,
Margrete Auken ,
Albert Deß ,
Bogdan Golik ,
Astrid Lulling ,
Katerina Batzeli ,
Maria Petre ,
Gábor Harangozó och
Béla Glattfelder .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Miroslav Mikolášik ,
Zdzisław Zbigniew Podkański ,
Friedrich-Wilhelm Graefe zu Baringdorf ,
Jim Allister ,
Mairead McGuinness ,
Neil Parish ,
Agnes Schierhuber och
Esther De Lange .
Talare: Iztok Jarc,
Mariann Fischer Boel och
Elisabeth Jeggle .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 5.4 i protokollet av den 12.03.2008
.
17
"Hälsokontroll" av den gemensamma jordbrukspolitiken (debatt)
Betänkande om "hälsokontroll" av den gemensamma jordbrukspolitiken [ 2007/2195(INI) ] - Utskottet för jordbruk och landsbygdens utveckling.
Föredragande: Lutz Goepel ( A6-0047/2008 )
Lutz Goepel redogjorde för sitt betänkande.
Talare:
Iztok Jarc (rådets tjänstgörande ordförande) och
Mariann Fischer Boel (ledamot av kommissionen) .
Talare:
Bart Staes (föredragande av yttrande från utskottet ENVI) och
Neil Parish för PPE-DE-gruppen .
ORDFÖRANDESKAP: Marek SIWIEC Vice talman
Talare:
Luis Manuel Capoulas Santos för PSE-gruppen,
Niels Busk för ALDE-gruppen,
Sergio Berlato för UEN-gruppen,
Friedrich-Wilhelm Graefe zu Baringdorf för Verts/ALE-gruppen,
Ilda Figueiredo för GUE/NGL-gruppen,
Witold Tomczak för IND/DEM-gruppen,
Peter Baco , grupplös,
Agnes Schierhuber ,
Bernadette Bourzai ,
Willem Schuth ,
Janusz Wojciechowski ,
Alyn Smith ,
Kartika Tamara Liotard ,
Vladimír Železný ,
Jean-Claude Martinez ,
Mairead McGuinness ,
María Isabel Salinas García ,
Jan Mulder ,
Andrzej Tomasz Zapałowski ,
Marie-Hélène Aubert ,
Bairbre de Brún ,
Derek Roland Clark ,
Jim Allister ,
Véronique Mathieu ,
Csaba Sándor Tabajdi ,
Anne Laperrouze ,
Liam Aylward ,
Carmen Fraga Estévez ,
Lily Jacobs ,
Kyösti Virrankoski ,
Zdzisław Zbigniew Podkański ,
Petya Stavreva ,
Bogdan Golik ,
Magor Imre Csibi ,
Zbigniew Krzysztof Kuźmiuk ,
Czesław Adam Siekierski ,
Katerina Batzeli ,
Francesco Ferrari och
Struan Stevenson .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Constantin Dumitriu ,
James Nicholson ,
Andrzej Jan Szejna ,
Markus Pieper och
Marian Harkin .
Talare:
Iztok Jarc ,
Mariann Fischer Boel och
Lutz Goepel .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 5.5 i protokollet av den 12.03.2008
.
18
Uppföljning efter översynen av Lamfalussyprocessen (debatt)
Muntlig fråga (
O-0015/2008 ) från
Pervenche Berès , för utskottet ECON, till rådet:
Uppföljning efter översynen av Lamfalussyprocessen ( B6-0011/2008 )
Muntlig fråga (
O-0016/2008 ) från
Pervenche Berès , för utskottet ECON, till kommissionen:
Uppföljning efter översynen av Lamfalussyprocessen ( B6-0012/2008 )
Pervenche Berès utvecklade de muntliga frågorna.
Janez Lenarčič (rådets tjänstgörande ordförande) besvarade frågan (
B6-0011/2008 ).
ORDFÖRANDESKAP: Diana WALLIS Vice talman
Joaquín Almunia (ledamot av kommissionen) besvarade frågan (
B6-0012/2008 ).
Talare:
Alexander Radwan för PPE-DE-gruppen,
Ieke van den Burg för PSE-gruppen,
Josu Ortuondo Larrea för ALDE-gruppen,
Piia-Noora Kauppi ,
Elisa Ferreira ,
Antolín Sánchez Presedo och
Harald Ettl .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Reinhard Rack .
Talare:
Joaquín Almunia .
Talmannen förklarade debatten avslutad.
19
Frågestund (frågor till kommissionen)
Parlamentet behandlade en rad frågor till kommissionen (
B6-0013/2008 ).
Talare:
Marian Harkin yttrade sig om organisationen av frågestunden.
Första delen
Fråga 32 (Stavros Arnaoutakis): Negativa konsekvenser av den internationella kreditkrisen inom handeln
H-0075/08 .
Stavros Arnaoutakis och
H-0086/08 .
Manolis Mavrommatis och
H-0090/08 .
Avril Doyle ,
Lambert van Nistelrooij och
Marian Harkin .
H-0092/08 .
Colm Burke ,
Avril Doyle och
H-0100/08 .
Bernd Posselt ,
Justas Vincas Paleckis och
Talare:
Jim Higgins yttrade sig om hur frågestunden genomfördes.
Fråga 41 (Georgios Papastamkos): Lösning av tvisten i Världshandelsorganisationen mellan EU och Förenta staterna om genetiskt förändrade organismer
H-0076/08 .
Georgios Papastamkos och
H-0079/08 .
H-0080/08 .
H-0085/08 .
H-0122/08 .
H-0124/08 .
H-0153/08 .
Bart Staes ,
Glenis Willmott ,
David Martin ,
Sarah Ludford och
Paul Rübig .
(
) .
ORDFÖRANDESKAP: Mario MAURO Vice talman
20
Kvinnornas situation i EU:s landsbygdsområden (debatt)
Betänkande om kvinnornas situation i EU:s landsbygdsområden [ 2007/2117(INI) ] - Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män.
Föredragande: Christa Klaß ( A6-0031/2008 )
Christa Klaß redogjorde för sitt betänkande.
Talare:
Mariann Fischer Boel (ledamot av kommissionen) .
Talare:
Edit Bauer för PPE-DE-gruppen,
Iratxe García Pérez för PSE-gruppen,
Jan Tadeusz Masiel för UEN-gruppen,
Raül Romeva i Rueda för Verts/ALE-gruppen,
Ilda Figueiredo för GUE/NGL-gruppen,
Urszula Krupa för IND/DEM-gruppen,
Rodi Kratsa-Tsagaropoulou ,
Christa Prets ,
Zdzisław Zbigniew Podkański ,
Eva-Britt Svensson ,
Rumiana Jeleva ,
Ewa Tomaszewska ,
Esther Herranz García ,
Corina Creţu och
Lidia Joanna Geringer de Oedenberg .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Mairead McGuinness ,
Silvia-Adriana Ţicău ,
Danutė Budreikaitė ,
Avril Doyle ,
Roberta Alma Anastase ,
Anna Záborská och
Monica Maria Iacob-Ridzi .
Talare:
Mariann Fischer Boel och
Christa Klaß .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 5.6 i protokollet av den 12.03.2008
.
21
Hållbart jordbruk och biogas: behov av översyn av EU-lagstiftningen (debatt)
Betänkande om hållbart jordbruk och biogas: behov av översyn av EU-lagstiftningen [ 2007/2107(INI) ] - Utskottet för jordbruk och landsbygdens utveckling.
Föredragande: Csaba Sándor Tabajdi ( A6-0034/2008 )
Csaba Sándor Tabajdi redogjorde för sitt betänkande.
Talare:
Mariann Fischer Boel (ledamot av kommissionen) .
ORDFÖRANDESKAP: Rodi KRATSA-TSAGAROPOULOU Vice talman
Talare:
Jens Holm (föredragande av yttrande från utskottet ENVI),
Werner Langen (föredragande av yttrande från utskottet ITRE),
Albert Deß för PPE-DE-gruppen,
Bogdan Golik för PSE-gruppen,
Willem Schuth för ALDE-gruppen,
Wiesław Stefan Kuc för UEN-gruppen,
Friedrich-Wilhelm Graefe zu Baringdorf för Verts/ALE-gruppen,
Derek Roland Clark för IND/DEM-gruppen,
Jim Allister , grupplös,
Mairead McGuinness ,
Gábor Harangozó ,
Anne Laperrouze ,
Leopold Józef Rutowicz ,
Nils Lundgren ,
Neil Parish ,
Cristian Silviu Buşoi och
Samuli Pohjamo .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Miroslav Mikolášik ,
Avril Doyle ,
James Nicholson ,
Czesław Adam Siekierski och
Claude Turmes .
Talare:
Mariann Fischer Boel och
Csaba Sándor Tabajdi .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 5.7 i protokollet av den 12.03.2008
.
22
Energistatistik ***I (debatt)
Betänkande om förslaget till Europaparlamentets och rådets förordning om energistatistik [ KOM(2006)0850 - C6-0035/2007 - 2007/0002(COD) ] - Utskottet för industrifrågor, forskning och energi.
Föredragande: Claude Turmes ( A6-0487/2007 )
Talare:
Joaquín Almunia (ledamot av kommissionen) .
Claude Turmes redogjorde för sitt betänkande.
Talare:
Eija-Riitta Korhola för PPE-DE-gruppen,
Catherine Trautmann för PSE-gruppen,
Fiona Hall för ALDE-gruppen,
Avril Doyle ,
Teresa Riera Madurell ,
Jerzy Buzek och
Silvia-Adriana Ţicău .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Paul Rübig .
Talare:
Claude Turmes .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 5.2 i protokollet av den 12.03.2008
.
23
Statistik om växtskyddsmedel ***I (debatt)
Betänkande om förslaget till Europaparlamentets och rådets förordning om statistik om växtskyddsmedel [ KOM(2006)0778 - C6-0457/2006 - 2006/0258(COD) ] - Utskottet för miljö, folkhälsa och livsmedelssäkerhet.
Föredragande: Bart Staes ( A6-0004/2008 )
Talare:
Joaquín Almunia (ledamot av kommissionen) .
Bart Staes redogjorde för sitt betänkande.
Talare:
Hartmut Nassauer för PPE-DE-gruppen,
Gyula Hegyi för PSE-gruppen,
Marios Matsakis för ALDE-gruppen,
Hiltrud Breyer för Verts/ALE-gruppen,
Jens Holm för GUE/NGL-gruppen,
Irena Belohorská , grupplös,
Christa Klaß och
Péter Olajos .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Paul Rübig ,
Czesław Adam Siekierski ,
Avril Doyle och
Marios Matsakis .
Talare:
Bart Staes .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 5.3 i protokollet av den 12.03.2008
.
24 Föredragningslista för nästa sammanträde
Föredragningslistan för nästa sammanträde fastställdes ("Föredragningslista" PE 403.203/OJME).
25 Avslutande av sammanträdet
Sammanträdet avslutades kl. 23.55.
Harald R
ømer
Rodi Kratsa-Tsagaropoulou
Generalsekreterare
Vice talman
NÄRVAROLISTA
Följande skrev på:
Agnoletto
Aita
Albertini
Allister
Alvaro
Anastase
Andersson
Andrejevs
Andria
Angelakas
Angelilli
Arif
Arnaoutakis
Ashworth
Atkins
Attard-Montalto
Attwooll
Aubert
Audy
Auken
Ayala Sender
Aylward
Ayuso
Baco
Badia i Cutchet
Baeva
Barón Crespo
Barsi-Pataky
Battilocchio
Batzeli
Bauer
Beazley
Becsey
Belder
Belet
Belohorská
Beňová
Berend
Berès
Berlato
Berlinguer
Berman
Binev
Blokland
Bobošíková
Bodu
Böge
Bösch
Bonde
Bonsignore
Borghezio
Borrell Fontelles
Bossi
Boştinaru
Botopoulos
Bourzai
Bowis
Bowles
Bozkurt
Bradbourn
Braghetto
Brejc
Breyer
Březina
Brie
Brok
Brunetta
Budreikaitė
van Buitenen
Bulfon
Bullmann
Bulzesc
van den Burg
Burke
Bushill-Matthews
Busk
Buşoi
Busquin
Buzek
Cabrnoch
Calabuig Rull
Callanan
Camre
Capoulas Santos
Cappato
Carlshamre
Carnero González
Carollo
Casaca
Casini
Caspary
Castex
del Castillo Vera
Cederschiöld
Cercas
Chatzimarkakis
Chichester
Chiesa
Chmielewski
Christensen
Chruszcz
Chukolov
Claeys
Clark
Cocilovo
Coelho
Cohn-Bendit
Corbett
Corda
Corlăţean
Cornillet
Paolo Costa
Coûteaux
Cramer
Corina Creţu
Gabriela Creţu
Crowley
Csibi
Marek Aleksander Czarnecki
Ryszard Czarnecki
Dăianu
Daul
Davies
De Blasio
de Brún
Degutis
Dehaene
De Keyser
Demetriou
De Michelis
Deprez
De Rossa
Descamps
Désir
Deß
Deva
De Veyrac
De Vits
Díaz de Mera García Consuegra
Dičkutė
Didžiokas
Dillen
Dimitrakopoulos
Dobolyi
Dombrovskis
Donnici
Doorn
Douay
Dover
Doyle
Drčar Murko
Duchoň
Duff
Duka-Zólyomi
Dumitriu
Ebner
Ehler
Ek
El Khadraoui
Elles
Esteves
Estrela
Ettl
Jonathan Evans
Robert Evans
Färm
Fajmon
Falbr
Farage
Fatuzzo
Fava
Fazakas
Ferber
Fernandes
Fernández Martín
Ferrari
Anne Ferreira
Elisa Ferreira
Figueiredo
Filip
Fjellner
Flasarová
Flautre
Florenz
Foglietta
Foltyn-Kubicka
Fontaine
Ford
Fouré
Fourtou
Fraga Estévez
França
Frassoni
Friedrich
Frunzăverde
Gacek
Gahler
Gál
Gaľa
Garcés Ramón
García-Margallo y Marfil
García Pérez
Gargani
Garriga Polledo
Gaubert
Gauzès
Gawronski
Gebhardt
Gentvilas
Georgiou
Geremek
Geringer de Oedenberg
Gewalt
Gibault
Gierek
Giertych
Gill
Gklavakis
Glante
Glattfelder
Gobbo
Goebbels
Goepel
Golik
Gollnisch
Gomes
Gomolka
Gottardi
Goudin
Grabowska
Grabowski
Graça Moura
Graefe zu Baringdorf
Gräßle
de Grandes Pascual
de Groen-Kouwenhoven
Groote
Grosch
Grossetête
Guardans Cambó
Guellec
Guerreiro
Guidoni
Gurmai
Gutiérrez-Cortines
Guy-Quint
Gyürk
Hänsch
Hall
Hammerstein
Hamon
Handzlik
Hannan
Harangozó
Harbour
Harkin
Harms
Hasse Ferreira
Hassi
Haug
Heaton-Harris
Hedh
Hegyi
Helmer
Hennicot-Schoepges
Hennis-Plasschaert
Herranz García
Herrero-Tejedor
Hieronymi
Higgins
Hökmark
Holm
Hołowczyc
Honeyball
Hoppenstedt
Horáček
Howitt
Hudacký
Hudghton
Hutchinson
Hyusmenova
Iacob-Ridzi
Ibrisagic
in 't Veld
Iotova
Irujo Amezaga
Isler Béguin
Itälä
Iturgaiz Angulo
Jackson
Jacobs
Jäätteenmäki
Jałowiecki
Janowski
Járóka
Jarzembowski
Jeggle
Jeleva
Jensen
Jöns
Jørgensen
Jonckheer
Jordan Cizelj
Jouye de Grandmaison
Juknevičienė
Kacin
Kaczmarek
Kallenbach
Kamall
Karas
Karim
Kasoulides
Kaufmann
Kauppi
Kazak
Tunne Kelam
Kilroy-Silk
Kindermann
Kinnock
Kirilov
Kirkhope
Klamt
Klaß
Klinz
Knapman
Koch
Kohlíček
Konrad
Koppa
Korhola
Kósáné Kovács
Koterec
Kozlík
Krahmer
Krasts
Kratsa-Tsagaropoulou
Krehl
Kreissl-Dörfler
Kristovskis
Krupa
Kuc
Kuhne
Kułakowski
Kušķis
Kusstatscher
Kuźmiuk
Lagendijk
Lamassoure
Lambert
Lambrinidis
Lang
De Lange
Langen
Langendries
Laperrouze
La Russa
Lauk
Lavarra
Lax
Lebech
Lechner
Le Foll
Lefrançois
Lehideux
Lehne
Lehtinen
Leichtfried
Leinen
Le Rachinel
Lévai
Lewandowski
Liberadzki
Libicki
Lichtenberger
Lienemann
Liotard
Lipietz
Losco
Louis
Lucas
Ludford
Lulling
Lundgren
Lyubcheva
Maaten
McAvan
McCarthy
McGuinness
McMillan-Scott
Madeira
Maldeikis
Manders
Mănescu
Maňka
Thomas Mann
Marinescu
Markov
Marques
Martens
David Martin
Hans-Peter Martin
Martinez
Martínez Martínez
Masiel
Masip Hidalgo
Maštálka
Mathieu
Matsakis
Matsis
Matsouka
Mauro
Mavrommatis
Mayer
Medina Ortega
Méndez de Vigo
Menéndez del Valle
Meyer Pleite
Miguélez Ramos
Mikko
Mikolášik
Millán Mon
Mitchell
Mladenov
Mölzer
Mohácsi
Moreno Sánchez
Morgantini
Morillon
Morin
Mote
Mulder
Musacchio
Muscardini
Myller
Napoletano
Nassauer
Nattrass
Nechifor
Newton Dunn
Neyts-Uyttebroeck
Nicholson
Niculescu
Niebler
van Nistelrooij
Novak
Obiols i Germà
Öger
Olbrycht
Ó Neachtain
Onesta
Onyszkiewicz
Oomen-Ruijten
Oprea
Ortuondo Larrea
Őry
Ouzký
Oviir
Paasilinna
Pack
Pahor
Paleckis
Panayotopoulos-Cassiotou
Panayotov
Panzeri
Papadimoulis
Paparizov
Papastamkos
Parish
Paşcu
Peillon
Pęk
Alojz Peterle
Petre
Pflüger
Piecyk
Pieper
Pīks
Pinheiro
Pinior
Piotrowski
Pirker
Piskorski
Pistelli
Pittella
Pleguezuelos Aguilar
Pleštinská
Plumb
Podestà
Podimata
Podkański
Pöttering
Pohjamo
Polfer
Pomés Ruiz
Mihaela Popa
Nicolae Vlad Popa
Posdorf
Posselt
Prets
Pribetich
Vittorio Prodi
Protasiewicz
Purvis
Queiró
Rack
Radwan
Raeva
Ransdorf
Rasmussen
Remek
Resetarits
Reul
Ribeiro e Castro
Riera Madurell
Ries
Riis-Jørgensen
Rivera
Rizzo
Rocard
Rogalski
Roithová
Romagnoli
Romeva i Rueda
Rosati
Roszkowski
Roth-Behrendt
Rouček
Roure
Rovsing
Rübig
Rühle
Rutowicz
Ryan
Sacconi
Saïfi
Sakalas
Saks
Salafranca Sánchez-Neyra
Salinas García
Sánchez Presedo
dos Santos
Sartori
Saryusz-Wolski
Savi
Sbarbati
Schaldemose
Scheele
Schierhuber
Schinas
Schlyter
Frithjof Schmidt
Olle Schmidt
Schmitt
Schnellhardt
Schöpflin
Jürgen Schröder
Schroedter
Schulz
Schuth
Schwab
Seeber
Segelström
Seppänen
Severin
Siekierski
Silva Peneda
Simpson
Sinnott
Siwiec
Skinner
Škottová
Smith
Sógor
Sommer
Søndergaard
Sonik
Sornosa Martínez
Sousa Pinto
Speroni
Staes
Staniszewska
Starkevičiūtė
Šťastný
Stauner
Stavreva
Sterckx
Stevenson
Stihler
Stockmann
Stolojan
Stoyanov
Strejček
Strož
Stubb
Sudre
Sumberg
Surján
Susta
Svensson
Swoboda
Szájer
Szejna
Szent-Iványi
Szymański
Tabajdi
Tajani
Takkula
Tarand
Tatarella
Thomsen
Thyssen
Ţicău
Titley
Toia
Tőkés
Tomaszewska
Tomczak
Toubon
Toussas
Trakatellis
Trautmann
Triantaphyllides
Turmes
Tzampazi
Uca
Ulmer
Urutchev
Vaidere
Vakalis
Vălean
Vanhecke
Van Hecke
Van Lancker
Van Orden
Varela Suanzes-Carpegna
Varvitsiotis
Vatanen
Vaugrenard
Ventre
Veraldi
Vergnaud
Vernola
Vidal-Quadras
Vigenin
de Villiers
Virrankoski
Visser
Vlasák
Wagenknecht
Wallis
Walter
Watson
Manfred Weber
Renate Weber
Weiler
Weisgerber
Westlund
Whittaker
Wieland
Wiersma
Wijkman
Willmott
Iuliu Winkler
Wise
von Wogau
Bernard Wojciechowski
Janusz Wojciechowski
Wortmann-Kool
Wurtz
Yañez-Barnuevo García
Záborská
Zahradil
Zaleski
Zapałowski
Zappalà
Zatloukal
Ždanoka
Zdravkova
Železný
Zieleniec
Zīle
Zimmer
Zlotea
Zvěřina
Zwiefka
-//EP//TEXT TA 20080424 ITEMS DOC XML V0//SV
Sanktioner till skydd för miljön
Miljö
2008-05-21 - 16:02
För att garantera att EU:s miljölagstiftning efterlevs, så blir det möjligt att utfärda straffrättsliga påföljder för miljöbrott.
Det är innebörden i en kompromiss som träffats mellan Europaparlamentet och rådet.
Kompromissen godkändes i plenum idag.
Syftet är ett effektivare miljöskydd och alla medlemsstater är överens om att ett antal handlingar som orsakar miljöskador skall vara kriminellt.
Efter att lagstiftningen träder i kraft blir de nationella regeringarna skyldiga att införa "effektiva, proportionerliga och avskräckande" straffrättsliga påföljder.
Europaparlamentet är också överens med rådet att direktivet endast ska omfatta brott mot gemenskapslagstiftningen om miljöskydd, enligt bilagan i betänkandet.
Svenska inlägg i debatten
Jens Holm (GUE/NGL) ansåg att straffrätten inte ska harmoniseras.
– Risken med harmoniseringslagstiftning är alltid att progressiva länder blir tvungna att sänka nivån på sin lagstiftning, menade Holm.
– Självklart ska EU verka för att medlemsstaterna ska bli bättre på att arbeta med miljölagstiftning.
Debatt: 19.5.2008
20080520IPR29449 Antagna texter (provisorisk utgåva)
SV
1
LINK
/activities/plenary/ta/calendar.do?language=SV
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//TEXT TA 20080522 ITEMS DOC XML V0//SV
Hög standard på livsmedelshygien
Livsmedelssäkerhet
2008-06-05 - 15:48
Det anser Europaparlamentet i ett betänkande som antogs idag.
Med rösterna 556 för, 67 emot och 19 nedlagda röster antog Europaparlamentet ett betänkande om livsmedelshygien av Horst SCHNELLHARDT (EPP-ED, DE).
Förslaget är en del av kommissionens åtgärdsprogram för minskning av de administrativa bördorna.
Förslaget ändrar den tidigare förordningen om livsmedelshygien från 2004.
Kommissionen föreslår att små livsmedelsföretag undantas från det så kallade HACCP-förfarandet.
Det är ett system för riskanalys och står för Hazard Analysis and Critical Control Point.
Undantaget ska gälla för mikroföretag som huvudsakligen säljer mat direkt till slutkund.
HACCP-förfarandet är ett arbetssätt för att ta reda på, bedöma och kontrollera alla faror i produktionen.
Farorna är ett hot mot livsmedelssäkerheten.
Utifrån flödesscheman över tillverkningsprocesserna sammanställer man alla faror som kan finnas.
Det kan vara mikrobiologiska, kemiska, allergena och fysikaliska faror.
Föredragande: Horst SCHNELLHARDT (EPP-ED,DE)
Debatt och omröstning: 5.6.2008
20080604IPR30762
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
Dag för dag: plenarsammanträdet i Bryssel 4-5 juni
Institutioner
2008-06-09 - 14:21
Ledamöterna röstade för ett betänkande som kräver åtgärder mot olagligt fiske och debatterade hur tvångsprostitution kan förhindras.
På dagordningen var dessutom EU:s säkerhets- och försvarspolitik som diskuterades med EU:s höge representant för utrikesfrågor Javier Solana.
Via länkarna nedan kan du läsa sammanfattningar, dag för dag, av frågorna som behandlades på minisessionen.
Nästa plenarsammanträde inleds den 16 juni i Strasbourg
20080605FCS30922
Onsdag i plenum: EU-USA, säkerhet och försvar
Javier Solana debatterar EU:s utrikespolitik med ledamöterna Inför toppmötet mellan EU-USA i Slovenien den 9-10 juni gav ledamöterna sina synpunkter på hur dialogen med Washington kan förbättras.
Ledamöterna debatterade också EU:s gemensamma utrikespolitik samt förvars- och säkerhetspolitik.
På dagordningen var också en muntlig fråga om kampen mot människohandel och tvångsprostitution.
Och ledamöterna diskuterade även ett initiativ mot tjuvfiske.
Årets gröna vecka var i fokus då talmannen Hans-Gert Pöttering öppnade plenarsammanträdet i Bryssel den 4–5 juni.
Han påminde om Europaparlamentets mål att minska koldioxidutsläppen från den egna verksamheten med trettio procent fram till 2020.
I år kommer toppmötet att fokusera på det bilaterala transatlantiska partnerskapet, aktuella globala utmaningar och säkerhetsfrågor.
Europaparlamentet debatterade innehållet i en resolution (omröstning torsdag) med deras prioriteringar inför mötet.
Även Cem Özdemir (De Gröna, Tyskland) betonade behovet av att stärka den parlamentariska dimensionen, och sade att det innebär att involvera den amerikanska kongressen och Europaparlamentet.
Europaparlamentet höll också en debatt om den gemensamma utrikespolitiken samt förvars- och säkerhetspolitiken.
Två betänkanden från utskottet för utrikesfrågor debatterades: Det ena om rådets årliga rapport om den gemensamma utrikes- och säkerhetspolitiken (GUSP) för 2006, av Jacek Saryusz-Wolski (EPP-ED, Polen), och det andra om genomförandet av europeiska säkerhetsstrategin (ESS) och den europeiska säkerhets- och försvarspolitiken (ESFP), av Helmut Kuhne (PSE, Tyskland).
Utvecklingen på västra Balkan och behovet att stärka den europeiska grannskapspolitiken är exempel på några av de frågor som lyftes fram i debatten.
Flera talare underströk dessutom förbättringarna som Lissabonfördraget kommer att föra med sig för EU på utrikesområdet.
Javier Solana, EU:s höge representant för utrikes- och säkerhetspolitiken, deltog i debatten och sade:
Den första prioriteten för oss alla är att fördraget ratificeras.
Solana instämde med Sayusz-Wolski och Kuhne att ny områden måste tas i beaktande, exempelvis klimatförändringens påverkan på internationell säkerhet, energisäkerhet, olaglig invandring och informationssäkerhet.
Toppmötet mellan EU och USA den 9–10 juni i Slovenien Toppmötet EU-USA Finansiella tjänster utan gränser?
Större parlamentarisk kontroll av utrikespolitiken Debatt om tvångsprostitution, människohandel och sexuellt utnyttjande Ledamöterna debatterar initiativ mot tjuvfiske EU-USA toppmötet (rådet och kommissionen) EU-USA toppmötet (politiska grupperna)
Torsdag i plenum: en union för Medelhavsområdet
Debatt om Medelhavsunionen Fred, säkerhet och välstånd för Medelhavsområdets invånare var i fokus när ledamöterna på torsdagen debatterade planen om en uppgradering av Barcelonaprocessen och skapandet av en union, för att stärka relationerna mellan länderna kring Medelhavet.
Frankrikes president Nicholas Sarkozy har varit pådrivande i frågan som troligen kommer att prioriteras när Frankrike tar över EU-ordförandeskapet i juli.
I den resolution om Medelhavsunionen som antogs på torsdagen understryker Europaparlamentet att samarbetets sekretariat ska fokusera på regionala projekt.
Ledamöterna nämner solenergiprojekt, motorvägsprojekt och projekt för att stoppa utsläpp i Medelhavet som viktiga regionala projekt för den nya unionen.
"Vi behöver inte nya institutioner och mer byråkrati", sade Martin Schulz (PSE, Tyskland).
Vito Bonsignore (Gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater, Italien) välkomnade den franske presidentens initiativ och sade att det är "värt en applåd".
Han betonade vikten av multilaterala projekt och sade att det behövs ett frihandelsområde senast 2010.
Utmaningar
Samarbetet står också inför utmaningar.
Martin Schulz (Socialdemokratiska gruppen, Tyskland) sade att "social stabilitet är en nödvändig förutsättning för fred".
Regionens uteblivna välstånd och den svåra situationen invandrare möter i Europa togs upp av Francis Wurtz (Gruppen Europeiska enade vänstern/Nordisk grön vänster, Frankrike).
Behovet av mekanismer för garanti av de mänskliga rättigheterna betonades av Hélène Flautre (De Gröna, Frankrike) som också talade om kärnenergisäkerhet i Medelhavsområdet.
Se länkarna nedan för omröstningsresultat och mer information om frågorna på plenarsammanträdets dagordning, den 4-5 juni.
SV
1
PHOTO
20080605PHT31007.jpg
SV
2
PHOTO
20080603PHT30732.jpg
SV
3
LINK
SV
6
LINK
//news/expert/briefing_page/29027-156-06-23-20080516BRI29012-04-06-2008-2008/default_p001c001_sv.htm
SV
7
PHOTO
-//EP//TEXT IM-PRESS 20080604IPR30761 0 NOT XML V0//SV
-//EP//TEXT MOTION P6-RC-2008-0281 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20070314STO04222 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 FCS DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 FCS DOC XML V0//EN
NÄRVAROLISTA
Följande skrev på:
Adamou
Agnoletto
Aita
Albertini
Allister
Alvaro
Andersson
Andrejevs
Andrikienė
Angelakas Emmanouil
Angelilli
Antinucci Rapisardo
Antoniozzi
Arnaoutakis
Ashworth
Assis
Atkins
Attard-Montalto
Attwooll
Aubert
Audy
Auken
Ayala Sender
Aylward
Ayuso
Baco
Badia i Cutchet
Baeva Mariela Velichkova
Barón Crespo
Barsi-Pataky
Basile Domenico Antonio
Batten
Battilocchio
Batzeli
Bauer
Beaupuy
Beazley
Becsey
Beer
Belet
Belohorská
Bennahmias
Beňová
Berend
Berès
Berlato
Berlinguer
Berman
Bielan
Binev Slavi
Birutis
Blokland
Bloom
Bobošíková
Böge
Bösch
Bono
Bonsignore
Borghezio
Borrell Fontelles
Boştinaru Victor
Botopoulos Costas
Boursier Catherine
Bourzai
Bova Giuseppe
Bowis
Bowles
Bozkurt
Myller
Braghetto
Brejc
Brepoels
Breyer
Březina
Brie
Budreikaitė
van Buitenen
Buitenweg
Bullmann
Bulzesc Nicodim
van den Burg
Burke Colm
Bushill-Matthews
Busk
Buşoi
Philippe Busquin
Busuttil
Buzek
Callanan
Camre
Capoulas Santos
Cappato
Carlotti
Carlshamre
Carnero González
Carollo
Casa
Casaca
Cashman
Casini
Caspary
Castex
del Castillo Vera
Catania
Cavada
Cederschiöld
Cercas
Chatzimarkakis
Chichester
Chiesa
Chmielewski
Christensen
Chruszcz
Chukolov Desislav
Philip Claeys
Clark
Cocilovo
Coelho
Cohn-Bendit
Corbett
Corbey
Corda Giovanna
Corlăţean
Cornillet
Cottigny
Coûteaux
Cramer
Cremers Jan
Corina Creţu
Gabriela Creţu
Crowley
Csibi Magor Imre
Marek Aleksander Czarnecki
Ryszard Czarnecki
Dahl Hanne
Dăianu Daniel
Daul
David Dragoş Florin
Davies
De Blasio
de Brún
Degutis
De Keyser
Demetriou
Breyer
De Rossa
De Sarnez
Descamps
Deß
De Veyrac
De Vits
Díaz de Mera García Consuegra
Dičkutė
Didžiokas
Dillen
Dimitrakopoulos
Dobolyi
Dombrovskis
Donnici
Doorn
Douay
Dover
Doyle
Drčar Murko
Droutsas Konstantinos
Duchoň
Dührkop Dührkop
Duff
Duka-Zólyomi
Dumitriu Constantin
Ehler
Ek
El Khadraoui
Elles
Esteves
Estrela
Ettl
Väyrynen
Jonathan Evans
Robert Evans
Färm
Fajmon
Falbr
Farage
Fatuzzo
Fava
Fazakas
Ferber
Fernandes
Fernández Martín
Ferrari Francesco
Panayotov
Elisa Ferreira
Figueiredo
Filip Petru
Fiore Roberto
Fjellner
Flasarová
Flautre
Florenz
Foglietta
Foltyn-Kubicka
Fontaine
Ford
Fouré Brigitte
Fourtou
Fraga Estévez
Fraile Cantón Juan
França Armando
Freitas
Friedrich
Gacek Urszula
Gahler
Gál
Gaľa
Galeote
Garcés Ramón Vicente Miguel
García-Margallo y Marfil
García Pérez
Gargani
Garriga Polledo
Gaubert
Gauzès
Gawronski
Gebhardt
Gentvilas
Georgiou Georgios
Geremek
Geringer de Oedenberg
Gewalt
Gibault
Gierek
Giertych
Gill
Gklavakis
Glattfelder
Désir
Konrad
Goepel
Golik
Gollnisch
Gomes
Gomolka
Gottardi
Goudin
Grabowska
Grabowski
Graça Moura
Graefe zu Baringdorf
Gräßle
de Grandes Pascual
Grau i Segú Martí
Grech
Griesbeck
Gröner
de Groen-Kouwenhoven
Groote
Grosch
Grossetête
Gruber
Guardans Cambó
Guellec
Guerreiro
Guidoni
Gurmai
Gutiérrez-Cortines
Guy-Quint
Gyürk
Hänsch
Hall
Hammerstein
Hamon
Handzlik
Harangozó
Harbour
Harkin
Harms
Hasse Ferreira
Hassi
Haug
Heaton-Harris
Hedh
Hegyi
Helmer
Henin
Hennicot-Schoepges
Hennis-Plasschaert
Herczog
Herranz García
Herrero-Tejedor
Hieronymi
Higgins
Hökmark
Holm
Honeyball
Hoppenstedt
Horáček
Howitt
Hudacký
Hudghton
Hughes
Hutchinson
Husmenova
Iacob-Ridzi
Ibrisagic
in 't Veld
Iotova Iliana Malinova
Irujo Amezaga Mikel
Isler Béguin
Itälä
Jackson
Jacobs Lily
Jäätteenmäki
Jałowiecki
Janowski
Járóka
Jarzembowski
Jeggle
Jeleva Rumiana
Jensen
Jöns
Jørgensen
Jonckheer
Jordan Cizelj
Jouye de Grandmaison Madeleine
Juknevičienė
Kacin
Kaczmarek
Kallenbach
Kamall
Karas
Karim
Kasoulides
Kaufmann
Kauppi
Kazak Metin
Tunne Kelam
Kindermann
Kinnock
Kirilov
Kirkhope
Klamt
Klaß
Klinz
Knapman
Koch
Koch-Mehrin
Kohlíček
Konrad
Koppa Maria Eleni
Korhola
Kósáné Kovács
Koterec
Kozlík
Krahmer
Krasts
Tajani
Krehl
Kreissl-Dörfler
Kristovskis
Krupa
Kuc
Kuhne
Kułakowski
Kušķis
Kusstatscher
Kuźmiuk
Lagendijk
Laignel
Lamassoure
Lambert
Lambrinidis
Landsbergis
Lang
De Lange
Langen
Laperrouze
La Russa
Lavarra
Lax
Lebech Johannes
Lechner
Le Foll
Lefrançois Roselyne
Lehideux
Lehne
Lehtinen
Leichtfried
Leinen
Jean-Marie Le Pen
Marine Le Pen
Le Rachinel
Lévai
Lewandowski
Liberadzki
Libicki
Lichtenberger
Lienemann
Liese
Liotard
Lipietz
Locatelli
López-Istúriz White
Losco
Louis
Lucas
Ludford
Lulling
Lundgren
Luque Aguilar Florencio
Lynne
Lyubcheva
McAvan
McCarthy
McGuinness
McMillan-Scott
Madeira
Maldeikis
Manders
Mănescu Ramona Nicole
Maňka
Erika Mann
Thomas Mann
Marinescu
Marini Catiuscia
Markov
Marques
Martens
David Martin
Hans-Peter Martin
Martinez
Martínez Martínez
Masiel
Maštálka
Mathieu
Matsakis
Matsouka
Mauro
Mavrommatis
Mayer
Mayor Oreja
Medina Ortega
Meijer
Méndez de Vigo
Menéndez del Valle
Meyer Pleite
Miguélez Ramos
Mikko
Mikolášik
Millán Mon
Mitchell
Mladenov Nickolay
Mölzer
Mohácsi
Moraes
Moreno Sánchez
Morgan
Morgantini
Morillon
Mote
Mulder
Musacchio
Muscardini
Grosch
Myller
Napoletano
Nassauer
Nattrass
Navarro
Nechifor Cătălin-Ioan
Neris Catherine
Newton Dunn
Nicholson
Nicholson of Winterbourne
Niculescu Rareş-Lucian
Niebler
van Nistelrooij
Novak
Obiols i Germà
Öger
Özdemir
Olbrycht
Ó Neachtain
Onesta
Onyszkiewicz
Ford
Ortuondo Larrea
Paasilinna
Pack
Pafilis
Pahor
Paleckis
Panayotopoulos-Cassiotou
Panayotov Vladko Todorov
Pannella
Panzeri
Papadimoulis
Paparizov
Papastamkos
Parish
Paşcu
Patriciello
Patrie
Peillon
Pęk
Alojz Peterle
Petre
Pflüger
Piecyk
Pieper
Pietikäinen Sirpa
Pīks
Pinheiro
Pinior
Piotrowski
Pirilli
Piskorski
Pittella
Pleguezuelos Aguilar
Pleštinská
Plumb
Podestà
Podimata Anni
Podkański
Pöttering
Pohjamo
Poignant
Polfer
Pomés Ruiz
Popa Mihaela
Popa
Portas
Posdorf
Posselt
Prets
Pribetich Pierre
Vittorio Prodi
Protasiewicz
Purvis
Queiró
Rack
Radwan
Raeva Bilyana Ilieva
Ransdorf
Rapkay
Remek
Reul
Mote
Riera Madurell
Ries
Riis-Jørgensen
Rivera
Rizzo
Robusti Giovanni
Rocard
Rogalski
Roithová
Romagnoli
Rosati
Roszkowski
Roth-Behrendt
Rothe
Rouček
Roure
Rovsing
Rübig
Rühle
Rutowicz
Ryan
Sacconi
Saïfi
Sakalas
Saks
Salafranca Sánchez-Neyra
Salinas García
Sánchez Presedo
dos Santos
Sanzarello Sebastiano
Sanz Palacio Salvador Domingo
Sartori
Saryusz-Wolski
Savary
Savi
Schaldemose
Schapira
Schenardi
Schierhuber
Schinas Margaritis
Schlyter
Frithjof Schmidt
Olle Schmidt
Schmitt
Schnellhardt
Schöpflin
Jürgen Schröder
Schroedter
Schuth
Schwab
Seeber
Segelström
Seppänen
Severin
Siekierski
Silva Peneda
Simpson
Sinnott
Siwiec
Skinner
Škottová
Smith
Sógor Csaba
Sommer
Søndergaard
Sonik
Sornosa Martínez
Sousa Pinto
Spautz
Speroni
Obiols i Germà
Staniszewska
Starkevičiūtė
Šťastný
Stauner
Stavreva Petya
Stevenson
Stihler
Stolojan Theodor Dumitru
Stoyanov
Strejček
Strož
Sturdy
Sudre
Sumberg
Surján
Susta
Svensson
Swoboda
Szájer
Szejna
Szent-Iványi
Szymański
Tabajdi
Takkula
Tannock
Tarand
Tatarella
Thomsen
Thyssen
Ţicău
Titford
Titley
Toia
Tőkés László
Tomaszewska Ewa
Tomczak
Toubon
Toussas
Trakatellis
Trautmann
Triantaphyllides
Trüpel
Turmes
Tzampazi
Uca
Ulmer
Urutchev Vladimir
Vakalis
Vălean
Vanhecke
Van Hecke
Van Lancker
Bösch
Varela Suanzes-Carpegna
Varvitsiotis
Vatanen
Vaugrenard
Veneto
Ventre
Veraldi
Vergnaud
Vernola
McCarthy
Vigenin
Virrankoski
Visser Cornelis
Vlasák
Zdravkova
Voggenhuber
Wagenknecht
Wallis
Walter
Watson
Henri Weber
Manfred Weber
Weber Renate
Weiler
Weisgerber
Westlund
Whittaker
Wiersma
Wijkman
Willmott
Winkler Iuliu
Wise
Wohlin
Bernard Wojciechowski
Janusz Wojciechowski
Wortmann-Kool
Wurtz
Yañez-Barnuevo García
Záborská
Zahradil
Zaleski
Zanicchi Iva
Zapałowski
Zappalà
Zatloukal
Ždanoka
Zdravkova Dushana
Zieleniec
Zīle
Zimmer
Zvěřina
Zwiefka
Inte bara politik
Kultur
2008-08-18 - 09:00
Inte bara politik EU:s 27 medlemsstaters befolkning på nästan en halv miljard med sina särskilda traditioner, vanor och kulturer skapar en av de mest färgstarka bilder man kan föreställa sig: Folkets Europa.
På vår webbplats har vi flera gånger skrivit om olika traditioner, vad européerna gör på sin fritid, kultur och evenemang.
Läs några av artiklarna här om fotboll, påsk, alla hjärtans dag och Europas kulturhuvudstäder.
Vi frågade några ledamöter om deras synpunkter.
Påsktraditioner i Europa
20080707FCS33614
Vi frågade några ledamöter om deras synpunkter.
– Fans från hela världen samlades för att njuta av sin favoritsport.
Han uppmärksammar att namnet på mästerskapets officiella boll är "Europass", det syftar på spelarnas och fansens samarbete och gruppanda.
– Det är en metafor för vårt arbete i Europaparlamentet.
Vi "passar" argument mellan oss, utbyter åsikter och erfarenheter för att uppnå ett gemensamt "mål".
Jan Andersson berättar att han ska åka till Salzburg för att se Sverige, och Henrik Larsson som inledde sin karriär i just Högaborg, spela mot Grekland.
För Ramona Mănescu (Gruppen Alliansen liberaler och demokrater för Europa, Rumänien) är sport ett sätt att mötas och på så sätt förenas människor.
Sportens värderingar är universella, och de är emot uppdelningar.
En fotbollsmatch är inte en kamp utan en möjlighet att jämföra sig i en ärlig match.
I Europa är vi ibland tillsammans och i andra fall var för sig.
Och så måste det fortsätta att vara.
Syftet är att bjuda in ungdomar för att delta i en europeisk kampanj mot våld och rasism inom idrotten.
Ett ungdomsforum kommer att hållas 18-20 september i italienska Bologna.
Påsk runt om i Europa För många är påsken en tid då man ser fram mot grönskan, ljuset och våren.
Påsken är en stor religiös högtid, men den handlar också om icke religiösa traditioner.
Läs mer om hur påsken firas i olika delar av Europa.
Också för Bastiaan Belder (gruppen Självständighet/Demokrati, IND/DEM) från Nederländerna är påsken en familjehögtid.
Han firade den med sin fru, barn och barnbarn.
Han säger att påsken också har en viktig religiös innebörd och att den "är inte bara en ledig dag".
Vi hade påskliljor på bordet som dekoration och en påskkärring i fönstret."
Tjeckiska ledamoten Jana Hybášková (EPP-ED) berättar att man, under mycket tjoande, på annandag påskmorgonen "piskar" varandra med vide i hennes familj.
Att måla påskägg är ytterligare en vanlig tradition."
Han berättar också att folk ger varandra videkvistar och att man frågar barnen "om solen dansar".
Nytt liv och ett nytt år
Hammerstein ska också fira den judiska påsken, som i år firas mellan den 20-26 april.
Och då kommer han särskilt att tänka på befrielsen av folk som lever under förtryck, som tibetanerna.
Tyska ledamoten Feleknas Uca (Gruppen Europeiska enade vänstern/Nordisk grön vänster) var i Turkiet för att fira newroz, det kurdiska nyåret som infaller på vårdagjämningen den 21 mars.
Vi lämnar ofta över det till poeter och musiker, men sällan till politiker.
Så vad passar bättre än att låta politikerna komma till tals idag på Alla hjärtans dag.
Vi tog mod till oss och talade med några ledamöter om kärlek.
Vad skulle en europeisk stadga om kärlek omfatta?
– Inga åldersbegränsningar eller sanktioner.
Den måste grundas på övertygelse och förtroende.
Katalin Lévai (PSE, Ungern) betonar vikten av ömsesidig förståelse och respekt.
Annars försvinner lusten.
– Kärlek misslyckas aldrig.
Om vi lyckas att genomföra den här idén, då skulle världen bli mycket trevligare.
Europeiska unionen är ett område där tankar, känslor, attityder uppmuntras att öppet blomstra.
Jag tror att den här stadgan redan existerar.
Vi har den inom oss, säger Roberta Alma Anastase (EPP-ED, Rumänien).
Den som spelar en roll misslyckas till sist, råder Katalin Lévai .
Astrid Lulling (EPP-ED, Luxemburg) menar att det inte går att organisera eller planera romantik och kärlek.
– Det finns inget värre gift för kärleken än leda.
– Ju mer du älskar desto mer utsätter du dig själv för lidande.
- Njut fullt ut av romantiken.
Men ta inga avgörande beslut innan du vet om det är kärlek eller något annat, säger Henrik Lax.
Men det viktigaste är att vara säker på att personen du älskar är där för dig, tycker Roberta Alma Anastase .
För Katalin Lévai är en bok är den mest värdefulla gåvan, men gärna ackompanjerat av blommor.
Medan Genowefa Grabowska skulle vilja få en röd ros.
Ge av tid, fantasi och sitt hjärta.
Har du planerat något speciellt för Alla hjärtans dag?
– Alla hjärtans dag blev på modet när jag redan var över fyrtio.
Men man kan ju alltid drömma, varför inte hoppas att en god vän tar initiativet till en fin överraskning, säger Astrid Lulling .
- Nej, jag kommer att vara i Kiev, Ukraina, långt från min hustru som jag träffade för fyrtiotre år sedan.
Teater- och filmvisningar, konserter, utställningar och andra kulturevenemang förväntas att locka besökare till de två städerna och placera dem på Europas kulturkarta.
EU:s kulturministrar i ministerrådet utser en eller flera europeiska kulturhuvudstäder.
Och Europaparlamentet deltar i urvalsprocessen.
Liverpool: Mer än Beatles
Liverpool är internationellt kanske mest berömd som Beatles hemstad och för fotbollslagen Everton och Liverpool.
Det är också en stor hamnstad, vars hamnområde 2004 upptogs på Unesco världsarvslista, och en mångkulturell mötesplats.
Uppskattningsvis talas ungefär 60 olika språk bland staden över 440 000 invånare.
Liverpool inledde året med en konsert: Liverpoolmusikalen med ex-beatlen Ringo Starr och Royal Liverpool Philharmonic Orchestra.
Men också teater, dans, bok- och poesifestivaler och fotoutställningar är på programmet.
Stavanger: "Open port"
Stavanger är liksom Liverpool en hamnstad.
Men är mer känd för sina ljusa sommarnätter och det vackra fjordlandskapet än fotboll och musik.
Stavangers gamla del består till stor del av vita trähus.
Oljeindustrin har bidragit till att göra Stavanger till en välmående stad.
Arbetslösheten är 1 procent.
Stavanger program som kulturhuvudstad är "Open port", och öppenhet och yttrandefrihet är viktiga delar.
Vissa ateljéer uppmuntrar exempelvis besökare att skapa sina egna alster, och internationella konstnärer kommer till Stavanger för att arbeta med lokala konstnärer.
Arkitektur, litteratur, musik och bildkonst är också del av evenemangsprogrammet.
SV
1
PHOTO
20080715PHT34210.jpg
SV
2
PHOTO
20080605PHT31009.jpg
SV
3
LINK
http://www.euro2008.uefa.com/
SV
4
LINK
/activities/committees/homeCom.do?body=CULT&language=SV
SV
5
LINK
/members.do?language=SV
SV
6
PHOTO
20080327PHT25026.jpg
SV
7
LINK
SV
9
PHOTO
20080211PHT20849.jpg
SV
10
LINK
-//EP//TEXT IM-PRESS 20070125STO02408 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 FEA DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 FEA DOC XML V0//EN
Föredragningslista
Onsdagen den 9 juli 2008
9:00 - 11:50 [LAGSTIFTNINGSDEBATT] Betänkande Olle Schmidt A6-0241/2008
ECB:s årsrapport för 2007
om ECB:s årsrapport för 2007
[ 2008/2107(INI) ]
Europeiska centralbankens ordförande Jean-Claude Trichet deltar i debatten
Gemensam debatt
Sociala trygghetssystem
Betänkande Jean Lambert A6-0251/2008
Samordning av socialförsäkringssystemen
om förslaget till Europaparlamentets och rådets förordning om tillämpningsbestämmelser till förordning (EG) nr 883/2004 om samordning av de sociala trygghetssystemen
[ KOM(2006)0016 - C6-0037/2006 - 2006/0006(COD) ]
Utskottet för sysselsättning och sociala frågor
Betänkande Emine Bozkurt A6-0229/2008
Samordning av socialförsäkringssystemen: bilaga XI
om förslaget till Europaparlamentets och rådets förordning om ändring av förordning (EG) nr 883/2004 om samordning av de sociala trygghetssystemen och om fastställande av innehållet i bilaga XI
[ KOM(2006)0007 - C6-0029/2006 - 2006/0008(COD) ]
Utskottet för sysselsättning och sociala frågor
Betänkande Jean Lambert A6-0209/2008
Utvidgning av bestämmelserna i förordning (EG) nr 883/2004 till att gälla de tredjelandsmedborgare som inte omfattas av dessa bestämmelser
om förslaget till rådets förordning om utvidgning av bestämmelserna i förordning (EG) nr 883/2004 och förordning (EG) nr […] till att gälla de medborgare i tredje land som enbart på grund av sitt medborgarskap inte omfattas av dessa bestämmelser
[ KOM(2007)0439 - C6-0289/2007 - 2007/0152(CNS) ]
Utskottet för sysselsättning och sociala frågor
Slut på den gemensamma debatten
12:00 - 13:00 Omröstning om begäran om brådskande förfarande ( artikel 134 i arbetsordningen)
Eventuellt: Omröstning
Resolutionsförslag B6-0336/2008
Årliga handlingsprogram för Brasilien och Argentina (2008)
om förslagen till kommissionens beslut om inrättande av årliga handlingsprogram för Brasilien 2008 och Argentina 2008
(CMTD 2008-0263) – D000422-01, CMTD-2008-0263 – D000421-01)
Utskottet för utveckling
Artikel 81 i arbetsordningen
Betänkande Alexander Graf Lambsdorff A6-0265/2008
Europaparlamentets rekommendationer till rådet om EU:s prioriteringar inför den 63:e sessionen i FN:s generalförsamling
om ett förslag till Europaparlamentets rekommendation till rådet om EU:s prioriteringar för FN:s generalförsamlings 63:e session
[ 2008/2111(INI) ]
Utskottet för utrikesfrågor
Artikel 90 i arbetsordningen
Betänkande Christoph Konrad A6-0240/2008
Program för modernisering av den europeiska företags- och handelsstatistiken (Meets-programmet)
om förslaget till Europaparlamentets och rådets beslut om ett program för modernisering av den europeiska företags- och handelsstatistiken (Meets-programmet)
[ KOM(2007)0433 - C6-0234/2007 - 2007/0156(COD) ]
Utskottet för ekonomi och valutafrågor
Betänkande Johannes Blokland A6-0244/2008
Batterier och ackumulatorer och förbrukade batterier och ackumulatorer
[ KOM(2008)0211 - C6-0165/2008 - 2008/0081(COD) ]
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Betänkande Miroslav Ouzký A6-0135/2008
Begränsning av användning och utsläppande på marknaden av vissa farliga ämnen och preparat (beredningar)
om förslaget till Europaparlamentets och rådets beslut om ändring av rådets direktiv 76/769/EEG om begränsning av användning och utsläppande på marknaden av vissa farliga ämnen och preparat (beredningar) 2 (2 metoxietoxi)etanol, 2-(2-butoxietoxi)etanol, metylendifenyldiisocyanat, cyklohexan och ammoniumnitrat
[ KOM(2007)0559 - C6-0327/2007 - 2007/0200(COD) ]
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Betänkande Diana Wallis A6-0224/2008
Den nationelle domarens roll i det europeiska rättssystemet
om den nationelle domarens roll i det europeiska rättssystemet
[ 2007/2027(INI) ]
Utskottet för rättsliga frågor
15:00 - 18:30 [DEBATT OM AKTUELLA ÄMNEN] Uttalanden av rådet och kommissionen
Situationen i Kina efter jordbävningen och inför de olympiska spelen
Betänkande Elmar Brok A6-0266/2008
Kommissionens strategidokument för utvidgningen
om kommissionens strategidokument för utvidgningen
[ 2007/2271(INI) ]
Utskottet för utrikesfrågor
Muntliga frågor
Palestinska fångar i israeliska fängelser
O-0040/2008 Luisa Morgantini Hélène Flautre Richard Howitt Thijs Berman Kyriacos Triantaphyllides Proinsias De Rossa Pasqualina Napoletano Margrete Auken Jean Lambert Marios Matsakis David Hammerstein Jill Evans Jamila Madeira Eugenijus Maldeikis Philippe Morillon Chris Davies Vincenzo Aita Françoise Castex Caroline Lucas Antonio Masip Hidalgo Alyn Smith Ana Maria Gomes Karin Scheele Alain Hutchinson Marco Cappato John Bowis Giovanni Berlinguer Giusto Catania Roberto Musacchio Vittorio Agnoletto Frieda Brepoels Mauro Zani Umberto Guidoni Luigi Cocilovo Linda McAvan Alessandro Battilocchio Baroness Nicholson of Winterbourne Francis Wurtz Tokia Saïfi Edward McMillan-Scott Emilio Menéndez del Valle Ioannis Kasoulides Véronique De Keyser Kader Arif Béatrice Patrie Rodi Kratsa-Tsagaropoulou B6-0166/2008 rådet Palestinska fångar i israeliska fängelser
O-0041/2008 Luisa Morgantini Hélène Flautre Richard Howitt Thijs Berman Kyriacos Triantaphyllides Proinsias De Rossa Pasqualina Napoletano Margrete Auken Jean Lambert Marios Matsakis David Hammerstein Jill Evans Jamila Madeira Eugenijus Maldeikis Philippe Morillon Chris Davies Vincenzo Aita Françoise Castex Caroline Lucas Antonio Masip Hidalgo Alyn Smith Ana Maria Gomes Karin Scheele Alain Hutchinson Marco Cappato John Bowis Giovanni Berlinguer Giusto Catania Roberto Musacchio Vittorio Agnoletto Frieda Brepoels Mauro Zani Umberto Guidoni Luigi Cocilovo Linda McAvan Alessandro Battilocchio Baroness Nicholson of Winterbourne Francis Wurtz Tokia Saïfi Edward McMillan-Scott Emilio Menéndez del Valle Ioannis Kasoulides Véronique De Keyser Kader Arif Béatrice Patrie Rodi Kratsa-Tsagaropoulou B6-0167/2008 kommissionen Palestinska fångar i israeliska fängelser
Situationen i Zimbabwe
18:30 - 20:00 Frågestund med frågor till kommissionen B6-0168/2008
21:00 - 24:00 Betänkande Karl von Wogau A6-0250/2008
Världsrymden och säkerheten
om världsrymden och säkerheten
[ 2008/2030(INI) ]
Utskottet för utrikesfrågor
Betänkande Carmen Fraga Estévez A6-0278/2008
Fiskemöjligheter och den ekonomiska ersättning som föreskrivs i partnerskapsavtalet om fiske mellan EG och Mauretanien
om förslaget till rådets förordning om ingående av protokollet om fastställande för perioden 1 augusti 2008–31 juli 2012 av de fiskemöjligheter och den ekonomiska ersättning som föreskrivs i partnerskapsavtalet om fiske mellan Europeiska gemenskapen och Islamiska republiken Mauretanien
[ KOM(2008)0243 - C6-0199/2008 - 2008/0093(CNS) ]
Fiskeriutskottet
Betänkande Sarah Ludford A6-0459/2007
Gemensamma konsulära instruktioner: biometriska kännetecken och visumansökningar
om förslaget till Europaparlamentets och rådets förordning om ändring av de gemensamma konsulära anvisningarna angående viseringar till diplomatiska beskickningar och karriärkonsulat i samband med införandet av biometri samt bestämmelser om organiseringen av mottagandet och behandlingen av viseringsansökningar
[ KOM(2006)0269 - C6-0166/2006 - 2006/0088(COD) ]
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Eventuellt: Betänkande upptaget i enlighet med artikel 134 i arbetsordningen
Talartid ( artikel 142 i arbetsordningen)
9:00 - 11:50 [LAGSTIFTNINGSDEBATT] Kommissionen (inklusive repliker)
Föredragande (3 x 6')
Föredragande av yttrande
Talarlistor Ledamöter
PPE-DE
24
PSE
18
ALDE
10
UEN
5
Verts/ALE
5
GUE/NGL
5
IND/DEM
4
NI
4
"Catch the eye" (2 x 5')
15:00 - 18:30 [DEBATT OM AKTUELLA ÄMNEN] Rådet (inklusive repliker)
Kommissionen (inklusive repliker)
Föredragande
Föredragande av yttrande
Frågeställare
Talarlistor Ledamöter
PPE-DE
29
PSE
22
ALDE
12
UEN
6
Verts/ALE
6
GUE/NGL
6
IND/DEM
4
NI
5
"Catch the eye" (4 x 5')
21:00 - 24:00 Kommissionen (inklusive repliker)
Föredragande (3 x 6')
Föredragande av yttrande (3 x 1')
Talarlistor Ledamöter
PPE-DE
24
PSE
18
ALDE
10
UEN
5
Verts/ALE
5
GUE/NGL
5
IND/DEM
4
NI
4
"Catch the eye"
Tidsfrister
Betänkande Olle Schmidt A6-0241/2008
ECB:s årsrapport för 2007
Ändringsförslag
har löpt ut
Betänkande Jean Lambert A6-0251/2008
Samordning av socialförsäkringssystemen
Ändringsförslag
har löpt ut
Betänkande Emine Bozkurt A6-0229/2008
Samordning av socialförsäkringssystemen: bilaga XI
Ändringsförslag
har löpt ut
Betänkande Jean Lambert A6-0209/2008
Utvidgning av bestämmelserna i förordning (EG) nr 883/2004 till att gälla de tredjelandsmedborgare som inte omfattas av dessa bestämmelser
Ändringsförslag
har löpt ut
Resolutionsförslag B6-0336/2008
Årliga handlingsprogram för Brasilien och Argentina (2008)
Ändringsförslag
Måndagen den 7 juli, 19:00
Betänkande Christoph Konrad A6-0240/2008
Program för modernisering av den europeiska företags- och handelsstatistiken (Meets-programmet)
Ändringsförslag
Måndagen den 7 juli, 19:00
Begäran om särskild omröstning, delad omröstning eller omröstning med namnupprop
Tisdagen den 8 juli, 19:00
Betänkande Johannes Blokland A6-0244/2008
Batterier och ackumulatorer och förbrukade batterier och ackumulatorer
Ändringsförslag
Måndagen den 7 juli, 19:00
Begäran om särskild omröstning, delad omröstning eller omröstning med namnupprop
Tisdagen den 8 juli, 19:00
Betänkande Miroslav Ouzký A6-0135/2008
Begränsning av användning och utsläppande på marknaden av vissa farliga ämnen och preparat (beredningar)
Ändringsförslag
Måndagen den 7 juli, 19:00
Begäran om särskild omröstning, delad omröstning eller omröstning med namnupprop
Tisdagen den 8 juli, 19:00
Betänkande Diana Wallis A6-0224/2008
Den nationelle domarens roll i det europeiska rättssystemet
Ändringsförslag
Måndagen den 7 juli, 19:00
Begäran om särskild omröstning, delad omröstning eller omröstning med namnupprop
Tisdagen den 8 juli, 19:00
Uttalanden av rådet och kommissionen
Situationen i Kina efter jordbävningen och inför de olympiska spelen
Resolutionsförslag
har löpt ut
Ändringsförslag och gemensamma resolutionsförslag
Måndagen den 7 juli, 19:00
Betänkande Elmar Brok A6-0266/2008
Kommissionens strategidokument för utvidgningen
Ändringsförslag
har löpt ut
Muntliga frågor
Palestinska fångar i israeliska fängelser
O-0040/2008 Luisa Morgantini Hélène Flautre Richard Howitt Thijs Berman Kyriacos Triantaphyllides Proinsias De Rossa Pasqualina Napoletano Margrete Auken Jean Lambert Marios Matsakis David Hammerstein Jill Evans Jamila Madeira Eugenijus Maldeikis Philippe Morillon Chris Davies Vincenzo Aita Françoise Castex Caroline Lucas Antonio Masip Hidalgo Alyn Smith Ana Maria Gomes Karin Scheele Alain Hutchinson Marco Cappato John Bowis Giovanni Berlinguer Giusto Catania Roberto Musacchio Vittorio Agnoletto Frieda Brepoels Mauro Zani Umberto Guidoni Luigi Cocilovo Linda McAvan Alessandro Battilocchio Baroness Nicholson of Winterbourne Francis Wurtz Tokia Saïfi Edward McMillan-Scott Emilio Menéndez del Valle Ioannis Kasoulides Véronique De Keyser Kader Arif Béatrice Patrie Rodi Kratsa-Tsagaropoulou B6-0166/2008 rådet Palestinska fångar i israeliska fängelser
O-0041/2008 Luisa Morgantini Hélène Flautre Richard Howitt Thijs Berman Kyriacos Triantaphyllides Proinsias De Rossa Pasqualina Napoletano Margrete Auken Jean Lambert Marios Matsakis David Hammerstein Jill Evans Jamila Madeira Eugenijus Maldeikis Philippe Morillon Chris Davies Vincenzo Aita Françoise Castex Caroline Lucas Antonio Masip Hidalgo Alyn Smith Ana Maria Gomes Karin Scheele Alain Hutchinson Marco Cappato John Bowis Giovanni Berlinguer Giusto Catania Roberto Musacchio Vittorio Agnoletto Frieda Brepoels Mauro Zani Umberto Guidoni Luigi Cocilovo Linda McAvan Alessandro Battilocchio Baroness Nicholson of Winterbourne Francis Wurtz Tokia Saïfi Edward McMillan-Scott Emilio Menéndez del Valle Ioannis Kasoulides Véronique De Keyser Kader Arif Béatrice Patrie Rodi Kratsa-Tsagaropoulou B6-0167/2008 kommissionen Palestinska fångar i israeliska fängelser
Resolutionsförslag
Onsdagen den 27 augusti, 12:00
Ändringsförslag och gemensamma resolutionsförslag
Måndagen den 1 september, 19:00
Uttalanden av rådet och kommissionen
Situationen i Zimbabwe
Resolutionsförslag
Måndagen den 7 juli, 19:00
Ändringsförslag och gemensamma resolutionsförslag
Tisdagen den 8 juli, 17:00
Begäran om särskild omröstning, delad omröstning eller omröstning med namnupprop
Onsdagen den 9 juli, 17:00
Betänkande Karl von Wogau A6-0250/2008
Världsrymden och säkerheten
Ändringsförslag
har löpt ut
Betänkande Carmen Fraga Estévez A6-0278/2008
Fiskemöjligheter och den ekonomiska ersättning som föreskrivs i partnerskapsavtalet om fiske mellan EG och Mauretanien
Ändringsförslag
har löpt ut
Betänkande Sarah Ludford A6-0459/2007
Gemensamma konsulära instruktioner: biometriska kännetecken och visumansökningar
Ändringsförslag
Måndagen den 7 juli, 19:00
Begäran om särskild omröstning, delad omröstning eller omröstning med namnupprop
Onsdagen den 9 juli, 17:00
Särskild omröstning - delad omröstning - omröstning med namnupprop Texter som kommer att gå till omröstning tisdag
Fredagen den 4 juli, 12:00
Texter som kommer att gå till omröstning onsdag
Måndagen den 7 juli, 19:00
Texter som kommer att gå till omröstning torsdag
Tisdagen den 8 juli, 19:00
Resolutionsförslag om debatter om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer ( artikel 115 i arbetsordningen)
Torsdagen den 10 juli, 10:00
Utskottet för utveckling
DEVE(2008)0901_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Måndagen den 1 september 2008 kl. 19.00–20.30
Bryssel
Lokal: ASP 1 G 3
1.
Godkännande av föredragningslistan
I närvaro av rådet och kommissionen
2.
Meddelanden från ordföranden
3.
Budgeten för 2009: Avsnitt III – kommissionen
DEVE/6/58984
2008/2026(BUD)
Föredragande:
Maria Martens (PPE-DE)
Ansv. utsk.:
BUDG
Jutta Haug (PSE)
· Antagande av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 19 augusti 2008 kl. 12.00
4.
Övriga frågor
5.
ARBETSORDNING
16:e upplagan
Oktober 2008
Anmärkning
till
läsaren
:
I enlighet med parlamentets beslut om användningen av könsneutralt språk i sina handlingar har arbetsordningen anpassats för att ta hänsyn till de riktlinjer beträffande denna fråga som antogs av högnivågruppen för jämställdhet mellan kvinnor och män samt mångfald den 13 februari 2008 och som godkändes av presidiet den 19 maj 2008.
Tolkningar till arbetsordningen återges (i enlighet med artikel 201) i kursiv stil.
INNEHÅLL
AVDELNING
I
LEDAMÖTER, PARLAMENTETS ORGAN OCH POLITISKA GRUPPER
KAPITEL
1
EUROPAPARLAMENTETS LEDAMÖTER
Artikel
1
Europaparlamentet
Artikel
2
Obundet mandat
Artikel
3
Valprövning
Artikel
4
Mandatets varaktighet
Artikel
5
Immunitet och privilegier
Artikel
6
Upphävande av immunitet
Artikel
7
Immunitetsförfaranden
Artikel
8
Kostnadsersättning och andra ersättningar
Artikel
9
Ledamöternas ekonomiska intressen, ordningsregler och tillträde till parlamentet
Artikel
10
Interna utredningar som utförs av Europeiska byrån för bedrägeribekämpning (OLAF)
KAPITEL
2
UPPDRAG
Artikel
11
Äldste ledamoten
Artikel
12
Nomineringar och allmänna bestämmelser
Artikel
13
Val av talman - öppningsanförande
Artikel
14
Val av vice talmän
Artikel
15
Val av kvestorer
Artikel
16
Mandattid
Artikel
17
Lediga poster
Artikel
18
Entledigande
KAPITEL
3
ORGAN OCH UPPGIFTER
Artikel
19
Talmannens uppgifter
Artikel
20
Vice talmännens uppgifter
Artikel
21
Presidiets sammansättning
Artikel
22
Presidiets uppgifter
Artikel
23
Talmanskonferensens sammansättning
Artikel
24
Talmanskonferensens uppgifter
Artikel
25
Kvestorernas uppgifter
Artikel
26
Utskottsordförandekonferensen
Artikel
27
Delegationsordförandekonferensen
Artikel
28
Offentlighet när det gäller presidiet och talmanskonferensen
KAPITEL
4
POLITISKA GRUPPER
Artikel
29
Bildande av politiska grupper
Artikel
30
De politiska gruppernas verksamhet och rättsliga ställning
Artikel
31
Grupplösa ledamöter
Artikel
32
Fördelning av platser i plenisalen
AVDELNING
II
LAGSTIFTNING, BUDGET OCH ANDRA FÖRFARANDEN
KAPITEL
1
LAGSTIFTNINGSFÖRFARANDEN - ALLMÄNNA BESTÄMMELSER
Artikel
33
Kommissionens lagstiftnings- och arbetsprogram
Artikel
34
Prövning av respekten för de grundläggande rättigheterna, subsidiaritets- och proportionalitetsprinciperna och rättsstatsprincipen samt av de ekonomiska konsekvenserna
Artikel
35
Prövning av den rättsliga grunden
Artikel
36
Prövning av ekonomisk förenlighet
Artikel
37
Parlamentets tillgång till handlingar och information till parlamentet
Artikel
38
Parlamentets företrädare vid rådsmöten
Artikel
38 a
Parlamentets initiativrätt enligt fördragen
Artikel
39
Initiativ enligt artikel 192 i EG-fördraget
Artikel
40
Beredning av lagstiftningsdokument
Artikel
41
Samråd om initiativ som läggs fram av en medlemsstat
KAPITEL
2
FÖRFARANDEN I UTSKOTTEN
Artikel
42
Betänkanden som avser lagstiftning
Artikel
43
Förenklat förfarande
Artikel
44
Betänkanden som inte avser lagstiftning
Artikel
45
Initiativbetänkanden
Artikel
46
Utskottsyttranden
Artikel
47
Förfarande med associerade utskott
Artikel
48
Utarbetande av betänkanden
KAPITEL
3
FÖRSTA BEHANDLINGEN
I utskotten
Artikel
49
Ändring av kommissionsförslag
Artikel
50
Kommissionens och rådets ståndpunkt vid ändringsförslag
I kammaren
Artikel
51
Avslutande av första behandlingen
Artikel
52
Förkastande av kommissionsförslag
Artikel
53
Antagande av ändringar till ett kommissionsförslag
Uppföljning
Artikel
54
Uppföljning av parlamentets yttranden
Artikel
55
Framläggande av ett nytt förslag för parlamentet
Artikel
56
Medlingsförfarandet enligt den gemensamma förklaringen från 1975
KAPITEL
4
ANDRA BEHANDLINGEN
I utskotten
Artikel
57
Mottagande av rådets gemensamma ståndpunkt
Artikel
58
Förlängning av tidsfrister
Artikel
59
Hänvisning till och förfarande i ansvarigt utskott
I kammaren
Artikel
60
Avslutande av andra behandlingen
Artikel
61
Avvisning av rådets gemensamma ståndpunkt
Artikel
62
Ändringsförslag till rådets gemensamma ståndpunkt
KAPITEL
5
TREDJE BEHANDLINGEN
Förlikning
Artikel
63
Sammankallande av förlikningskommittén
Artikel
64
Delegationen till förlikningskommittén
I kammaren
Artikel
65
Gemensamt utkast
KAPITEL
6
LAGSTIFTNINGSFÖRFARANDET - AVSLUTANDE
Artikel
66
Överenskommelse vid första behandlingen
Artikel
67
Överenskommelse vid andra behandlingen
Artikel
68
Undertecknande av antagna rättsakter
KAPITEL
7
BUDGETFÖRFARANDEN
Artikel
69
Allmänna budgeten
Artikel
70
Ansvarsfrihet för kommissionen beträffande genomförandet av budgeten
Artikel
71
Andra förfaranden för beviljande av ansvarsfrihet
Artikel
72
Parlamentets kontroll över genomförandet av budgeten
KAPITEL
8
INTERNA BUDGETFÖRFARANDEN
Artikel
73
Parlamentets budgetberäkning
Artikel
74
Ekonomiska åtaganden och reglering av utgifter
KAPITEL
9
SAMTYCKESFÖRFARANDET
Artikel
75
Samtyckesförfarandet
KAPITEL
10
NÄRMARE SAMARBETE
Artikel
76
Förfaranden i parlamentet
KAPITEL
11
ÖVRIGA FÖRFARANDEN
Artikel
77
Yttranden i enlighet med artikel 122 i EG-fördraget
Artikel
78
Förfaranden som rör dialogen mellan arbetsmarknadens parter
Artikel
79
Förfaranden för kontroll av frivilliga överenskommelser
Artikel
80
Kodifiering
Artikel
80 a
Omarbetning
Artikel
81
Genomförandeåtgärder
KAPITEL
12
FÖRDRAG OCH INTERNATIONELLA AVTAL
Artikel
82
Anslutningsfördrag
Artikel
83
Internationella avtal
Artikel
84
Förfaranden enligt artikel 300 i EG-fördraget när det gäller provisorisk tillämpning eller tillfälligt upphävande av internationella avtal eller fastställande av gemenskapens ståndpunkt i ett organ som inrättats genom ett internationellt avtal
KAPITEL
13
UNIONENS EXTERNA REPRESENTATION OCH DEN GEMENSAMMA UTRIKES- OCH SÄKERHETSPOLITIKEN
Artikel
85
Utnämning av den höge representanten för den gemensamma utrikes- och säkerhetspolitiken
Artikel
86
Utnämning av särskilda representanter inom ramen för den gemensamma utrikes- och säkerhetspolitiken
Artikel
87
Uttalanden av den höge representanten för den gemensamma utrikes- och säkerhetspolitiken och andra särskilda representanter
Artikel
88
Internationell representation
Artikel
89
Samråd med och underrättande av parlamentet inom ramen för den gemensamma utrikes- och säkerhetspolitiken
Artikel
90
Rekommendationer inom ramen för den gemensamma utrikes- och säkerhetspolitiken
Artikel
91
Kränkningar av de mänskliga rättigheterna
KAPITEL
14
POLISSAMARBETE OCH STRAFFRÄTTSLIGT SAMARBETE
Artikel
92
Information till parlamentet när det gäller polissamarbete och straffrättsligt samarbete
Artikel
93
Samråd med parlamentet när det gäller polissamarbete och straffrättsligt samarbete
Artikel
94
Rekommendationer när det gäller polissamarbete och straffrättsligt samarbete
KAPITEL
15
EN MEDLEMSSTATS ÅSIDOSÄTTANDE AV GRUNDLÄGGANDE PRINCIPER
Artikel
95
Fastslående av åsidosättande
AVDELNING
III
ÖPPENHET OCH INSYN
Artikel
96
Insyn i parlamentets verksamhet
Artikel
97
Allmänhetens tillgång till handlingar
AVDELNING
IV
FÖRBINDELSER MED ANDRA ORGAN
KAPITEL
1
NOMINERINGAR OCH UTNÄMNINGAR
Artikel
98
Val av kommissionens ordförande
Artikel
99
Val av kommissionen
Artikel
100
Misstroendeförklaring mot kommissionen
Artikel
101
Utnämning av revisionsrättens ledamöter
Artikel
102
Utnämning av direktionsledamöter i Europeiska centralbanken
KAPITEL
2
UTTALANDEN
Artikel
103
Uttalanden av kommissionen, rådet och Europeiska rådet
Artikel
104
Förklaringar av kommissionens beslut
Artikel
105
Uttalanden av revisionsrätten
Artikel
106
Uttalanden av Europeiska centralbanken
Artikel
107
Rekommendation om de allmänna riktlinjerna för den ekonomiska politiken
KAPITEL
3
FRÅGOR TILL RÅDET, KOMMISSIONEN OCH EUROPEISKA CENTRALBANKEN
Artikel
108
Frågor för muntligt besvarande med debatt
Artikel
109
Frågestund
Artikel
110
Frågor till rådet och kommissionen för skriftligt besvarande
Artikel
111
Frågor till Europeiska centralbanken för skriftligt besvarande
KAPITEL
4
RAPPORTER FRÅN ANDRA INSTITUTIONER
Artikel
112
Årsrapporter och andra rapporter från andra institutioner
KAPITEL
5
RESOLUTIONER OCH REKOMMENDATIONER
Artikel
113
Resolutionsförslag
Artikel
114
Rekommendationer till rådet
Artikel
115
Debatter om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer
Artikel
116
Skriftliga förklaringar
Artikel
117
Samråd med Europeiska ekonomiska och sociala kommittén
Artikel
118
Samråd med Regionkommittén
Artikel
119
Begäran till EU-organ
KAPITEL
6
INTERINSTITUTIONELLA AVTAL
Artikel
120
Interinstitutionella avtal
KAPITEL
7
FÖRFARANDEN VID DOMSTOLEN
Artikel
121
Förfaranden vid domstolen
Artikel
122
Följder av rådets underlåtenhet att agera efter det att dess gemensamma ståndpunkt har godkänts enligt samarbetsförfarandet
AVDELNING
V
FÖRBINDELSER MED NATIONELLA PARLAMENT
Artikel
123
Utbyte av uppgifter samt kontakter och ömsesidiga resurser
Artikel
124
Konferensen mellan organ för EG- och EU-frågor (COSAC)
Artikel
125
Parlamentariska konferenser
AVDELNING
VI
SESSIONER
KAPITEL
1
PARLAMENTETS SESSIONER
Artikel
126
Parlamentets valperiod, sessioner, sammanträdesperioder, sammanträden
Artikel
127
Sammankallande av parlamentet
Artikel
128
Plats för sammanträden
Artikel
129
Deltagande i sammanträden
KAPITEL
2
PARLAMENTETS ARBETSGÅNG
Artikel
130
Förslag till föredragningslista
Artikel
131
Förfarande i kammaren utan ändringsförslag och debatt
Artikel
131 a
Kortfattad redogörelse
Artikel
132
Godkännande och ändring av föredragningslistan
Artikel
133
Särskild debatt
Artikel
134
Brådskande debatt
Artikel
135
Gemensam debatt
Artikel
136
Tidsfrister
KAPITEL
3
ALLMÄNNA BESTÄMMELSER FÖR PLENARSAMMANTRÄDEN
Artikel
137
Tillträde till plenisalen
Artikel
138
Språk
Artikel
139
Övergångsbestämmelser
Artikel
140
Utdelning av handlingar
Artikel
141
Tilldelning av ordet och anförandens innehåll
Artikel
142
Fördelning av talartid
Artikel
143
Talarlista
Artikel
144
Anföranden på en minut
Artikel
145
Personliga uttalanden
KAPITEL
4
ÅTGÄRDER VID LEDAMÖTERS ÖVERTRÄDELSE AV ORDNINGSREGLERNA
Artikel
146
Omedelbara åtgärder
Artikel
147
Påföljder
Artikel
148
Internt förfarande för överklagande
KAPITEL
5
BESLUTFÖRHET OCH OMRÖSTNING
Artikel
149
Beslutförhet
Artikel
150
Ingivande och framläggande av ändringsförslag
Artikel
151
Ändringsförslags tillåtlighet
Artikel
152
Omröstningar
Artikel
153
Lika röstetal
Artikel
154
Grundläggande principer för omröstningen
Artikel
155
Omröstningsordning vid ändringsförslag
Artikel
156
Behandling i utskott av ändringsförslag ingivna för behandling i plenum
Artikel
157
Delad omröstning
Artikel
158
Rösträtt
Artikel
159
Omröstning
Artikel
160
Omröstning med namnupprop
Artikel
161
Elektronisk omröstning
Artikel
162
Sluten omröstning
Artikel
163
Röstförklaringar
Artikel
164
Invändningar beträffande omröstningar
KAPITEL
6
PROCEDURFRÅGOR
Artikel
165
Förslag som rör förfaranden
Artikel
166
Ordningsfrågor
Artikel
167
Avvisning av ett ärende som otillåtligt
Artikel
168
Återförvisning till utskott
Artikel
169
Avslutande av debatt
Artikel
170
Uppskjutande av debatt och omröstning
Artikel
171
Avbrytande eller avslutande av sammanträde
KAPITEL
7
DOKUMENTATION AV SAMMANTRÄDEN
Artikel
172
Protokoll
Artikel
173
Fullständigt förhandlingsreferat
Artikel
173 a
Audiovisuell upptagning av förhandlingar
AVDELNING
VII
UTSKOTT, UNDERSÖKNINGSKOMMITTÉER OCH DELEGATIONER
KAPITEL
1
UTSKOTT OCH UNDERSÖKNINGSKOMMITTÉER - TILLSÄTTNING OCH BEHÖRIGHETSOMRÅDEN
Artikel
174
Tillsättning av ständiga utskott
Artikel
175
Tillsättning av tillfälliga utskott
Artikel
176
Undersökningskommittéer
Artikel
177
Utskottens och undersökningskommittéernas sammansättning
Artikel
178
Suppleanter
Artikel
179
Utskottens behörighetsområden
Artikel
180
Utskott med ansvar för valprövning
Artikel
181
Underutskott
Artikel
182
Utskottspresidium
KAPITEL
2
UTSKOTT OCH UNDERSÖKNINGSKOMMITTÉER - ARBETSSÄTT
Artikel
183
Utskottssammanträden
Artikel
184
Protokoll från utskottssammanträden
Artikel
185
Omröstningar i utskott
Artikel
186
Bestämmelser för plenarsammanträden som även ska gälla utskottssammanträden
Artikel
187
Frågestund i utskott
KAPITEL
3
INTERPARLAMENTARISKA DELEGATIONER
Artikel
188
Tillsättning av interparlamentariska delegationer och delegationernas uppgifter
Artikel
189
Samarbete med Europarådets parlamentariska församling
Artikel
190
Gemensamma parlamentarikerkommittéer
AVDELNING
VIII
FRAMSTÄLLNINGAR
Artikel
191
Rätt att inge framställningar
Artikel
192
Prövning av framställningar
Artikel
193
Tillkännagivande av framställningar
AVDELNING
IX
OMBUDSMANNEN
Artikel
194
Utnämning av ombudsmannen
Artikel
195
Ombudsmannens verksamhet
Artikel
196
Avsättning av ombudsmannen
AVDELNING
X
PARLAMENTETS GENERALSEKRETARIAT
Artikel
197
Generalsekretariat
AVDELNING
XI
BEFOGENHETER GÄLLANDE POLITISKA PARTIER PÅ EUROPEISK NIVÅ
Artikel
198
Talmannens befogenheter
Artikel
199
Presidiets befogenheter
Artikel
200
Ansvarigt utskotts och plenums befogenheter
AVDELNING
XII
TILLÄMPNING OCH ÄNDRING AV ARBETSORDNINGEN
Artikel
201
Tillämpning av arbetsordningen
Artikel
202
Ändring av arbetsordningen
AVDELNING
XIII
DIVERSE BESTÄMMELSER
Artikel
203
Oavslutade ärenden
Artikel
204
Bilagor till arbetsordningen
Artikel
204 a
Rättelser
BILAGA
I
BILAGA
II
Genomförande av frågestunden i artikel 109
BILAGA
II a
Riktlinjer för frågor för skriftligt besvarande enligt artiklarna 110 och 111
BILAGA
III
Riktlinjer och allmänna principer för att fastställa vilka frågor som ska tas upp på föredragningslistan till debatter om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer enligt artikel 115
BILAGA
IV
Genomförandebestämmelser för behandling av Europeiska unionens allmänna budget och tilläggsbudgetar
BILAGA
V
Förfarande för överläggningar om och antagande av beslut om beviljande av ansvarsfrihet
BILAGA
VI
Ständiga utskotts behörighetsområden
I.
Utskottet för utrikesfrågor
II.
Utskottet för utveckling
III.
Utskottet för internationell handel
IV.
Budgetutskottet
V.
Budgetkontrollutskottet
VI.
Utskottet för ekonomi och valutafrågor
VII.
Utskottet för sysselsättning och sociala frågor
VIII.
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
IX.
Utskottet för industrifrågor, forskning och energi
X.
Utskottet för den inre marknaden och konsumentskydd
XI.
Utskottet för transport och turism
XII.
Utskottet för regional utveckling
XIII.
Utskottet för jordbruk och landsbygdens utveckling
XIV.
Fiskeriutskottet
XV.
Utskottet för kultur och utbildning
XVI.
Utskottet för rättsliga frågor
XVII.
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
XVIII.
Utskottet för konstitutionella frågor
XIX.
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
XX.
Utskottet för framställningar
BILAGA
VII
Sekretessbelagda handlingar och känslig information
BILAGA
VIII
Närmare föreskrifter för utövandet av Europaparlamentets undersökningsrätt
BILAGA
IX
BILAGA
X
Ombudsmannens ämbetsutövning
BILAGA
XI
Villkor och närmare bestämmelser för interna utredningar för att bekämpa bedrägerier, korruption och all annan olaglig verksamhet som kan skada gemenskapernas intressen
BILAGA
XII
Överenskommelse mellan Europaparlamentet och kommissionen om tillämpningsföreskrifter till rådets beslut 1999/468/EG, om de förfaranden som ska tillämpas vid utövandet av kommissionens genomförandebefogenheter, ändrat genom beslut 2006/512/EG
BILAGA
XIII
Ramavtal om förbindelserna mellan Europaparlamentet och kommissionen
BILAGA
XIV
(utgår)
BILAGA
XV
Förteckning över de handlingar som allmänheten ges direkt tillgång till via register över parlamentshandlingar
BILAGA
XVI
Förordning (EG) nr 1049/2001 om allmänhetens tillgång till handlingar
BILAGA
XVI a
Riktlinjer för tolkning av ordningsreglerna för ledamöterna
BILAGA
XVI b
Riktlinjer för godkännande av kommissionen
BILAGA
XVI c
Förfarandet för att bevilja tillstånd att utarbeta initiativbetänkanden
AVDELNING
I
LEDAMÖTER, PARLAMENTETS ORGAN OCH POLITISKA GRUPPER
KAPITEL
1
EUROPAPARLAMENTETS LEDAMÖTER
Artikel
1
Europaparlamentet
1.
Europaparlamentet är den församling som är vald i överensstämmelse med fördragen, akten av den 20 september 1976 om allmänna direkta val av ledamöter av Europaparlamentet samt den från fördragen härledda nationella lagstiftningen.
2.
Europaparlamentets valda företrädare benämns:
"Членове на Европейския парламент" på bulgariska,
"Diputados al Parlamento Europeo" på spanska,
"Poslanci Evropského parlamentu" på tjeckiska,
"Medlemmer af Europa-Parlamentet" på danska,
"Mitglieder des Europäischen Parlaments" på tyska,
"Euroopa Parlamendi liikmed" på estniska,
"Βoυλευτές τoυ Ευρωπαϊκoύ Κoιvoβoυλίoυ" på grekiska,
"Members of the European Parliament" på engelska,
"Deputés au Parlement européen" på franska,
"Feisirí de Pharlaimint na hEorpa" på iriska,
"Deputati al Parlamento europeo" på italienska,
"Eiropas Parlamenta deputāti" på lettiska,
"Europos Parlamento nariai" på litauiska,
"Európai Parlamenti Képviselők" på ungerska,
"Membru tal-Parlament Ewropew" på maltesiska,
"Leden van het Europees Parlement" på nederländska,
"Posłowie do Parlamentu Europejskiego" på polska,
"Deputados ao Parlamento Europeu" på portugisiska,
"Deputaţi în Parlamentul European" på rumänska,
"Poslanci Európskeho parlamentu" på slovakiska,
"Poslanci Evropskega parlamenta" på slovenska,
"Euroopan parlamentin jäsenet" på finska samt
"Ledamöter av Europaparlamentet" på svenska.
Artikel
2
Obundet mandat
Europaparlamentets ledamöter har ett obundet mandat.
De får inte bindas av instruktioner eller uppdrag.
Artikel
3
Valprövning
1.
Efter val till Europaparlamentet ska dess ordförande (härefter kallad talman) uppmana de behöriga myndigheterna i medlemsstaterna att utan dröjsmål meddela parlamentet namnen på de valda ledamöterna, så att alla ledamöter kan tillträda sitt uppdrag i parlamentet från och med öppnandet av det första sammanträdet efter valet.
Samtidigt ska talmannen göra dessa myndigheter uppmärksamma på de relevanta bestämmelserna i akten av den 20 september 1976 och uppmana dem att vidta de åtgärder som är nödvändiga för att undvika oförenlighet med uppdraget som ledamot av Europaparlamentet.
2.
Efter allmänna val ska denna förklaring om möjligt avges senast sex dagar före parlamentets konstituerande sammanträde.
Fram till dess att bevis om val av ledamöter har granskats eller beslut fattats beträffande en eventuell tvist, förutsatt att han undertecknat den ovannämnda skriftliga förklaringen, ska ledamoten tillträda sina uppdrag i parlamentet och i dess organ, varvid han ska ha alla de rättigheter som följer av uppdragen.
3.
Med utgångspunkt i ett betänkande från behörigt utskott ska parlamentet omgående granska bevisen om val av ledmöter och avgöra varje enskild ny ledamots mandat, samt eventuella tvister som uppkommer till följd av bestämmelserna i akten av den 20 september 1976 med undantag av invändningar som grundar sig på nationella vallagar.
4.
Behörigt utskotts betänkande ska grunda sig på de officiella kungörelserna från de enskilda medlemsstaterna om det samlade valresultatet, vilka innehåller namnen på de valda kandidaterna och deras ersättare samt en rangordning baserad på valresultatet.
Giltigheten av en ledamots mandat får inte bekräftas förrän ledamoten har avgivit de skriftliga förklaringar som följer av denna artikel och bilaga I till arbetsordningen.
Parlamentet kan när som helst på grundval av ett betänkande från sitt behöriga utskott yttra sig om varje invändning mot ett mandats giltighet.
5.
6.
När behöriga myndigheter i medlemsstaterna inleder ett förfarande som kan leda till att en ledamot skiljs från sitt uppdrag, ska talmannen begära regelbunden information från dem om hur förfarandet framskrider.
Talmannen ska hänvisa ärendet till behörigt utskott, och parlamentet kan yttra sig på förslag av detta utskott.
Artikel
4
Mandatets varaktighet
1.
Mandatet börjar och slutar i enlighet med akten av den 20 september 1976.
Det upphör också när en ledamot avlider eller begär entledigande.
2.
Alla ledamöter har kvar sina uppdrag till dess att parlamentets första sammanträde efter valet öppnas.
3.
Varje ledamot som begär entledigande ska anmäla detta till talmannen tillsammans med angivande av det datum då avgången ska gälla, vilket inte får vara senare än tre månader efter anmälan.
Anser det behöriga utskottet att begäran om entledigande strider mot andan eller bokstaven i akten av den 20 september 1976, ska parlamentet underrättas om detta, så att parlamentet kan avgöra om platsen ska förklaras vakant eller inte.
I annat fall konstateras platsen vakant från och med det datum som den avgående ledamoten har angivit i det skriftliga protokollet.
Det sker ingen omröstning i parlamentet i detta fall.
4.
5.
Medlemsstaternas eller unionens myndigheter ska underrätta talmannen om varje uppdrag som de ämnar anförtro en ledamot.
Talmannen ska hänvisa frågan om huruvida uppdraget är förenligt med andan och bokstaven i akten av den 20 september 1976 till det behöriga utskottet.
Talmannen ska underrätta kammaren, den berörde ledamoten och de berörda myndigheterna om utskottets slutsatser.
6.
Mandatet ska anses ha upphört och platsen vara vakant från och med följande tidpunkter:
-
Vid tilldelning av ett uppdrag eller val till ett ämbete (se artikel 4.4 andra stycket) som inte är förenligt med uppdraget som ledamot av Europaparlamentet enligt vad som avses i artikel 7.1 eller 7.2 i akten av den 20 september 1976: från och med den dag som ledamoten eller medlemsstaternas eller unionens behöriga myndigheter angivit.
7.
När parlamentet fastställt att en plats är vakant ska det underrätta berörd medlemsstat om detta och uppmana den att utan dröjsmål tillsätta den vakanta platsen.
8.
Alla tvister rörande giltigheten av mandatet för en ledamot vars bevis redan granskats ska hänvisas till behörigt utskott, som omgående och senast vid början av nästföljande sammanträdesperiod ska underrätta parlamentet.
9.
Parlamentet förbehåller sig rätten att ogiltigförklara det mandat som är under prövning eller att inte fastställa att platsen (se t.ex. punkt 9) är vakant, då det i förbindelse med godkännandet eller upphävandet av mandatet konstateras att felaktigheter eller brister föreligger.
Artikel
5
Immunitet och privilegier
1.
Ledamöterna åtnjuter immunitet och privilegier i enlighet med protokollet om Europeiska gemenskapernas immunitet och privilegier.
2.
Passerkort som tillåter ledamöterna att fritt röra sig i medlemsstaterna ska utfärdas av parlamentets talman så snart talmannen meddelats vilka ledamöter som valts.
3.
Ledamöterna har rätt att ta del av alla handlingar som parlamentets eller ett utskott innehar, med undantag av personakter och personliga räkenskaper, vilka endast de berörda ledamöterna har rätt att ta del av.
I bilaga VII till denna arbetsordning finns bestämmelser om undantag från denna princip när det gäller hantering av sådana handlingar som allmänheten kan nekas tillgång till i enlighet med Europaparlamentets och rådets förordning (EG) nr 1049/2001 om allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar.
Artikel
6
Upphävande av immunitet
1.
Parlamentet ska vid utövandet av sina befogenheter i frågor som rör immunitet och privilegier i första hand försöka upprätthålla parlamentets integritet som en demokratisk lagstiftande församling och befästa ledamöternas oberoende när dessa fullgör sina åligganden.
2.
Varje begäran ställd till talmannen från en i en medlemsstat behörig myndighet om upphävande av en ledamots immunitet ska tillkännages i kammaren och hänvisas till behörigt utskott.
3.
Varje begäran om fastställelse av immunitet och privilegier som en ledamot eller före detta ledamot lämnar in till talmannen ska tillkännages i kammaren och hänvisas till behörigt utskott.
Ledamoten eller den före detta ledamoten kan representeras av en annan ledamot.
En begäran kan inte lämnas in av en annan ledamot utan den berörde ledamotens samtycke.
4.
Om en ledamot grips eller får sin rörelsefrihet begränsad på ett sätt som förmodas kränka ledamotens immunitet och privilegier kan talmannen, i brådskande fall och efter samråd med det behöriga utskottets ordförande och föredragande, själv ta initiativ till att bekräfta ledamotens immunitet och privilegier.
Talmannen ska meddela utskottet detta och informera parlamentet.
Artikel
7
Immunitetsförfaranden
1.
Behörigt utskott ska utan dröjsmål, och i den ordning de inkommit, pröva varje begäran om upphävande av immunitet och varje begäran om fastställelse av immunitet eller privilegier.
2.
Utskottet ska lägga fram ett förslag till beslut, i vilket utskottet endast ska rekommendera huruvida en begäran om upphävande av immuniteten eller en begäran om fastställelse av immunitet och privilegier ska bifallas eller avslås.
3.
Utskottet kan uppmana den berörda myndigheten att förse utskottet med alla upplysningar och preciseringar som det anser sig behöva för att kunna ta ställning till om immuniteten bör upphävas eller fastställas.
De har rätt att låta sig företrädas av en annan ledamot.
4.
Om en begäran om upphävande av immunitet hänför sig till flera gärningar kan upphävande av immuniteten beträffande var och en av dessa gärningar bli föremål för ett enskilt beslut.
I utskottets betänkande kan det i undantagsfall föreslås att upphävandet av immuniteten endast ska beröra åtalet och att ledamoten, så länge som det inte finns någon lagakraftvunnen dom varken kan gripas, anhållas, häktas eller utsättas för någon annan åtgärd som skulle förhindra ledamoten att utföra sina åligganden i enlighet med uppdraget som ledamot av Europaparlamentet.
5.
När en ledamot anmodas att vittna eller framträda som sakkunnig behöver ingen begäran om upphävande av immuniteten inges, under förutsättning att
ledamoten inte är skyldig att avlägga vittnesmål som omfattar sådana sekretessbelagda uppgifter som erhållits under utövandet av uppdraget som ledamot och som ledamoten inte anser sig kunna röja.
6.
7.
Utskottet får emellertid under inga omständigheter uttala sig i skuldfrågan, eller på annat sätt yttra sig över ledamoten eller om det riktiga i att väcka åtal för de uttalanden eller handlingar som tillskrivs ledamoten, inte ens vid tillfällen där utskottet genom prövning av en begäran erhåller detaljerad kunskap i fallet.
8.
Utskottets betänkande ska tas upp som första punkt på föredragningslistan till det första sammanträdet efter det att betänkandet har getts in.
Det är inte tillåtet att lägga fram ändringsförslag till förslaget eller förslagen till beslut.
Det är endast tillåtet att debattera grunderna för och emot varje enskilt förslag om att upphäva eller upprätthålla immunitet eller fastställa immunitet eller privilegier.
Utan att det påverkar tillämpningen av artikel 145 får den ledamot vars immunitet eller privilegier det är fråga om inte yttra sig i debatten.
Omröstning om betänkandets förslag till beslut ska ske vid det första omröstningstillfället efter det att debatten avslutats.
Efter behandling i kammaren ska särskild omröstning ske om varje enskilt förslag i betänkandet.
Om ett förslag förkastas ska motsatt beslut anses fattat.
9.
Talmannen ska omedelbart meddela parlamentets beslut till ledamoten i fråga och till behörig myndighet i berörd medlemsstat och begära att talmannen hålls underrättad om hur de relevanta förfarandena fortskrider och om eventuella beslut i samband därmed.
När talmannen erhåller denna information, ska parlamentet, vid behov efter samråd med behörigt utskott, underrättas på det sätt talmannen finner mest lämpligt.
10.
Om utskottet anser det nödvändigt kan det lägga fram ett betänkande till parlamentet.
11.
Utskottet ska vid behandlingen av dessa ärenden och eventuella handlingar det tar emot iaktta strikt sekretess.
12.
Efter att ha hört medlemsstaterna kan utskottet utarbeta en vägledande förteckning över de myndigheter i de olika medlemsstaterna som är behöriga att inkomma med en begäran om upphävande av en ledamots immunitet.
13.
Alla förfrågningar som en behörig myndighet gör beträffande omfattningen av ledamöternas immunitet och privilegier ska behandlas i enlighet med bestämmelserna ovan.
Artikel
8
Kostnadsersättning och andra ersättningar
Presidiet ska fastställa bestämmelser om kostnadsersättning och andra ersättningar till ledamöterna.
Artikel
9
Ledamöternas ekonomiska intressen, ordningsregler och tillträde till parlamentet
1.
Parlamentet kan fastställa regler om öppenhet i fråga om ledamöternas ekonomiska intressen, vilka fogas som bilaga till arbetsordningen
Se bilaga I.
.
Dessa regler får på intet sätt hindra eller begränsa en ledamots utövande av sitt mandat, politisk verksamhet eller annan verksamhet i förbindelse härmed.
2.
Ledamöternas uppträdande ska präglas av ömsesidig respekt baserad på de värderingar och principer som fastställs i Europeiska unionens grundläggande rättsakter, ledamöterna ska slå vakt om parlamentets värdighet, samt uppträda på ett sätt som inte stör parlamentets arbete eller ordningen i någon av parlamentets byggnader.
Om dessa principer inte respekteras kan de åtgärder som föreskrivs i artiklarna 146, 147 och 148 komma att tillämpas.
3.
Tillämpningen av denna artikel ska inte ligga till hinder för en livlig debatt i parlamentet eller begränsa ledamöternas yttrandefrihet.
Artikeln ska tillämpas med fullt iakttagande av ledamöternas befogenheter, i enlighet med vad som fastställs i primärrätten och i ledamotsstadgan.
Artikeln ska tillämpas med iakttagande av öppenhetsprincipen och på ett sätt som medför att ledamöterna underrättas om alla gällande bestämmelser om öppenhet samt informeras personligen om sina rättigheter och skyldigheter.
4.
Kvestorerna ska ansvara för utfärdandet av personliga passerkort med en giltighet på högst ett år till personer som regelbundet vill ha tillträde till parlamentets lokaler för att i eget eller tredje mans intresse förse ledamöter med information inom ramen för ledamöternas mandat.
Dessa personer ska i gengäld
-
följa de ordningsregler som anges i en bilaga till arbetsordningen
Se bilaga IX.
,
-
skriva in sig i ett register som förs av kvestorerna.
Allmänheten kan på begäran få ta del av detta register på alla parlamentets arbetsorter och på parlamentets informationskontor i medlemsstaterna på det sätt som kvestorerna fastställer.
Närmare föreskrifter för tillämpningen av denna punkt ska anges i en bilaga till arbetsordningen
Se bilaga IX.
.
5.
Ordningsregler, rättigheter och privilegier för före detta ledamöter ska fastställas genom ett beslut av presidiet.
Alla före detta ledamöter ska behandlas lika.
Artikel
10
Interna utredningar som utförs av Europeiska byrån för bedrägeribekämpning (OLAF)
Se bilaga XI.
.
KAPITEL
2
UPPDRAG
Artikel
11
Äldste ledamoten
1.
2.
Under den äldste ledamotens ledning får inga andra frågor behandlas än sådana som rör val av talman eller granskning av bevis om val av ledamöter.
Övriga frågor som rör granskning av bevis om val av ledamöter och som tas upp under den ledamotens ledning av sammanträdet ska hänvisas till utskottet med behörighet i frågor som rör valprövning.
Artikel
12
Nomineringar och allmänna bestämmelser
1.
Talman, vice talmän och kvestorer väljs genom sluten omröstning i enlighet med vad som föreskrivs i artikel 162.
Nominering kan endast ske med de berörda parternas samtycke.
Nomineringar kan endast göras av politiska grupper eller minst 40 ledamöter.
Om antalet kandidater inte överstiger antalet lediga platser, kan emellertid kandidaterna väljas med acklamation.
2.
Vid val av talman, vice talmän och kvestorer bör hänsyn tas till behovet av en för medlemsstaterna och de politiska åsiktsriktningarna övergripande rättvis representation.
Artikel
13
Val av talman - öppningsanförande
1.
Talmannen ska väljas först.
Före varje omröstning ska nomineringarna föreläggas ålderspresidenten, som ska underrätta parlamentet.
Har ingen kandidat erhållit absolut majoritet av de avgivna rösterna efter tre valomgångar, begränsas den fjärde valomgången till de två kandidater som i den tredje valomgången erhöll flest antal röster.
Vid lika röstetal förklaras den äldste kandidaten vald.
2.
Så snart talmannen är vald ska ålderspresidenten överlämna ordförandeposten till talmannen.
Endast den nyvalde talmannen får hålla ett öppningsanförande.
Artikel
14
Val av vice talmän
1.
Därefter ska 14 vice talmän väljas från en enda valsedel.
Är antalet valda kandidater lägre än antalet personer som ska väljas, hålls en andra valomgång under samma betingelser för att fylla de återstående platserna.
Blir en tredje valomgång nödvändig, betraktas de kandidater som får flest röster som valda till de återstående platserna.
Vid lika röstetal förklaras de äldsta kandidaterna valda.
2.
När val inte har förrättats genom sluten omröstning är rangordningen den ordning i vilken talmannen läst upp namnen.
Artikel
15
Val av kvestorer
Efter valet av vice talmän ska parlamentet välja fem kvestorer.
Kvestorerna väljs enligt samma förfarande som de vice talmännen.
Trots vad som sägs i första stycket ska parlamentet för perioden januari 2007 till juli 2009 utse sex kvestorer.
Artikel
16
Mandattid
1.
Mandattiden för talmannen, vice talmännen och kvestorerna är två och ett halvt år.
Även om en ledamot ändrar sin grupptillhörighet, ska ledamoten under den resterande delen av sin mandattid på två och ett halvt år behålla sin eventuella plats i presidiet eller kvestorskollegiet.
2.
Blir en av dessa poster vakant före denna periods utgång, ska den ledamot som då väljs endast inneha sitt uppdrag till och med utgången av företrädarens mandattid.
Artikel
17
Lediga poster
1.
Om det blir nödvändigt att ersätta talmannen, en vice talman eller en kvestor ska ersättare väljas i enlighet med bestämmelserna ovan.
En nyvald vice talman intar sin företrädares plats enligt rangordningen för vice talmän.
2.
Blir talmansposten ledig ska förste vice talmannen utföra talmannens uppgifter till dess att en ny talman valts.
Artikel
18
Entledigande
Talmanskonferensen får med en majoritet av tre femtedelar av de avgivna rösterna, som ska företräda minst tre politiska grupper, föreslå parlamentet att entlediga talmannen, en vice talman, en kvestor, en ordförande eller vice ordförande i ett utskott, en ordförande eller vice ordförande i en interparlamentarisk delegation, eller någon annan befattningshavare som utsetts av parlamentet, om talmanskonferensen anser att ledamoten i fråga har gjort sig skyldig till allvarlig försummelse.
För att godkänna ett sådant förslag krävs två tredjedelar av de avgivna rösterna och en majoritet av parlamentets samtliga ledamöter.
KAPITEL
3
ORGAN OCH UPPGIFTER
Artikel
19
Talmannens uppgifter
1.
Talmannen leder i enlighet med de i arbetsordningen fastställda reglerna allt arbete i parlamentet och dess organ.
I de befogenheter som följer av denna artikel ingår även att låta textdelar gå till omröstning i en annan ordning än den ordning i vilken de förekommer i den handling som omröstningen avser.
2.
Talmannen ska avgöra huruvida ändringsförslag ska förklaras tillåtliga, avgöra ärenden som rör frågor till rådet och kommissionen samt avgöra huruvida betänkanden uppfyller arbetsordningens bestämmelser.
Talmannen ska se till att arbetsordningen efterlevs, upprätthålla ordningen, ge talare ordet, förklara debatter avslutade, förrätta omröstningar och tillkännage omröstningsresultat.
3.
Talmannen får endast yttra sig i en debatt för att sammanfatta debatten och för att upprätthålla ordningen.
Om talmannen önskar delta i en debatt ska ordförandeskapet överlåtas, och talmannen får inte återta ordförandeskapet förrän debatten i fråga är avslutad.
4.
Artikel
20
Vice talmännens uppgifter
1.
2.
3.
Artikel
21
Presidiets sammansättning
1.
Presidiet består av talmannen och parlamentets 14 vice talmän.
2.
Kvestorerna är medlemmar av presidiet med rådgivande funktion.
3.
Talmannen har utslagsröst vid lika röstetal vid omröstningar i presidiet.
Artikel
22
Presidiets uppgifter
1.
Presidiet ska utföra de uppgifter det tilldelas enligt arbetsordningen.
2.
Presidiet ska avgöra ekonomiska, organisatoriska och administrativa ärenden som rör ledamöterna, parlamentets interna organisation, dess sekretariat och dess organ.
3.
Presidiet ska avgöra frågor som rör sammanträdesordningen.
Begreppet sammanträdesordning inbegriper frågor som rör ledamöternas uppträdande i parlamentets samtliga lokaler.
4.
Presidiet ska fastställa föreskrifter för grupplösa ledamöter i enlighet med artikel 31.
5.
Presidiet ska fastställa generalsekretariatets tjänsteförteckning samt föreskrifter för tjänstemäns och övriga anställdas rättsliga ställning och ekonomiska situation.
6.
Presidiet ska utarbeta parlamentets preliminära budgetberäkning.
7.
Presidiet ska fastställa riktlinjer för kvestorerna i enlighet med artikel 25.
8.
Presidiet är det organ som godkänner utskottssammanträden utanför de vanliga arbetsorterna, utskottsutfrågningar samt studie- och informationsresor för föredragande.
När sådana sammanträden eller sammankomster godkänns ska det fastställas vilka språkregler som ska gälla med utgångspunkt i de officiella språk som ledamöterna och suppleanterna i utskottet i fråga använder och begär.
Detsamma ska gälla för delegationerna, om inte berörda ledamöter och suppleanter beslutar annat.
9.
Presidiet ska utse en generalsekreterare i enlighet med artikel 197.
10.
Presidiet ska fastställa tillämpningsföreskrifter till Europaparlamentets och rådets förordning (EG) nr 2004/2003 om regler för och finansiering av politiska partier på europeisk nivå, och i samband med genomförandet av den förordningen utföra de uppgifter det tilldelas i arbetsordningen.
11.
Talmannen eller presidiet kan tilldela en eller flera medlemmar av presidiet allmänna eller specifika uppgifter som ligger inom talmannens eller presidiets behörighetsområde.
Samtidigt ska det fastställas hur dessa uppgifter ska genomföras.
12.
Vid nyval till parlamentet ska det avgående presidiet ha kvar sina uppgifter fram till dess att det nya parlamentet sammanträder för första gången.
Artikel
23
Talmanskonferensens sammansättning
1.
Talmanskonferensen består av talmannen och ordförandena i de politiska grupperna.
En ordförande i en politisk grupp kan låta sig företrädas av en medlem av sin grupp.
2.
De grupplösa ledamöterna ska ge en av sina ledamöter i uppdrag att delta vid talmanskonferensens sammanträden.
Denna ledamot har inte rösträtt.
3.
Talmanskonferensen ska anstränga sig för att nå konsensus i frågor som föreläggs den.
I fall där konsensus inte kan nås ska frågan gå till omröstning, i vilken gruppernas röster räknas i förhållande till antalet medlemmar i respektive grupp.
Artikel
24
Talmanskonferensens uppgifter
1.
Talmanskonferensen ska utföra de uppgifter den tilldelas enligt arbetsordningen.
2.
Talmanskonferensen ska fatta beslut om parlamentets arbetsorganisation och ärenden som rör planering av lagstiftningsarbete.
3.
Talmanskonferensen ska ansvara för frågor som rör förbindelserna med Europeiska unionens övriga organ och institutioner och med medlemsstaternas nationella parlament.
Presidiet ska utse två vice talmän som ska ansvara för förbindelserna med de nationella parlamenten.
Dessa ska regelbundet rapportera till talmanskonferensen om sin verksamhet i detta avseende.
4.
Talmanskonferensen ska ansvara för frågor som rör förbindelser med tredje land samt med institutioner och organisationer utanför Europeiska unionen.
5.
Talmanskonferensen ska utarbeta förslag till föredragningslista till parlamentets sammanträdesperioder.
6.
Talmanskonferensen ska ansvara för sammansättning av och befogenheter för utskott, undersökningskommittéer, gemensamma parlamentarikerkommittéer, ständiga delegationer och ad hoc-delegationer.
7.
Talmanskonferensen ska i enlighet med artikel 32 avgöra platsfördelningen i plenisalen.
8.
Talmanskonferensen är det organ som har behörighet att ge tillstånd att utarbeta initiativbetänkanden.
9.
Talmanskonferensen ska lämna in förslag till presidiet angående administrativa frågor och budgetfrågor som rör de olika politiska grupperna.
Artikel
25
Kvestorernas uppgifter
Kvestorerna ska ha ansvaret för administrativa och ekonomiska ärenden som direkt berör ledamöterna enligt riktlinjer fastställda av presidiet.
Artikel
26
Utskottsordförandekonferensen
1.
2.
Utskottsordförandekonferensen kan utfärda rekommendationer till talmanskonferensen angående utskottens arbete och upprättandet av föredragningslista till sammanträdesperioderna.
3.
Presidiet och talmanskonferensen kan ge utskottsordförandekonferensen i uppdrag att utföra vissa uppgifter.
Artikel
27
Delegationsordförandekonferensen
1.
2.
Delegationsordförandekonferensen kan utfärda rekommendationer till talmanskonferensen angående delegationernas arbete.
3.
Presidiet och talmanskonferensen kan ge delegationsordförandekonferensen i uppdrag att utföra vissa uppgifter.
Artikel
28
Offentlighet när det gäller presidiet och talmanskonferensen
1.
2.
Varje ledamot kan ställa frågor som rör presidiets, talmanskonferensens eller kvestorernas arbete.
Sådana frågor ska inges skriftligen till talmannen och tillsammans med de avgivna svaren offentliggöras i parlamentets bulletin inom trettio dagar från det att de ingavs.
KAPITEL
4
POLITISKA GRUPPER
Artikel
29
Bildande av politiska grupper
1.
Ledamöter får bilda grupper efter politisk samhörighet.
Parlamentet behöver i normala fall inte bedöma gruppledamöters politiska samhörighet.
Ledamöter som tillsammans bildar en grupp i enlighet med denna artikel ska per definition acceptera att de har politisk samhörighet.
Endast då de berörda ledamöterna förnekar detta blir det nödvändigt för parlamentet att utvärdera huruvida gruppen har bildats i överensstämmelse med arbetsordningens bestämmelser.
2.
En politisk grupp ska omfatta ledamöter som valts i minst en femtedel av medlemsstaterna.
För att bilda en politisk grupp fordras minst 20 ledamöter.
3.
En ledamot får inte tillhöra flera än en politisk grupp.
4.
Bildandet av en politisk grupp ska anmälas till talmannen.
Anmälan ska omfatta gruppens namn, dess medlemmar och dess ledning.
5.
Anmälan ska offentliggöras i Europeiska unionens officiella tidning.
Artikel
30
De politiska gruppernas verksamhet och rättsliga ställning
1.
De politiska grupperna ska utföra sina uppgifter inom ramen för unionens verksamhet, även de arbetsuppgifter som tillkommer dem genom arbetsordningen.
De politiska grupperna ska inom ramen för generalsekretariatets tjänsteförteckning förfoga över ett sekretariat, administrativa faciliteter och de anslag som förs upp i parlamentets budget.
2.
Presidiet ska fastställa bestämmelser om hur dessa faciliteter och anslag ska tillhandahållas, utnyttjas och kontrolleras samt om de härtill hörande delegeringarna av befogenheter att genomföra budgeten.
3.
I dessa bestämmelser ska anges de administrativa och ekonomiska konsekvenserna i händelse av att en politisk grupp upplöses.
Artikel
31
Grupplösa ledamöter
1.
Ledamöter som inte tillhör någon politisk grupp ska ha tillgång till ett sekretariat.
Närmare regler ska fastställas av presidiet på förslag av generalsekreteraren.
2.
Presidiet ska även avgöra sådana ledamöters ställning och parlamentariska rättigheter.
3.
Presidiet ska också fastställa bestämmelser om tillhandahållande, utnyttjande och kontroll av anslag som förs upp i parlamentets budget för att täcka de grupplösa ledamöternas utgifter för sekretariat och administrativa faciliteter.
Artikel
32
Fördelning av platser i plenisalen
Talmanskonferensen ska avgöra fördelningen av platser i plenisalen för de politiska grupperna, de grupplösa ledamöterna och Europeiska unionens institutioner.
AVDELNING
II
LAGSTIFTNING, BUDGET OCH ANDRA FÖRFARANDEN
KAPITEL
1
LAGSTIFTNINGSFÖRFARANDEN - ALLMÄNNA BESTÄMMELSER
Artikel
33
Kommissionens lagstiftnings- och arbetsprogram
1.
Parlamentet ska tillsammans med kommissionen och rådet utforma Europeiska unionens lagstiftningsprogram.
Parlamentet och kommissionen ska samarbeta under förberedelserna av kommissionens lagstiftnings- och arbetsprogram i enlighet med den tidsplan och de närmare föreskrifter som de två institutionerna kommit överens om och som fogats som bilaga till arbetsordningen
Se bilaga XIV.
.
2.
Vid brådskande och oförutsedda omständigheter har en institution rätt att på eget initiativ, och i enlighet med de förfaranden som föreskrivs i fördragen, föreslå lagstiftningsåtgärder utöver dem som föreslås i lagstiftningsprogrammet.
3.
Talmannen ska översända den av parlamentet antagna resolutionen till de andra institutionerna som deltar i Europeiska unionens lagstiftningsprocess och till medlemsstaternas parlament.
Talmannen ska uppmana rådet att yttra sig över kommissionens årliga lagstiftningsprogram samt över parlamentets resolution.
4.
Om en av institutionerna inte kan följa den fastställda tidsplanen ska den underrätta de andra institutionerna om skälen till förseningen och föreslå en ny tidsplan.
Artikel
34
Prövning av respekten för de grundläggande rättigheterna, subsidiaritets- och proportionalitetsprinciperna och rättsstatsprincipen samt av de ekonomiska konsekvenserna
Vid prövning av ett förslag till rättsakt ska parlamentet ta särskild hänsyn till huruvida förslaget respekterar de grundläggande rättigheterna och framför allt att rättsakten står i överensstämmelse med Europeiska unionens stadga om de grundläggande rättigheterna, subsidiaritets- och proportionalitetsprinciperna samt rättsstatsprincipen.
Har ett förslag ekonomiska konsekvenser ska parlamentet fastställa huruvida tillräckliga finansiella medel har föreslagits.
Artikel
35
Prövning av den rättsliga grunden
1.
Innan kommissionsförslag och andra dokument som avser lagstiftning behandlas, ska ansvarigt utskott först göra en bedömning av den rättsliga grund som valts.
2.
Om ansvarigt utskott anser att den rättsliga grunden är inkorrekt eller olämplig– inbegripet prövning i enlighet med artikel 5 i EG-fördraget – ska det begära att utskottet med behörighet i rättsliga frågor yttrar sig.
3.
Utskottet med behörighet i rättsliga frågor kan också på eget initiativ behandla frågor som rör den rättsliga grunden för förslag som kommissionen lagt fram.
I sådana fall ska ansvarigt utskott underrättas.
4.
Om utskottet med behörighet i rättsliga frågor anser att den rättsliga grunden är inkorrekt eller olämplig, ska det underrätta parlamentet om sina slutsatser.
Parlamentet ska rösta om dessa slutsatser innan det röstar om innehållet i förslaget.
5.
Ändringsförslag som läggs fram i parlamentet i syfte att ändra den rättsliga grunden för en av kommissionen föreslagen rättsakt är tillåtliga endast om ansvarigt utskott eller utskottet med behörighet i rättsliga frågor anser att den rättsliga grunden är inkorrekt eller olämplig.
6.
Om kommissionen inte är villig att ändra sitt förslag i överensstämmelse med den rättsliga grund som parlamentet har godkänt, kan föredraganden eller ordföranden i utskottet med behörighet i rättsliga frågor eller i det ansvariga utskottet föreslå att omröstningen om innehållet i förslaget ska skjutas upp till ett senare sammanträde.
Artikel
36
Prövning av ekonomisk förenlighet
1.
Utan att det påverkar tillämpningen av artikel 40 ska ansvarigt utskott i samband med alla kommissionsförslag och alla övriga handlingar som avser lagstiftning pröva om en rättsakts finansiering är förenlig med budgetplanen.
2.
Om ansvarigt utskott ändrar några uppgifter i anslagstilldelningen i den berörda rättsakten ska utskottet begära att utskottet med behörighet i budgetfrågor yttrar sig.
3.
Utskottet med behörighet i budgetfrågor kan även på eget initiativ studera den ekonomiska förenligheten i ett förslag som kommissionen lagt fram.
I så fall ska behörigt utskott underrättas.
4.
Om utskottet med behörighet i budgetfrågor anser att förslaget inte är ekonomiskt förenligt, ska utskottet översända sina slutsatser till parlamentet som ska låta dessa gå till omröstning.
5.
Parlamentet får med budgetmyndighetens medgivande anta en rättsakt som förklarats oförenlig.
Artikel
37
Parlamentets tillgång till handlingar och information till parlamentet
1.
Genom hela lagstiftningsförfarandet ska parlamentet och dess utskott begära att på samma villkor som rådet och dess arbetsgrupper få tillgång till alla handlingar som rör kommissionsförslag.
2.
Vid beredning av ett kommissionsförslag ska ansvarigt utskott uppmana kommissionen och rådet att hålla utskottet underrättat om hur arbetet med detta förslag fortskrider i rådet och rådets arbetsgrupper, i synnerhet när det gäller kompromisser som i väsentlig grad ändrar kommissionens ursprungliga förslag, eller meddela om kommissionen har för avsikt att dra tillbaka förslaget.
Artikel
38
Parlamentets företrädare vid rådsmöten
När rådet inbjuder parlamentet att delta vid ett rådsmöte där rådet handlar i sin egenskap av lagstiftare, ska talmannen uppdra åt ordföranden för det ansvariga utskottet, föredraganden eller någon annan ledamot som utsetts av det ansvariga utskottet att företräda parlamentet.
Artikel
38 a
Parlamentets initiativrätt enligt fördragen
I fall där fördragen ger parlamentet initiativrätt får det ansvariga utskottet besluta att utarbeta ett initiativbetänkande.
Betänkandet ska innehålla följande:
a)
Ett resolutionsförslag.
b)
När det är lämpligt ett förslag till beslut eller ett utkast till förslag.
c)
En motivering inklusive när det är lämpligt en finansieringsöversikt.
Om parlamentets antagande av en rättsakt kräver godkännande eller samtycke från rådet och yttrande eller samtycke från kommissionen får parlamentet, efter omröstningen om den föreslagna rättsakten och på förslag från föredraganden, besluta att skjuta upp omröstningen om resolutionsförslaget fram till det att rådet eller kommissionen har framfört sin ståndpunkt.
Artikel
39
Initiativ enligt artikel 192 i EG-fördraget
1.
Resolutionen ska antas av en majoritet av parlamentets samtliga ledamöter.
Parlamentet kan samtidigt fastställa en frist för att lägga fram ett sådant förslag.
2.
Parlamentets resolutioner ska ange den relevanta rättsliga grunden och omfatta detaljerade rekommendationer angående innehållet i förslaget i fråga, vilket ska respektera de grundläggande rättigheterna och subsidiaritetsprincipen.
3.
Om ett förslag har ekonomiska konsekvenser, ska parlamentet ange hur tillräcklig ekonomisk täckning kan garanteras.
4.
Ansvarigt utskott ska följa utvecklingen när det gäller varje förslag till rättsakt som utarbetas till följd av en särskild uppmaning från parlamentet.
Artikel
40
Beredning av lagstiftningsdokument
1.
Kommissionens förslag och andra dokument som avser lagstiftning ska av talmannen hänvisas till behörigt utskott för beredning.
När ett förslag är upptaget i lagstiftningsprogrammet, kan ansvarigt utskott besluta att utse en föredragande som ska följa utarbetandet av förslaget.
När rådet eller kommissionen begär att parlamentet ska yttra sig, ska talmannen vidarebefordra denna begäran till det utskott som ansvarar för beredningen av förslaget i fråga.
Bestämmelserna om första behandlingen i artiklarna 34-37, 49-56 och 66 ska tillämpas på lagstiftningsförslag, oavsett om det krävs en, två eller tre behandlingar.
2.
Rådets gemensamma ståndpunkter ska hänvisas för beredning till det utskott som var ansvarigt vid första behandlingen.
Bestämmelserna om andra behandlingen i artiklarna 57-62 och 67 ska tillämpas på gemensamma ståndpunkter.
3.
Under det förlikningsförfarande mellan parlamentet och rådet som följer på andra behandlingen får ingen återförvisning till utskott äga rum.
Bestämmelserna om tredje behandlingen i artiklarna 63, 64 och 65 ska tillämpas vid förlikningsförfarandet.
4.
5.
Om en bestämmelse i arbetsordningen som rör andra och tredje behandlingen strider mot någon annan bestämmelse i arbetsordningen, ska de bestämmelser som rör andra och tredje behandlingen ha företräde.
Artikel
41
Samråd om initiativ som läggs fram av en medlemsstat
1.
2.
Ansvarigt utskott kan inbjuda en företrädare för den medlemsstat som lagt fram initiativet till utskottet för att redogöra för initiativet.
Företrädaren för medlemsstaten kan åtföljas av företrädare för rådets ordförandeskap.
3.
Innan ansvarigt utskott påbörjar sin omröstning, ska utskottet fråga kommissionen om den har förberett en ståndpunkt om initiativet och om så är fallet uppmana kommissionen att tillkännage ståndpunkten inför det ansvariga utskottet.
4.
Om parlamentet samtidigt eller inom en kort tidsperiod föreläggs två eller flera förslag, med samma lagstiftningssyfte, från kommissionen och/eller medlemsstaterna, ska parlamentet behandla dessa i ett enda betänkande.
Ansvarigt utskott ska i betänkandet ange till vilken text det föreslår ändringar och i lagstiftningsresolutionen hänvisa till de övriga texterna.
5.
KAPITEL
2
FÖRFARANDEN I UTSKOTTEN
Artikel
42
Betänkanden som avser lagstiftning
1.
Ordföranden för det utskott till vilket ett kommissionsförslag har hänvisats ska föreslå utskottet vilket förfarande som ska tillämpas.
2.
Efter ett beslut om vilket förfarande som ska tillämpas, och om artikel 43 inte ska tillämpas, ska utskottet bland sina ledamöter eller ständiga suppleanter utse en föredragande för kommissionens förslag, om detta inte redan har skett på grundval av det lagstiftningsprogram som avses i artikel 33.
3.
Utskottets betänkande ska omfatta följande delar:
a)
b)
c)
Vid behov en motivering, inklusive en finansieringsöversikt som anger omfattningen av betänkandets eventuella ekonomiska konsekvenser och överensstämmelsen med budgetplanen.
Artikel
43
Förenklat förfarande
1.
Efter en första diskussion om ett förslag till rättsakt får utskottsordföranden föreslå att förslaget godkänns utan ändringsförslag.
2.
Ordföranden kan i stället föreslå att ordföranden själv eller föredraganden utarbetar ett antal ändringsförslag som återger diskussionen i utskottet.
Om utskottet går med på detta, ska dessa ändringsförslag sändas till utskottets ledamöter.
Betänkandet ska anses ha blivit antaget i utskottet såvida inte minst en tiondel av utskottets ledamöter har framfört invändningar före en fastställd tidpunkt, som inte får infalla tidigare än 21 dagar efter det att förslaget sänts ut.
3.
Om minst en tiondel av ledamöterna framför invändningar ska ändringsförslagen tas upp till omröstning vid nästföljande utskottssammanträde.
4.
Första och andra meningen i punkt 1, första, andra och tredje meningen i punkt 2 samt punkt 3 ska också gälla i tillämpliga delar på utskottsyttranden i den mening som avses i artikel 46.
Artikel
44
Betänkanden som inte avser lagstiftning
1.
Utarbetar ett utskott ett betänkande som inte avser lagstiftning, ska det bland sina ledamöter eller ständiga suppleanter utse en föredragande.
2.
Utskottets föredragande är ansvarig för utarbetandet av utskottets betänkande och för att detta på utskottets vägnar läggs fram i kammaren.
3.
Utskottets betänkande ska omfatta följande delar:
a)
Ett resolutionsförslag.
b)
En motivering, inklusive en finansieringsöversikt som anger omfattningen av betänkandets eventuella ekonomiska konsekvenser och överensstämmelsen med budgetplanen.
c)
Artikel
45
Initiativbetänkanden
1.
Ett eventuellt avslag på en sådan begäran ska alltid åtföljas av en motivering.
Talmanskonferensen ska fatta beslut om en begäran om tillstånd att utarbeta ett betänkande enligt punkt 1 på grundval av bestämmelser som talmanskonferensen själv fastställer.
Om ett utskotts befogenhet att utarbeta ett betänkande för vilket tillstånd har begärts ifrågasätts, ska talmanskonferensen inom sex veckor fatta ett beslut på grundval av en rekommendation från utskottsordförandekonferensen, eller, om ingen sådan rekommendation föreligger, från utskottsordförandekonferensens ordförande.
Om inget beslut har fattats av talmanskonferensen inom denna period, ska rekommendationen anses ha blivit godkänd.
2.
Resolutionsförslag i initiativbetänkanden ska behandlas av parlamentet i enlighet med det förfarande för kortfattad redogörelse som fastställs i artikel 131a.
Se talmanskonferensens relevanta beslut, som återges i bilaga ... till arbetsordningen.
.
3.
Om ämnet för betänkandet omfattas av den initiativrätt som avses i artikel 38a får medgivande vägras endast om villkoren i fördragen inte är uppfyllda.
4.
I de fall som avses i artiklarna 38a och 39 ska talmanskonferensen fatta ett beslut inom två månader.
Artikel
46
Utskottsyttranden
1.
2.
Föredraganden ska ansvara för motiveringarna, vilka inte ska gå till omröstning.
Om det behövs kan det rådgivande utskottet lämna in en kortfattad skriftlig motivering som omfattar hela yttrandet.
När det rör sig om texter som inte avser lagstiftning ska yttrandet innehålla förslag till delar av det ansvariga utskottets resolutionsförslag.
Det ansvariga utskottet ska rösta om dessa ändringsförslag eller förslag till nya punkter.
Yttrandet ska enbart omfatta sådana frågor som faller inom det rådgivande utskottets behörighetsområde.
3.
Det ansvariga utskottet ska fastställa när det rådgivande utskottet måste avge sina yttranden för att det ansvariga utskottet ska kunna ta hänsyn till dem.
Det ansvariga utskottet ska omedelbart meddela rådgivande utskott alla ändringar av denna frist.
Ansvarigt utskott ska inte fatta beslut innan tidsfristen har löpt ut.
4.
Alla antagna yttranden ska återges i det ansvariga utskottets betänkande.
5.
Endast det ansvariga utskottet har rätt att lägga fram ändringsförslag i kammaren.
6.
Ordföranden och föredraganden i det rådgivande utskottet ska inbjudas att i en rådgivande roll delta i det ansvariga utskottets sammanträden om det rör sig om ett ärende av gemensamt intresse.
Artikel
47
Förfarande med associerade utskott
-
De berörda utskotten ska gemensamt komma överens om tidsplanen.
-
Föredraganden och föredragandena av yttrande ska hålla varandra underrättade och sträva efter att komma överens om den text de lägger fram för sina respektive utskott och hur de ställer sig till eventuella ändringsförslag.
-
De ordförande, den föredragande och de föredragande av yttrande som berörs ska sträva efter att tillsammans fastställa vilka delar av texten som faller inom respektive utskotts exklusiva behörighetsområde och vilka delar av texten som faller inom ett gemensamt behörighetsområde samt komma överens om hur samarbetet dem emellan ska bedrivas.
-
Det ansvariga utskottet ska utan omröstning godta ändringsförslag från ett associerat utskott om förslagen rör frågor som det ansvariga utskottets ordförande, på grundval av bilaga VI och efter samråd med det associerade utskottets ordförande, anser falla inom det associerade utskottets exklusiva behörighetsområde, och som inte strider mot andra delar av betänkandet.
Det ansvariga utskottets ordförande ska ta hänsyn till alla eventuella överenskommelser som uppnåtts i enlighet med den tredje strecksatsen.
-
Om ett förlikningsförfarande inleds om förslaget ska de associerade utskottens föredragande ingå i parlamentets delegation.
I denna artikel föreskrivs ingen begränsning av tillämpningsområdet.
Artikel
48
Utarbetande av betänkanden
2.
I betänkandet ska resultatet från omröstningen om betänkandet i sin helhet anges.
3.
Denna ska anmälas i samband med omröstningen om hela texten och kan på författarnas begäran utgöra en skriftlig reservation på högst 200 ord, som fogas som bilaga till motiveringen.
Utskottsordföranden ska avgöra alla tvister som kan uppkomma till följd av dessa bestämmelser.
4.
Ett utskott kan på förslag av sitt presidium fastställa en tidsfrist för när utskottets föredragande ska lägga fram sitt förslag till betänkande.
Tidsfristen kan förlängas, och en ny föredragande kan även utses.
5.
Debatter kan i så fall äga rum på grundval av en muntlig rapport från utskottet i fråga.
KAPITEL
3
FÖRSTA BEHANDLINGEN
I utskotten
Artikel
49
Ändring av kommissionsförslag
1.
Om kommissionen underrättar parlamentet om att kommissionen har för avsikt att ändra sitt förslag, eller om ansvarigt utskott på annat sätt får kännedom om detta, ska detta utskott skjuta upp sin beredning av ärendet till dess att utskottet har mottagit det nya förslaget eller kommissionens ändringar.
2.
Om rådet väsentligt ändrar kommissionens förslag, ska bestämmelserna i artikel 55 tillämpas.
Artikel
50
Kommissionens och rådets ståndpunkt vid ändringsförslag
1.
Innan ansvarigt utskott övergår till slutomröstningen om ett kommissionsförslag, ska kommissionen uppmanas att tillkännage sin ståndpunkt angående alla de ändringsförslag till kommissionens förslag som utskottet antagit, och rådet ska uppmanas att ge en kommentar.
2.
Utskottet kan skjuta upp slutomröstning om kommissionen inte har möjlighet att tillkännage sin ståndpunkt, eller om kommissionen förklarar att den inte är beredd att godta alla de ändringsförslag som utskottet antagit.
3.
Kommissionens ståndpunkt ska vid behov ingå i betänkandet.
I kammaren
Artikel
51
Avslutande av första behandlingen
1.
Parlamentet ska behandla ett förslag till rättsakt på grundval av ett betänkande som ansvarigt utskott utarbetat i enlighet med artikel 42.
2.
Samrådsförfarandet är avslutat om förslaget till lagstiftningsresolution antas.
Om parlamentet inte antar lagstiftningsresolutionen, ska förslaget återförvisas till det ansvariga utskottet.
Alla betänkanden som läggs fram i enlighet med lagstiftningsförfarandet måste följa bestämmelserna i artiklarna 35, 40 och 42.
Alla resolutionsförslag som ett utskott lägger fram, och som inte avser lagstiftning, måste följa de särskilda förfaranden som anges i artikel 45 eller 179.
3.
Förslaget, så som det godkänts av parlamentet, och tillhörande resolution ska av talmannen såsom parlamentets yttrande översändas till rådet och kommissionen.
Artikel
52
Förkastande av kommissionsförslag
1.
Om ett kommissionsförslag inte får en majoritet av de avgivna rösterna ska talmannen, innan parlamentet röstar om förslaget till lagstiftningsresolution, uppmana kommissionen att dra tillbaka förslaget.
2.
Drar kommissionen tillbaka sitt förslag, ska talmannen fastslå att samrådsförfarandet är överflödigt och underrätta rådet om detta.
3.
Drar kommissionen inte tillbaka sitt förslag, ska parlamentet återförvisa frågan till ansvarigt utskott utan att rösta om förslaget till lagstiftningsresolution.
I sådana fall ska ansvarigt utskott, muntligen eller skriftligen, rapportera till parlamentet före utgången av en av parlamentet fastställd tidsfrist som inte får överstiga två månader.
4.
Artikel
53
Antagande av ändringar till ett kommissionsförslag
1.
Godkänns kommissionens förslag i sin helhet, men med antagna ändringar, ska omröstningen om förslaget till lagstiftningsresolution skjutas upp till dess att kommissionen redogjort för sin ståndpunkt beträffande var och en av parlamentets ändringar.
Om kommissionen vid avslutandet av parlamentets omröstning om kommissionens förslag inte har möjlighet att lämna en sådan redogörelse, ska kommissionen meddela talmannen eller ansvarigt utskott när den kommer att kunna göra detta.
2.
Meddelar kommissionen att den inte har för avsikt att godta alla parlamentets ändringar, ska ansvarigt utskotts föredragande eller, om föredraganden inte är närvarande, utskottets ordförande lägga fram ett formellt förslag till parlamentet om huruvida förslaget till lagstiftningsresolution ska gå till omröstning.
Utskottets föredragande eller ordförande kan före framläggandet av det formella förslaget uppmana talmannen att avbryta ärendets behandling.
Beslutar parlamentet att skjuta upp omröstningen, ska ärendet anses återförvisat till ansvarigt utskott för ytterligare beredning.
Endast ändringsförslag som ingivits av ansvarigt utskott, och som syftar till att få till stånd en kompromiss med kommissionen, ska tillåtas i detta skede.
3.
Vad som sägs i punkt 2 utesluter inte att andra ledamöter kan begära återförvisning i enlighet med artikel 168.
Om ett ärende återförvisas i enlighet med punkt 2, är ansvarigt utskott i enlighet med vad som fastställs vid återförvisningen skyldigt att lägga fram ett nytt betänkande före utgången av den fastställda tidsfristen.
Eftersom endast kompromissändringsförslag från utskottet är tillåtliga och för att kammarens suveränitet ska bevaras, måste det i sådana fall i det betänkande som avses i punkt 2 klart och tydligt framgå vilka redan godkända delar av förslaget som bortfaller om ändringsförslagen antas.
Uppföljning
Artikel
54
Uppföljning av parlamentets yttranden
1.
När parlamentet har yttrat sig om ett kommissionsförslag, ska ansvarigt utskotts ordförande och föredragande följa hur arbetet med förslaget fortskrider till dess att det har antagits av rådet, särskilt för att försäkra sig om att rådets och kommissionen verkligen respekterar sina åtaganden gentemot parlamentet när det gäller parlamentets ändringar.
2.
Ansvarigt utskott kan bjuda in kommissionen och rådet för att diskutera ärendet med utskottet.
3.
Ansvarigt utskott kan enligt denna artikel, om det anser det nödvändigt, när som helst under uppföljningsförfarandet lägga fram ett resolutionsförslag i vilket det rekommenderas att parlamentet
-
uppmanar kommissionen att dra tillbaka sitt förslag,
-
uppmanar kommissionen eller rådet att på nytt höra parlamentet i enlighet med artikel 55 eller uppmana kommissionen att lägga fram ett nytt förslag,
-
beslutar att vidta andra åtgärder som det finner lämpligt.
Detta förslag ska tas upp på förslaget till föredragningslista till den sammanträdesperiod som följer på utskottets beslut.
Artikel
55
Framläggande av ett nytt förslag för parlamentet
Medbeslutandeförfarandet
1.
Talmannen ska på begäran av ansvarigt utskott uppmana kommissionen att på nytt höra parlamentet om kommissionens förslag
-
om kommissionen, efter det att parlamentet har antagit sin ståndpunkt, drar tillbaka sitt ursprungliga förslag för att ersätta det, såvida detta inte sker i syfte att föra in parlamentets ändringar,
-
om kommissionen väsentligt ändrar eller har för avsikt att ändra sitt ursprungliga förslag, såvida detta inte sker i syfte att föra in parlamentets ändringar,
-
om problemställningen som förslaget avser väsentligt har förändrats på grund av tidens gång eller ändrade förhållanden,
-
om ett nytt val till parlamentet har ägt rum sedan parlamentet antog sin ståndpunkt och om talmanskonferensen anser att så är önskvärt.
2.
Parlamentet ska på ansvarigt utskotts begäran uppmana rådet att på nytt höra parlamentet om ett förslag som kommissionen lagt fram i enlighet med artikel 251 i EG-fördraget, om rådet har för avsikt att ändra förslagets rättsliga grund och det får till följd att förfarandet i artikel 251 i EG-fördraget inte längre är tillämpligt.
Andra förfaranden
3.
På begäran av ansvarigt utskott ska talmannen uppmana rådet att höra parlamentet på nytt under samma förutsättningar och på samma villkor som anges i punkt 1, och dessutom om rådet väsentligen ändrar eller har för avsikt att avsevärt ändra det ursprungliga förslag som parlamentet har yttrat sig över, såvida detta inte sker i syfte att föra in parlamentets ändringar.
4.
Talmannen ska även begära att parlamentet hörs på nytt om ett förslag till rättsakt under de förutsättningar som fastställs i denna artikel, om parlamentet så beslutar på förslag av en politisk grupp eller minst 40 ledamöter.
Artikel
56
Medlingsförfarandet enligt den gemensamma förklaringen från 1975
1.
När rådet i samband med vissa viktiga gemenskapsrättsakter har för avsikt att avvika från parlamentets yttrande, kan parlamentet med aktivt deltagande från kommissionen inleda ett medlingsförfarande med rådet i samband med att parlamentet avger sitt yttrande.
2.
Detta förfarande ska inledas av parlamentet antingen på eget eller på rådets initiativ.
3.
Vid sammansättningen av delegationen till medlingskommittén och när det gäller hur kommittén ska arbeta och meddela parlamentet sina resultat ska bestämmelserna i artikel 64 tillämpas.
4.
Ansvarigt utskott ska meddela resultatet av medlingen i ett betänkande.
Detta betänkande ska vara föremål för debatt och omröstning i kammaren.
KAPITEL
4
ANDRA BEHANDLINGEN
I utskotten
Artikel
57
Mottagande av rådets gemensamma ståndpunkt
1.
Parlamentet ska anses ha blivit delgiven rådets gemensamma ståndpunkt i enlighet med artiklarna 251 och 252 i EG-fördraget när talmannen tillkännager mottagandet i kammaren.
Talmannen ska tillkännage detta efter att ha mottagit de handlingar som innehåller den gemensamma ståndpunkten, alla förklaringar som fogats till rådets protokoll när det antog den gemensamma ståndpunkten, skälen till antagandet av denna samt kommissionens ståndpunkt, allt vederbörligen översatt till Europeiska unionens officiella språk.
Detta tillkännagivande ska göras vid den sammanträdesperiod som följer på mottagandet av dessa handlingar.
Före tillkännagivandet, men efter att ha hört ansvarigt utskotts ordförande och/eller föredragande, ska talmannen fastställa att den mottagna texten verkligen är en gemensam ståndpunkt och att sådana omständigheter som avses i artikel 55 inte föreligger.
Om detta inte kan fastställas ska talmannen tillsammans med ansvarigt utskott och om möjligt i samförstånd med rådet försöka hitta en lämplig lösning.
2.
En förteckning över sådana delgivna handlingar ska tillsammans med namnet på ansvarigt utskott offentliggöras i sammanträdesprotokollet.
Artikel
58
Förlängning av tidsfrister
1.
2.
3.
Artikel
59
Hänvisning till och förfarande i ansvarigt utskott
1.
2.
Den gemensamma ståndpunkten ska tas upp som första punkt på föredragningslistan till ansvarigt utskotts första sammanträde efter tidpunkten för mottagandet.
Rådet kan uppmanas att redogöra för den gemensamma ståndpunkten.
3.
Beslutas inte annorlunda ska föredraganden vid andra behandlingen vara densamme som vid första behandlingen.
4.
Endast detta utskotts ledamöter eller ständiga suppleanter har rätt att lägga fram förslag om avvisning eller ändringsförslag.
Utskottets beslut ska fattas med en majoritet av de avgivna rösterna.
5.
Utskottet kan före omröstningen begära att utskottsordföranden och föredraganden tillsammans med rådets ordförande eller företrädaren för rådets ordförande och i närvaro av ansvarig kommissionsledamot diskuterar ändringsförslag som lagts fram i utskottet.
Föredraganden kan lägga fram kompromissändringsförslag till följd av en sådan diskussion.
6.
Ansvarigt utskott ska avge en andrabehandlingsrekommendation där det föreslås att rådets gemensamma ståndpunkt godkänns, ändras eller avvisas.
Rekommendationen ska innehålla en kort motivering till föreslaget beslut.
I kammaren
Artikel
60
Avslutande av andra behandlingen
1.
Rådets gemensamma ståndpunkt, och i förekommande fall ansvarigt utskotts andrabehandlingsrekommendation, ska utan föregående beslut tas upp på förslaget till föredragningslista till den sammanträdesperiod vars onsdag infaller närmast före utgången av tidsfristen på tre eller, om denna förlängts i enlighet med artikel 58, fyra månader, såvida inte ärendet har behandlats vid en tidigare sammanträdesperiod.
Utskottens andrabehandlingsrekommendationer är likvärdiga med en motivering i vilken utskottet redogör för sin ståndpunkt i förhållande till rådets gemensamma ståndpunkt.
Andrabehandlingsrekommendationer ska därför inte gå till omröstning.
2.
Andra behandlingen avslutas när parlamentet, inom de tidsfrister och i enlighet med de villkor som fastställs i artiklarna 251 och 252 i EG-fördraget, godkänner, avvisar eller ändrar den gemensamma ståndpunkten.
Artikel
61
Avvisning av rådets gemensamma ståndpunkt
1.
Ansvarigt utskott, en politisk grupp eller minst 40 ledamöter kan skriftligen och före utgången av en av talmannen fastställd tidsfrist lägga fram ett förslag om avvisning av rådets gemensamma ståndpunkt.
För att ett sådant förslag ska antas krävs en majoritet av parlamentets samtliga ledamöter.
Omröstningen om förslag till avvisning av rådets gemensamma ståndpunkt ska äga rum före omröstningen om eventuella ändringsförslag.
2.
3.
Avvisas rådets gemensamma ståndpunkt ska talmannen tillkännage i kammaren att lagstiftningsförfarandet är avslutat.
4.
Med avvikelse från punkt 3 ska talmannen uppmana kommissionen att dra tillbaka sitt förslag om parlamentets avvisning omfattas av bestämmelserna i artikel 252 i EG-fördraget.
Drar kommissionen tillbaka sitt förslag ska talmannen tillkännage i kammaren att lagstiftningsförfarandet är avslutat.
Artikel
62
Ändringsförslag till rådets gemensamma ståndpunkt
1.
Ansvarigt utskott, en politisk grupp eller minst 40 ledamöter har rätt att inge ändringsförslag till rådets gemensamma ståndpunkt för behandling i kammaren.
2.
Ett ändringsförslag till den gemensamma ståndpunkten är tillåtligt endast om det är förenligt med bestämmelserna i artiklarna 150 och 151 samt om det syftar till att
a)
helt eller delvis återinföra den ståndpunkt som parlamentet intog vid första behandlingen,
b)
nå en kompromiss mellan rådet och parlamentet,
c)
ändra sådana delar av den gemensamma ståndpunkten som inte ingick i eller som innehållsmässigt skiljer sig från det vid första behandlingen framlagda förslaget, och som inte medför en väsentlig förändring av förslaget enligt vad som avses i artikel 55,
d)
beakta ett faktum eller ett nytt rättsligt läge som uppstått sedan första behandlingen.
Talmannens beslut om huruvida ett ändringsförslag är tillåtligt eller otillåtligt kan inte överklagas.
3.
Om ett nytt val har ägt rum sedan första behandlingen och artikel 55 inte har åberopats kan talmannen besluta att göra undantag från begränsningarna beträffande tillåtlighet i punkt 2.
4.
Ett ändringsförslag kan antas endast om det får en majoritet av rösterna från parlamentets samtliga ledamöter.
5.
Innan ändringsförslagen går till omröstning kan talmannen uppmana kommissionen att tillkännage sin ståndpunkt och rådet att ge en kommentar.
KAPITEL
5
TREDJE BEHANDLINGEN
Förlikning
Artikel
63
Sammankallande av förlikningskommittén
Om rådet meddelar parlamentet att det inte kan godkänna alla parlamentets ändringar i den gemensamma ståndpunkten ska talmannen tillsammans med rådet komma överens om tid och plats för ett första sammanträde i förlikningskommittén.
Artikel
64
Delegationen till förlikningskommittén
1.
Parlamentets delegation till förlikningskommittén ska bestå av samma antal ledamöter som rådets delegation.
2.
Delegationens politiska sammansättning ska motsvara parlamentets sammansättning av politiska grupper.
Talmanskonferensen ska fastställa det exakta antalet ledamöter från varje politisk grupp.
3.
Med undantag av tre ledamöter som för en tid av tolv månader utses som ständiga ledamöter av olika delegationer, ska delegationens ledamöter utses av de politiska grupperna för varje enskild förlikning, företrädesvis bland de berörda utskottens ledamöter.
De tre ständiga ledamöterna ska utses av de politiska grupperna bland de vice talmännen och ska företräda minst två olika politiska grupper.
Ansvarigt utskotts ordförande och föredragande ska alltid ingå i delegationen.
4.
De i delegationen företrädda grupperna ska utse suppleanter.
5.
Politiska grupper och grupplösa som inte är företrädda i delegationen har rätt att sända var sin företrädare till alla delegationens interna förberedande sammanträden.
6.
Delegationen leds av talmannen eller en av de tre ständiga ledamöterna.
7.
Delegationen ska fatta beslut med en majoritet av sina ledamöter.
Delegationens överläggningar är inte offentliga.
Talmanskonferensen får fastställa ytterligare procedurregler för arbetet i delegationen till förlikningskommittén.
8.
Delegationen ska meddela parlamentet resultatet av förlikningen.
I kammaren
Artikel
65
Gemensamt utkast
1.
Uppnås enighet i förlikningskommittén om ett gemensamt utkast ska ärendet tas upp på föredragningslistan i så god tid att det kan behandlas i kammaren inom sex eller, vid en förlängning av tidsfristen, åtta veckor från dagen för förlikningskommitténs godkännande av det gemensamma utkastet.
2.
Ordföranden eller någon annan utsedd medlem av parlamentets delegation till förlikningskommittén ska göra ett uttalande om det gemensamma utkastet vilket ska åtföljas av ett betänkande.
3.
Inga ändringsförslag får läggas fram till det gemensamma utkastet.
4.
Det gemensamma utkastet i sin helhet ska vara föremål för en enda omröstning.
Det gemensamma utkastet godkänns om det får en majoritet av de avgivna rösterna.
5.
Uppnås ingen enighet om ett gemensamt utkast i förlikningskommittén, ska ordföranden eller någon annan utsedd medlem av parlamentets delegation till förlikningskommittén göra ett uttalande.
Detta uttalande ska följas av en debatt.
KAPITEL
6
LAGSTIFTNINGSFÖRFARANDET - AVSLUTANDE
Artikel
66
Överenskommelse vid första behandlingen
1.
2.
Före detta tillkännagivande ska talmannen kontrollera att inga tekniska förändringar av förslaget som rådet gjort påverkar innehållet i förslaget.
I tveksamma fall ska talmannen samråda med ansvarigt utskott.
Om de ändringar som gjorts anses påverka innehållet, ska talmannen underrätta rådet om att parlamentet kommer att gå vidare med en andra behandling så snart villkoren i artikel 57 har uppfyllts.
3.
Efter tillkännagivandet i punkt 1 ska talmannen tillsammans med rådets ordförande underteckna den föreslagna rättsakten och i enlighet med artikel 68 se till att den offentliggörs i Europeiska unionens officiella tidning.
Artikel
67
Överenskommelse vid andra behandlingen
Antas inte något förslag om avvisning av den gemensamma ståndpunkten eller något ändringsförslag enligt artiklarna 61 och 62 före utgången av tidsfristen för att inge och rösta om ändringsförslag eller förslag om avvisning, ska talmannen tillkännage i kammaren att den föreslagna rättsakten är slutgiltigt antagen.
Talmannen ska tillsammans med rådets ordförande underteckna den föreslagna rättsakten och i enlighet med artikel 68 se till att den offentliggörs i Europeiska unionens officiella tidning.
Artikel
68
Undertecknande av antagna rättsakter
1.
Texten till sådana rättsakter som antas av parlamentet och rådet ska undertecknas av talmannen och av generalsekreteraren efter att dessa har kontrollerat att alla förfaranden vederbörligen avslutats.
2.
I rättsakter som antas av parlamentet och rådet gemensamt inom ramen för förfarandet i artikel 251 i EG-fördraget ska anges vilken typ av rättsakt det rör sig om, ordningsnumret, dagen för dess antagande och en uppgift om innehållet.
3.
Rättsakter som antas av parlamentet och rådet gemensamt ska innehålla följande:
a)
Formuleringen "Europaparlamentet och Europeiska unionens råd".
b)
En uppgift om de bestämmelser på grundval av vilka rättsakten antas, föregången av orden "med beaktande av".
c)
En hänvisning till framlagda förslag, avgivna yttranden och hållna samråd.
d)
Skälen till rättsakten.
e)
En formulering såsom "härigenom föreskrivs följande" eller "har beslutat följande" följd av bestämmelserna i rättsakten.
4.
Rättsakter ska delas in i artiklar som får grupperas i kapitel och avsnitt.
5.
Sista artikeln i en rättsakt ska bestämma dagen för ikraftträdandet, om denna dag inträffar före eller efter den tjugonde dagen efter det att rättsakten offentliggjorts.
6.
Sista artikeln i en rättsakt ska följas av
-
en lämplig slutformulering, i enlighet med relevant artikel i fördraget, beträffande rättsaktens tillämplighet,
-
"Utfärdad i/Utfärdat i..." följt av dagen för antagandet av rättsakten,
-
formuleringen "På Europaparlamentets vägnar Ordförande", "På rådets vägnar Ordförande" med namnet på talmannen och namnet på ordföranden i rådet vid tidpunkten för antagandet av rättsakten infört före ordet "Ordförande".
7.
De rättsakter som avses ovan ska offentliggöras i Europeiska unionens officiella tidning på initiativ av parlamentets och rådets generalsekreterare.
KAPITEL
7
BUDGETFÖRFARANDEN
Artikel
69
Allmänna budgeten
Genomförandebestämmelser för granskning av Europeiska unionens allmänna budget och tilläggsbudgetar, i enlighet med de finansiella bestämmelserna i fördragen om upprättandet av Europeiska gemenskaperna, ska antas av parlamentet i form av en resolution och fogas som bilaga till arbetsordningen
Se bilaga IV.
.
Artikel
70
Ansvarsfrihet för kommissionen beträffande genomförandet av budgeten
Bestämmelser för beviljande av ansvarsfrihet för kommissionen beträffande genomförandet av budgeten, i enlighet med de finansiella bestämmelserna i fördragen om upprättandet av Europeiska gemenskaperna och budgetförordningen, ska fogas som bilaga till arbetsordningen
Se bilaga V.
.
Artikel
71
Andra förfaranden för beviljande av ansvarsfrihet
Bestämmelserna angående förfarandet för beviljande av ansvarsfrihet för kommissionen vad gäller genomförandet av budgeten gäller på motsvarande sätt för följande förfaranden:
-
Förfarandet för beviljande av ansvarsfrihet för Europaparlamentets talman vad gäller genomförandet av Europaparlamentets budget.
-
Förfarandet för beviljande av ansvarsfrihet för de personer som är ansvariga för genomförandet av budgetarna för Europeiska unionens övriga institutioner och organ, exempelvis rådet (i fråga om rådets verkställande verksamhet), EG-domstolen, revisionsrätten, Europeiska ekonomiska och sociala kommittén och Regionkommittén.
-
Förfarandet för beviljande av ansvarsfrihet för kommissionen vad gäller genomförandet av Europeiska utvecklingsfondens budget.
-
Förfarandet för beviljande av ansvarsfrihet för de organ som ansvarar för genomförandet av budgeten för juridiskt oberoende enheter vilka sköter uppgifter åt gemenskapen, i den mån de bestämmelser som reglerar deras verksamhet föreskriver att ansvarsfrihet ska beviljas av Europaparlamentet.
Artikel
72
Parlamentets kontroll över genomförandet av budgeten
1.
Parlamentet ska övervaka genomförandet av den löpande budgeten.
Parlamentet ska överlåta denna uppgift till utskotten med behörighet i frågor som rör budget och budgetkontroll samt övriga berörda utskott.
2.
Varje år ska parlamentet, före första behandlingen av budgetförslaget för det följande budgetåret, behandla problem i samband med genomförandet av den löpande budgeten, eventuellt på grundval av ett resolutionsförslag från behörigt utskott.
KAPITEL
8
INTERNA BUDGETFÖRFARANDEN
Artikel
73
Parlamentets budgetberäkning
1.
På grundval av en rapport från generalsekreteraren ska presidiet upprätta ett preliminärt förslag till budgetberäkning.
2.
Talmannen ska översända det preliminära förslaget till budgetberäkning till behörigt utskott, som ska utarbeta ett förslag till budgetberäkning och rapportera till parlamentet.
3.
Talmannen ska fastställa en tidsfrist för ingivande av ändringsförlag till förslaget till budgetberäkning.
Behörigt utskott ska yttra sig över dessa ändringsförslag.
4.
Parlamentet ska anta budgetberäkningen.
5.
Talmannen ska översända budgetberäkningen till kommissionen och rådet.
6.
Ovanstående bestämmelser ska även tillämpas vid tilläggsbudgetberäkningar.
7.
Genomförandebestämmelser för upprättandet av parlamentets budgetberäkning ska antas med en majoritet av de avgivna rösterna och fogas som bilaga till arbetsordningen
Se bilaga IV.
.
Artikel
74
Ekonomiska åtaganden och reglering av utgifter
1.
Talmannen ska göra de ekonomiska åtaganden och reglera de utgifter - eller se till att så sker - som omfattas av de interna finansbestämmelser som presidiet fastställt efter att ha hört behörigt utskott.
2.
Talmannen ska översända förslaget till avslutande av räkenskaperna till behörigt utskott.
3.
På grundval av ett betänkande från behörigt utskott ska parlamentet fastställa avslutandet av räkenskaperna och besluta om beviljande av ansvarsfrihet.
KAPITEL
9
SAMTYCKESFÖRFARANDET
Artikel
75
Samtyckesförfarandet
1.
När parlamentet uppmanas att ge sitt samtycke till ett förslag till rättsakt ska det fatta beslut med utgångspunkt i en rekommendation från det ansvariga utskottet om att godkänna eller förkasta rättsakten.
Den för samtycke nödvändiga majoriteten ska vara den majoritet som anges i den artikel i EG-fördraget eller EU-fördraget som utgör den rättsliga grunden för förslaget till rättsakt.
2.
Vid anslutningsfördrag och internationella avtal samt när det gäller att slå fast att en medlemsstat allvarligt och ihållande åsidosätter gemensamma principer ska artiklarna 82, 83 och 95 i arbetsordningen tillämpas.
Vid närmare samarbete på ett område som omfattas av det förfarande som fastställs i artikel 251 i EG-fördraget ska artikel 76 i denna arbetsordning tillämpas.
3.
När parlamentets samtycke krävs i samband med ett förslag till rättsakt kan ansvarigt utskott, för att förfarandet ska leda till ett positivt resultat, besluta att förelägga parlamentet ett interimsbetänkande om kommissionens förslag med ett resolutionsförslag som innehåller rekommendationer om ändring eller genomförande av förslaget till rättsakt.
Om parlamentet antar minst en rekommendation ska talmannen anhålla om ytterligare diskussioner med rådet.
Ansvarigt utskott ska lämna sin slutgiltiga rekommendation angående parlamentets samtycke på grundval av resultatet av diskussionerna med rådet.
KAPITEL
10
NÄRMARE SAMARBETE
Artikel
76
Förfaranden i parlamentet
1.
Artiklarna 35, 36, 37, 40, 49-56 och 75 i arbetsordningen ska tillämpas på lämpligt sätt.
2.
Behörigt utskott ska kontrollera om förslaget är förenligt med artikel 11 i EG-fördraget samt artiklarna 27a, 27b, 40, 43, 44 och 44a i EU-fördraget.
3.
Förslag till rättsakter som därefter läggs fram inom ramen för det närmare samarbetet, när detta väl upprättats, ska behandlas i parlamentet på samma sätt som när det inte förekommer något närmare samarbete.
KAPITEL
11
ÖVRIGA FÖRFARANDEN
Artikel
77
Yttranden i enlighet med artikel 122 i EG-fördraget
1.
2.
Artikel
78
Förfaranden som rör dialogen mellan arbetsmarknadens parter
1.
2.
3.
Artikel
79
Förfaranden för kontroll av frivilliga överenskommelser
1.
Om kommissionen meddelar parlamentet att den avser att undersöka möjligheten att som ett alternativ till lagstiftning använda sig av frivilliga överenskommelser, får det ansvariga utskottet utarbeta ett betänkande om själva sakfrågan i enlighet med artikel 45.
2.
När kommissionen uppger att den har för avsikt att ingå en frivillig överenskommelse, ska det ansvariga utskottet inge ett förslag till resolution som rekommenderar huruvida förslaget ska antas eller förkastas, och på vilka villkor.
Artikel
80
Kodifiering
1.
När ett kommissionsförslag om kodifiering av gemenskapslagstiftning föreläggs parlamentet, ska det hänvisas till utskottet med behörighet i rättsliga frågor.
Utskottet ska behandla förslaget i enlighet med de förfaranden som överenskommits på interinstitutionell nivå
2.
för att se till att förslaget inskränker sig till en enkel kodifiering som inte i sak ändrar innehållet.
2.
3.
Om utskottet med behörighet i rättsliga frågor anser att förslaget inte innebär någon ändring i sak av gemenskapslagstiftningen ska det förelägga parlamentet förslaget för godkännande.
Om utskottet anser att förslaget innebär en ändring i sak, ska det föreslå att parlamentet förkastar förslaget.
I båda dessa fall ska parlamentet fatta beslut genom en enkel omröstning utan vare sig ändringsförslag eller debatt.
Artikel
80 a
Omarbetning
1.
När ett kommissionsförslag om omarbetning av gemenskapslagstiftning föreläggs parlamentet, ska det hänvisas till utskottet med behörighet i rättsliga frågor och till det ansvariga utskottet.
2.
Utskottet med behörighet i rättsliga frågor ska behandla förslaget i enlighet med de förfaranden som överenskommits på interinstitutionell nivå
Interinstitutionellt avtal av den 28 november 2001 om en mer strukturerad användning av omarbetningstekniken för rättsakter, punkt 9 (EGT C 77, 28.3.2002, s.
1).
för att se till att förslaget inte innebär några andra ändringar i sak än dem som angivits som sådana.
3.
Om utskottet med behörighet i rättsliga frågor anser att förslaget inte innebär några andra ändringar i sak än dem som angivits som sådana, ska det informera det ansvariga utskottet om detta.
Det ansvariga utskottet kan i så fall bara behandla ändringsförslag om de berör de delar av förslaget som innehåller ändringar och uppfyller villkoren i artiklarna 150 och 151.
Ändringsförslag till de oförändrade delarna kan emellertid tillåtas undantagsvis och från fall till fall av ordföranden i det utskottet om han eller hon anser att detta är nödvändigt för att texten ska bli logisk eller för att det finns ett samband med andra tillåtliga ändringsförslag.
En skriftlig motivering som rättfärdigar dessa undantag ska upprättas för dessa ändringsförslag.
4.
Om utskottet med behörighet i rättsliga frågor anser att förslaget innebär andra ändringar i sak än dem som har angivits som sådana, ska det föreslå att parlamentet förkastar förslaget och underrätta det ansvariga utskottet om detta.
I detta fall ska talmannen uppmana kommissionen att dra tillbaka sitt förslag.
Om kommissionen drar tillbaka sitt förslag ska talmannen slå fast att förfarandet är överflödigt och underrätta rådet om detta.
Om kommissionen inte drar tillbaka sitt förslag ska parlamentet hänvisa det till det ansvariga utskottet, som ska ta upp det till förnyad behandling i enlighet med det gängse förfarandet.
Artikel
81
Genomförandeåtgärder
2.
Ordföranden för det ansvariga utskottet ska fastställa en tidsfrist inom vilken ledamöterna kan föreslå att utskottet motsätter sig förslaget till åtgärder.
Om utskottet finner det lämpligt kan det besluta att utse en föredragande bland sina ledamöter eller ständiga suppleanter.
3.
Om det inte hålls någon sammanträdesperiod före tidsfristens utgång ska rätten att svara anses ha delegerats till ansvarigt utskott.
Svaret ska vara i form av en skrivelse från utskottets ordförande till ansvarig kommissionsledamot.
Samtliga ledamöter ska informeras om detta.
4.
a)
I detta fall ska artikel 138 inte tillämpas.
b)
Parlamentet kan med en majoritet av sina ledamöter motsätta sig att ett förslag till åtgärder antas, samtidigt som det motiverar sina invändningar genom att ange att förslaget till åtgärder överskrider de genomförandebefogenheter som fastställs i den grundläggande rättsakten eller att utkastet inte är förenligt med syftet med eller innehållet i den grundläggande rättsakten eller att det inte respekterar subsidiaritets- eller proportionalitetsprincipen.
c)
KAPITEL
12
FÖRDRAG OCH INTERNATIONELLA AVTAL
Artikel
82
Anslutningsfördrag
1.
Varje ansökan från en europeisk stat om medlemskap i Europeiska unionen ska hänvisas till behörigt utskott för beredning.
2.
Parlamentet kan på förslag av behörigt utskott, en politisk grupp eller minst 40 ledamöter besluta att uppmana kommissionen och rådet att delta i en debatt innan förhandlingarna med den ansökande staten inleds.
3.
4.
Parlamentet har rätt att när som helst under förhandlingarna, på grundval av ett betänkande från ansvarigt utskott, anta rekommendationer och kräva att dessa beaktas innan ett fördrag om en ansökande stats anslutning till Europeiska unionen ingås.
För antagandet av sådana rekommendationer fordras samma majoritet som vid samtycke.
5.
När förhandlingarna slutförts, men innan något avtal undertecknas, ska förslaget till fördrag föreläggas parlamentet för samtycke.
6.
Parlamentet ska på grundval av ett betänkande från ansvarigt utskott och med en majoritet av samtliga sina ledamöter ge sitt samtycke till en ansökan från en europeisk stat om medlemskap i Europeiska unionen.
Artikel
83
Internationella avtal
1.
2.
Parlamentet kan på förslag av ansvarigt utskott, en politisk grupp eller minst 40 ledamöter uppmana rådet att inte tillåta att förhandlingar inleds förrän parlamentet, med ett betänkande från ansvarigt utskott som grund, har yttrat sig om det föreslagna förhandlingsmandatet.
3.
När avsikten är att inleda förhandlingar, ska ansvarigt utskott se till att kommissionen angett en rättslig grund för att ingå de internationella avtal som avses i punkt 1.
Ansvarigt utskott ska granska den valda rättsliga grunden i enlighet med artikel 35.
Om kommissionen inte har angett en rättslig grund eller om dess lämplighet kan ifrågasättas, ska artikel 35 tillämpas.
4.
5.
Parlamentet har rätt att när som helst under förhandlingarna, på grundval av ett betänkande från ansvarigt utskott och efter att ha prövat eventuella förslag som lagts fram i enlighet med artikel 114, anta rekommendationer och begära att dessa beaktas innan det internationella avtalet i fråga ingås.
6.
När förhandlingarna slutförts, men innan något avtal undertecknas, ska förslaget till avtal föreläggas parlamentet för yttrande eller samtycke.
När det gäller samtyckesförfarandet ska artikel 75 tillämpas.
7.
8.
Om parlamentet avstyrker, ska talmannen uppmana rådet att inte ingå avtalet i fråga.
9.
Om parlamentet med en majoritet av de avgivna rösterna inte ger sitt samtycke till ett internationellt avtal, ska talmannen meddela rådet att avtalet inte kan ingås.
Artikel
84
Förfaranden enligt artikel 300 i EG-fördraget när det gäller provisorisk tillämpning eller tillfälligt upphävande av internationella avtal eller fastställande av gemenskapens ståndpunkt i ett organ som inrättats genom ett internationellt avtal
Parlamentet kan utfärda rekommendationer i enlighet med artikel 83 eller 90 i arbetsordningen.
KAPITEL
13
UNIONENS EXTERNA REPRESENTATION OCH DEN GEMENSAMMA UTRIKES- OCH SÄKERHETSPOLITIKEN
Artikel
85
Utnämning av den höge representanten för den gemensamma utrikes- och säkerhetspolitiken
1.
Före utnämningen av den höge representanten för den gemensamma utrikes- och säkerhetspolitiken, ska talmannen uppmana rådets tjänstgörande ordförande att inför parlamentet göra ett uttalande i enlighet med artikel 21 i EU-fördraget.
Talmannen ska uppmana kommissionens ordförande att uttala sig vid samma tillfälle.
2.
3.
Uttalandet och svaren i punkterna 1 och 2 kan följas av rekommendationer från parlamentet på initiativ från behörigt utskott eller i enlighet med artikel 114.
Artikel
86
Utnämning av särskilda representanter inom ramen för den gemensamma utrikes- och säkerhetspolitiken
1.
2.
När den särskilde representanten har utsetts, men ännu inte tillträtt, kan han eller hon uppmanas att inför det behöriga utskottet göra ett uttalande och besvara frågor.
3.
Inom tre månader från utfrågningen kan utskottet föreslå en rekommendation enligt artikel 114 som direkt hänför sig till uttalandet och svaren.
4.
Den särskilde representanten ska uppmanas att utförligt och regelbundet hålla parlamentet informerat om det praktiska genomförandet av representantens mandat.
Artikel
87
Uttalanden av den höge representanten för den gemensamma utrikes- och säkerhetspolitiken och andra särskilda representanter
1.
Den höge representanten ska inbjudas att minst fyra gånger om året uttala sig i kammaren.
Artikel 103 ska tillämpas.
2.
Den höge representanten ska minst fyra gånger om året inbjudas att närvara vid det behöriga utskottets sammanträden för att där göra ett uttalande och besvara frågor.
Den höge representanten kan bjudas in vid andra tillfällen när utskottet anser det vara nödvändigt eller på representantens egen begäran.
3.
När en särskild representant med mandat för en särskild politisk fråga utses av rådet, ska han eller hon på parlamentets eller på eget initiativ inbjudas för att göra ett uttalande inför behörigt utskott.
Artikel
88
Internationell representation
2.
Artikel
89
Samråd med och underrättande av parlamentet inom ramen för den gemensamma utrikes- och säkerhetspolitiken
1.
2.
De berörda utskotten ska sträva efter att förmå den höge representanten för den gemensamma utrikes- och säkerhetspolitiken, rådet och kommissionen att förse dem med regelbunden och aktuell information om utvecklingen och genomförandet av den gemensamma utrikes- och säkerhetspolitiken, den beräknade kostnaden för varje beslut på detta område som har ekonomiska konsekvenser och om övriga finansiella aspekter som rör genomförandet av den gemensamma utrikes- och säkerhetspolitiken.
På begäran av kommissionen, rådet eller den höge representanten kan ett utskott i undantagsfall besluta att hålla sina sammanträden inom stängda dörrar.
3.
En gång om året ska det hållas en debatt om det samrådsdokument som rådet utarbetat om de viktigaste aspekterna och de grundläggande valmöjligheterna när det gäller den gemensamma utrikes- och säkerhetspolitiken, inbegripet konsekvenserna för unionens budget.
Förfarandet i artikel 103 ska tillämpas.
(Se även tolkningen till artikel 114.)
4.
Rådet och/eller den höge representanten och kommissionen ska inbjudas till alla plenardebatter som rör utrikes-, säkerhets- eller försvarspolitik.
Artikel
90
Rekommendationer inom ramen för den gemensamma utrikes- och säkerhetspolitiken
1.
Utskottet med behörighet i frågor som rör den gemensamma utrikes- och säkerhetspolitiken kan, efter att ha beviljats tillstånd av talmanskonferensen eller på grundval av ett förslag i enlighet med artikel 114, utarbeta rekommendationer till rådet inom sitt behörighetsområde.
2.
I brådskande fall kan det tillstånd som avses i punkt 1 beviljas av talmannen, som även kan ge utskottet tillstånd att hålla ett brådskande sammanträde.
3.
Undantaget beträffande tillämpningen av artikel 138 gäller endast utskott och i brådskande fall.
Bestämmelserna i artikel 138 ska tillämpas vid utskottssammanträden som inte har förklarats som brådskande och vid plenarsammanträden.
Bestämmelsen om att muntliga ändringsförslag får läggas fram innebär att ledamöter inte kan motsätta sig att muntliga ändringsförslag går till omröstning i utskottet.
4.
De på detta sätt utarbetade rekommendationerna ska föras upp på föredragningslistan till nästföljande sammanträdesperiod.
I brådskande fall, som fastställs av talmannen, kan rekommendationer föras upp på föredragningslistan till en pågående sammanträdesperiod.
Rekommendationer ska anses antagna om inte minst 40 ledamöter före sammanträdesperiodens början inger en skriftlig invändning.
I sådana fall ska var och en av utskottets rekommendationer föras upp på föredragningslistan för debatt och omröstning vid ett plenarsammanträde under denna sammanträdesperiod.
En politisk grupp eller minst 40 ledamöter kan inge ändringsförslag.
Artikel
91
Kränkningar av de mänskliga rättigheterna
KAPITEL
14
POLISSAMARBETE OCH STRAFFRÄTTSLIGT SAMARBETE
Artikel
92
Information till parlamentet när det gäller polissamarbete och straffrättsligt samarbete
1.
2.
På kommissionens eller rådets begäran kan ett utskott i undantagsfall besluta att hålla sina sammanträden inom stängda dörrar.
3.
Artikel
93
Samråd med parlamentet när det gäller polissamarbete och straffrättsligt samarbete
När parlamentet hörs om rådets förslag till beslut om utnämning av Europols direktör och styrelse ska artikel 101 i arbetsordningen gälla i tillämpliga delar.
Artikel
94
Rekommendationer när det gäller polissamarbete och straffrättsligt samarbete
1.
Utskottet med behörighet i frågor som rör polissamarbete och straffrättsligt samarbete kan, efter att ha inhämtat talmanskonferensens tillstånd eller på grundval av ett förslag i enlighet med artikel 114, utarbeta rekommendationer till rådet inom sitt behörighetsområde inom det område som faller inom avdelning VI i EU-fördraget.
2.
I brådskande fall kan det tillstånd som avses i punkt 1 beviljas av talmannen, som även kan bevilja utskottet tillstånd att hålla ett brådskande sammanträde.
3.
(Se även tolkningen till artikel 114.)
KAPITEL
15
EN MEDLEMSSTATS ÅSIDOSÄTTANDE AV GRUNDLÄGGANDE PRINCIPER
Artikel
95
Fastslående av åsidosättande
1.
Parlamentet kan, på grundval av ett särskilt betänkande från det ansvariga utskottet i enlighet med artikel 45,
a)
b)
c)
2.
Parlamentet ska fatta beslut på grundval av ett förslag från det ansvariga utskottet, utom i brådskande fall och om det finns goda skäl.
3.
Beslut i enlighet med punkterna 1 och 2 kräver två tredjedelars majoritet av de avgivna rösterna och en majoritet av parlamentets samtliga ledamöter.
4.
Behörigt utskott kan lägga fram ett kompletterande resolutionsförslag i de fall då parlamentet uppmanas att ge sitt samtycke i enlighet med punkt 2.
Ett sådant resolutionsförslag ska innehålla parlamentets synpunkter på en medlemsstats allvarliga åsidosättande på lämpliga åtgärder och på förutsättningarna för att ändra eller upphöra med dessa åtgärder.
5.
Behörigt utskott ska se till att parlamentet hålls fullständigt informerat och vid behov hörs om alla åtgärder som vidtas efter det att parlamentet gett sitt samtycke i enlighet med punkt 3.
Rådet ska uppmanas att informera om utvecklingen på lämpligt sätt.
På förslag av behörigt utskott, utarbetat med talmanskonferensens medgivande, kan parlamentet anta rekommendationer till rådet.
AVDELNING
III
ÖPPENHET OCH INSYN
Artikel
96
Insyn i parlamentets verksamhet
1.
2.
Parlamentets överläggningar ska vara offentliga.
3.
Parlamentets utskott ska normalt hålla offentliga sammanträden.
Om tystnadsplikten inte respekteras ska artikel 147 tillämpas.
4.
Behandlingen i behörigt utskott av begäran som berör förfarandet om upphävande av immunitet i enlighet med artikel 7 ska alltid äga rum inom stängda dörrar.
Artikel
97
Allmänhetens tillgång till handlingar
1.
Varje unionsmedborgare och varje fysisk eller juridisk person som är bosatt eller har sitt säte i en medlemsstat ska ha rätt till tillgång till parlamentets handlingar i enlighet med artikel 255 i EG-fördraget, med beaktande av de principer, villkor och gränser som fastställs i Europaparlamentets och rådets förordning (EG) nr 1049/2001 och i enlighet med de särskilda bestämmelser som ingår i arbetsordningen.
Andra fysiska och juridiska personer ska i den mån det är möjligt ha tillgång till parlamentets handlingar på samma sätt.
Förordning (EG) nr 1049/2001 ska offentliggöras för kännedom vid sidan om arbetsordningen.
2.
Handlingar som utarbetats av enskilda ledamöter eller politiska grupper ska i frågor som berör tillgången till handlingar anses som parlamentets handlingar, om de framlagts i enlighet med arbetsordningen.
Presidiet ska fastställa bestämmelser för att säkerställa att alla parlamentets handlingar registreras.
3.
Parlamentet ska inrätta ett register över parlamentets handlingar.
Lagstiftningshandlingar och andra handlingar som anges i en bilaga till arbetsordningen
Se bilaga XV.
ska göras direkt tillgängliga i enlighet med förordning (EG) nr 1049/2001 via parlamentets register.
Hänvisningar till andra av parlamentets handlingar ska i största möjliga utsträckning tas med i registret.
De handlingar som är direkt tillgängliga ska tas upp i en förteckning som ska godkännas av parlamentet och bifogas arbetsordningen
Se bilaga XV.
som bilaga.
Detta innebär inte att tillgången till handlingar av typer som inte finns med i förteckningen begränsas.
De av parlamentets handlingar som inte är direkt tillgängliga via registret ska tillhandahållas efter skriftlig begäran.
Presidiet kan anta bestämmelser, som är i överensstämmelse med förordning (EG) nr 1049/2001, om hur tillgången praktiskt ska organiseras, och som ska offentliggöras i Europeiska unionens officiella tidning.
4.
Presidiet ska fastställa vilka myndigheter som ska ansvara för behandling av ursprungliga ansökningar (artikel 7 i förordning (EG) nr 1049/2001) samt anta beslut om bekräftande ansökningar (artikel 8 i nämnda förordning) och ansökningar om känsliga handlingar (artikel 9 i nämnda förordning).
5.
6.
Tillsynen över hur ansökningar om tillgång till handlingar behandlas ska en av de vice talmännen vara ansvarig för.
7.
Ansvarigt parlamentsutskott ska, på grundval av upplysningar från presidiet och andra källor, utarbeta den årsrapport som avses i artikel 17 i förordning (EG) nr 1049/2001 och lägga fram den för kammaren.
Ansvarigt utskott ska också granska och utvärdera de rapporter som i enlighet med artikel 17 i nämnda förordning antas av andra institutioner och organ.
AVDELNING
IV
FÖRBINDELSER MED ANDRA ORGAN
KAPITEL
1
NOMINERINGAR OCH UTNÄMNINGAR
Artikel
98
Val av kommissionens ordförande
1.
När rådet har enats om nomineringen av en kandidat till ämbetet som kommissionens ordförande, ska talmannen uppmana kandidaten att göra ett uttalande och redogöra för sitt politiska program inför parlamentet.
Uttalandet ska följas av en debatt.
Rådet ska uppmanas att delta i debatten.
2.
Parlamentet ska godkänna eller avslå nomineringen med en majoritet av de avgivna rösterna.
Omröstningen ska vara sluten.
3.
Om kandidaten blir vald, ska talmannen underrätta rådet och uppmana rådet och den person som valts till kommissionens ordförande att i samförstånd nominera de övriga personer som de vill utse till ledamöter av kommissionen.
4.
Om parlamentet inte godkänner nomineringen, ska talmannen uppmana rådet att nominera en ny kandidat.
Artikel
99
Val av kommissionen
1.
Talmannen ska, efter att ha hört kommissionens nyvalde ordförande, uppmana dem som den nyvalde ordföranden och rådet nominerat till ledamöter av kommissionen att framträda inför lämpligt utskott i enlighet med sina framtida ansvarsområden.
Dessa utfrågningar ska vara offentliga.
2.
Behörigt eller behöriga utskott ska uppmana den nominerade kommissionsledamoten att göra ett uttalande och besvara frågor.
Utfrågningarna ska anordnas på sådant sätt att de nominerade kommissionsledamöterna får möjlighet att lämna alla relevanta upplysningar till parlamentet.
Bestämmelser om anordnandet av utfrågningarna ska fastställas i en bilaga till arbetsordningen
Se bilaga XVI b.
.
3.
Den nyvalde ordföranden ska presentera kollegiet och dess program vid ett plenarsammanträde, där hela rådet inbjuds att delta.
Programförklaringen ska följas av en debatt.
4.
Som avslutning på debatten har varje politisk grupp eller minst 40 ledamöter rätt att lägga fram ett resolutionsförslag.
Efter omröstningen om resolutionsförslaget ska parlamentet välja eller avvisa kommissionen med en majoritet av de avgivna rösterna.
Omröstningen ska förrättas med namnupprop.
Parlamentet kan skjuta upp omröstningen till nästföljande sammanträde.
5.
Talmannen ska underrätta rådet om huruvida kommissionen har valts eller avvisats.
6.
Om det under mandatperioden sker en avsevärd förändring beträffande ansvarsområden inom kommissionen, om det utnämns en ersättare eller om det utses en ny kommissionsledamot till följd av anslutning av en ny medlemsstat, ska berörda kommissionsledamöter bjudas in till det utskott som ansvarar för deras behörighetsområde i enlighet med punkt 2.
Artikel
100
Misstroendeförklaring mot kommissionen
1.
En tiondel av parlamentsledamöterna kan förelägga talmannen ett förslag till misstroendeförklaring mot kommissionen.
2.
Förslaget ska betecknas "förslag till misstroendeförklaring" och vara försett med motivering.
Det ska översändas till kommissionen.
3.
Så snart talmannen mottagit ett förslag till misstroendeförklaring, ska talmannen underrätta ledamöterna om att ett sådant förslag har ingivits.
4.
Debatten om misstroendeförklaringen ska äga rum tidigast 24 timmar efter det att ledamöterna underrättats om förslaget till misstroendeförklaring.
5.
Omröstningen om förslaget ska förrättas med namnupprop och ska hållas tidigast 48 timmar efter debattens början.
6.
Debatten och omröstningen ska äga rum senast under den sammanträdesperiod som följer på ingivandet av förslaget.
7.
Förslaget till misstroendeförklaring antas om det erhåller en majoritet av två tredjedelar av de avgivna rösterna och en majoritet av parlamentets samtliga ledamöter.
Rådets ordförande och kommissionens ordförande ska underrättas om omröstningsresultatet.
Artikel
101
Utnämning av revisionsrättens ledamöter
1.
Kandidater som har nominerats till ledamöter av revisionsrätten ska uppmanas att göra ett uttalande inför behörigt utskott samt besvara frågor från dess ledamöter.
Utskottet ska genom sluten omröstning rösta om varje enskild nominering.
2.
3.
Omröstningen i kammaren ska förrättas inom två månader från det att nomineringen mottagits, såvida inte parlamentet på begäran av behörigt utskott, en politisk grupp eller minst 40 ledamöter beslutar annorlunda.
Omröstningen ska vara sluten och parlamentet ska rösta separat om varje nominering och fatta sitt beslut med majoritet av de avgivna rösterna.
4.
Om parlamentet avstyrker en enskild nominering ska talmannen uppmana rådet att dra tillbaka sitt förslag och förelägga parlamentet ett nytt.
Artikel
102
Utnämning av direktionsledamöter i Europeiska centralbanken
1.
Den kandidat som nomineras till Europeiska centralbankens ordförande ska uppmanas att göra ett uttalande inför behörigt utskott samt besvara frågor från dess ledamöter.
2.
Utskottet ska till parlamentet lämna en rekommendation av vilken det framgår huruvida det tillstyrker utnämningen av den nominerade kandidaten.
3.
Omröstningen ska förrättas inom två månader från det att nomineringen mottagits, såvida inte parlamentet på begäran av behörigt utskott, en politisk grupp eller minst 40 ledamöter beslutar annorlunda.
4.
Om parlamentet avstyrker nomineringen ska talmannen uppmana rådet att dra tillbaka sitt förslag och förelägga parlamentet ett nytt.
5.
Samma förfarande ska tillämpas vid nomineringar till vice ordförande och andra direktionsledamöter i Europeiska centralbanken.
KAPITEL
2
UTTALANDEN
Artikel
103
Uttalanden av kommissionen, rådet och Europeiska rådet
1.
Ledamöter av kommissionen, rådet och Europeiska rådet kan när som helst anhålla om talmannens tillstånd att göra ett uttalande.
Talmannen avgör när ett uttalande får göras och huruvida ett sådant uttalande ska följas av en fullständig debatt eller endast 30 minuters frågestund med korta och koncisa frågor från ledamöterna.
2.
När ett uttalande med debatt har förts upp på föredragningslistan, ska kammaren besluta om debatten ska avslutas med att en resolution antas.
Om inte talmannen på grund av särskilda omständigheter beslutar annorlunda, ska debatten inte avslutas med att en resolution antas om ett betänkande om samma ämne ska tas upp under samma eller nästkommande sammanträdesperiod.
Om kammaren beslutar att en debatt ska avslutas med antagandet av en resolution får ett utskott, en politisk grupp eller minst 40 ledamöter lägga fram ett resolutionsförslag.
3.
Ett sådant resolutionsförslag ska gå till omröstning samma dag.
Talmannen ska fatta beslut om eventuella undantag.
Röstförklaringar ska tillåtas.
4.
Ett gemensamt resolutionsförslag kan ersätta de resolutionsförslag som förslagsställarna ingivit tidigare, men inte dem som ingivits av andra utskott, politiska grupper eller ledamöter.
5.
När en resolution har antagits får inga andra resolutionsförslag gå till omröstning om inte talmannen i undantagsfall beslutar annorlunda.
Artikel
104
Förklaringar av kommissionens beslut
Talmannen kan efter samråd med talmanskonferensen uppmana kommissionens ordförande, den kommissionsledamot som ansvarar för förbindelserna med parlamentet, eller enligt överenskommelse någon annan kommissionsledamot, att uttala sig inför parlamentet efter vart och ett av kommissionens sammanträden för att förklara de viktigaste besluten.
Uttalandet ska följas av en minst 30 minuter lång debatt, under vilken ledamöterna får ställa korta och koncisa frågor.
Artikel
105
Uttalanden av revisionsrätten
1.
Revisionsrättens ordförande kan, som ett led i ansvarsfrihetsförfarandet eller parlamentets verksamhet inom budgetkontrollområdet, uppmanas att presentera kommentarerna i revisionsrättens årsrapport, särskilda rapporter eller yttranden, eller att förklara rättens arbetsprogram.
2.
Parlamentet kan besluta att i närvaro av kommissionen och rådet hålla en särskild debatt om varje fråga som tas upp i ett sådant uttalande, särskilt om oegentligheter i budgetförvaltningen har påvisats.
Artikel
106
Uttalanden av Europeiska centralbanken
1.
Europeiska centralbankens ordförande ska förelägga parlamentet bankens årsrapport om verksamheten inom Europeiska centralbankssystemet och om den monetära politiken under det föregående och det innevarande året.
2.
Därefter ska parlamentet hålla en allmän debatt.
3.
Europeiska centralbankens ordförande ska uppmanas att närvara vid sammanträden i behörigt utskott åtminstone fyra gånger om året för att göra ett uttalande och besvara frågor.
4.
Europeiska centralbankens ordförande, vice ordförande och övriga direktionsledamöter ska inbjudas att närvara vid ytterligare sammanträden, om de själva eller parlamentet begär detta.
5.
Ett fullständigt förhandlingsreferat från de sammanträden som hålls i enlighet med punkterna 3 och 4 ska upprättas på de officiella språken.
Artikel
107
Rekommendation om de allmänna riktlinjerna för den ekonomiska politiken
1.
Kommissionens rekommendation om de allmänna riktlinjerna för medlemsstaternas och gemenskapens ekonomiska politik ska hänvisas till behörigt utskott, som ska förelägga kammaren ett betänkande.
2.
Rådet ska uppmanas att informera parlamentet om innehållet i sin rekommendation och om den ståndpunkt som intagits av Europeiska rådet.
KAPITEL
3
FRÅGOR TILL RÅDET, KOMMISSIONEN OCH EUROPEISKA CENTRALBANKEN
Artikel
108
Frågor för muntligt besvarande med debatt
1.
Ett utskott, en politisk grupp eller minst 40 ledamöter får ställa frågor till rådet och kommissionen och begära att de ska föras upp på parlamentets föredragningslista.
Sådana frågor ska skriftligen inges till talmannen som utan dröjsmål ska hänskjuta dem till talmanskonferensen.
Talmanskonferensen ska avgöra om och i vilken ordning frågor ska föras upp på föredragningslistan.
Frågor som inte förts upp på parlamentets föredragningslista inom tre månader efter det att de ingivits ska utgå.
2.
Frågor till kommissionen ska vidarebefordras till denna institution minst en vecka före det sammanträde då frågorna enligt föredragningslistan ska behandlas.
3.
4.
En av frågeställarna har högst fem minuter till förfogande för att utveckla frågan.
En ledamot av den berörda institutionen ska besvara frågan.
Frågeställaren har rätt att utnyttja hela sin talartid.
5.
Artikel
109
Frågestund
1.
Frågestund för frågor till rådet och kommissionen ska hållas under varje sammanträdesperiod vid tidpunkter som bestäms av parlamentet på förslag av talmanskonferensen.
Särskild tid kan avsättas för frågor till kommissionens ordförande och enskilda ledamöter av kommissionen.
2.
Under en och samma sammanträdesperiod får ingen ledamot ställa mer än en fråga till rådet och kommissionen.
3.
Frågor ska inges skriftligen till talmannen, som avgör deras tillåtlighet och den ordning i vilken de ska behandlas.
Frågeställaren ska omgående underrättas om beslutet.
4.
Närmare bestämmelser om förfarandet ska fastställas genom riktlinjer som ingår i en bilaga till arbetsordningen
Se bilaga II.
.
Artikel
110
Frågor till rådet och kommissionen för skriftligt besvarande
1.
Alla ledamöter får ställa frågor för skriftligt besvarande till rådet och kommissionen i enlighet med riktlinjerna
Se bilaga IIa.
.
Frågeställaren får själv avgöra vad frågorna ska handla om.
2.
Sådana frågor ska skriftligen inges till talmannen, som ska vidarebefordra dem till berörd institution.
I tveksamma fall ska talmannen avgöra om en fråga är tillåtlig eller inte.
Talmannens beslut ska meddelas frågeställaren.
3.
Om en fråga inte kan besvaras inom utsatt tid, ska den på frågeställarens begäran föras upp på föredragningslistan till nästa sammanträde i behörigt utskott.
Artikel 109 ska gälla i tillämpliga delar.
4.
Frågor som kräver ett omedelbart svar, men inte någon ingående undersökning (prioriterade frågor), ska besvaras inom tre veckor.
Varje ledamot har rätt att ställa en prioriterad fråga per månad.
Andra frågor (icke-prioriterade frågor) ska besvaras senast sex veckor efter det att de ingivits till den berörda institutionen.
Ledamöter ska ange vilken typ av fråga det rör sig om.
Det slutgiltiga avgörandet träffas av talmannen.
5.
Frågor och svar ska offentliggöras i Europeiska unionens officiella tidning.
Artikel
111
Frågor till Europeiska centralbanken för skriftligt besvarande
1.
Alla ledamöter får ställa frågor för skriftligt besvarande till Europeiska centralbanken i enlighet med riktlinjerna
Se bilaga IIa.
.
2.
3.
Frågor och svar ska offentliggöras i Europeiska unionens officiella tidning.
4.
Om en fråga inte har besvarats inom den fastställda tidsfristen ska den på frågeställarens begäran föras upp på föredragningslistan för det ansvariga utskottets närmast påföljande sammanträde med ordföranden för Europeiska centralbanken.
KAPITEL
4
RAPPORTER FRÅN ANDRA INSTITUTIONER
Artikel
112
Årsrapporter och andra rapporter från andra institutioner
1.
Årsrapporter och andra rapporter från andra institutioner som parlamentet enligt fördragen eller enligt andra rättsliga bestämmelser ska höras om, ska behandlas genom ett betänkande som ska läggas fram för kammaren.
2.
Årsrapporter och andra rapporter från andra institutioner vilka inte omfattas av vad som sägs i punkt 1 ska hänvisas till behörigt utskott som sedan får föreslå att ett betänkande ska utarbetas i enlighet med artikel 45.
KAPITEL
5
RESOLUTIONER OCH REKOMMENDATIONER
Artikel
113
Resolutionsförslag
1.
Varje ledamot får inge ett resolutionsförslag i ett ämne som faller inom Europeiska unionens verksamhetsområde.
Förslaget får omfatta högst 200 ord.
2.
Ansvarigt utskott ska avgöra vilket förfarande som ska tillämpas.
Utskottet kan sammanfoga ett resolutionsförslag med andra resolutionsförslag eller betänkanden.
Utskottet kan besluta att avge ett yttrande, eventuellt i form av en skrivelse.
Utskottet kan besluta att utarbeta ett betänkande i enlighet med artikel 45.
3.
Författarna till ett resolutionsförslag ska underrättas om utskottets och talmanskonferensens beslut.
4.
Betänkandet ska innehålla resolutionsförslagets text.
5.
Yttranden i form av skrivelser adresserade till andra institutioner inom Europeiska unionen ska översändas av talmannen.
6.
7.
Ett resolutionsförslag som lagts fram i enlighet med punkt 1 kan dras tillbaka av författaren, författarna eller den förste som undertecknat förslaget om detta görs innan ansvarigt utskott i enlighet med punkt 2 har beslutat att utarbeta ett betänkande om förslaget.
När ett förslag på detta sätt har övertagits av utskottet har endast utskottet självt rätt att dra tillbaka det fram till dess att slutomröstningen om förslaget inleds.
8.
Ett resolutionsförslag som dragits tillbaka kan omgående övertas och inges på nytt av en grupp, ett utskott eller samma antal ledamöter som ursprungligen hade rätt att inge förslaget.
Utskotten är skyldiga att se till att alla resolutionsförslag som lagts fram i enlighet med denna artikel, och som uppfyller de krav som fastställts, följs upp och nämns i de handlingar som utarbetas i samband med uppföljandet.
Artikel
114
Rekommendationer till rådet
1.
En politisk grupp eller minst 40 ledamöter kan förelägga rådet ett förslag till rekommendation om frågor som behandlas i avdelningarna V och VI i EU-fördraget eller, när parlamentet inte har hörts, om internationella avtal som omfattas av artikel 83 eller 84 i arbetsordningen.
2.
Sådana förslag ska hänvisas till behörigt utskott för beredning.
I förekommande fall ska behörigt utskott överlämna ärendet till kammaren i enlighet med bestämmelserna i denna arbetsordning.
3.
När behörigt utskott avger ett betänkande ska det förelägga parlamentet ett förslag till rekommendation till rådet, tillsammans med en kortfattad motivering och eventuella yttranden från de utskott som har hörts.
Tillämpning av punkt 3 kräver inte förhandsgodkännande av talmanskonferensen.
4.
Bestämmelserna i artikel 90 eller 94 ska tillämpas.
Artikel
115
Debatter om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer
1.
2.
På grundval av en sådan begäran som avses i punkt 1, och i enlighet med bestämmelserna i bilaga III, ska talmanskonferensen upprätta en förteckning över de ämnen som ska föras upp i det slutgiltiga förslaget till föredragningslista inför nästa debatt om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer.
Högst tre ämnen, inklusive underavdelningar, får föras upp på föredragningslistan.
Parlamentet kan i enlighet med artikel 132 besluta att ett ämne som ska debatteras ska utgå och ersättas med ett debattämne som inte finns på föredragningslistan.
Resolutionsförslag om de ämnen som valts ska inges senast på kvällen den dag då föredragninglistan godkänns.
Talmannen ska fastställa den exakta tidsfristen för ingivande av sådana resolutionsförslag.
3.
När den tid som beräknats för redogörelse för och omröstning om resolutionsförslag liksom även den talartid som eventuellt tilldelats rådet eller kommissionen räknats bort, ska återstående talartid fördelas mellan de politiska grupperna och de grupplösa ledamöterna.
4.
Omröstning ska förrättas omedelbart efter debattens slut.
Artikel 163 ska inte tillämpas.
Omröstningar som förrättas i överensstämmelse med denna artikel får efter talmannens och talmanskonferensens beslut anordnas som en enda omröstning.
5.
6.
Talmannen och ordförandena i de politiska grupperna får besluta att låta ett resolutionsförslag gå till omröstning utan debatt.
För ett sådant beslut fordras enhällighet bland ordförandena i samtliga politiska grupper.
Bestämmelserna i artiklarna 167, 168 och 170 ska inte tillämpas på resolutionsförslag som tagits upp på föredragningslistan till en debatt om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer.
Resolutionsförslag till en debatt om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer ska läggas fram först efter det att förteckningen över ämnen har godkänts.
Alla resolutionsförslag som inte hinner behandlas inom den tidsram som avsatts för debatten bortfaller.
Ledamöter har naturligtvis rätt att åter lägga fram sådana förslag, antingen för beredning i utskott i enlighet med artikel 113 eller till debatten om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer vid nästföljande sammanträdesperiod.
Ett ämne kan inte tas upp på föredragningslistan till en debatt om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer, om det redan förekommer på föredragningslistan till den sammanträdesperioden.
Artikel
116
Skriftliga förklaringar
1.
En skriftlig förklaring på högst 200 ord om ett ämne som faller inom Europeiska unionens verksamhetsområde kan inges av upp till fem ledamöter.
Skriftliga förklaringar ska tryckas på de officiella språken och delas ut.
De ska tillsammans med namnen på undertecknarna finnas i ett register.
Detta register ska vara offentligt och ska under sammanträdesperioderna placeras utanför ingången till plenisalen, medan det mellan sammanträdesperioderna ska placeras på en lämplig plats som bestäms av kvestorskollegiet.
Innehållet i en skriftlig förklaring ska inte överskrida den sedvanliga formen för en förklaring och, i synnerhet, inte innehålla beslut om frågor för vars antagande det i arbetsordningen anges särskilda förfaranden och behörigheter.
2.
Varje ledamot har rätt att underteckna en skriftlig förklaring som införts i registret.
3.
När en majoritet av parlamentets samtliga ledamöter har undertecknat en förklaring ska talmannen underrätta parlamentet om detta och i protokollet offentliggöra namnen på undertecknarna.
4.
En sådan förklaring ska efter sammanträdesperioden översändas till de institutioner som anges i förklaringen, tillsammans med namnen på undertecknarna.
Förklaringen ska ingå i protokollet från det sammanträde där förklaringen tillkännagavs.
När förklaringen på detta sätt har offentliggjorts är förfarandet avslutat.
5.
En skriftlig förklaring bortfaller om den har varit införd i registret längre än tre månader och inte har undertecknats av minst hälften av parlamentets samtliga ledamöter.
Artikel
117
Samråd med Europeiska ekonomiska och sociala kommittén
1.
Ett utskott kan begära att Europeiska ekonomiska och sociala kommittén hörs i allmänna eller särskilda frågor.
Utskottet ska ange när Europeiska ekonomiska och sociala kommittén ska ha yttrat sig.
2.
En begäran om att höra Europeiska ekonomiska och sociala kommittén ska godkännas av kammaren utan debatt.
Artikel
118
Samråd med Regionkommittén
1.
Ett utskott kan begära att Regionkommittén hörs i allmänna eller särskilda frågor.
Utskottet ska ange när Regionkommittén ska ha yttrat sig.
2.
En begäran om att höra Regionkommittén ska godkännas av kammaren utan debatt.
Artikel
119
Begäran till EU-organ
1.
I de fall parlamentet har rätt att rikta en begäran till ett EU-organ har varje ledamot möjlighet att lämna in en sådan begäran i form av en skrivelse till parlamentets talman.
En begäran ska gälla frågor som faller inom ifrågavarande EU-organs uppdrag och åtföljas av bakgrundsinformation som förklarar den fråga som ska beaktas och gemenskapens intresse däri.
2.
Efter att ha rådfrågat ansvarigt utskott ska talmannen antingen vidarebefordra en inlämnad begäran till organet eller vidta annan lämplig åtgärd.
Den ledamot som inlämnat en begäran ska omedelbart underrättas om talmannens åtgärder.
I samband med varje begäran som talmannen översänder till ett organ ska även tidsfrist för det begärda svaret anges.
3.
Om organet anser att det inte har möjlighet att yttra sig över en begäran såsom den framställts, eller anser att den bör omformuleras, ska det omgående meddela talmannen, som ska vidta lämpliga åtgärder efter att vid behov ha rådfrågat ansvarigt utskott.
KAPITEL
6
INTERINSTITUTIONELLA AVTAL
Artikel
120
Interinstitutionella avtal
1.
Parlamentet kan ingå avtal med andra institutioner om fördragens tillämpning och om förbättring eller förtydligande av olika förfaranden.
Sådana avtal kan utgöras av gemensamma uttalanden, skriftväxlingar, förhållningsregler eller andra lämpliga instrument.
De ska efter behandling i utskottet med behörighet i konstitutionella frågor och efter parlamentets godkännande undertecknas av talmannen.
De kan för kännedom fogas som bilagor till arbetsordningen.
2.
KAPITEL
7
FÖRFARANDEN VID DOMSTOLEN
Artikel
121
Förfaranden vid domstolen
1.
Före utgången av de tidsfrister för att väcka talan som gäller för Europeiska unionens institutioner och för fysiska och juridiska personer i enlighet med fördragen och domstolens stadgar, ska parlamentet granska gemenskapslagstiftningen och genomförandebestämmelserna för att försäkra sig om att fördragen till fullo respekteras, framför allt vad gäller parlamentets rättigheter.
2.
Ansvarigt utskott ska underrätta parlamentet, vid behov muntligen, om det misstänker en överträdelse av gemenskapsrätten.
3.
Talmannen ska i enlighet med en rekommendation från det behöriga utskottet väcka talan på parlamentets vägnar.
I början av nästföljande sammanträdesperiod kan talmannen förelägga kammaren ett beslut om att vidhålla talan.
Om kammaren med en majoritet av de avgivna rösterna fattar ett beslut som går emot talan, ska talmannen dra tillbaka denna.
Om talmannen väcker talan i strid med rekommendationen från det behöriga utskottet, ska han eller hon i början av nästföljande sammanträdesperiod förelägga kammaren ett beslut om att vidhålla talan.
4.
Talmannen ska efter att ha hört ansvarigt utskott avge yttranden eller agera på parlamentets vägnar i domstolsförfaranden.
Om talmannen avser att avvika från det ansvariga utskottets rekommendation ska han eller hon informera utskottet om detta samt hänskjuta frågan till talmanskonferensen med angivande av sina skäl.
Om talmanskonferensen anser att parlamentet undantagsvis inte bör inkomma med inlagor eller skriftliga yttranden till domstolen i mål där giltigheten av en rättsakt som parlamentet antagit ifrågasätts, ska ärendet utan dröjsmål föreläggas kammaren.
I brådskande fall får talmannen vidta förebyggande åtgärder för att den berörda domstolens tidsfrister ska respekteras.
I sådana fall ska det förfarande som anges i denna punkt genomföras så snart som möjligt.
Inget i arbetsordningen hindrar det ansvariga utskottet från att i brådskande fall fatta beslut om lämpliga förfaranden för att kunna översända rekommendationen i rätt tid.
Artikel
122
Följder av rådets underlåtenhet att agera efter det att dess gemensamma ståndpunkt har godkänts enligt samarbetsförfarandet
Har parlamentet inom tre eller, med rådets samtycke, fyra månader efter mottagandet av den gemensamma ståndpunkten i enlighet med artikel 252 i EG-fördraget varken avvisat eller ändrat den gemensamma ståndpunkten och rådet underlåter att anta den föreslagna rättsakten i enlighet med den gemensamma ståndpunkten, får talmannen på parlamentets vägnar och efter att ha hört utskottet med behörighet i rättsliga frågor väcka talan vid domstolen mot rådet i enlighet med artikel 232 i EG-fördraget.
AVDELNING
V
FÖRBINDELSER MED NATIONELLA PARLAMENT
Artikel
123
Utbyte av uppgifter samt kontakter och ömsesidiga resurser
1.
Parlamentet ska regelbundet informera medlemsstaternas nationella parlament om parlamentets verksamhet.
2.
Talmanskonferensen kan ge talmannen mandat att förhandla om resurser som på ömsesidig grund ska ställas till medlemsstaternas nationella parlaments förfogande och föreslå andra åtgärder för att underlätta kontakterna med de nationella parlamenten.
Artikel
124
Konferensen mellan organ för EG- och EU-frågor (COSAC)
1.
Talmanskonferensen ska på förslag av talmannen utse och ge mandat åt ledamöterna i parlamentets delegation till COSAC.
Delegationen ska ledas av en av de vice talmännen med ansvar för förbindelserna med de nationella parlamenten.
2.
De övriga delegationsledamöterna ska utses med hänsyn till de ämnen som ska behandlas vid COSAC:s sammanträde och med beaktande av den övergripande politiska jämvikten i parlamentet.
Delegationen ska lämna en rapport efter varje sammanträde.
Artikel
125
Parlamentariska konferenser
Delegationerna ska själva utse ordförande och i förekommande fall en eller flera vice ordförande.
AVDELNING
VI
SESSIONER
KAPITEL
1
PARLAMENTETS SESSIONER
Artikel
126
Parlamentets valperiod, sessioner, sammanträdesperioder, sammanträden
1.
Parlamentets valperiod sammanfaller med ledamöternas mandattid enligt akten av den 20 september 1976.
2.
Session är den årslånga period som föreskrivs i ovannämnda akt och i fördragen.
3.
Sammanträdesperioder är de perioder - som regel varje månad - då parlamentet sammanträder.
Plenarsammanträden som hålls samma dag betraktas som ett enda sammanträde.
Artikel
127
Sammankallande av parlamentet
1.
Parlamentet sammanträder utan att kallelse krävs den andra tisdagen i mars varje år och avgör då de sammanträdesfria periodernas längd under sessionen.
2.
3.
4.
Talmannen ska, efter att ha hört talmanskonferensen, sammankalla parlamentet till ett extra sammanträde om en majoritet av parlamentets samtliga ledamöter, kommissionen eller rådet begär detta.
I undantagsfall kan talmannen med talmanskonferensens samtycke i brådskande fall sammankalla parlamentet till ett extra sammanträde.
Artikel
128
Plats för sammanträden
1.
Parlamentet ska hålla sina plenarsammanträden och utskottssammanträden i enlighet med vad som föreskrivs i fördragen.
Förslag om extra sammanträdesperioder i Bryssel och ändringsförslag till dessa behöver endast majoritet av de avgivna rösterna för att antas.
2.
Alla utskott kan begära att ett eller flera sammanträden hålls på annan ort.
En begäran försedd med motivering ska överlämnas till talmannen som ska lägga fram den för presidiet.
I brådskande fall kan talmannen själv fatta beslut i frågan.
Om presidiet eller talmannen avslår begäran ska skälen till detta redovisas.
Artikel
129
Deltagande i sammanträden
1.
Vid varje sammanträde ska det finnas en närvarolista som ledamöterna ska skriva på.
2.
Namnen på de ledamöter som är närvarande enligt närvarolistan ska föras till protokollet från varje sammanträde.
KAPITEL
2
PARLAMENTETS ARBETSGÅNG
Artikel
130
Förslag till föredragningslista
1.
Före varje sammanträdesperiod ska talmanskonferensen upprätta ett förslag till föredragningslista på grundval av utskottsordförandekonferensens rekommendationer och med beaktande av det antagna lagstiftningsprogram som avses i artikel 33.
Kommissionen och rådet har rätt att på talmannens inbjudan delta i talmanskonferensens överläggningar om förslag till föredragningslista.
2.
I förslaget till föredragningslista kan tider för omröstningar fastställas för enskilda punkter på föredragningslistan.
3.
I förslaget till föredragningslista kan en eller två perioder på sammanlagt högst 60 minuter avsättas för debatter om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer i enlighet med artikel 115.
4.
Det slutgiltiga förslaget till föredragningslista ska delas ut till ledamöterna senast tre timmar före sammanträdesperiodens början.
Artikel
131
Förfarande i kammaren utan ändringsförslag och debatt
1.
Lagstiftningsförslag (första behandlingen) och resolutionsförslag som inte avser lagstiftning och som har antagits av utskottet varvid färre än en tiondel av utskottsledamöterna röstat emot, ska föras upp på parlamentets förslag till föredragningslista för omröstning utan ändringsförslag.
Ärendet ska sedan vara föremål för en enda omröstning, såvida inte politiska grupper eller enskilda ledamöter som tillsammans utgör en tiondel av parlamentets ledamöter före upprättandet av det slutgiltiga förslaget till föredragningslistan skriftligen begär att ärendet ska vara föremål för ändringsförslag.
I så fall ska talmannen fastställa en tidsfrist för att inge ändringsförslag.
2.
Ärenden som har förts upp på det slutgiltiga förslaget till föredragningslista för omröstning utan ändringsförslag ska även avgöras utan debatt, såvida inte parlamentet, på förslag av talmanskonferensen eller på begäran av en politisk grupp eller minst 40 ledamöter, beslutar annorlunda då föredragningslistan godkänns vid sammanträdesperiodens inledning.
3.
När talmanskonferensen upprättar det slutgiltiga förslaget till föredragningslista för en sammanträdesperiod får den föreslå att andra ärenden ska behandlas utan ändringsförslag eller debatt.
När parlamentet godkänner föredragningslistan får det inte godkänna något sådant förslag om en politisk grupp eller minst 40 ledamöter skriftligen har motsatt sig detta minst en timme innan sammanträdesperioden inleds.
4.
När ett ärende avgörs utan debatt får föredraganden eller ordföranden i behörigt utskott omedelbart före omröstningen göra ett kort uttalande på högst två minuter.
Artikel
131 a
Kortfattad redogörelse
På begäran av föredraganden eller på förslag från talmanskonferensen får parlamentet också besluta att en fråga som inte behöver tas upp i en omfattande debatt ska behandlas genom att föredraganden gör en kortfattad redogörelse i kammaren.
Artikel
132
Godkännande och ändring av föredragningslistan
1.
Parlamentet ska vid början av varje sammanträdesperiod fatta beslut om det slutgiltiga förslaget till föredragningslista.
Ändringsförslag kan läggas fram av ett utskott, en politisk grupp eller minst 40 ledamöter.
Alla sådana förslag ska vara talmannen tillhanda senast en timme före sammanträdesperiodens början.
Talmannen kan ge ordet till förslagsställaren, en talare som är för förslaget och en talare som är emot förslaget.
Talartiden får inte överstiga en minut.
2.
När föredragningslistan väl har godkänts kan den inte ändras, förutom i enlighet med artiklarna 134 och 167-171 eller på förslag av talmannen.
Förkastas ett förslag om att ändra föredragningslistan, kan detta förslag inte läggas fram på nytt vid samma sammanträdesperiod.
3.
Innan talmannen avslutar sammanträdet ska datum, tidpunkt och föredragningslista för nästa sammanträde meddelas.
Artikel
133
Särskild debatt
1.
En politisk grupp eller minst 40 ledamöter kan begära att en särskild debatt om ett ämne av större vikt med anknytning till Europeiska unionens politik ska föras upp på parlamentets föredragningslista.
Under varje sammanträdesperiod ska det i regel endast hållas en särskild debatt.
2.
En sådan begäran ska inges skriftligen till talmannen senast tre timmar före inledningen av den sammanträdesperiod under vilken den särskilda debatten ska äga rum.
Omröstningen om ett sådant förslag ska genomföras vid sammanträdesperiodens inledning i samband med godkännandet av föredragningslistan.
3.
För att kunna reagera på händelser som inträffar efter godkännandet av föredragningslistan för en sammanträdesperiod kan talmannen, efter samråd med de politiska gruppernas ordförande, föreslå en särskild debatt.
4.
Talmannen ska fastställa tidpunkten för en särskild debatt.
Den sammanlagda tiden för en sådan debatt får inte överstiga 60 minuter.
5.
Debatten ska avslutas utan att någon resolution antas.
Artikel
134
Brådskande debatt
1.
Denna begäran ska inges skriftligen och vara försedd med motivering.
2.
Så snart talmannen har mottagit en begäran om brådskande debatt ska talmannen underrätta parlamentet om detta.
Omröstning om en sådan begäran ska hållas vid inledningen av det sammanträde som följer på det sammanträde då tillkännagivandet gjordes, förutsatt att det förslag som begäran avser har delats ut på de officiella språken.
Finns det flera än en begäran om brådskande debatt som rör samma ämne, ska bifall respektive avslag på en begäran om brådskande debatt gälla varje begäran som rör detta ämne.
3.
Före omröstningen kan endast den som inkommit med en begäran, en talare för, en talare emot samt ansvarigt utskotts ordförande eller föredragande tilldelas ordet i högst tre minuter var.
4.
De ärenden om vilka kammaren beslutar att tillämpa brådskande debatt ska ges företräde framför andra punkter på föredragningslistan.
Talmannen fastställer tidpunkten för debatt och omröstning.
5.
En brådskande debatt kan hållas utan betänkande eller i undantagsfall på grundval av en muntlig rapport från ansvarigt utskott.
Artikel
135
Gemensam debatt
Beslut kan när som helst fattas om att vid ett och samma tillfälle debattera liknande ärenden eller ärenden som hör ihop.
Artikel
136
Tidsfrister
Förutom i de brådskande fall som avses i artiklarna 115 och 134, får en debatt eller omröstning om en text endast inledas om texten delats ut minst 24 timmar tidigare.
KAPITEL
3
ALLMÄNNA BESTÄMMELSER FÖR PLENARSAMMANTRÄDEN
Artikel
137
Tillträde till plenisalen
1.
Tillträde till plenisalen har endast parlamentsledamöter, ledamöter av kommissionen och rådet, parlamentets generalsekreterare, parlamentspersonal vars uppgifter kräver närvaro där samt unionens experter och tjänstemän.
2.
Endast innehavare av ett av talmannen eller parlamentets generalsekreterare vederbörligen utställt tillträdeskort har rätt att vistas på åhörarläktaren.
3.
Åhörare som vistas på åhörarläktaren måste förbli sittande och vara tysta.
Åhörare som uttrycker bifall eller ogillande ska genast föras ut av vaktmästarna.
Artikel
138
Språk
1.
Samtliga parlamentets handlingar ska avfattas på de officiella språken.
2.
Samtliga ledamöter ska ha rätt att hålla sina anföranden i parlamentet på det officiella språk de önskar.
Anföranden på ett av de officiella språken ska simultantolkas till övriga officiella språk och till varje annat språk som presidiet anser nödvändigt.
3.
Vid varje utskotts- och delegationssammanträde ska tolkning finnas tillgänglig från och till de officiella språk som ledamöterna och suppleanterna i utskottet eller delegationen i fråga använder och begär.
4.
Vid utskotts- och delegationssammanträden utanför de vanliga arbetsorterna ska tolkning finnas tillgänglig från och till de språk som används av de ledamöter som bekräftat att de kommer att delta i sammanträdet.
Avsteg från dessa regler får göras undantagsvis med godkännande från ledamöterna i utskottet eller delegationen.
Om en överenskommelse inte kan uppnås ska presidiet avgöra frågan.
Originalversionen kan inte alltid betraktas som den officiella texten, eftersom en situation kan uppstå där alla de övriga språken avviker från originalversionen.
Artikel
139
Övergångsbestämmelser
1.
Under en övergångsperiod fram till sjätte valperiodens utgång ska det vara tillåtet att göra undantag från bestämmelserna i artikel 138, om och i den utsträckning det för ett officiellt språk inte finns tillräckligt många tolkar eller översättare trots att lämpliga åtgärder vidtagits.
2.
På förslag från generalsekreteraren ska presidiet fastställa om villkoren i punkt 1 är uppfyllda för vart och ett av de berörda officiella språken, och var sjätte månad ska det se över sitt beslut på grundval av en rapport från generalsekreteraren om de framsteg som gjorts.
Presidiet ska anta de genomförandebestämmelser som behövs.
3.
De särskilda tidsbegränsade bestämmelser som rör utarbetandet av rättsakter och som rådet utfärdat med stöd av fördragen ska tillämpas; med undantag för förordningar som Europaparlamentet och rådet antar gemensamt.
4.
Parlamentet kan efter det att presidiet lämnat en motiverad rekommendation när som helst besluta att upphäva denna artikel i förtid, eller att förlänga giltighetstiden för densamma vid utgången av den frist som anges i punkt 1.
Artikel
140
Utdelning av handlingar
Handlingar som utgör underlag för parlamentets debatter och beslut ska tryckas och delas ut till ledamöterna.
En förteckning över dessa handlingar ska offentliggöras i protokollen från parlamentets sammanträden.
Utan att det påverkar tillämpningen av första stycket, ska ledamöter och politiska grupper ha direkt tillgång till parlamentets interna datasystem för att konsultera alla förberedande handlingar som inte är sekretessbelagda (förslag till betänkanden, förslag till rekommendationer, förslag till yttranden, arbetsdokument och ändringsförslag som lagts fram i utskott).
Artikel
141
Tilldelning av ordet och anförandens innehåll
1.
Ingen ledamot har rätt att yttra sig om inte talmannen tilldelat ledamoten ordet.
2.
Om en talare avviker från ämnet, ska talmannen återkalla talaren till ordningen.
Har talaren vid samma debatt redan återkallats till ordningen två gånger, har talmannen rätt att den tredje gången frånta talaren ordet för återstoden av den debatt som rör detta ämne.
3.
Utan att det påverkar talmannens övriga disciplinära befogenheter, kan talmannen från det fullständiga förhandlingsreferatet avföra anföranden och inlägg från ledamöter som inte tilldelats ordet eller som överskridit den tilldelade talartiden.
4.
En talare får endast avbrytas av talmannen.
Talaren kan dock med talmannens medgivande själv avbryta sitt anförande för att låta en annan ledamot, kommissionen eller rådet ställa en fråga angående en bestämd punkt i anförandet.
Artikel
142
Fördelning av talartid
1.
Talmanskonferensen kan föreslå parlamentet att talartid fördelas för en bestämd debatt.
Parlamentet ska utan debatt fatta beslut om ett sådant förslag.
2.
Talartiden ska fördelas i enlighet med följande kriterier:
a)
En första del av talartiden ska fördelas lika mellan alla politiska grupper.
b)
En andra del ska fördelas mellan de politiska grupperna i proportion till deras sammanlagda antal ledamöter.
c)
De grupplösa ledamöterna ska tilldelas en sammanlagd talartid som baseras på de delar som respektive politisk grupp tilldelas enligt a och b ovan.
3.
Avsätts en gemensam talartid för flera punkter på föredragningslistan, ska de politiska grupperna underrätta talmannen om hur stor del av talartiden som de avser att använda för varje enskild punkt.
Talmannen ska se till att dessa talartider respekteras.
4.
Talartiden för inlägg om sammanträdesprotokollen, arbetsordningen, ändringar till det slutgiltiga förslaget till föredragningslista eller till föredragningslistan får inte överstiga en minut.
5.
Kommissionen och rådet ska som regel ha rätt att yttra sig i en debatt om ett betänkande direkt efter det att betänkandet har lagts fram av föredraganden.
Kommissionen, rådet och föredraganden får höras igen, särskilt för att bemöta uttalanden från Europaparlamentets ledamöter.
6.
Utan att det påverkar tillämpningen av artikel 197 i EG-fördraget ska talmannen försöka komma överens med kommissionen och rådet om en lämplig fördelning av talartiden för dessa institutioner.
7.
Ledamöter som inte yttrat sig under en debatt kan, högst en gång per sammanträdesperiod, lämna in en skriftlig förklaring på högst 200 ord som ska bifogas protokollet från debatten.
Artikel
143
Talarlista
1.
Namnen på de ledamöter som begär ordet ska föras upp på talarlistan i den ordning deras begäran togs emot.
2.
Talmannen tilldelar ledamöter ordet och ska så långt det är möjligt se till att talare från olika politiska åsiktsriktningar och talare som talar olika språk växelvis tilldelas ordet.
3.
Ansvarigt utskotts föredragande, politiska gruppers ordförande som önskar tala på gruppens vägnar, eller talare som ersätter dessa, kan på begäran ges företräde framför andra talare.
4.
Ingen ledamot får utan talmannens medgivande yttra sig mer än två gånger om samma ämne.
Berörda utskotts ordförande och föredragande ska dock på egen begäran få tala under en tid som bestäms av talmannen.
Artikel
144
Anföranden på en minut
Under högst trettio minuter vid varje sammanträdesperiods första sammanträde ska talmannen tilldela de ledamöter ordet som önskar göra anföranden för att uppmärksamma parlamentet på en fråga av politisk vikt.
Talartiden för var och en av ledamöterna får inte överskrida en minut.
Talmannen kan besluta att tillåta ytterligare en sådan period senare under samma sammanträdesperiod.
Artikel
145
Personliga uttalanden
1.
En ledamot som begär att få göra ett personligt uttalande ska tilldelas ordet i slutet av debatten om den punkt på föredragningslistan som behandlas, eller när protokollet från det sammanträde begäran av ordet avser ska justeras.
Ledamoten i fråga får inte yttra sig i sakfrågan utan ska begränsa sitt inlägg till att bemöta yttranden som under debattens gång fällts om ledamotens person eller påståenden om ledamotens åsikter eller för att tillrättalägga sina egna tidigare yttranden.
2.
Ett personligt uttalande får inte överstiga tre minuter om inte kammaren beslutar annorlunda.
KAPITEL
4
ÅTGÄRDER VID LEDAMÖTERS ÖVERTRÄDELSE AV ORDNINGSREGLERNA
Artikel
146
Omedelbara åtgärder
1.
Varje ledamot som uppträder störande under ett sammanträde eller uppträder på ett sätt som strider mot tillämpliga bestämmelser i artikel 9 ska kallas till ordningen av talmannen.
2.
Upprepas förseelsen ska talmannen återigen kalla ledamoten till ordningen, och saken ska föras till sammanträdesprotokollet.
3.
Vid upprepat störande uppträdande eller om ytterligare förseelser begås kan talmannen förbjuda ledamoten att ta till orda eller uppmana ledamoten att lämna plenisalen för återstoden av sammanträdet.
Vid synnerligen grova ordningsförseelser kan talmannen omedelbart uppmana ledamoten att lämna plenisalen utan att dessförinnan än en gång ha återkallat till ordningen.
Generalsekreteraren ska utan dröjsmål se till att denna disciplinära åtgärd verkställs med hjälp av vaktmästarna och vid behov med hjälp av parlamentets säkerhetstjänst.
4.
Om ett störande uppträdande hotar att förhindra överläggningarna får talmannen, för att återställa ordningen, avbryta sammanträdet under en viss tid eller avsluta detsamma.
Kan talmannen inte göra sig hörd ska talmannen lämna ordförandeplatsen, vilket avslutar sammanträdet.
Talmannen är den som kallar till fortsatt sammanträde.
5.
De befogenheter som fastställs i punkterna 1-4 ska i tillämpliga delar tillkomma organens, utskottens och delegationernas mötesordförande enligt den definition som ges i arbetsordningen.
6.
I förekommande fall och beroende på hur allvarlig överträdelsen av ordningsreglerna är kan mötesordföranden senast vid nästkommande sammanträdesperiod eller berörda organs, utskotts eller delegations nästkommande sammanträde uppmana talmannen att tillämpa artikel 147.
Artikel
147
Påföljder
1.
2.
Sådana påföljder kan bestå av en eller flera av följande åtgärder:
a)
prickning
b)
indragning av dagtraktamentet under två till tio dagar,
c)
utan att det inverkar på rätten att rösta i kammaren, och under förutsättning att ordningsreglerna följs strikt, tidsbegränsad avstängning från deltagande i samtliga eller vissa av parlamentets eller något av dess organs, utskotts eller delegationers verksamhet under 2 till 10 på varandra följande sammanträdesdagar,
d)
framläggande till talmanskonferensen, i enlighet med artikel 18, av ett förslag om avstängning eller entledigande från ett eller flera av de uppdrag till vilka ledamoten har valts.
Artikel
148
Internt förfarande för överklagande
Presidiet kan senast fyra veckor efter att överklagandet inkommit upphäva, fastställa eller reducera påföljden, utan att detta påverkar ledamotens externa överklaganderättigheter.
Om presidiet inte fattar beslut inom angiven tid betraktas påföljden som ogiltig.
KAPITEL
5
BESLUTFÖRHET OCH OMRÖSTNING
Artikel
149
Beslutförhet
1.
Parlamentet har rätt att hålla överläggningar, fastställa föredragningslista och justera sammanträdesprotokoll oavsett antalet närvarande ledamöter.
2.
Beslutförhet föreligger om en tredjedel av parlamentets samtliga ledamöter är närvarande i plenisalen.
3.
Alla omröstningar är giltiga oavsett antalet deltagare i en omröstning, såvida inte talmannen i samband med omröstningen, till följd av en begäran gjord av minst 40 ledamöter innan omröstningen inletts, förklarar att beslutförhet inte föreligger.
Om omröstningen visar att beslutförhet inte föreligger, ska omröstningen tas upp på föredragningslistan till nästföljande sammanträde.
En begäran om fastställandet av huruvida beslutförhet föreligger måste göras av minst 40 ledamöter.
En begäran på en politisk grupps vägnar är inte tillåtlig.
När omröstningsresultatet fastställs ska hänsyn tas dels till antalet närvarande ledamöter i kammaren enligt punkt 2, dels till antalet ledamöter som begärt ett fastställande av beslutförhet enligt punkt 4.
Det elektroniska omröstningssystemet får inte användas för detta syfte.
Plenisalens dörrar får inte stängas.
Om antalet närvarande ledamöter inte uppgår till det antal som krävs för beslutförhet, ska talmannen inte tillkännage omröstningsresultatet utan förklara att beslutförhet inte föreligger.
Punkt 3 sista meningen ska inte tillämpas vid omröstningar om procedurfrågor utan endast vid omröstningar om sakfrågor.
4.
Ledamöter som begärt ett fastställande av beslutförhet ska räknas som närvarande enligt punkt 2, även om de inte längre befinner sig i plenisalen.
5.
Är färre än 40 ledamöter närvarande, har talmannen rätt att förklara att beslutförhet inte föreligger.
Artikel
150
Ingivande och framläggande av ändringsförslag
1.
Ansvarigt utskott, en politisk grupp eller minst 40 ledamöter kan inge ändringsförslag för behandling i kammaren.
Ändringsförslag ska inges skriftligen och vara undertecknade av författarna.
Ändringsförslag till handlingar som avser lagstiftning enligt artikel 40.1 kan förses med en kort motivering.
2.
Utan att det påverkar tillämpningen av artikel 151 kan ett ändringsförslag syfta till att ändra vilken del som helst av en text och till att stryka, tillföra eller ersätta ord eller siffror.
Med "text" avses i denna artikel och i artikel 151 hela den samlade textmassan i ett resolutionsförslag, förslag till lagstiftningsresolution, förslag till beslut eller kommissionsförslag.
3.
Talmannen ska fastställa en tidsfrist för ingivande av ändringsförslag.
4.
Ett ändringsförslag kan under debatten läggas fram av förslagsställaren eller av varje annan ledamot som förslagsställaren utsett till ersättare.
5.
Om en förslagsställare drar tillbaka sitt ändringsförslag ska detta bortfalla, såvida det inte genast övertas av en annan ledamot.
6.
Ändringsförslag ska gå till omröstning först efter det att de tryckts och delats ut på alla officiella språk, såvida inte kammaren beslutar annorlunda.
Kammaren kan inte fatta ett sådant beslut om minst 40 ledamöter motsätter sig detta.
Artikel 139 ska gälla i tillämpliga delar på denna punkt.
Muntliga ändringsförslag som läggs fram i ett utskott kan gå till omröstning, såvida inte någon av utskottets ledamöter motsätter sig detta.
Artikel
151
Ändringsförslags tillåtlighet
1.
Ett ändringsförslag är otillåtligt om
a)
det inte har något direkt samband med den text som det syftar till att ändra,
b)
det avser att stryka eller ersätta texten i sin helhet,
c)
det avser att ändra fler än en av de enskilda artiklarna eller punkterna i den text som avses.
Denna bestämmelse ska inte tillämpas vid kompromissändringsförslag eller ändringsförslag som avser att ändra ett visst ord eller en viss formulering på exakt samma sätt genom hela texten,
d)
2.
Ett ändringsförslag bortfaller om det är oförenligt med tidigare fattade beslut om samma text vid samma omröstning.
3.
Talmannen ska avgöra om ett ändringsförslag är tillåtligt.
Talmannens beslut i punkt 3 angående ändringsförslags tillåtlighet ska inte uteslutande grundas på bestämmelserna i punkt 1 och 2 i denna artikel utan på bestämmelserna i arbetsordningen i allmänhet.
4.
En politisk grupp eller minst fyrtio ledamöter får inge ett alternativt resolutionsförslag till ett resolutionsförslag i ett utskottsbetänkande som inte avser lagstiftning.
I så fall får gruppen eller de berörda ledamöterna inte inge ändringsförslag till utskottets resolutionsförslag.
Ett sådant alternativt resolutionsförslag får inte vara längre än utskottets resolutionsförslag.
Resolutionsförslaget ska gå till omröstning genom en enda omröstning och utan ändringsförslag.
Artikel
152
Omröstningar
1.
Vid betänkanden ska följande omröstningsordning tillämpas:
a)
Omröstning om eventuella ändringsförslag till det förslag som tas upp i ansvarigt utskotts betänkande.
b)
Omröstning om hela förslaget - ändrat eller inte.
c)
Omröstning om ändringsförslag till resolutionsförslag eller till förslag till lagstiftningsresolutioner.
d)
Omröstning om resolutionsförslag eller förslag till lagstiftningsresolutioner i sin helhet (slutomröstning).
Parlamentet ska inte rösta om betänkandets motivering.
2.
Följande omröstningsordning ska tillämpas vid andra behandlingen:
a)
Har inget förslag om att avvisa eller ändra rådets gemensamma ståndpunkt lagts fram, ska den gemensamma ståndpunkten anses godkänd, i enlighet med artikel 67.
b)
c)
Har flera ändringsförslag till den gemensamma ståndpunkten lagts fram, ska omröstning om dessa förrättas i den ordning som fastställs i artikel 155.
d)
3.
Förfarandet i artikel 65 ska tillämpas vid tredje behandlingen.
4.
Vid omröstningar om lagstiftningstexter och resolutionsförslag som inte avser lagstiftning, ska de delar som rör det egentliga innehållet gå till omröstning först.
Om ett ändringsförslag står i strid med ett tidigare omröstningsresultat ska det bortfalla.
5.
Utskottets föredragande är den ende ledamot som får yttra sig i samband med omröstningen och endast för att kortfattat redovisa sitt utskotts ståndpunkter angående de ändringsförslag som omröstningen gäller.
Artikel
153
Lika röstetal
1.
2.
Uppkommer lika röstetal vid en omröstning om föredragningslistan i sin helhet (artikel 132), protokollet i sin helhet (artikel 172) eller vid en delad omröstning enligt artikel 157, ska texten anses antagen.
3.
I alla övriga fall av lika röstetal, utan att det påverkar tillämpningen av de artiklar som föreskriver kvalificerad majoritet ska texter eller förslag som gått till omröstning anses förkastade.
Artikel
154
Grundläggande principer för omröstningen
1.
Omröstning om ett betänkande ska förrättas på grundval av en rekommendation från ansvarigt utskott.
Utskottet kan delegera denna uppgift till sin ordförande eller föredragande.
2.
Utskottet kan rekommendera att en gemensam omröstning förrättas om alla eller flera av ändringsförslagen och att dessa ska antas, förkastas eller utgå.
Utskottet kan även lägga fram kompromissändringsförslag.
3.
Rekommenderar ansvarigt utskott en gemensam omröstning om ändringsförslag, ska den gemensamma omröstningen förrättas först.
4.
Om ansvarigt utskott lägger fram ett kompromissändringsförslag, ska omröstning om detta förrättas först.
5.
Omröstning om ändringsförslag för vilka namnupprop har begärts, ska förrättas separat.
6.
Delad omröstning ska inte tillåtas vid en gemensam omröstning eller en omröstning om ett kompromissändringsförslag.
Artikel
155
Omröstningsordning vid ändringsförslag
1.
Ändringsförslag har företräde framför den text de avser och ska gå till omröstning före den texten.
2.
Har två eller flera ändringsförslag, som ömsesidigt utesluter varandra, lagts fram till samma textavsnitt, ska det ändringsförslag som avviker mest från den ursprungliga texten ha företräde och vara det som först går till omröstning.
Antas det ändringsförslaget ska de övriga ändringsförslagen anses ha förkastats.
Förkastas det ska omröstning förrättas om det ändringsförslag som står närmast i tur och på samma sätt för vart och ett av de återstående ändringsförslagen.
Råder det tvekan om den inbördes ordningen, ska denna avgöras av talmannen.
Förkastas samtliga ändringsförslag ska den ursprungliga texten anses antagen om inte särskild omröstning begärts inom föreskriven tid.
3.
Talmannen kan låta den ursprungliga texten gå till omröstning först, eller låta ett ändringsförslag, som står närmare den ursprungliga texten än det ändringsförslag som avviker mest gå till omröstning före detta förslag.
Erhåller endera av dessa majoritet bortfaller alla övriga ändringsförslag som avser samma text.
4.
I undantagsfall kan det på förslag av talmannen förrättas omröstning om ändringsförslag som lagts fram efter det att debatten avslutats, om ändringsförslagen är kompromissändringsförslag eller om tekniska problem föreligger.
Talmannen ska inhämta kammarens samtycke till att låta sådana ändringsförslag gå till omröstning.
Vid kompromissändringsförslag som lagts fram efter en debatts avslutande i enlighet med denna punkt, ska talmannen i varje enskilt fall avgöra ändringsförslagens tillåtlighet med hänsyn till deras kompromisskaraktär.
Följande allmänna kriterier för tillåtlighet kan tillämpas:
-
Kompromissändringsförslag får normalt inte avse de delar av texten som när fr
i
sten för att inge ändringsförslag löpt ut inte varit föremål för ändringsförslag.
-
Kompromissändringsförslag ska
Endast talmannen kan föreslå att ett kompromissändringsförslag ska behandlas.
För att ett kompromissändringsförslag ska gå till omröstning, måste talmannen inhämta kammarens samtycke genom att fråga om det finns några invändningar mot en sådan omröstning.
Framförs invändningar ska kammaren avgöra frågan med majoritet av de avgivna rösterna.
5.
När ansvarigt utskott har lagt fram en rad ändringsförslag som avser samma text som betänkandet, ska talmannen låta dem gå till gemensam omröstning, såvida inte en politisk grupp eller minst 40 ledamöter begärt särskild omröstning eller andra ändringsförslag lagts fram.
6.
Talmannen kan låta andra ändringsförslag gå till gemensam omröstning om de kompletterar varandra.
I så fall ska talmannen tillämpa förfarandet i punkt 5.
Författarna till ändringsförslag som kompletterar varandra har rätt att föreslå en gemensam omröstning.
7.
Efter det att ett visst ändringsförslag har antagits eller förkastats, kan talmannen besluta att flera andra ändringsförslag med liknande innehåll eller liknande syften ska gå till gemensam omröstning.
Talmannen kan i förväg inhämta kammarens medgivande.
Sådana grupper av ändringsförslag kan avse olika delar av den ursprungliga texten.
8.
Om två eller flera identiska ändringsförslag läggs fram av olika personer, ska de gå till omröstning som ett enda ändringsförslag.
Artikel
156
Behandling i utskott av ändringsförslag ingivna för behandling i plenum
Om flera än 50 ändringsförslag har ingetts till ett betänkande för behandling i plenum får talmannen, efter samråd med utskottsordföranden, uppmana det ansvariga utskottet att hålla ett sammanträde för att behandla ändringsförslagen.
Endast ändringsförslag som då stöds av minst en tiondel av utskottets ledamöter ska tas upp till omröstning i plenum.
Artikel
157
Delad omröstning
1.
En politisk grupp eller minst 40 ledamöter kan begära delad omröstning om ett textavsnitt som ska gå till omröstning innehåller två eller flera bestämmelser, syftar på två eller flera punkter eller kan indelas i två eller flera delar som var och en har en egen logisk betydelse eller ett eget normativt värde.
2.
Begäran om delad omröstning ska göras kvällen före omröstningen, såvida inte talmannen fastställer en ny tidsfrist.
Talmannen ska fatta beslut om en sådan begäran.
Artikel
158
Rösträtt
Rösträtten är personlig.
Ledamöter ska avge sina röster personligen och var för sig.
Artikel
159
Omröstning
1.
Parlamentet röstar normalt med handuppräckning.
2.
Finner talmannen att resultatet av omröstningen är oklart ska en ny omröstning äga rum med hjälp av det elektroniska omröstningssystemet eller, om detta är ur funktion, genom att ledamöterna reser sig upp.
3.
Omröstningsresultaten ska registreras.
Artikel
160
Omröstning med namnupprop
1.
2.
Namnuppropet ska ske i bokstavsordning och börja med namnet på en ledamot som tas fram genom lottdragning.
Talmannen ska rösta sist.
Omröstningen sker genom att varje ledamot högt och tydligt säger "ja", "nej" eller "avstår".
Vid rösträkningen ska hänsyn endast tas till de röster som avgivits för eller emot ett förslag.
Talmannen ska fastställa omröstningsresultatet och tillkännage detta.
Artikel
161
Elektronisk omröstning
1.
Talmannen kan när som helst besluta att de omröstningar som avses i artiklarna 159, 160 och 162 ska förrättas med elektroniskt omröstningssystem.
Tekniska instruktioner för användningen av det elektroniska omröstningssystemet ska fastställas av presidiet.
2.
Används det elektroniska omröstningssystemet ska resultatet registreras endast i siffror.
3.
Det förfarande som beskrivs i punkt 1 i denna artikel kan användas för att avgöra om en sådan majoritet föreligger.
Artikel
162
Sluten omröstning
1.
Endast röstsedlar med nominerade ledamöters namn ska beaktas vid räkningen av antalet avgivna röster.
2.
Sluten omröstning kan även förrättas om minst en femtedel av parlamentets samtliga ledamöter så begär.
En sådan begäran måste framställas innan omröstningen inleds.
Parlamentet ska förrätta sluten omröstning om en begäran om sluten omröstning framställs av minst en femtedel av parlamentets samtliga ledamöter innan omröstningen inleds.
3.
En begäran om sluten omröstning har företräde framför en begäran om omröstning med namnupprop.
4.
Två till sex genom lottdragning framtagna ledamöter ska räkna de röster som avges i en sluten omröstning.
Vid omröstning enligt punkt 1 får nominerade kandidater inte vara rösträknare.
Namnen på de ledamöter som deltagit i en sluten omröstning ska föras till protokollet från det sammanträde då omröstningen ägde rum.
Artikel
163
Röstförklaringar
1.
När den allmänna debatten har avslutats, har varje ledamot rätt att i samband med slutomröstningen avge en muntlig röstförklaring på högst en minut eller en skriftlig röstförklaring på högst 200 ord, vilka ska ingå i det fullständiga förhandlingsreferatet.
Varje politisk grupp har rätt att avge en röstförklaring på högst två minuter.
När den första röstförklaringen har påbörjats ska ingen ytterligare begäran om att få avge röstförklaringar beviljas.
Röstförklaringar till slutomröstning kan avges om alla frågor som tagits upp i kammaren.
Termen "slutomröstning" anger inte vilken typ av omröstning det gäller, utan avser den sista omröstningen beträffande en fråga.
2.
Röstförklaringar ska inte tillåtas vid omröstning om procedurfrågor.
3.
Är ett kommissionsförslag eller ett betänkande uppfört på föredragningslistan enligt artikel 131, kan ledamöter inge en skriftlig röstförklaring i enlighet med punkt 1.
Såväl muntliga som skriftliga röstförklaringar måste ha ett direkt samband med den text som är föremål för omröstning.
Artikel
164
Invändningar beträffande omröstningar
1.
Talmannen ska vid varje enskild omröstning förklara omröstningen påbörjad och avslutad.
2.
När talmannen har förklarat en omröstning påbörjad, har endast talmannen rätt att göra inlägg innan omröstningen är avslutad.
3.
Ordningsfrågor beträffande en omröstnings giltighet kan tas upp efter det att talmannen har förklarat omröstningen avslutad.
4.
När resultatet av en omröstning med handuppräckning har tillkännagivits, kan en ledamot begära att resultatet ska kontrolleras med hjälp av det elektroniska omröstningssystemet.
5.
Talmannen avgör om det tillkännagivna resultatet är giltigt.
Talmannens beslut kan inte ifrågasättas.
KAPITEL
6
PROCEDURFRÅGOR
Artikel
165
Förslag som rör förfaranden
1.
En begäran om följande förslag som rör förfaranden ska ha företräde framför varje annan begäran om att tilldelas ordet:
a)
Förslag om avvisning av ett ärende som otillåtligt (artikel 167).
b)
Förslag om återförvisning till utskott (artikel 168).
c)
Förslag om avslutande av debatt (artikel 169).
d)
Förslag om uppskjutande av debatt och omröstning (artikel 170).
e)
Förslag om avbrytande eller avslutande av sammanträde (artikel 171).
Endast förslagsställaren samt en talare för, en talare emot och ansvarigt utskotts ordförande eller föredragande har rätt att yttra sig om sådana förslag.
2.
Talartiden får inte överstiga en minut.
Artikel
166
Ordningsfrågor
1.
En ledamot kan tilldelas ordet för att göra talmannen uppmärksam på eventuella överträdelser av parlamentets arbetsordning.
Ledamoten ska först ange vilken artikel som åsyftas.
2.
En begäran om att ta upp en sådan ordningsfråga ska ha företräde framför varje annan begäran om att tilldelas ordet.
3.
Talartiden får inte överstiga en minut.
4.
Talmannen ska omedelbart fatta beslut i ordningsfrågor i enlighet med arbetsordningen och ska meddela sitt beslut omedelbart efter det att ordningsfrågan har tagits upp.
Det ska inte förrättas någon omröstning om detta.
5.
Talmannen kan i undantagsfall förklara att beslutet kommer att tillkännages senare, dock senast 24 timmar efter det att ordningsfrågan togs upp.
Skjuts beslutet upp medför detta emellertid inte att debatten skjuts upp.
Talmannen kan hänvisa ärendet till behörigt utskott.
En begäran om att ta upp en ordningsfråga ska röra den punkt på föredragningslistan som just då behandlas.
En ledamot kan tilldelas ordet för att ta upp en ordningsfråga avseende ett annat ämne vid lämplig tidpunkt, exempelvis när behandlingen av den aktuella punkten på föredragningslistan avslutats eller innan sammanträdet avbryts.
Artikel
167
Avvisning av ett ärende som otillåtligt
1.
När en debatt om en bestämd punkt på föredragningslistan inleds kan förslag väckas om att avvisa denna punkt som otillåtlig.
Ett sådant förslag ska omedelbart gå till omröstning.
2.
Godkänns förslaget ska kammaren genast fortsätta till nästa punkt på föredragningslistan.
Artikel
168
Återförvisning till utskott
1.
En politisk grupp eller minst 40 ledamöter kan begära återförvisning till utskott när föredragningslistan ska fastställas eller innan debatten inleds.
2.
En politisk grupp eller minst 40 ledamöter kan även begära återförvisning till utskott före eller under en omröstning.
En sådan begäran ska tas upp till omröstning omedelbart.
3.
En sådan begäran kan endast göras en gång vid var och en av dessa olika etapper i förfarandet.
4.
Återförvisning till utskott innebär att debatten av punkten i fråga skjuts upp.
5.
Kammaren kan fastställa en tidpunkt före vilken utskottet ska redogöra för sina slutsatser.
Artikel
169
Avslutande av debatt
1.
Kammaren kan på förslag av talmannen eller på begäran av en politisk grupp eller minst 40 ledamöter avsluta en debatt innan samtliga talare på talarlistan tilldelats ordet.
Ett sådant förslag eller en sådan begäran ska genast gå till omröstning.
2.
Om förslaget godkänns eller begäran beviljas har endast en ledamot från varje politisk grupp som ännu inte haft ordet rätt att göra inlägg.
3.
Efter de inlägg som avses i punkt 2 ska debatten avslutas och kammaren övergå till omröstning om punkten i fråga, såvida det inte i förväg har fastställts en tidpunkt för omröstning.
4.
Ett förslag eller en begäran som förkastats respektive avslagits kan endast läggas fram på nytt vid samma debatt av talmannen.
Artikel
170
Uppskjutande av debatt och omröstning
1.
Vid inledandet av en debatt om en punkt på föredragningslistan kan en politisk grupp eller minst 40 ledamöter begära att debatten skjuts upp till en viss bestämd tidpunkt.
Ett sådant förslag ska omedelbart gå till omröstning.
2.
Om begäran bifalls ska kammaren gå vidare till nästa punkt på föredragningslistan.
Den uppskjutna debatten ska återupptas vid den tidpunkt som angivits.
3.
Om begäran avslås kan den inte läggas fram på nytt under samma sammanträdesperiod.
4.
Före eller under en omröstning kan en politisk grupp eller minst 40 ledamöter begära att omröstningen ska skjutas upp.
Omröstning om en sådan begäran ska ske omedelbart.
Beslutar parlamentet att skjuta upp en debatt till en senare sammanträdesperiod ska beslutet ange den sammanträdesperiod på vars föredragningslista debatten ska tas upp, varvid föredragningslistan till den sammanträdesperioden ovillkorligen ska upprättas i enlighet med artiklarna 130 och 132 i arbetsordningen.
Artikel
171
Avbrytande eller avslutande av sammanträde
Ett sammanträde kan avbrytas eller avslutas under en debatt eller omröstning, om parlamentet på förslag av talmannen eller på begäran av en politisk grupp eller minst 40 ledamöter så beslutar.
Ett sådant förslag eller en sådan begäran ska omedelbart gå till omröstning.
KAPITEL
7
DOKUMENTATION AV SAMMANTRÄDEN
Artikel
172
Protokoll
1.
Protokollet från varje sammanträde, innehållande parlamentets beslut och namnen på talarna, ska delas ut minst en halvtimme före inledningen av det därpå följande sammanträdets eftermiddagsblock.
2.
Vid inledningen av varje sammanträdes eftermiddagsblock ska talmannen förelägga kammaren protokollet från föregående sammanträde för justering.
3.
Framförs invändningar mot protokollet ska kammaren avgöra huruvida de föreslagna ändringarna ska beaktas.
Ingen ledamot får yttra sig om protokollet i mer än en minut.
4.
Protokollet ska undertecknas av talmannen och generalsekreteraren och förvaras i parlamentets arkiv.
Det ska inom en månad offentliggöras i Europeiska unionens officiella tidning.
Artikel
173
Fullständigt förhandlingsreferat
1.
För varje sammanträde ska ett fullständigt förhandlingsreferat upprättas på alla officiella språk.
2.
Talare är skyldiga att återlämna rättelser av utskrifter av sina anföranden till sekretariatet inom en vecka.
3.
Det fullständiga förhandlingsreferatet ska offentliggöras som bilaga till Europeiska unionens officiella tidning.
4.
Ledamöter kan kräva att utdrag från det fullständiga förhandlingsreferatet ska översättas med kort varsel.
Artikel
173 a
Audiovisuell upptagning av förhandlingar
Omedelbart efter sammanträdet ska en audiovisuell upptagning av förhandlingarna, inklusive ljudinspelningar från alla tolkbås, produceras och göras tillgänglig via Internet.
AVDELNING
VII
UTSKOTT, UNDERSÖKNINGSKOMMITTÉER OCH DELEGATIONER
KAPITEL
1
UTSKOTT OCH UNDERSÖKNINGSKOMMITTÉER - TILLSÄTTNING OCH BEHÖRIGHETSOMRÅDEN
Artikel
174
Tillsättning av ständiga utskott
Parlamentet ska på förslag från talmanskonferensen tillsätta ständiga utskott vars behörighetsområden fastställs i en bilaga till denna arbetsordning
Val av utskottsledamöter ska äga rum vid den första sammanträdesperioden efter nyval till parlamentet och på nytt två och ett halvt år därefter.
Ständiga utskotts behörighetsområden kan fastställas vid en annan tidpunkt än när dessa utskott tillsätts.
Artikel
175
Tillsättning av tillfälliga utskott
Eftersom tillfälliga utskotts behörighetsområden, sammansättning och mandatperioder fastställs vid samma tidpunkt som dessa utskott tillsätts, kan parlamentet inte vid en senare tidpunkt besluta att ändra behörighetsområdena genom att begränsa eller utvidga dessa.
Artikel
176
Undersökningskommittéer
1.
Parlamentet kan på begäran av en fjärdedel av ledamöterna tillsätta en undersökningskommitté för att utreda påstådda överträdelser av gemenskapsrätten eller fall av missförhållanden vid tillämpningen av gemenskapsrätten, oavsett om den som har gjort sig skyldig till överträdelsen är en gemenskapsinstitution, ett gemenskapsorgan, en offentlig myndighet i en medlemsstat eller en person som enligt gemenskapsrätten har befogenhet att tillämpa denna.
Beslut om att tillsätta en undersökningskommitté ska inom en månad offentliggöras i Europeiska unionens officiella tidning.
2.
Undersökningskommitténs arbetssätt ska regleras av de bestämmelser i denna arbetsordning som rör utskott, om inte annat följer av denna artikel och Europaparlamentets, rådets och kommissionens beslut av den 19 april 1995 om närmare föreskrifter för utövandet av Europaparlamentets undersökningsrätt
3.
I en begäran om att en undersökningskommitté ska tillsättas ska det anges vad som ska utredas och den ska innehålla en detaljerad redogörelse för de skäl som motiverar undersökningen.
På förslag av talmanskonferensen ska kammaren fatta beslut om huruvida undersökningskommittén ska tillsättas och hur den i så fall ska vara sammansatt.
Beslut om sammansättning ska fattas i enlighet med bestämmelserna i artikel 177.
4.
Undersökningskommittén ska avsluta sitt arbete genom att lägga fram en rapport inom tolv månader.
Parlamentet kan två gånger besluta att förlänga denna tidsfrist med ytterligare tre månader.
Endast ordinarie ledamöter, eller i deras frånvaro de ständiga suppleanterna, har rösträtt i en undersökningskommitté.
5.
Undersökningskommittén ska välja sin ordförande och två vice ordförande samt en eller flera föredragande.
6.
När en undersökningskommitté anser att någon av dess rättigheter inte har respekterats, kan den föreslå talmannen att vidta lämpliga åtgärder.
7.
Kostnader för resa och uppehälle för andra personer som hörs av en undersökningskommitté ska ersättas av Europaparlamentet enligt gällande villkor för utfrågning av sakkunniga.
De ska informeras om dessa rättigheter innan de hörs av undersökningskommittén.
8.
Ordföranden i en undersökningskommitté ska i samarbete med presidiet se till att eventuell sekretess respekteras och att ledamöterna vederbörligen informeras om detta.
Ordföranden ska dessutom uttryckligen hänvisa till bestämmelserna i artikel 2.2 i ovannämnda beslut.
Bestämmelserna i bilaga VII, del A i arbetsordningen ska tillämpas.
9.
När sekretessbelagda handlingar, som har vidarebefordrats, behandlas ska sådana tekniska hjälpmedel användas som kan garantera att endast de ledamöter som är ansvariga för ärendet i fråga får tillgång till dessa handlingar.
Sammanträden ska hållas i lokaler som utrustats på ett sådant sätt att ingen obehörig har möjlighet till avlyssning.
10.
Denna rapport ska offentliggöras.
På begäran av undersökningskommittén ska kammaren hålla en debatt om denna rapport under den sammanträdesperiod som följer på dess framläggande.
Inga ändringsförslag får inges vad beträffar ämnet för undersökningen såsom det har fastställts av en fjärdedel av parlamentets samtliga ledamöter (punkt 3) och inte heller till den tidsfrist inom vilken en rapport ska läggas fram i enlighet med punkt 4.
Artikel
177
Val av ledamöter till utskott
2.
Ändringsförslag till talmanskonferensens förslag är endast tillåtliga om de inges av minst 40 ledamöter.
Kammaren ska förrätta sluten omröstning om sådana förslag.
3.
4.
Om en politisk grupp underlåter att inom en av talmanskonferensen fastställd tidsfrist inge nomineringar till ledamöter av en undersökningskommitté i enlighet med punkt 1, ska talmanskonferensen endast förelägga parlamentet de nomineringar som ingivits före utgången av denna tidsfrist.
5.
Talmanskonferensen kan, med de berörda ledamöternas samtycke och med beaktande av punkt 1 ovan, besluta att tillfälligt fylla en vakant plats.
6.
Artikel
178
Suppleanter
1.
De politiska grupperna och de grupplösa ledamöterna kan till varje utskott utse ett antal ständiga suppleanter, vars antal ska svara mot det antal ordinarie ledamöter som företräder de olika grupperna och de grupplösa ledamöterna i respektive utskott.
Talmannen ska underrättas om detta.
Ständiga suppleanter har rätt att närvara och yttra sig vid utskottssammanträden och, i en ordinarie ledamots frånvaro, delta i omröstningar.
2.
Är en ordinarie ledamot frånvarande och inga ständiga suppleanter har utsetts, eller om även suppleanterna är frånvarande, kan den ordinarie ledamoten välja att låta sig företrädas av en annan ledamot från samma politiska grupp, vilken har rätt att rösta på den ledamotens vägnar.
Namnet på företrädaren ska anmälas till utskottsordföranden före omröstningen.
Punkt 2 ska i tillämpliga delar gälla även för de grupplösa ledamöterna.
a
a
-
a
t
-
Under inga omständigheter får en utskottsledamot vara suppleant för en ledamot som tillhör en annan politisk grupp.
Artikel
179
Utskottens behörighetsområden
1.
Ständiga utskott ska behandla ärenden som hänvisas till dem av kammaren eller, under ett sessionsuppehåll, av talmannen på talmanskonferensens vägnar.
(Se tolkningen till artikel 175.)
2.
Om ett ständigt utskott förklarar sig obehörigt att behandla ett ärende, eller om en behörighetstvist uppstår mellan två eller flera ständiga utskott, ska frågan om behörighet hänskjutas till talmanskonferensen senast fyra arbetsveckor efter det att ärendets hänvisning till utskott har tillkännagivits i kammaren.
Utskottsordförandekonferensen ska underrättas, vilken kan utfärda rekommendationer till talmanskonferensen.
Talmanskonferensen ska fatta beslut senast sex arbetsveckor efter det att ärendet hänskjutits till konferensen.
Annars ska ärendet tas upp till beslut på föredragningslistan för påföljande sammanträdesperiod.
3.
Om två eller flera ständiga utskott är behöriga att bereda ett ärende ska ett utskott utses till ansvarigt utskott och de övriga till rådgivande utskott.
Ett ärende får dock inte samtidigt hänvisas till fler än tre utskott, såvida det inte på goda grunder beslutas att denna regel ska frångås i enlighet med bestämmelserna i punkt 1.
4.
Två eller flera utskott eller underutskott kan gemensamt bereda ärenden som hör till deras behörighetsområden, men de har inte rätt att fatta beslut.
5.
Alla utskott kan med presidiets samtycke ge en eller flera av sina ledamöter ett studie- eller informationsuppdrag.
Artikel
180
Utskott med ansvar för valprövning
Bland de utskott som tillsatts i överensstämmelse med bestämmelserna i denna arbetsordning ska ett utskott ha ansvaret för att granska bevis om val av ledamöter och bereda beslut om alla invändningar om huruvida ett val är giltigt.
Artikel
181
Underutskott
1.
Efter att först ha inhämtat talmanskonferensens medgivande kan ett ständigt eller tillfälligt utskott, om dess arbete så kräver, tillsätta ett eller flera underutskott och samtidigt fastställa dessa underutskotts sammansättning (se artikel 177) och behörighetsområden.
Underutskott ska inge rapporter till det utskott som tillsatt dem.
2.
Det förfarande som gäller för utskott ska även gälla för underutskott.
3.
Suppleanter har rätt att närvara vid underutskottssammanträden på samma villkor som vid utskottssammanträden.
4.
Denna artikel ska tillämpas på ett sådant sätt att beroendeförhållandet mellan ett underutskott och det utskott som tillsatt det garanteras.
Därför ska alla ordinarie ledamöter i ett underutskott väljas bland de ledamöter som sitter i huvudutskottet.
Artikel
182
Utskottspresidium
1.
Vid det första utskottssammanträdet efter det att val av utskottsledamöter har förrättats i enlighet med artikel 177, ska utskottet i separata omröstningar välja ett presidium bestående av en ordförande och en, två eller tre vice ordförande.
Trots vad som sägs i första stycket ska fyra vice ordförande ingå i varje utskottspresidium under perioden januari 2007 till juli 2009.
Denna bestämmelse utgör inte hinder för ordföranden för huvudutskottet att låta ordförandena för underutskotten delta i arbetet i presidiet, eller att tillåta att de är ordförande vid debatter om de särskilda frågor som behandlas av de berörda underutskotten, förutsatt att detta sätt att förfara i sin helhet granskas och godkänns av presidiet.
2.
Om antalet kandidater svarar mot antalet lediga platser, kan valet ske med acklamation.
Om detta inte är fallet, eller på begäran av en sjättedel av utskottets ledamöter, ska valet ske med sluten omröstning.
Om det finns fler än en kandidat i den första valomgången, ska den kandidat väljas som erhåller en absolut majoritet av de avgivna rösterna, i enlighet med föregående stycke.
Vid den andra valomgången ska den kandidat som erhåller flest röster väljas.
Vid lika antal röster ska den äldste kandidaten anses vald.
Om en andra valomgång krävs kan nya kandidater utses.
KAPITEL
2
UTSKOTT OCH UNDERSÖKNINGSKOMMITTÉER - ARBETSSÄTT
Artikel
183
Utskottssammanträden
1.
ska sammanträda på kallelse av sin ordförande eller på uppmaning av talmannen.
2.
Kommissionen och rådet får delta i utskottssammanträden, om de av utskottets ordförande på utskottets vägnar inbjuds att delta.
Ett utskott får efter särskilt beslut inbjuda vem som helst att närvara och yttra sig vid ett sammanträde.
Beslut om huruvida en ledamots personliga assistenter ska få närvara vid utskottssammanträden ska på samma sätt överlåtas till varje enskilt utskott.
Ett ansvarigt utskott får med presidiets medgivande anordna en utfrågning av sakkunniga om det anser att en sådan utfrågning är nödvändig för att på ett effektivt sätt kunna utföra sitt arbete i ett bestämt ärende.
Rådgivande utskott har rätt att närvara vid utfrågningen om de så önskar.
3.
Sådana ledamöter kan emellertid av utskottet bemyndigas att i en rådgivande roll delta i utskottets arbete.
Artikel
184
Protokoll från utskottssammanträden
Protokoll från varje utskottssammanträde ska delas ut till utskottets samtliga ledamöter och föreläggas utskottet för justering vid det därpå följande sammanträdet.
Artikel
185
Omröstningar i utskott
1.
Alla ledamöter har rätt att inge ändringsförslag för beredning i utskott.
2.
I ett utskott föreligger beslutförhet endast när minst en fjärdedel av ledamöterna är närvarande.
Om en sjättedel av utskottets ledamöter innan omröstningen inleds så kräver, ska emellertid omröstningen anses giltig endast om en majoritet av utskottets samtliga ledamöter har deltagit i den.
3.
4.
Utskottets ordförande har rätt att delta i överläggningar och omröstningar, men har inte utslagsröst.
5.
Med beaktande av de ingivna ändringsförslagen kan utskottet, i stället för att låta förslagen gå till omröstning, uppmana föredraganden att inkomma med ett nytt förslag i vilket så många ändringsförslag som möjligt beaktas.
En ny tidsfrist ska därefter fastställas för ändringsförslag till detta förslag.
Artikel
186
Bestämmelser för plenarsammanträden som även ska gälla utskottssammanträden
Artikel
187
Frågestund i utskott
Ett utskott kan hålla en frågestund om utskottet så beslutar.
Varje utskott fastställer självt regler för frågestundens genomförande.
KAPITEL
3
INTERPARLAMENTARISKA DELEGATIONER
Artikel
188
Tillsättning av interparlamentariska delegationer och delegationernas uppgifter
1.
På talmanskonferensens förslag ska parlamentet tillsätta ständiga interparlamentariska delegationer samt besluta om deras utformning och antalet ledamöter med hänsyn till delegationernas uppgifter.
Val av ledamöter i delegationerna för hela valperioden ska förrättas vid den första eller andra sammanträdesperioden efter nyval till parlamentet.
2.
Val av ledamöter förrättas efter att de politiska grupperna och de grupplösa parlamentsledamöterna ingivit nomineringar till talmanskonferensen.
3.
Sammansättningen av delegationernas presidier ska fastställas enligt det förfarande som gäller för de ständiga utskotten enligt artikel 182.
4.
Kammaren ska fastställa de enskilda delegationernas allmänna befogenheter.
Den får när som helst besluta att utvidga eller inskränka dessa befogenheter.
5.
De genomförandebestämmelser som krävs för att delegationerna ska kunna utföra sitt arbete ska antas av talmanskonferensen på förslag av delegationsordförandekonferensen.
6.
Delegationsordföranden ska överlämna en rapport om delegationens verksamhet till utskottet med behörighet i utrikes- och säkerhetsfrågor.
Artikel
189
Samarbete med Europarådets parlamentariska församling
1.
Parlamentets organ, framförallt utskotten, ska samarbeta med motsvarande organ i Europarådets parlamentariska församling på de områden som är av gemensamt intresse för att på så sätt effektivisera arbetet och undvika dubbelarbete.
2.
Talmanskonferensen ska i samförstånd med behöriga organ vid Europarådets parlamentariska församling fastställa närmare föreskrifter för genomförandet av dessa bestämmelser.
Artikel
190
Gemensamma parlamentarikerkommittéer
1.
Europaparlamentet kan tillsätta gemensamma parlamentarikerkommittéer tillsammans med parlamenten i stater associerade med gemenskapen eller stater med vilka anslutningsförhandlingar har inletts.
Sådana kommittéer har rätt att utarbeta rekommendationer till de deltagande parlamenten.
När det gäller Europaparlamentet ska dessa rekommendationer hänvisas till behörigt utskott, vilket ska lägga fram förslag om åtgärder som bör vidtas.
2.
De gemensamma parlamentarikerkommittéernas allmänna befogenheter ska fastställas av Europaparlamentet och genom avtal med berört tredje land.
3.
Gemensamma parlamentarikerkommittéer ska lyda under de bestämmelser som fastställs i själva avtalet i fråga.
Dessa bestämmelser ska baseras på principen om jämlikhet mellan Europaparlamentets delegation och det berörda parlamentets delegation.
4.
5.
Val av ledamöter till Europaparlamentets delegationer till gemensamma parlamentarikerkommittéer och tillsättning av delegationernas presidier ska ske enligt det förfarande som fastställts för interparlamentariska delegationer.
AVDELNING
VIII
FRAMSTÄLLNINGAR
Artikel
191
Rätt att inge framställningar
1.
Alla medborgare i Europeiska unionen och alla fysiska och juridiska personer som är bosatta i eller har sin hemvist eller säte i en medlemsstat har rätt att ensamma eller tillsammans med andra medborgare eller personer göra en framställning till parlamentet i en fråga som hör till Europeiska unionens verksamhetsområde och som direkt berör framställaren.
2.
Framställningar till parlamentet ska vara försedda med namn, nationalitet och hemvist för varje framställare.
3.
Framställningar ska vara avfattade på ett av Europeiska unionens officiella språk.
Framställningar som är avfattade på ett annat språk ska endast behandlas om framställaren bifogar en översättning eller en sammanfattning av innehållet på ett av Europeiska unionens officiella språk.
Översättningen eller sammanfattningen ska utgöra parlamentets arbetsunderlag.
Parlamentets korrespondens med framställaren ska ske på det officiella språk som översättningen eller sammanfattningen avfattats på.
4.
5.
Framställningar som upptagits i registret, ska av talmannen hänvisas till behörigt utskott, som ska bedöma huruvida de faller inom Europeiska unionens verksamhetsområde.
6.
7.
Det ansvariga utskottet kan i sådana fall föreslå framställaren att vända sig till behörig myndighet i den berörda medlemsstaten eller till behörig myndighet i Europeiska unionen.
8.
Såvida inte framställaren begär att sekretess ska gälla vid behandlingen av framställningen, ska den tas upp i ett offentligt register.
9.
Om utskottet anser det lämpligt kan det hänvisa ärendet till ombudsmannen.
10.
Framställningar till parlamentet som ingivits av fysiska eller juridiska personer som varken är medborgare i Europeiska unionen, bosatta i en medlemsstat eller har sin hemvist eller säte i en medlemsstat, ska registreras och arkiveras separat.
En gång i månaden ska talmannen översända en förteckning över de framställningar som mottagits under föregående månad, med angivande av vilket ämne de behandlar, till utskottet med behörighet i frågor som rör prövning av framställningar.
Artikel
192
Prövning av framställningar
1.
Ansvarigt utskott kan besluta att utarbeta ett betänkande eller på annat sätt yttra sig över de framställningar som det har förklarat tillåtliga.
Utskottet kan, speciellt vid framställningar som söker ändra gällande lagstiftning, begära yttranden från andra utskott i enlighet med artikel 46.
2.
Det ska inrättas ett elektroniskt register i vilket medborgarna kan ge sitt stöd till framställaren genom att med sin egen elektroniska underskrift skriva på en framställning som har förklarats tillåtlig och som har upptagits i registret.
3.
Vid prövningen av framställningar eller för att utreda sakförhållanden kan utskottet höra framställare, anordna allmänna utfrågningar eller skicka ut ledamöter för att på ort och ställe orientera sig om sakförhållanden.
4.
Som ett led i förberedandet av sitt yttrande kan utskottet uppmana kommissionen att inkomma med handlingar, lämna upplysningar och ge utskottet tillgång till dess tjänster.
5.
Utskottet kan eventuellt förelägga parlamentet resolutionsförslag om framställningar som det har behandlat.
Utskottet kan även uppmana talmannen att vidarebefordra utskottets yttrande till kommissionen eller rådet.
6.
En gång varje halvår ska utskottet underrätta parlamentet om resultatet av sina överläggningar.
Utskottet ska i synnerhet underrätta parlamentet om åtgärder som kommissionen eller rådet vidtagit beträffande framställningar som parlamentet vidarebefordrat till dem.
7.
Talmannen ska underrätta framställarna om fattade beslut och skälen till dessa.
Artikel
193
Tillkännagivande av framställningar
1.
Sådana tillkännagivanden ska föras till protokollet från sammanträdet.
2.
Titel på och sammanfattning av texterna till de i registret upptagna framställningarna samt de yttranden som översänts och de viktigaste beslut som fattats i samband med behandlingen av framställningarna ska med framställarens medgivande göras tillgängliga för allmänheten i en databas.
Sekretessbelagda framställningar ska förvaras i parlamentets arkiv, där de ska vara tillgängliga för alla ledamöter.
AVDELNING
IX
OMBUDSMANNEN
Artikel
194
Utnämning av ombudsmannen
1.
Omedelbart efter valet av talman vid början av varje valperiod eller vid de fall som avses i punkt 8 ska talmannen begära nomineringar till ämbetet som ombudsman samt fastställa en tidsfrist för ingivandet av dessa nomineringar.
Denna begäran ska offentliggöras i Europeiska unionens officiella tidning.
2.
Nomineringar måste ha stöd av minst 40 av parlamentets ledamöter som ska komma från minst två medlemsstater.
Varje ledamot kan endast stödja en nominering.
Nomineringarna ska innehålla alla de handlingar som krävs för att styrka att kandidaten uppfyller villkoren i föreskrifterna för utövandet av ämbetet som ombudsman.
3.
Utfrågningarna ska vara öppna för parlamentets samtliga ledamöter.
4.
En alfabetisk förteckning över godkända nomineringar föreläggs sedan parlamentet för omröstning.
5.
Omröstningen ska vara sluten, och en majoritet av de avgivna rösterna krävs.
Om ingen kandidat har valts efter de två första valomgångarna, får endast de två kandidater som erhöll flest antal röster vid andra valomgången kvarstå som kandidater.
Vid lika röstetal ges företräde åt den äldste kandidaten.
6.
Talmannen ska innan omröstningen inleds försäkra sig om att minst hälften av parlamentets samtliga ledamöter är närvarande.
7.
Den utnämnda ombudsmannen ska omedelbart avlägga en ed inför domstolen.
8.
Ombudsmannen ska, såvida han eller hon inte avsätts eller avlider, utföra sina uppgifter till dess att en efterträdare övertar ämbetet.
Artikel
195
Ombudsmannens verksamhet
1.
Beslutet om de föreskrifter och allmänna villkor för ombudsmannens ämbetsutövning samt bestämmelserna för genomförandet av detta beslut, sådana de antagits av ombudsmannen, bifogas parlamentets arbetsordning
Se bilaga X.
2.
Ombudsmannen ska i enlighet med artikel 3.6 och 3.7 i ovannämnda beslut underrätta parlamentet om fel och försummelser som upptäckts, och det behöriga utskottet kan utarbeta ett betänkande om dessa.
Det behöriga utskottet ska utarbeta ett betänkande om denna rapport, vilket ska läggas fram för debatt i kammaren.
3.
Ombudsmannen kan också underrätta behörigt utskott på begäran av detta eller på eget initiativ höras av behörigt utskott.
Artikel
196
Avsättning av ombudsmannen
1.
En tiondel av parlamentets ledamöter kan begära att ombudsmannen ska avsättas, om ombudsmannen inte längre uppfyller de krav som ställs för att utföra uppgifterna eller om ombudsmannen gjort sig skyldig till allvarlig försummelse.
2.
En sådan begäran ska översändas till ombudsmannen och till behörigt utskott som, om en majoritet av dess ledamöter anser skälen vara välgrundade, ska förelägga parlamentet ett betänkande.
Ombudsmannen ska, om han eller hon så begär, höras innan betänkandet går till omröstning.
Parlamentet ska efter en debatt fatta beslut med sluten omröstning.
3.
Innan omröstningen inleds ska talmannen förvissa sig om att minst hälften av parlamentets samtliga ledamöter är närvarande.
4.
Om parlamentet antar förslaget om avsättning av ombudsmannen och ombudsmannen därefter inte avgår frivilligt ska talmannen, senast vid den sammanträdesperiod som följer på den vid vilken omröstningen ägde rum, vända sig till domstolen med en hemställan om att utan dröjsmål förklara ombudsmannen avsatt.
Avgår ombudsmannen på egen begäran inställs detta förfarande.
AVDELNING
X
PARLAMENTETS GENERALSEKRETARIAT
Artikel
197
Generalsekretariat
1.
Parlamentet ska biträdas av en generalsekreterare som utses av presidiet.
Generalsekreteraren ska inför presidiet avge en högtidlig försäkran om att utföra sina uppgifter samvetsgrant och helt opartiskt.
2.
Generalsekreteraren ska leda ett sekretariat, vars sammansättning och organisation ska fastställas av presidiet.
3.
Presidiet ska fastställa generalsekretariatets tjänsteförteckning och föreskrifter för tjänstemäns och övriga anställdas rättsliga ställning och ekonomiska situation.
Presidiet ska också fastställa vilka kategorier av tjänstemän och övriga anställda som helt eller delvis omfattas av artiklarna 12-14 i Europeiska gemenskapernas protokoll om immunitet och privilegier.
Talmannen ska vederbörligen underrätta Europeiska unionens berörda institutioner.
AVDELNING
XI
BEFOGENHETER GÄLLANDE POLITISKA PARTIER PÅ EUROPEISK NIVÅ
Artikel
198
Talmannens befogenheter
Artikel
199
Presidiets befogenheter
1.
Presidiet ska besluta om en ansökan om finansiering som lämnats in av ett politiskt parti på europeisk nivå och om fördelningen av anslagen mellan de stödmottagande partierna.
Presidiet ska upprätta en förteckning över stödmottagare och beviljade belopp.
2.
Presidiet ska besluta om eventuell indragning eller minskning av finansieringen och eventuellt återbetalning av belopp som erhållits felaktigt.
3.
Efter budgetåret ska presidiet godkänna den slutliga verksamhetsrapporten och den ekonomiska redovisningen från de politiska partier som har erhållit stöd.
4.
Presidiet får enligt de villkor som fastställs i Europaparlamentets och rådets förordning (EG) nr 2004/2003 ge tekniskt stöd till politiska partier på europeisk nivå i överensstämmelse med deras förslag.
Vissa beslut om att ge tekniskt stöd får presidiet delegera till generalsekreteraren.
5.
I alla de fall som avses i föregående punkter ska presidiet agera på förslag av generalsekreteraren.
Utom i de fall som avses i punkterna 1 och 4, ska presidiet innan det fattar beslut höra företrädare för det berörda politiska partiet.
Presidiet får när som helst begära att talmanskonferensen yttrar sig.
6.
Om parlamentet efter kontroll konstaterar att ett politiskt parti på europeisk nivå inte längre respekterar principerna om frihet, demokrati och respekt för de mänskliga rättigheterna och de grundläggande friheterna samt rättsstatsprincipen ska presidiet besluta att detta parti ska uteslutas från finansiering.
Artikel
200
Ansvarigt utskotts och plenums befogenheter
1.
På begäran av en fjärdedel av parlamentets ledamöter, vilka ska företräda minst tre politiska grupper, ska talmannen efter diskussion med talmanskonferensen ge ansvarigt utskott i uppdrag att kontrollera om ett politiskt parti på europeisk nivå fortfarande respekterar (i synnerhet i sitt program och i sin verksamhet) de principer på vilka Europeiska unionen grundas, nämligen principerna om frihet, demokrati och respekt för de mänskliga rättigheterna och de grundläggande friheterna samt rättsstatsprincipen.
2.
Det ansvariga utskottet ska, innan det lägger fram ett förslag till beslut för parlamentet, höra företrädarna för det berörda politiska partiet på europeisk nivå, begära att den kommitté bestående av oavhängiga personer, som avses i Europaparlamentets och rådets förordning (EG) nr 2004/2003, yttrar sig i frågan samt behandla kommitténs yttrande.
3.
Om förslaget till beslut inte antas med en majoritet av de avgivna rösterna ska motsatt beslut anses antaget.
4.
Parlamentets beslut gäller från den dag då den begäran som avses i punkt 1 ingavs.
5.
Talmannen ska företräda parlamentet i kommittén bestående av oavhängiga personer.
6.
Det ansvariga utskottet ska utarbeta den i Europaparlamentets och rådets förordning (EG) nr 2004/2003 angivna rapporten om tillämpningen av den förordningen och de finansierade verksamheterna och lägga fram rapporten för kammaren.
AVDELNING
XII
TILLÄMPNING OCH ÄNDRING AV ARBETSORDNINGEN
Artikel
201
Tillämpning av arbetsordningen
1.
Uppstår tveksamheter vid tillämpningen eller tolkningen av denna arbetsordning kan talmannen hänvisa frågan till behörigt utskott för beredning.
En utskottsordförande kan göra detta när sådana tveksamheter uppstår i utskottets arbete och har samband med detta arbete.
2.
Utskottet ska avgöra om det är nödvändigt att föreslå en ändring av arbetsordningen.
I så fall ska förfarandet i artikel 202 tillämpas.
3.
Beslutar utskottet att en tolkning av gällande arbetsordning är tillräcklig, ska det översända sin tolkning till talmannen som ska underrätta parlamentet under den påföljande sammanträdesperioden.
4.
Om en politisk grupp eller minst 40 ledamöter framför invändningar mot utskottets tolkning, ska frågan gå till omröstning i parlamentet.
Texten ska antas med majoritet av de avlagda rösterna, under förutsättning att minst en tredjedel av samtliga ledamöter är närvarande.
Vid avslag ska frågan återförvisas till utskottet.
5.
Tolkningar som inte bestrids och tolkningar som antas av parlamentet ska i kursiv stil fogas som förklarande kommentarer till berörda artiklar i arbetsordningen.
6.
Dessa tolkningar ska utgöra prejudikat för framtida tillämpning och tolkning av de berörda artiklarna.
7.
Ansvarigt utskott ska regelbundet se över tolkningar och arbetsordningens artiklar.
8.
När arbetsordningen ger ett bestämt antal ledamöter vissa rättigheter, ska detta antal automatiskt justeras till det närmaste hela antal som svarar mot samma procentandel av parlamentets ledamöter om parlamentets totala antal ledamöter ökar, t.ex. efter en utvidgning av Europeiska unionen.
Artikel
202
Ändring av arbetsordningen
1.
Alla ledamöter har rätt att föreslå ändringar av arbetsordningen och dess bilagor.
Sådana ändringsförslag ska översättas, tryckas, delas ut och hänvisas till behörigt utskott, som bereder dem och avgör om de ska föreläggas parlamentet.
Då artiklarna 150, 151 och 155 tillämpas vid behandlingen i kammaren av ändringsförslag till arbetsordningen, ska benämningarna "den ursprungliga texten" och "ett kommissionsförslag" i dessa artiklar betraktas som hänvisningar till gällande bestämmelser.
2.
Ändringsförslag till denna arbetsordning ska endast antas om de erhåller en majoritet av rösterna från parlamentets samtliga ledamöter.
3.
Såvida det inte vid omröstningstillfället beslutas annorlunda, ska ändringar till denna arbetsordning och dess bilagor träda i kraft den första dagen under den sammanträdesperiod som följer på deras antagande.
AVDELNING
XIII
DIVERSE BESTÄMMELSER
Artikel
203
Oavslutade ärenden
Vid slutet av den sista sammanträdesperioden före val till parlamentet, ska samtliga oavslutade ärenden, som förelagts parlamentet, anses ha bortfallit, om inte annat följer av bestämmelserna i andra stycket.
I början på varje valperiod ska talmanskonferensen fatta beslut om varje motiverad begäran från utskott och övriga institutioner om att återuppta eller fortsätta behandlingen av dessa ärenden.
Dessa bestämmelser gäller inte framställningar och texter om vilka beslut inte ska fattas.
Artikel
204
Bilagor till arbetsordningen
Bilagor till arbetsordningen ska ha följande indelning:
a)
Genomförandebestämmelser för arbetsordningens förfaranden, antagna med en majoritet av de avgivna rösterna (bilaga VI).
b)
Bestämmelser antagna enligt särskilda föreskrifter i arbetsordningen och enligt de förfaranden och majoritetsregler som anges i dessa föreskrifter (bilagorna I, II, III, IV, V, VII del A och del C, IX och XV).
c)
Interinstitutionella avtal och andra bestämmelser som utfärdats enligt fördragen och som gäller i parlamentet eller är av intresse för parlamentets verksamhet.
De sistnämnda bestämmelserna kan fogas som bilagor till arbetsordningen efter ett beslut av kammaren med en majoritet av de avgivna rösterna och på förslag av behörigt utskott (bilagorna VII del B, VIII, X, XI, XII, XIII, XIV och XVI.).
Artikel
204 a
Rättelser
1.
Om ett fel upptäcks i en text som antagits av parlamentet ska talmannen, när så är lämpligt, till det ansvariga utskottet lämna ett förslag till rättelse.
2.
Om ett fel upptäcks i en text som antagits av parlamentet och överenskommits med en annan institution ska talmannen inhämta denna institutions samtycke till de nödvändiga rättelserna och därefter tillämpa punkt 1.
3.
Det ansvariga utskottet ska behandla förslaget till rättelse och inge det till kammaren om det konstaterar att det begåtts ett fel som kan rättas på föreslaget sätt.
4.
Rättelsen ska tillkännages vid följande sammanträdesperiod.
Den ska anses ha godkänts om det inte senast 48 timmar efter tillkännagivandet inkommit en begäran från en politisk grupp eller minst 40 ledamöter om att rättelsen ska bli föremål för omröstning.
Om rättelsen inte godkänns ska den återförvisas till det ansvariga utskottet, som kan föreslå en ändrad rättelse eller avsluta förfarandet.
5.
BILAGA
I
Artikel
1
1.
Varje ledamot som har direkta ekonomiska intressen i en fråga som debatteras ska muntligen uppge dessa intressen om denne föreslås som föredragande samt innan denne yttrar sig i kammaren eller i något av parlamentets organ.
2.
Artikel
2
Kvestorerna ska föra ett register dit samtliga ledamöter personligen lämnar detaljerade upplysningar angående:
a)
Yrkesmässig verksamhet och alla övriga relevanta uppdrag eller all annan verksamhet som de utför mot ersättning.
b)
Ledamöterna har inte rätt att ta emot andra gåvor eller förmåner vid utövande av sitt mandat.
Varje ledamot har ett personligt ansvar för de upplysningar som lämnas till registret, vilka ska uppdateras årligen.
Presidiet kan regelbundet ange de uppgifter det anser bör ingå i registret.
Om en ledamot efter vederbörlig uppmaning inte lämnar uppgifter enligt led a och b ovan ska talmannen på nytt uppmana ledamoten att lämna dessa uppgifter inom två månader.
Löper denna tidsfrist ut utan att uppgifterna lämnats ska ledamotens namn, med uppgift om överträdelsen, offentliggöras genom en anteckning i protokollet från det första sammanträdet under varje sammanträdesperiod sedan tidsfristen löpt ut.
Vägrar ledamoten även sedan överträdelsen offentliggjorts att lämna dessa uppgifter ska talmannen tillämpa bestämmelserna i artikel 147 i arbetsordningen och avstänga ledamoten i fråga.
Ordförandena för de olika grupperingarna inom parlamentet, både tvärpolitiska grupper och andra inofficiella grupperingar av ledamöter, ska redogöra för alla bidrag, både ekonomiska och andra (exempelvis sekreterarhjälp), som, om de hade erbjudits ledamöterna personligen, skulle ha uppgivits i enlighet med denna artikel.
Kvestorerna ska ansvara för att ett register förs och ska fastställa detaljerade bestämmelser för hur grupperingarna ska redogöra för bidrag från utomstående.
Artikel
3
Registret ska vara offentligt.
Registret kan vara tillgängligt för allmänheten på elektronisk väg.
Artikel
4
I avvaktan på att en stadga införs för ledamöter av Europaparlamentet, som kan ersätta det stora antalet nationella bestämmelser, omfattas ledamöterna när det gäller deklaration av förmögenhet av lagstiftningen i den medlemsstat där de valts.
BILAGA
II
Genomförande av frågestunden i artikel 109
A.
Riktlinjer
1.
Frågor är tillåtliga endast om de
-
är kortfattade och formulerade på ett sådant sätt att ett kort svar kan lämnas,
-
faller inom kommissionens och rådets behörighets- och ansvarsområden och är av allmänt intresse,
-
inte kräver omfattande förstudier eller efterforskningar för berörd institution,
-
är klart formulerade och avser en konkret punkt,
-
inte innehåller påståenden eller omdömen,
-
inte avser rent personliga angelägenheter,
-
inte syftar till att skaffa fram handlingar eller statistiska upplysningar,
-
är formulerade som frågor.
2.
Frågor är inte tillåtliga om de avser ärenden som redan är upptagna på föredragningslistan och om vilka överläggningar med deltagande av berörd institution redan har fastställts.
3.
Frågor är inte tillåtliga om identiska eller liknande frågor har ställts och besvarats under de närmast föregående tre månaderna, såvida det inte har skett en förändring av situationen eller frågeställaren vill ha ytterligare information.
I det första fallet ska en kopia av frågan och svaret överlämnas till frågeställaren.
Följdfrågor
4.
Varje ledamot har rätt att till varje fråga följa upp svaret med en följdfråga.
Ledamoten får endast ställa två följdfrågor.
5.
De bestämmelser om frågors tillåtlighet som fastställs i dessa riktlinjer ska även gälla följdfrågor.
6.
Talmannen avgör följdfrågors tillåtlighet och ska begränsa antalet så att varje ledamot som har ställt en fråga kan få den besvarad.
Även om en följdfråga uppfyller ovannämnda villkor är talmannen inte skyldig att förklara följdfrågan tillåtlig
a)
om det är sannolikt att den kommer att störa frågestundens normala förlopp,
b)
om den huvudfråga som följdfrågan avser redan har belysts tillräckligt av andra följdfrågor, eller
c)
om det inte finns något direkt samband med huvudfrågan.
Besvarande av frågor
7.
Berörd institution ska se till att svaren är kortfattade och av relevans för frågans ämne.
8.
Om innehållet i flera frågor så tillåter kan talmannen, efter att ha hört frågeställarna, besluta att berörd institution ska besvara dem tillsammans.
9.
En fråga får endast besvaras om frågeställaren är närvarande eller om frågeställaren före frågestundens inledande skriftligen underrättat ordföranden om namnet på sin ersättare.
10.
Om varken frågeställaren eller frågeställarens ersättare är närvarande bortfaller frågan.
11.
Om en ledamot inger en fråga, men varken ledamoten själv eller ledamotens ersättare är närvarande vid frågestunden, ska talmannen skriftligen påminna ledamoten om att det är hans eller hennes skyldighet att antingen närvara själv eller se till att det finns en ersättare.
Om talmannen tre gånger inom loppet av en tolvmånadersperiod är tvungen att sända en sådan skrivelse, ska ledamoten i fråga för en tid av sex månader förlora sin rätt att inge frågor.
12.
13.
Tidsfrister
14.
Frågor ska inges senast en vecka innan frågestunden inleds.
Frågor som inte ingivits inom denna tid får behandlas under frågestunden om berörd institution ger sitt samtycke.
Frågor som förklarats tillåtliga ska delas ut till ledamöterna och översändas till berörda institutioner.
Uppläggning
15.
Frågestunden med frågor till kommissionen kan med kommissionens samtycke delas upp i separata frågestunder med frågor till enskilda ledamöter av kommissionen.
Frågestunden med frågor till rådet kan med rådets samtycke delas upp i frågestunder med frågor till ordförandeskapet, frågor till den höge representanten för utrikes- och säkerhetspolitiken eller frågor till ordföranden för eurogruppen.
Den kan också delas in ämnesvis.
B.
Rekommendationer
(Utdrag ur parlamentets resolution av den 13 november 1986)
Europaparlamentet
1.
ser gärna att det sker en strängare tillämpning av riktlinjerna för genomförandet av frågestunden i artikel 43
Nu artikel 109.
i arbetsordningen, i synnerhet av punkt 1 i riktlinjerna beträffande tillåtlighet,
2.
i arbetsordningen, för att indela frågor för frågestunden efter ämne, men menar dock att endast de frågor på första halvan av den förteckning över frågor som ingivits till en viss sammanträdesperiod bör underkastas en sådan ämnesindelning,
3.
rekommenderar vad gäller följdfrågor, att talmannen som en allmän regel ska tillåta en följdfråga från frågeställaren och en eller högst två följdfrågor från andra ledamöter, vilka helst ska tillhöra en annan politisk grupp eller komma från en annan medlemsstat än huvudfrågeställaren; betonar att följdfrågor måste vara kortfattade och i form av frågor samt föreslår att deras längd bör begränsas till 30 sekunder,
4.
uppmanar kommissionen och rådet att i enlighet med punkt 7 i riktlinjerna se till att svaren är kortfattade och av relevans för frågans ämne.
BILAGA
II a
Riktlinjer för frågor för skriftligt besvarande enligt artiklarna 110 och 111
Punkterna 2 och 3 ska träda i kraft den första sammanträdesperiodens första dag under parlamentets sjunde valperiod.
1.
Frågor för skriftligt besvarande ska
-
falla inom den berörda institutionens kompetens- och ansvarsområde och vara av allmänt intresse,
-
vara korta och koncisa och innehålla en begriplig fråga,
-
vara skrivna på ett språk som inte innehåller stötande formuleringar,
-
beröra ämnen som inte är rent personliga.
2.
Om en fråga inte är förenlig med dessa riktlinjer ska generalsekretariatet informera frågeställaren om hur frågan kan formuleras för att den ska vara tillåtlig.
3.
Om en identisk eller liknande fråga har ingivits och besvarats under de närmast föregående sex månaderna ska generalsekretariatet till berörd institution översända en kopia av den tidigare frågan och det tillhörande svaret till frågeställaren.
Den nya frågan ska inte översändas såvida inte frågeställaren hänvisar till en betydande förändring av situationen eller efterfrågar ytterligare information.
4.
Om det i en fråga begärs fakta- eller statistikuppgifter som redan är tillgängliga för parlamentets bibliotek ska biblioteket informera ledamoten om detta; ledamoten har då möjlighet att dra tillbaka frågan.
5.
Frågor som rör relaterade ämnen får besvaras gemensamt.
BILAGA
III
Riktlinjer och allmänna principer för att fastställa vilka frågor som ska tas upp på föredragningslistan till debatter om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer enligt artikel 115
Grundläggande kriterier
1.
2.
Resolutionsförslag får omfatta högst 500 ord.
3.
De frågor ska ha företräde som avser befogenheter som Europeiska unionen har i enlighet med fördraget, under förutsättning att frågorna är av större vikt.
4.
Praktiska detaljer
5.
De grundläggande kriterier som har tillämpats för att bestämma valet av frågor som ska tas upp i debatten om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer ska meddelas parlamentet och de politiska grupperna.
Begränsning och tilldelning av talartid
6.
För att bättre utnyttja den tid som avsatts ska talmannen, efter att ha hört de politiska gruppernas ordförande, träffa en överenskommelse med rådet och kommissionen om en begränsning av talartiden för dessa två institutioners eventuella yttranden under debatten om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer.
Tidsfrist för ingivande av ändringsförslag
7.
Tidsfristen för ingivandet av ändringsförslag ska fastställas så att tillräckligt med tid finns från det att ändringsförslagen delas ut på de officiella språken till den tidpunkt som är fastställd för debatten om resolutionsförslagen, för att möjliggöra för ledamöter och politiska grupper att noggrant överväga dem.
BILAGA
IV
Genomförandebestämmelser för behandling av Europeiska unionens allmänna budget och tilläggsbudgetar
Artikel
1
Sammanträdeshandlingar
1.
Följande handlingar ska tryckas och delas ut:
a)
b)
Kommissionens eller rådets förslag om fastställandet av en ny sats.
c)
En sammanfattning av rådets överläggningar om de ändringar och ändringsförslag till budgetförslaget som parlamentet antagit.
d)
De modifieringar rådet företagit av de ändringar av budgetförslaget som parlamentet antagit.
e)
Rådets ståndpunkt beträffande fastställandet av en ny maximal procentsats.
f)
g)
2.
Dessa handlingar ska hänvisas till ansvarigt utskott.
Alla berörda utskott har rätt att yttra sig.
3.
Önskar andra utskott yttra sig ska talmannen fastställa när dessa yttranden ska ha inkommit till ansvarigt utskott.
Artikel
2
Maximal procentsats
1.
Varje ledamot kan, under förutsättning att nedanstående villkor beaktas, lägga fram och motivera förslag till beslut om fastställandet av en ny maximal procentsats.
2.
Sådana förslag är tillåtliga endast om de inges skriftligen och är undertecknade av minst 40 ledamöter, eller inges på en politisk grupps eller ett utskotts vägnar.
3.
Talmannen ska fastställa en tidsfrist för ingivandet av sådana förslag.
4.
Ansvarigt utskott ska avge ett betänkande om dessa förslag innan de behandlas i kammaren.
5.
Parlamentet ska därefter låta förslagen gå till omröstning.
Parlamentet ska fatta beslut med en majoritet av samtliga ledamöter och med en majoritet av tre femtedelar av de avgivna rösterna.
Har rådet meddelat parlamentet att det samtycker till fastställandet av en ny sats ska talmannen i kammaren förklara den nya satsen antagen.
Om så inte är fallet ska rådets ståndpunkt återförvisas till ansvarigt utskott.
Artikel
3
Behandling av budgetförslaget - första etappen
1.
Med de begränsningar som anges nedan får varje ledamot inge och framlägga:
-
Förslag till ändring av budgetförslaget.
-
Ändringsförslag till budgetförslaget.
2.
Förslag till ändringar ska för att kunna antas inges skriftligen, vara undertecknade av minst 40 ledamöter eller ingivna på en politisk grupps eller ett utskotts vägnar, ange den punkt i budgeten som de avser och respektera upprätthållandet av en balans mellan inkomster och utgifter.
Förslagen till ändringar ska omfatta alla relevanta uppgifter vad gäller de anmärkningar som berör den avsedda punkten i budgeten
Samma bestämmelser gäller för ändringsförslag.
Alla förslag till ändringar av och alla ändringsförslag till budgetförslaget måste åtföljas av en skriftlig motivering.
3.
Talmannen ska fastställa tidsfrister för ingivandet av förslag till ändringar och ändringsförslag.
Talmannen ska fastställa två tidsfrister för ingivande av förslag till ändringar och ändringsförslag: en före och en efter antagandet av betänkandet i ansvarigt utskott.
4.
Ansvarigt utskott ska yttra sig om de ingivna förslagen innan de behandlas i kammaren.
5.
Förslag till ändring av parlamentets budgetberäkning vars innehåll liknar de förslag som parlamentet redan förkastade när budgetberäkningen upprättades, ska endast behandlas om ansvarigt utskott ger sitt samtycke till detta.
6.
-
varje förslag till ändring och varje ändringsförslag,
-
varje avsnitt av budgetförslaget,
-
ett resolutionsförslag om detta budgetförslag.
7.
De artiklar, kapitel, avdelningar och avsnitt i budgetförslaget till vilka inga förslag till ändringar eller ändringsförslag har lagts fram ska anses antagna.
8.
För att godkännas måste ett förslag till ändring erhålla en majoritet av parlamentets samtliga ledamöter.
För att godkännas måste ett ändringsförslag erhålla en majoritet av de avgivna rösterna.
9.
Parlamentet ska fatta beslut med en majoritet av samtliga ledamöter och en majoritet av tre femtedelar av de avgivna rösterna.
Förkastas förslaget ska budgetförslaget i sin helhet återförvisas till ansvarigt utskott.
10.
Har parlamentet företagit ändringar av budgetförslaget eller godkänt ändringsförslag, ska det ändrade budgetförslaget eller ändringsförslagen översändas till rådet och kommissionen tillsammans med motiveringar.
Har parlamentet företagit ändringar av budgetförslaget eller godkänt ändringsförslag, ska det ändrade budgetförslaget eller ändringsförslagen översändas till rådet och kommissionen.
11.
Protokollet från det sammanträde vid vilket parlamentet yttrade sig över budgetförslaget ska översändas till rådet och kommissionen.
Artikel
4
Slutgiltigt antagande av budgeten efter första behandlingen
Artikel
5
Beaktande av rådets överläggningar - andra etappen
1.
Har rådet modifierat en eller flera av de av parlamentet antagna ändringarna ska den av rådet på detta sätt modifierade texten hänvisas till ansvarigt utskott.
2.
Varje ledamot kan, med de begränsningar som anges nedan, inge och lägga fram förslag till ändring av den av rådet modifierade texten.
3.
För att vara tillåtliga ska sådana förslag till ändringar inges skriftligen, vara undertecknade av minst 40 ledamöter eller ingivna på ett utskotts vägnar samt respektera upprätthållandet av balansen mellan inkomster och utgifter.
Förslag till ändringar är tillåtliga endast om de avser den av rådet modifierade texten.
4.
Talmannen ska fastställa en tidsfrist för ingivande av förslag till ändringar.
5.
Ansvarigt utskott ska ta ställning till den av rådet modifierade texten och yttra sig om förslagen till ändring av denna text.
6.
Parlamentet ska fatta beslut med en majoritet av samtliga ledamöter och tre femtedelar av de avgivna rösterna.
Antas förslagen till ändringar ska den av rådet modifierade texten anses förkastad.
Förkastas de ska den av rådet modifierade texten anses antagen.
7.
Rådets sammanfattning av resultatet av överläggningarna om de ändringsförslag som parlamentet har godkänt ska bli föremål för en debatt, vilken kan avslutas med omröstning om ett resolutionsförslag.
8.
Artikel
6
Avslag på hela budgetförslaget
1.
Ett utskott eller minst 40 ledamöter har rätt att, om synnerliga skäl föreligger, lägga fram ett förslag om att budgetförslaget ska avslås i sin helhet.
Ett sådant förslag är tillåtligt endast om det åtföljs av en skriftlig motivering och inges inom en av talmannen fastställd tid.
Skälen för avslag får inte vara inbördes oförenliga.
2.
Ansvarigt utskott ska yttra sig om ett sådant förslag innan det går till omröstning i kammaren.
Parlamentet ska fatta beslut med en majoritet av samtliga ledamöter och två tredjedelar av de avgivna rösterna.
Antas förslaget ska budgetförslaget i sin helhet återförvisas till rådet.
Artikel
7
Systemet med de provisoriska tolftedelarna
1.
Varje ledamot kan, med de begränsningar som anges nedan, lägga fram ett förslag till beslut som skiljer sig från det som rådet har fattat och som godkänner utgifter som överstiger den provisoriska tolftedelen, för utgifter utöver de som är en nödvändig följd av fördraget eller av rättsakter antagna på grundval av fördraget.
2.
För att vara tillåtliga ska sådana förslag till beslut inges skriftligen, vara undertecknade av minst 40 ledamöter eller ingivna av en politisk grupp eller ett utskott samt åtföljas av en motivering.
3.
Ansvarigt utskott ska yttra sig över de ingivna förslagen innan de behandlas i kammaren.
4.
Parlamentet ska fatta beslut med en majoritet av samtliga ledamöter och tre femtedelar av de avgivna rösterna.
Artikel
8
Förfarande för upprättandet av parlamentets budgetberäkning
1.
2.
3.
Detta ska i enlighet med artikel 73 i arbetsordningen ske etappvis på följande sätt:
a)
Presidiet ska upprätta ett preliminärt förslag till budgetberäkning av inkomster och utgifter (punkt 1).
b)
Utskottet med behörighet i frågor som rör budgetska upprätta ett förslag till budgetberäkning av inkomster och utgifter (punkt 2).
c)
Överläggningar ska hållas om ståndpunkterna från utskottet med behörighet i frågor som rör budget och presidiet kraftigt avviker från varandra.
BILAGA
V
Förfarande för överläggningar om och antagande av beslut om beviljande av ansvarsfrihet
Artikel
1
Handlingar
1.
Följande handlingar ska tryckas och delas ut:
a)
Resultaträkningen, analysen av den ekonomiska förvaltningen samt balansräkningen, som kommissionen översänder.
b)
Revisionsrättens årsrapport och särskilda rapporter, tillsammans med institutionernas yttranden.
c)
Revisionsrättens förklaring om räkenskapernas tillförlitlighet och de underliggande transaktionernas laglighet och korrekthet, i enlighet med artikel 248 i EG-fördraget.
d)
Rådets rekommendation.
2.
Dessa handlingar ska hänvisas till ansvarigt utskott.
Alla berörda utskott har rätt att yttra sig.
3.
Önskar andra utskott yttra sig ska talmannen fastställa när dessa yttranden ska ha inkommit till ansvarigt utskott.
Artikel
2
Behandling av betänkanden
1.
Parlamentet ska i enlighet med budgetförordningen senast den 30 april året efter det att revisionsrättens årsrapport har antagits behandla ett betänkande från ansvarigt utskott om ansvarsfrihet.
2.
Såvida annat inte föreskrivs i denna bilaga ska de bestämmelser i parlamentets arbetsordning som avser ändringsförslag och omröstningar tillämpas.
Artikel
3
Betänkandets innehåll
1.
Betänkandet om beviljande av ansvarsfrihet från ansvarigt utskott ska innehålla följande:
a)
Ett förslag till beslut om att bevilja ansvarsfrihet eller om att uppskjuta beslutet om beviljande av ansvarsfrihet (omröstning under sammanträdesperioden i april) eller ett förslag till beslut om att bevilja eller inte bevilja ansvarsfrihet (omröstning under sammanträdesperioden i oktober).
b)
Ett förslag till beslut om att avsluta räkenskaperna för gemenskapens samtliga inkomster, utgifter, tillgångar och skulder.
c)
Ett resolutionsförslag med kommentarer till det förslag till beslut som avses i punkt a ovan, däribland såväl en bedömning av kommissionens budgetförvaltning under räkenskapsåret som kommentarer beträffande effektueringen av framtida utgifter.
d)
En bilaga med en förteckning över de handlingar som erhållits från kommissionen respektive de handlingar som begärts av kommissionen, men som inte erhållits.
e)
Yttrandena från de berörda utskotten.
2.
Om ansvarigt utskott föreslår att beslutet om beviljande av ansvarsfrihet ska uppskjutas, ska i det tillhörande förslaget till resolution särskilt anges bland annat följande:
a)
anledningen till att beslutet föreslås bli uppskjutet,
b)
de ytterligare åtgärder som det förväntas att kommissionen vidtar, inbegripet en tidsfrist för dessa,
c)
de handlingar som parlamentet behöver ta del av för att på sakliga grunder kunna fatta sitt beslut.
Artikel
4
Behandling och omröstning i parlamentet
1.
Samtliga betänkanden från ansvarigt utskott som rör ansvarsfrihet ska tas upp på föredragningslistan till den sammanträdesperiod som följer på ingivandet.
2.
3.
Omröstning om förslag till beslut och förslag till resolution ska, såvida inget annat anges i artikel 5, ske i den ordning som anges i artikel 3.
4.
Parlamentet ska besluta med en majoritet av de avgivna rösterna, i enlighet med artikel 198 i EG-fördraget.
Artikel
5
Möjliga förfaranden
1.
Omröstning under sammanträdesperioden i april
I detta första skede ska betänkandet om beviljande av ansvarsfrihet innehålla ett förslag om att ansvarsfrihet beviljas eller att beslutet om beviljande av ansvarsfrihet uppskjuts.
a)
Om ett förslag om att bevilja ansvarsfrihet erhåller majoritet, innebär detta att ansvarsfrihet beviljas.
Om ett förslag om att bevilja ansvarsfrihet inte erhåller majoritet, innebär det att beviljandet av ansvarsfrihet uppskjuts och att ansvarigt utskott inom sex månader ska lägga fram ett nytt betänkande, som innehåller ett nytt förslag om att bevilja eller inte bevilja ansvarsfrihet.
b)
Om ett förslag om att uppskjuta beviljandet av ansvarsfrihet antas, ska ansvarigt utskott inom sex månader lägga fram ett nytt betänkande, som innehåller ett nytt förslag om att bevilja eller inte bevilja ansvarsfrihet.
Om ett förslag om att uppskjuta beviljandet av ansvarsfrihet inte erhåller majoritet, innebär det att ansvarsfrihet beviljas.
I detta fall ska beslutet även innebära att räkenskaperna avslutas.
Förslaget till resolution kan fortfarande gå till omröstning.
2.
Omröstning under sammanträdesperioden i oktober
I detta andra skede ska betänkandet om beviljande av ansvarsfrihet innehålla ett förslag om att bevilja eller inte bevilja ansvarsfrihet.
a.
Om ett förslag om att bevilja ansvarsfrihet erhåller majoritet, innebär detta att ansvarsfrihet beviljas.
Om ett förslag om att bevilja ansvarsfrihet inte erhåller majoritet, innebär detta att ansvarsfrihet inte beviljas.
Ett formellt förslag om avslutning av räkenskaperna för året i fråga ska läggas fram vid en senare sammanträdesperiod, då kommissionen också ska uppmanas att göra ett uttalande.
b.
Om ett förslag om att inte bevilja ansvarsfrihet erhåller majoritet, ska ett formellt förslag om avslutning av räkenskaperna för året i fråga läggas fram vid en senare sammanträdesperiod, då kommissionen också ska uppmanas att göra ett uttalande.
I detta fall ska beslutet även innebära att räkenskaperna avslutas.
Förslaget till resolution kan fortfarande gå till omröstning.
3.
Om förslaget till resolution eller förslaget om avslutning av räkenskaperna innehåller något som verkar stå i strid med parlamentets omröstning om ansvarsfrihet, får talmannen efter samråd med ordföranden i ansvarigt utskott uppskjuta omröstningen och fastställa en ny tidsfrist för ingivande av ändringsförslag.
Artikel
6
Genomförande av beslut om ansvarsfrihet
1.
Talmannen ska i enlighet med artikel 3 översända alla parlamentets beslut eller resolutioner till kommissionen och till var och en av de övriga institutionerna.
Talmannen ska se till att de offentliggörs i serien för bindande rättsakter (L-serien) i Europeiska unionens officiella tidning.
2.
Ansvarigt utskott ska minst en gång om året underrätta parlamentet om de åtgärder som institutionerna har vidtagit till följd av de i beslutet om ansvarsfrihet åtföljande kommentarerna och andra i parlamentets resolutioner ingående kommentarer som rör utgifter.
3.
På grundval av ett betänkande från utskottet med behörighet i frågor som rör budgetkontroll kan talmannen, på parlamentets vägnar och i enlighet med artikel 232 i EG-fördraget, väcka talan inför domstolen mot berörd institution för underlåtenhet att utföra de förpliktelser som anges i kommentarerna till beslutet om ansvarsfrihet eller andra resolutioner som avser genomförande av utgifter.
BILAGA
VI
Ständiga utskotts behörighetsområden
Antagen genom parlamentets beslut av den 29 januari 2004.
I.
Utskottet för utrikesfrågor
Utskottet är behörigt i frågor som rör följande områden:
1.
Den gemensamma utrikes- och säkerhetspolitiken (GUSP) och den europeiska säkerhets- och försvarspolitiken (ESFP).
Utskottet biträds i detta sammanhang av ett underutskott för säkerhet och försvar.
2.
Förbindelser med andra EU-institutioner, organ, FN och andra internationella organisationer och interparlamentariska församlingar när det gäller frågor som hör till utskottets behörighetsområde.
3.
Fördjupning av de politiska förbindelserna med tredje land, särskilt länderna i unionens omedelbara närhet, med hjälp av omfattande samarbets- och stödprogram eller internationella avtal, till exempel associerings- och partnerskapsavtal.
4.
Inledande, genomförande och avslutande av förhandlingar om europeiska staters anslutning till Europeiska unionen.
5.
Mänskliga rättigheter, skydd av minoriteter och främjandet av demokratiska värden i tredje land.
Utskottet biträds i detta sammanhang av ett underutskott för mänskliga rättigheter.
Utan att det påverkar tillämpningen av relevanta bestämmelser ska ledamöter från andra utskott och organ med ansvar på detta område inbjudas att delta i underutskottets sammanträden.
Utskottet ska samordna arbetet i de gemensamma parlamentariska kommittéerna, de parlamentariska samarbetskommittéerna och de interparlamentariska delegationerna samt i de ad hoc-delegationer och valövervakningsdelegationer som faller inom dess behörighetsområde.
II.
Utskottet för utveckling
Utskottet är behörigt i frågor som rör följande områden:
1.
2.
Partnerskapsavtal inom ramen för AVS-EU och förbindelser med relevanta organ.
3.
Utskottet ska samordna arbetet i de interparlamentariska delegationer och de ad hoc-delegationer som hör till utskottets behörighetsområde.
III.
Utskottet för internationell handel
Utskottet är behörigt i frågor som rör följande områden:
Inrättandet och genomförandet av unionens gemensamma handelspolitik och unionens externa ekonomiska förbindelser, särskilt inom följande områden:
1.
Finansiella, ekonomiska och handelsmässiga förbindelser med tredje land och regionala organisationer.
2.
Åtgärder beträffande teknisk harmonisering och standardisering på områden som omfattas av instrument inom folkrätten.
3.
Förbindelser med berörda internationella organisationer och med organisationer som främjar regional och handelsmässig integration utanför unionen.
4.
Förbindelser med Världshandelsorganisationen (WTO), däribland dess parlamentariska dimension.
Utskottet ska hålla kontakt med berörda interparlamentariska delegationer och ad hoc-delegationer när det gäller de ekonomiska och handelsmässiga aspekterna av förbindelserna med tredje land.
IV.
Budgetutskottet
Utskottet är behörigt i frågor som rör följande områden:
1.
Den fleråriga finansieringsramen för unionens inkomster och utgifter samt unionens system med egna medel.
2.
Parlamentets budgetbefogenheter, det vill säga unionens budget samt förhandling om och genomförande av interinstitutionella avtal på detta område.
3.
Parlamentets budgetberäkning i enlighet med det förfarande som fastställs i arbetsordningen.
4.
Budgeten för de decentraliserade organen.
5.
Europeiska investeringsbankens finansiella verksamhet.
6.
7.
8.
9.
Budgetförordningen, med undantag av frågor som rör budgetgenomförande, budgetförvaltning och budgetkontroll.
V.
Budgetkontrollutskottet
Utskottet är behörigt i frågor som rör följande områden:
1.
Kontroll av genomförandet av unionens och Europeiska utvecklingsfondens budget samt beslut om ansvarsfrihet som ska fattas av parlamentet, inklusive det interna förfarandet för ansvarsfrihet och alla andra åtgärder som följer av dessa beslut eller deras genomförande.
2.
Avslutande av räkenskaperna, framläggande av räkenskaperna och revision av räkenskaper och balansräkningar för Europeiska unionen, dess institutioner och alla organ som finansieras av Europeiska unionen, däribland uppförandet av de avsatta medel som ska överföras samt reglerandet av konton.
3.
Kontroll av Europeiska investeringsbankens finansiella verksamhet.
4.
Kontroll av kostnadseffektiviteten av gemenskapens olika finansieringsåtgärder vid genomförandet av unionens olika politikområden.
5.
Granskning av bedrägerier och oegentligheter vid genomförandet av unionens budget, åtgärder i syfte att förebygga och åtala sådana fall och ett allmänt tillvaratagande av unionens ekonomiska intressen.
6.
Förbindelser med revisionsrätten, utnämning av dess ledamöter och granskning av dess rapporter.
7.
Budgetförordningen, när det gäller frågor som rör budgetgenomförande, budgetförvaltning och budgetkontroll.
VI.
Utskottet för ekonomi och valutafrågor
Utskottet är behörigt i frågor som rör följande områden:
1.
Unionens ekonomiska politik och penningpolitik, Ekonomiska och monetära unionens funktion och det europeiska valuta- och finanssystemet (inklusive förbindelserna med berörda institutioner och organisationer).
2.
Den fria rörligheten för kapital och betalningar (gränsöverskridande betalningar, enhetligt betalningsområde, betalningsbalans, kapitalrörelser och in- och utlåningspolitik, kontroll av kapitalrörelser som har sitt ursprung i tredje land, åtgärder i syfte att främja unionens kapitalutförsel).
3.
Internationella valuta- och finanssystemet (inklusive förbindelserna med finansiella och monetära institutioner och organisationer).
4.
Bestämmelserna om konkurrens och statligt eller offentligt stöd.
5.
Skattebestämmelser.
6.
Reglering och övervakning av finansiella tjänster, institutioner och marknader, inklusive finansiell rapportering, revision, bokföringsbestämmelser, bolagsförvaltning och andra bolagsrättsliga frågor som särskilt rör finansiella tjänster.
VII.
Utskottet för sysselsättning och sociala frågor
Utskottet är behörigt i frågor som rör följande områden:
1.
Sysselsättningspolitik och alla aspekter av socialpolitik, exempelvis arbetsvillkor, social trygghet och socialt skydd.
2.
Åtgärder beträffande arbetsmiljö.
3.
Europeiska socialfonden.
4.
Yrkesutbildningspolitik, inklusive yrkeskvalifikationer.
5.
Fri rörlighet för arbetstagare och pensionärer.
6.
Dialogen mellan arbetsmarknadens parter.
7.
Alla former av diskriminering på arbetsplatsen och arbetsmarknaden, med undantag av könsdiskriminering.
8.
Förbindelser med följande organ:
-
Europeiskt centrum för utveckling av yrkesutbildning (Cedefop)
-
Europeiska fonden för förbättring av arbets- och levnadsvillkor
-
Europeiska yrkesutbildningsstiftelsen
-
Europeiska arbetsmiljöbyrån
Förbindelser med andra berörda EU-organ och internationella organisationer.
VIII.
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Utskottet är behörigt i frågor som rör följande områden:
1.
Miljöpolitik och miljöskyddsåtgärder, särskilt inom följande områden:
a)
Luft-, jord- och vattenföroreningar, avfallshantering och återvinning, farliga ämnen och beredningar, bullernivåer, klimatförändring och skydd av den biologiska mångfalden.
b)
En hållbar utveckling.
c)
Internationella och regionala åtgärder och avtal i syfte att skydda miljön.
d)
Återställande av miljöskador.
e)
Civilskydd.
f)
Europeiska miljöbyrån.
2.
Folkhälsa, särskilt inom följande områden:
a)
Program för särskilda åtgärder på folkhälsoområdet.
b)
Läkemedel och kosmetika.
c)
Hälsoaspekter av bioterrorism.
d)
Europeiska läkemedelsmyndigheten och Europeiska centrumet för förebyggande och kontroll av sjukdomar.
3.
Livsmedelssäkerhet, särskilt inom följande områden:
a)
Märkning av livsmedel och livsmedelssäkerhet.
b)
Veterinärlagstiftning som avser skydd mot hälsorisker för människor, kontroll av livsmedelsprodukter och system för livsmedelsproduktion med avseende på folkhälsan.
c)
Europeiska myndigheten för livsmedelssäkerhet och Kontoret för livsmedels- och veterinärfrågor.
IX.
Utskottet för industrifrågor, forskning och energi
Utskottet är behörigt i frågor som rör följande områden:
1.
Unionens industripolitik och tillämpning av ny teknik, bland annat åtgärder som rör små och medelstora företag.
2.
Unionens forskningspolitik, bland annat spridning och utnyttjande av forskningsresultat.
3.
Rymdpolitik.
4.
Verksamhet vid det gemensamma forskningscentrumet och centralbyrån för åtgärder inom kärnfysikområdet liksom JET, ITER och andra projekt inom samma område.
5.
Gemenskapsåtgärder som rör energipolitik i allmänhet, säkerhet när det gäller energiförsörjning och energieffektivitet, bland annat upprättande och utveckling av transeuropeiska nät för infrastruktur inom energisektorn.
6.
Euratomfördraget och Euratoms försörjningsbyrå, kärnsäkerhet, avveckling och avfallshantering inom kärnkraftsområdet.
7.
Informationssamhället och informationsteknik, bland annat upprättande och utveckling av transeuropeiska nät för infrastruktur inom telekommunikationssektorn.
X.
Utskottet för den inre marknaden och konsumentskydd
Utskottet är behörigt i frågor som rör följande områden:
1.
2.
Åtgärder som syftar till att identifiera och undanröja potentiella hinder för att den inre marknaden ska fungera.
3.
XI.
Utskottet för transport och turism
Utskottet är behörigt i frågor som rör följande områden:
1.
Utveckling av en gemensam politik för transporter på järnväg, landsväg och inre vattenväg samt sjöfart och luftfart, särskilt inom följande områden:
a)
3.
Posttjänster.
4.
Turism.
XII.
Utskottet för regional utveckling
Utskottet är behörigt i frågor som rör följande områden:
Regionalpolitik och sammanhållningspolitik, framför allt följande:
a)
Europeiska fonden för regional utveckling, Sammanhållningsfonden och andra instrument för Europeiska gemenskapens regionalpolitik.
b)
Bedömning av hur övrig EU-politik påverkar den ekonomiska och sociala sammanhållningen.
c)
Samordning av unionens strukturinstrument.
d)
De yttersta randområdena och öregionerna samt gränsöverskridande och interregionalt samarbete.
e)
Förbindelser med Regionkommittén, organisationer för interregionalt samarbete och med lokala och regionala myndigheter.
XIII.
Utskottet för jordbruk och landsbygdens utveckling
Utskottet är behörigt i frågor som rör följande områden:
1.
Genomförande och utveckling av den gemensamma jordbrukspolitiken.
2.
Landsbygdens utveckling, däribland verksamhet som bedrivs med hjälp av relevanta finansiella instrument.
3.
Lagstiftning om
a)
veterinärmedicinska frågor och växtskyddsfrågor samt djurfoder, förutsatt att åtgärderna inte syftar till att skydda mot risker för människans hälsa,
b)
djuruppfödning och djurskydd.
4.
Förbättring av kvaliteten på jordbruksprodukter.
5.
Tillgång på jordbruksråvaror.
6.
Gemenskapens växtsortsmyndighet.
7.
Skogsbruk.
XIV.
Fiskeriutskottet
Utskottet är behörigt i frågor som rör följande områden:
1.
Den gemensamma fiskeripolitiken, dess utveckling och förvaltning.
2.
Bevarande av fiskbestånden.
3.
Den gemensamma organisationen av marknaden för fiskeriprodukter.
4.
Strukturpolitik inom fiskeri- och vattenbrukssektorerna, däribland de finansiella instrumenten för utveckling av fisket.
5.
Internationella fiskeriavtal.
XV.
Utskottet för kultur och utbildning
Utskottet är behörigt i frågor som rör följande områden:
1.
Europeiska unionens kulturella aspekter, framför allt
a)
förbättring av kunskaperna om och spridning av kultur,
b)
skydd och främjande av kulturell och språklig mångfald,
c)
bevarande och skydd av kulturarvet, kulturutbyte och konstnärligt skapande.
2.
Unionens utbildningspolitik, däribland den högre Europautbildningen, främjande av systemet med Europaskolor och livslångt lärande.
3.
Audiovisuell politik och informationssamhällets kultur- och utbildningsaspekter.
4.
Ungdomspolitik och utveckling av en politik för idrott och fritid.
5.
Informations- och mediepolitik.
6.
Samarbete med tredje land på kultur- och utbildningsområdena och förbindelser med berörda internationella organisationer och institutioner.
XVI.
Utskottet för rättsliga frågor
Utskottet är behörigt i frågor som rör följande områden:
1.
Tolkning och tillämpning av EU-rätten, unionens rättsakters överensstämmelse med primärrätten, inbegripet valet av rättslig grund för rättsakterna och respekten för subsidiaritets- och proportionalitetsprinciperna.
2.
Tolkning och tillämpning av folkrätten, i den utsträckning Europeiska unionen berörs.
3.
Förenkling av gemenskapsrätten, särskilt förslag till kodifiering av gemenskapslagstiftningen.
4.
Rättsligt skydd för parlamentets rättigheter och befogenheter, särskilt vid parlamentets deltagande i processer inför domstolen och förstainstansrätten.
5.
6.
Miljöansvar och påföljder vid miljöbrott.
7.
Etiska frågor i samband med ny teknik vid tillämpning av förfarandet med associerade utskott med berörda utskott.
8.
Ledamotsstadgan och tjänsteföreskrifterna för Europeiska gemenskapernas personal.
9.
Privilegier och immunitet samt granskning av bevis för nyvalda ledamöter.
10.
Domstolens organisation och ställning.
11.
XVII.
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Utskottet är behörigt i frågor som rör följande områden:
1.
Skyddet inom unionens territorium av de medborgarliga rättigheter, de mänskliga rättigheter och de grundläggande rättigheter, inklusive skydd av minoriteter, som slås fast i fördragen och Europeiska unionens stadga om de grundläggande rättigheterna.
2.
Åtgärder som krävs för att bekämpa alla former av diskriminering, med undantag av diskriminering på grund av kön eller diskriminering på arbetsplatsen och på arbetsmarknaden.
3.
Lagstiftning om öppenhet och skydd för enskilda när det gäller behandling av personuppgifter.
4.
Förverkligande och fördjupning av ett område med frihet, säkerhet och rättvisa, framför allt följande:
5.
Europeiska centrumet för kontroll av narkotika och narkotikamissbruk och Europeiska centrumet för övervakning av rasism och främlingsfientlighet, Europol, Eurojust och Cepol och andra organ och kontor inom samma område.
6.
XVIII.
Utskottet för konstitutionella frågor
Utskottet är behörigt i frågor som rör följande områden:
1.
Institutionella aspekter av den europeiska integrationen, särskilt i samband med förberedande och genomförande av konvent och regeringskonferenser.
2.
Genomförande av EU-fördraget och utvärdering av hur det fungerar.
3.
De institutionella konsekvenserna av unionens utvidgningsförhandlingar.
4.
5.
Enhetlig valordning.
6.
7.
Fastslående av att det finns en klar risk för att en medlemsstat allvarligt och ihållande åsidosätter principer som är gemensamma för medlemsstaterna.
8.
Tolkning och tillämpning av arbetsordningen och förslag till ändring av denna.
XIX.
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
Utskottet är behörigt i frågor som rör följande områden:
1.
Fastställande, främjande och skydd av kvinnors rättigheter i unionen och gemenskapsåtgärder i samband med detta.
2.
Främjande av kvinnors rättigheter i tredje land.
3.
Politik för lika möjligheter, däribland lika möjlighet för kvinnor och män på arbetsmarknaden och lika behandling av kvinnor och män på arbetsplatsen.
4.
Undanröjande av alla former av könsdiskriminering.
5.
Genomförande och vidareutveckling av jämställdhetsperspektivet i alla sektorer (”gender mainstreaming”).
6.
Uppföljning och genomförande av internationella avtal och konventioner om kvinnors rättigheter.
7.
Informationspolitik med avseende på kvinnor.
XX.
1.
Framställningar.
2.
Förbindelser med Europeiska ombudsmannen.
BILAGA
VII
Sekretessbelagda handlingar och känslig information
A
Behandling av sekretessbelagda handlingar som förelagts parlamentet
Förfarande för behandling av sekretessbelagda handlingar som förelagts Europaparlamentet
1.
Som sekretessbelagda handlingar betraktas handlingar och upplysningar som kan undantas från allmänhetens tillgång av skäl som anges i artikel 4 i Europaparlamentets och rådets förordning (EG) nr 1049/2001, inklusive känsliga handlingar enligt artikel 9 i nämnda förordning.
När sekretessbelagda handlingar föreläggs parlamentet under skydd av sekretess, skall behörigt parlamentsutskotts ordförande omedelbart tillämpa sekretessförfarandet i punkt 3 nedan.
Närmare bestämmelser om skyddet av sekretessbelagda handlingar skall antas i kammaren på grundval av ett förslag från presidiet och skall fogas till arbetsordningen som bilaga.
Bestämmelserna skall beakta kontakter med kommissionen och rådet.
2.
Alla parlamentets utskott har rätt att på skriftlig eller muntlig begäran av en av sina ledamöter tillämpa sekretessförfarandet beträffande upplysningar eller handlingar ledamoten angivit.
En majoritet av två tredjedelar av de närvarande ledamöterna krävs för ett beslut om att tillämpa sekretessförfarande.
3.
Har utskottets ordförande väl förklarat att sekretessförfarandet skall tillämpas har endast utskottets ledamöter samt ett strängt begränsat antal tjänstemän och sakkunniga, vilka på förhand utsetts av ordföranden, rätt att närvara vid förhandlingarna.
Handlingarna skall numreras och delas ut vid sammanträdets början och samlas in vid dess slut.
Inga anteckningar får föras och fotokopiering är inte tillåten.
Protokollet från sammanträdet skall inte redogöra för behandlingen av en punkt som behandlas under sekretess.
Endast ett eventuellt beslut får föras till protokollet.
4.
Tre ledamöter av ett utskott som tillämpat sekretessförfarandet kan begära en prövning av brott mot tystnadsplikten samt att detta tas upp på föredragningslistan.
En majoritet av utskottets ledamöter kan besluta att brott mot tystnadsplikten skall tas upp på föredragningslistan till det första sammanträde som följer på att ordföranden mottagit en sådan begäran.
5.
Påföljder: Vid fall av överträdelser skall utskottets ordförande, efter att ha hört vice ordförandena, fastställa ett motiverat beslut om lämpliga påföljder (prickning, tillfällig uteslutning ur utskottet, förlängd eller permanent uteslutning ur utskottet).
Berörd ledamot har rätt att inkomma med besvär mot detta beslut utan att det har upphävande verkan.
Detta besvär skall gemensamt prövas av talmanskonferensen och berört utskotts presidium.
Beslut skall fattas med majoritet av de avlagda rösterna och kan inte överklagas.
Kan det styrkas att en tjänsteman inte har respekterat tystnadsplikten skall de i tjänsteföreskrifterna fastställda påföljderna tillämpas.
B
Parlamentets tillgång till känslig information om säkerhets- och försvarspolitiken
Interinstitutionellt avtal av den 20 november 2002 mellan Europaparlamentet och rådet om Europaparlamentets tillgång till känslig information i rådet om säkerhets- och försvarspolitiken
EGT C 298, 30.11.2002, s.
1.
I artikel 21 i Fördraget om Europeiska unionen anges det att rådets ordförandeskap skall höra Europaparlamentet om de viktigaste aspekterna och de grundläggande valmöjligheterna när det gäller den gemensamma utrikes- och säkerhetspolitiken och se till att vederbörlig hänsyn tas till Europaparlamentets synpunkter.
I samma artikel anges det också att rådets ordförandeskap och kommissionen regelbundet skall hålla Europaparlamentet informerat om utvecklingen av den gemensamma utrikes- och säkerhetspolitiken.
En mekanism bör införas för att se till att dessa principer tillämpas på detta område.
(2)
Enligt artikel 9.7 i Europaparlamentets och rådets förordning (EG) nr 1049/2001 av den 30 maj 2001 om allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar
EGT L 145, 31.5.2001, s.
43.
skall rådet informera Europaparlamentet om känsliga handlingar som avses i artikel 9.1 i den förordningen, i enlighet med en ordning om vilken institutionerna skall komma överens.
(4)
Genom detta interinstitutionella avtal bör Europaparlamentet få en behandling som överensstämmer med bästa praxis i medlemsstaterna.
EUROPAPARLAMENTET OCH RÅDET HAR ENATS OM FÖLJANDE.
1.
Räckvidd
1.1
Detta interinstitutionella avtal rör Europaparlamentets tillgång till känslig information, dvs. information som klassificeras TRÈS SECRET/TOP SECRET, SECRET eller CONFIDENTIEL, oberoende av dess ursprung, medium eller hur slutförd den är, som innehas av rådet inom säkerhets- och försvarspolitiken samt hantering av handlingar med denna klassificering.
1.2
Information med ursprung i en tredje stat eller en internationell organisation skall överlämnas efter godkännande från den staten eller organisationen.
Om information med ursprung i en medlemsstat överlämnas till rådet utan annan uttrycklig begränsning av dess spridande till andra institutioner än dess klassificering skall bestämmelserna i avsnitt 2 och 3 i detta interinstitutionella avtal tillämpas.
I övrigt skall sådan information överlämnas med godkännande av medlemsstaten i fråga.
I fall då överlämnande av information från en tredje stat, en internationell organisation eller en medlemsstat vägras, skall rådet ange skälen till detta.
1.3
Bestämmelserna i detta interinstitutionella avtal skall tillämpas i enlighet med tillämplig lag och utan att det påverkar tillämpningen av Europaparlamentets, rådets och kommissionens beslut 95/167/EG, Euratom, EKSG av den 19 april 1995 om närmare föreskrifter för utövandet av Europaparlamentets undersökningsrätt
EGT L 113, 19.5.1995, s.
2.
och utan att det påverkar tillämpningen av befintliga bestämmelser, särskilt det interinstitutionella avtalet av den 6 maj 1999 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och förbättring av budgetförfarandet
EGT C 172, 18.6.1999, s.
1.
.
2.
Allmänna bestämmelser
2.1
De två institutionerna skall agera i enlighet med sina ömsesidiga skyldigheter om lojalt samarbete och i en anda av ömsesidigt förtroende samt i enlighet med relevanta fördragsbestämmelser.
Vid överlämnande och hantering av den information som omfattas av detta interinstitutionella avtal måste hänsyn tas till de intressen som klassificeringen är avsedd att skydda och i synnerhet allmänhetens intresse beträffande säkerheten och försvaret av Europeiska unionen eller en eller flera av dess medlemsstater eller militär och icke-militär krishantering.
2.2
Rådets ordförandeskap eller generalsekreteraren/höge representanten skall på begäran av en av de personer som avses i punkt 3.1 nedan med all nödvändig skyndsamhet informera om innehållet i varje känslig information som krävs för utövande av de befogenheter som har tilldelats Europaparlamentet genom fördraget om Europeiska unionen på det område som omfattas av detta interinstitutionella avtal, med beaktande av allmänhetens intresse i frågor som rör säkerheten för och försvaret av Europeiska unionen eller en eller flera av dess medlemsstater eller militär och icke-militär krishantering samt i enlighet med bestämmelserna i avsnitt 3 nedan.
3.
Bestämmelser om tillgång till och hantering av känslig information
3.1
Inom ramen för detta interinstitutionella avtal får Europaparlamentets ordförande eller ordföranden för Europaparlamentets utskott för utrikesfrågor, mänskliga rättigheter, gemensam säkerhet och försvarspolitik begära att rådets ordförandeskap eller generalsekreteraren/höge representanten skall lämna information till detta utskott om utvecklingen av den europeiska säkerhets- och försvarspolitiken, inklusive känslig information, vilken omfattas av punkt 3.3.
3.2
I händelse av en kris eller på begäran av Europaparlamentets ordförande eller av ordföranden för utskottet för utrikesfrågor, mänskliga rättigheter, gemensam säkerhet och försvarspolitik skall denna information lämnas snarast möjligt.
3.3
Europaparlamentets ordförande och en särskild kommitté under ordförandeskap av ordföranden för utskottet för utrikesfrågor, mänskliga rättigheter, gemensam säkerhet och försvarspolitik, sammansatt av fyra medlemmar utsedda av talmanskonferensen, skall inom denna ram informeras av rådets ordförandeskap eller generalsekreteraren/höge representanten om innehållet i den känsliga informationen om detta krävs för utövande av de befogenheter som har tilldelats Europaparlamentet enligt fördraget om Europeiska unionen inom det område som omfattas av detta interinstitutionella avtal.
Europaparlamentets ordförande och den särskilda kommittén får begära att få del av dokumenten i fråga i rådets lokaler.
Om det är lämpligt och möjligt med beaktande av informationens eller dokumentens art och innehåll, skall dessa göras tillgängliga för Europaparlamentets ordförande som skall välja ett av följande alternativ:
a)
Information till ordföranden för utskottet för utrikesfrågor, mänskliga rättigheter, gemensam säkerhet och försvarspolitik.
b)
Tillgång till information som begränsas till endast medlemmar av utskottet för utrikesfrågor, mänskliga rättigheter, gemensam säkerhet och försvarspolitik.
c)
Behandling inom lyckta dörrar i utskottet för utrikesfrågor, mänskliga rättigheter, gemensam säkerhet och försvarspolitik i enlighet med bestämmelser som kan variera beroende på sekretessgraden i fråga.
d)
Överlämnande av dokument i vilka information har strukits med hänsyn till den sekretessgrad som krävs.
Dessa alternativ skall inte tillämpas om känslig information är klassificerad som TRÈS SECRET/TOP SECRET.
När det gäller dokument som klassificerats som SECRET eller CONFIDENTIEL skall Europaparlamentets ordförandes val av ett av dessa alternativ i förväg överenskommas med rådet.
Informationen eller dokumenten i fråga får inte offentliggöras eller lämnas vidare till någon annan mottagare.
4.
Slutbestämmelser
4.1
Europaparlamentet och rådet skall vart för sig vidta alla nödvändiga åtgärder för att säkerställa tillämpningen av detta interinstitutionella avtal, inklusive de åtgärder som krävs för säkerhetsundersökningen av de berörda personerna.
4.2
De två institutionerna är villiga att diskutera jämförbara interinstitutionella avtal om sekretessbelagd information inom andra av rådets verksamhetsområden, varvid skall gälla att bestämmelserna i detta interinstitutionella avtal inte blir prejudicerande för unionens eller gemenskapens andra verksamhetsområden och inte påverkar innehållet i några andra interinstitutionellt avtal.
4.3
Detta interinstitutionella avtal skall ses över efter två år på begäran av endera av de två institutionerna med beaktande av de erfarenheter som erhållits vid tillämpningen av detsamma.
Bilaga
Det interinstitutionella avtalet skall tillämpas i enlighet med relevanta tillämpliga bestämmelser, särskilt i överensstämmelse med principen att upphovsmannens samtycke krävs för överlämnande av sekretessbelagd information enligt punkt 1.2.
När medlemmarna i Europaparlamentets särskilda kommitté får tillgång till känsliga handlingar skall detta ske i en säkrad lokal på rådet.
Det interinstitutionella avtalet skall träda i kraft efter det att Europaparlamentet har antagit interna säkerhetsåtgärder som överensstämmer med de principer som anges i punkt 2.1 och som är jämförbara med de åtgärder som tillämpas på de andra institutionerna, i syfte att garantera en likvärdig skyddsnivå för den känsliga informationen i fråga.
C
Genomförandet av det interinstitutionella avtalet om Europaparlamentets tillgång till känslig information om säkerhets- och försvarspolitiken
Europaparlamentets beslut av den 23 oktober 2002 om genomförandet av det interinstitutionella avtalet om Europaparlamentets tillgång till känslig information i rådet om säkerhets- och försvarspolitiken
EGT C 298, 30.11.2002, s.
4.
.
EUROPAPARLAMENTET HAR BESLUTAT FÖLJANDE
med beaktande av artikel 9, särskilt punkterna 6 och 7, i Europaparlamentets och rådets förordning (EG) nr 1049/2001 av den 30 maj 2001 om allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar
EGT L 145, 31.5.2001, s.
43.
,
med beaktande av arbetsordningens bilaga VII, del A, punkt 1,
med beaktande av artikel 20 i presidiets beslut av den 28 november 2001 om allmänhetens tillgång till Europaparlamentets handlingar
EGT C 374, 29.12.2001, s.
1.
,
med beaktande av det interinstitutionella avtalet mellan Europaparlamentet och rådet om Europaparlamentets tillgång till känslig information från rådet på säkerhets- och försvarspolitikens område,
med beaktande av presidiets förslag och av följande skäl:
Viss information om säkerhets- och försvarspolitiken som är belagd med sträng sekretess är av särskild natur och har ett särskilt känsligt innehåll.
Rådet är förpliktigat att tillhandahålla Europaparlamentet information om känsliga handlingar i enlighet med vad som överenskommits mellan institutionerna.
De av Europaparlamentets ledamöter som ingår i den särskilda kommitté som inrättas genom det interinstitutionella avtalet bör genomgå en säkerhetsprövning för att få tillgång till känslig information i enlighet med principen att de behöver ha tillgång till uppgifterna för tjänsteutövningen.
Det är nödvändigt att införa särskilda arrangemang för att ta emot, hantera och kontrollera känslig information från rådet, medlemsstaterna, tredje länder eller internationella organisationer.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Syftet med detta beslut är att anta kompletterande åtgärder som är nödvändiga för att genomföra det interinstitutionella avtalet om Europaparlamentets tillgång till känslig information från rådet på säkerhets- och försvarspolitikens område.
Artikel 2
Europaparlamentets begäran om tillgång till känslig information från rådet skall behandlas av rådet i enlighet med dess bestämmelser.
När de begärda handlingarna har upprättats av andra institutioner, medlemsstater, tredje länder eller internationella organisationer, översänds handlingarna när dessa gett sitt medgivande.
Artikel 3
Europaparlamentets talman skall ansvara för genomförandet av detta interinstitutionella avtal inom parlamentet.
Talmannen skall för detta ändamål vidta alla nödvändiga åtgärder för att se till att den information som mottas direkt från rådets ordförande eller generalsekreterare/höge representant eller som inhämtas i samband med att känsliga handlingar konsulteras i rådets lokaler omfattas av sekretess.
Artikel 4
När Europaparlamentets talman eller ordföranden för utskottet för utrikesfrågor, mänskliga rättigheter, gemensam säkerhet och försvarspolitik uppmanar rådets ordförandeskap eller generalsekreterare/höge representant att tillhandahålla känslig information till den särskilda kommitté som inrättas genom det interinstitutionella avtalet, skall denna information tillhandahållas snarast.
Europaparlamentet skall utrusta ett rum särskilt för detta ändamål.
Valet av rum skall göras så att en likvärdig skyddsnivå garanteras som den som fastställs för denna typ av möten i rådets beslut 2001/264/EG av den 19 mars 2001 om antagande av rådets säkerhetsbestämmelser
EGT L 101, 11.4.2001, s.
1.
.
Artikel 5
Informationsmötet, som leds av Europaparlamentets talman eller av ovannämnda utskottsordförande, skall hållas inom stängda dörrar.
Med undantag för de fyra ledamöter som utses av talmanskonferensen skall enbart de tjänstemän som på grund av sina arbetsuppgifter eller tjänsteåligganden genomgått säkerhetsprövning och beviljats tillstånd, få tillträde till möteslokalen under förutsättning att de behöver ha tillgång till uppgifterna för tjänsteutövningen.
Artikel 6
När Europaparlamentets talman eller ordföranden i ovannämnda utskott beslutar att begära att få konsultera handlingar med känslig information, skall handlingarna i enlighet med punkt 3.3 i ovannämnda interinstitutionella avtal konsulteras i rådets lokaler.
Handlingarna skall konsulteras på plats i de versioner som finns tillgängliga.
Artikel 7
De ledamöter av Europaparlamentet som skall delta i informationsmöten eller ta del av känsliga handlingar skall genomgå ett liknande säkerhetsprövningsförfarande som medlemmarna av rådet och ledamöterna av kommissionen.
I detta avseende skall Europaparlamentets talman vidta nödvändiga åtgärder vid de behöriga nationella myndigheterna.
Artikel 8
De tjänstemän som skall få kännedom om känslig information skall genomgå säkerhetsprövning i enlighet med de bestämmelser som fastställts för övriga institutioner.
De tjänstemän som genomgått en sådan säkerhetsprövning, under förutsättning att de behöver ha tillgång till uppgifterna för tjänsteutövningen, skall kunna få delta i ovannämnda informationsmöten eller få kännedom om deras innehåll.
Generalsekreteraren skall bevilja tillstånd till detta efter att ha inhämtat yttranden från de nationella behöriga myndigheterna i medlemsstaterna och på grundval av de säkerhetsprövningar som samma myndigheter genomfört.
Artikel 9
Den information som erhålls vid dessa möten eller när handlingar konsulteras i rådets lokaler får inte röjas, spridas eller mångfaldigas, vare sig fullständigt eller delvis, i någon som helst form.
Det är inte heller tillåtet att göra någon form av upptagning av den känsliga information som rådet tillhandahållit.
Artikel 10
De ledamöter av Europaparlamentet som av talmanskonferensen utsetts för att få tillgång till känslig information skall ha tystnadsplikt.
Vid brott mot tystnadsplikten skall ledamöterna i den särskilda kommittén bytas ut mot en annan ledamot som talmanskonferensen utser.
En ledamot som brutit mot tystnadsplikten kan, innan han eller hon utesluts från den särskilda kommittén, höras av talmanskonferensen som då skall hålla ett särskilt sammanträde inom stängda dörrar.
Den ledamot som gjort sig skyldig till informationsläckan kan, i förekommande fall, förutom att bli utesluten ur den särskilda kommittén, även bli föremål för rättsliga åtgärder i enlighet med gällande lagstiftning.
Artikel 11
De tjänstemän som på vederbörligt sätt genomgått säkerhetsprövning och som skall få tillgång till känslig information på grundval av principen att de behöver ha tillgång till uppgifterna för tjänsteutövningen skall ha tystnadsplikt.
Eventuella brott mot tystnadsplikten skall bli föremål för en utredning som leds av Europaparlamentets talman och, i förekommande fall, ett disciplinförfarande i enlighet med tjänsteföreskrifterna.
Om det blir fråga om rättsliga åtgärder skall talmannen vidta de åtgärder som krävs för att de behöriga nationella myndigheterna skall kunna inleda lämpliga förfaranden.
Artikel 12
Presidiet skall vara behörigt att genomföra de eventuella anpassningar, ändringar eller tolkningar som kan bli nödvändiga för att tillämpa detta beslut.
Artikel 13
Detta beslut återges i Europaparlamentets arbetsordning och träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
BILAGA
VIII
Närmare föreskrifter för utövandet av Europaparlamentets undersökningsrätt
Europaparlamentets, rådets och kommissionens beslut av den 19 april 1995 om närmare föreskrifter för utövandet av Europaparlamentets undersökningsrätt
EGT L 113, 19.5.1995, s.
2.
Europaparlamentet, rådet och kommissionen har i samförstånd fattat detta beslut
med beaktande av Fördraget om upprättandet av Europeiska kol- och stålgemenskapen, särskilt artikel 20b,
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 193,
Det bör fastställas närmare föreskrifter för Europaparlamentets utövande av undersökningsrätten med hänsyn till bestämmelserna i Fördragen om upprättandet av Europeiska gemenskaperna.
De tillfälliga undersökningskommittéerna måste ha nödvändiga medel för att fullgöra sina uppgifter; i detta avseende är det viktigt att medlemsstaterna samt Europeiska gemenskapernas institutioner och organ vidtar alla åtgärder som kan underlätta fullgörandet av dessa uppgifter.
Sekretess och konfidentiell behandling i samband med de tillfälliga undersökningskommittéernas arbete måste säkerställas.
Föreskrifterna för utövandet av undersökningsrätten kan på begäran av en av de tre institutionerna ses över efter utgången av Europaparlamentets valperiod mot bakgrund av gjorda erfarenheter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE
Artikel
1
Närmare föreskrifter om utövandet av Europaparlamentets undersökningsrätt skall fastställas i detta beslut i enlighet med artikel 20b i EKSG-fördraget, artikel 193 i EG-fördraget och artikel 107b i Euratomfördraget.
Artikel
2
1.
Europaparlamentet kan vid fullgörandet av sina uppgifter på de villkor och inom de gränser som fastställs i de fördrag som anges i artikel 1 på begäran av en fjärdedel av sina ledamöter tillsätta en tillfällig undersökningskommitté för att undersöka påstådda fel eller missförhållanden vid tillämpningen av gemenskapsrätten, oavsett om dessa skulle ha begåtts av en gemenskapsinstitution, ett gemenskapsorgan, en offentlig myndighet i en medlemsstat eller av personer som enligt gemenskapsrätten är bemyndigade att tillämpa denna.
Europaparlamentet skall fastställa de tillfälliga undersökningskommittéernas sammansättning samt närmare regler för deras arbetssätt.
Beslutet om att tillsätta en tillfällig undersökningskommitté, i vilket särskilt skall anges kommitténs syfte och tidsfristen för att överlämna dess rapport, skall offentliggöras i Europeiska gemenskapernas officiella tidning.
2.
Den tillfälliga undersökningskommittén skall fullgöra sina uppgifter i enlighet med de befogenheter fördragen tilldelat gemenskapsinstitutionerna och gemenskapsorganen.
Medlemmarna av den tillfälliga undersökningskommittén och varje annan person som i sin tjänsteutövning får kännedom om sakförhållanden, information, kunskap, dokument eller annat där sekretess gäller i enlighet med en medlemsstats eller gemenskapsinstitutions bestämmelser är skyldig att bibehålla denna sekretess gentemot obehöriga personer och allmänheten, även efter att deras tjänsteutövning har upphört.
Förhör och avgivande av vittnesmål skall vara offentliga.
På begäran av en fjärdedel av medlemmarna i den tillfälliga undersökningskommittén, eller på begäran av gemenskapernas myndigheter eller nationella myndigheter, eller om den tillfälliga undersökningkommittén har förelagts uppgifter för vilka sekretess gäller, skall förhandlingarna ske bakom stängda dörrar.
Vittnen och sakkunniga har rätt att avge utlåtande eller vittnesmål bakom stängda dörrar.
3.
En tillfällig undersökningskommitté får inte utreda en sak som är föremål för rättslig prövning vid en gemenskapsinstans eller en nationell instans, så länge som den rättsliga prövningen inte är avslutad.
Inom en tidsfrist på två månader, antingen efter offentliggörandet i enlighet med punkt 1, eller efter att kommissionen har informerats om att undersökningskommittén har förelagts ett påstående om att en medlemsstat har överträtt gemenskapsrätten, får kommissionen underrätta Europaparlamentet om att en sak som är hänskjuten till en tillfällig undersökningskommitté är underkastad ett förberedande gemenskapsförfarande; i detta fall skall den tillfälliga undersökningskommittén vidta alla nödvändiga åtgärder för att kommissionen fullt ut skall kunna utöva de befogenheter den tilldelats i enlighet med fördragen.
4.
Den tillfälliga undersökningskommittén skall upplösas när den har överlämnat sin rapport inom den tidsfrist som fastställdes när den tillsattes, eller senast vid utgången av en tidsfrist på maximalt tolv månader från den dag då den tillsattes, eller, under alla omständigheter, vid utgången av valperioden.
Europaparlamentet kan efter ett motiverat beslut två gånger förlänga tolvmånadersfristen med tre månader.
Detta beslut skall offentliggöras i Europeiska gemenskapernas officiella tidning.
5.
En tillfällig undersökningskommitté får inte tillsättas eller tillsättas på nytt angående en sak som redan varit föremål för undersökning av en tillfällig undersökningskommitté förrän det har gått minst tolv månader efter överlämnandet av denna undersöknings rapport, eller efter det att uppgiften har avslutats, och endast under förutsättning att nya omständigheter har framkommit.
Artikel
3
1.
Den tillfälliga undersökningskommittén skall företa de undersökningar som är nödvändiga för att undersöka påstådda överträdelser eller missförhållanden vid tillämpningen av gemenskapsrätten enligt nedanstående villkor.
2.
Den tillfälliga undersökningskommittén kan anmoda en gemenskapsinstitution, ett gemenskapsorgan eller en medlemsstats regering att utse en av sina ledamöter eller medlemmar att delta i kommitténs arbete.
3.
På motiverad begäran av den tillfälliga undersökningskommittén skall berörda medlemsstater och gemenskapsinstitutioner eller gemenskapsorgan utse en tjänsteman eller annan anställd som de bemyndigar att uppträda inför den tillfälliga undersökningskommittén, såvida inte sekretess eller hänsyn till nationell och allmän säkerhet på grund av nationell lagstiftning eller gemenskapslagstiftning utgör hinder för detta.
De aktuella tjänstemännen eller andra anställda skall yttra sig på sin regerings eller institutions vägnar och efter instruktion från dessa.
De skall fortsätta att vara bundna av de förpliktelser som följer av de för dem gällande föreskrifterna.
4.
Medlemsstaternas myndigheter och gemenskapsinstitutionerna eller gemenskapsorganen skall, antingen på begäran av den tillfälliga undersökningskommittén eller på eget initiativ, tillhandahålla den tillfälliga undersökningskommittén de handlingar som är nödvändiga för att den skall kunna utföra sitt arbete om de inte på grund av sekretess eller av hänsyn till allmän och nationell säkerhet är förhindrade att göra detta på grund av medlemstaternas och gemenskapernas lagar och föreskrifter.
5.
Bestämmelserna i punkterna 3 och 4 skall inte påverka andra nationella bestämmelser som hindrar en tjänsteman att uppträda eller utlämning av handlingar.
Hinder som uppstår med hänsyn till sekretess, offentlig eller nationell säkerhet eller på grund av bestämmelserna i första stycket, skall anmälas till Europaparlamentet av en företrädare som är behörig att binda den berörda medlemsstatens regering eller institution.
6.
Gemenskapsinstitutionerna eller gemenskapsorganen får inte tillhandahålla den tillfälliga undersökningskommittén handlingar från en medlemsstat utan att först ha informerat den berörda medlemsstaten om detta.
De får inte överlämna handlingar som omfattas av punkt 5 till den tillfälliga undersökningskommittén utan att först ha inhämtat den berörda medlemsstatens samtycke.
7.
Bestämmelserna i punkterna 3-5 skall tillämpas på fysiska och juridiska personer som är bemyndigade enligt gemenskapsrätten att tillämpa denna.
8.
Den tillfälliga undersökningskommittén kan begära att varje annan person avlägger vittnesmål inför kommittén i den mån det är nödvändigt för fullgörandet av dess uppgifter.
Om omnämnandet av en person i förbindelse med en undersökning kan åsamka skada skall den tillfälliga undersökningskommittén underrätta personen om detta samt höra personen ifall denne så begär.
Artikel
4
1.
De upplysningar som den tillfälliga undersökningskommittén samlar in får endast användas för att fullgöra dess uppgifter.
Upplysningarna får inte offentliggöras om de innehåller sekretessbelagda uppgifter eller uppgifter av konfidentiell natur eller om personer härigenom namnges.
Europaparlamentet skall anta de administrativa och reglementariska bestämmelser som behövs för att säkerställa sekretess och konfidentiell behandling i förbindelse med de tillfälliga undersökningskommittéernas arbete.
2.
Den tillfälliga undersökningskommitténs rapport skall föreläggas Europaparlamentet som kan bestämma att rapporten skall offentliggöras, om inte annat följer av bestämmelserna i punkt 1.
3.
Europaparlamentet får överlämna de rekommendationer som det har antagit på grundval av den tillfälliga undersökningskommitténs rapport till gemenskapsinstitutionerna eller gemenskapsorganen eller medlemsstaterna.
Dessa skall dra de slutsatser därav som de anser lämpliga.
Artikel
5
Alla meddelanden till medlemsstaternas nationella myndigheter för genomförandet av detta beslut skall gå via medlemsstaternas fasta representationer vid Europeiska unionen.
Artikel
6
På begäran av Europaparlamentet, rådet eller kommissionen kan ovanstående bestämmelser ses över mot bakgrund av gjorda erfarenheter, från det att Europaparlamentets valperiod har löpt ut.
Artikel
7
Detta beslut skall träda i kraft den dag det offentliggörs i Europeiska gemenskapernas officiella tidning.
BILAGA
IX
Artikel
1
Passerkort
1.
Passerkortet ska utgöras av ett inplastat kort med ett fotografi av innehavaren, innehavarens för- och efternamn samt namnet på det företag, den organisation eller den person som innehavaren arbetar för.
Innehavare av passerkort ska alltid bära kortet synligt inom alla parlamentets lokaler.
Underlåtenhet att göra detta kan leda till att kortet dras in.
Passerkortet ska särskiljas i form och färg från de passerkort som utfärdas till tillfälliga besökare.
2.
I det fall en ledamot ifrågasätter en representants eller en lobbygrupps verksamhet ska frågan hänvisas till kvestorerna, som ska göra en utredning och avgöra om passerkortet ifråga får behållas eller ska dras in.
3.
Passerkort ger under inga omständigheter innehavaren rätt att närvara vid andra av parlamentets eller dess organs sammanträden än de som förklarats öppna för allmänheten och ger i detta fall inte innehavaren rätt till undantag från de regler om tillträde som gäller för alla övriga unionsmedborgare.
Artikel
2
Assistenter
1.
Vid början av varje mandatperiod ska kvestorerna besluta om det högsta antal assistenter som kan registreras av varje ledamot.
Registrerade assistenter ska när de tillträder sin tjänst avge en skriftlig förklaring beträffande sin yrkesverksamhet och andra uppdrag och verksamheter som de utför mot ersättning.
2.
Assistenterna ska ha tillträde till parlamentet enligt samma villkor som personal vid generalsekretariatet eller de politiska grupperna.
3.
Artikel
3
Ordningsregler
1.
a)
rätta sig efter bestämmelserna i artikel 9 i arbetsordningen och denna bilaga,
b)
uppge vems eller vilkas intressen de företräder vid kontakt med parlamentets ledamöter, ledamöternas medarbetare eller tjänstemän vid parlamentet,
c)
inte försöka få tag i information på ett oärligt sätt,
d)
inte uppge någon formell anknytning till parlamentet i sina förbindelser med tredje man,
e)
inte i vinstsyfte sprida handlingar som erhållits från parlamentet till tredje man,
f)
g)
h)
rätta sig efter bestämmelserna i tjänsteföreskrifterna vid anställning av före detta tjänstemän från institutionerna,
i)
rätta sig efter alla bestämmelser som parlamentet fastställer om före detta ledamöters rättigheter och skyldigheter,
j)
2.
Brott mot dessa ordningsregler kan medföra att passerkortet dras in för berörda personer, och eventuellt för deras företag.
BILAGA
X
Ombudsmannens ämbetsutövning
A.
Europaparlamentets beslut om föreskrifter och allmänna villkor för ombudsmannens ämbetsutövning
Antaget av parlamentet den 9 mars 1994 (EGT L 113, 4.5.1994, s.
15) och ändrat genom parlamentets beslut av den 14 mars 2002 (EGT L 92, 9.4.2002, s.
13) och den 18 juni 2008 (EUT L 189, 17.7.2008, s.
25).
Europaparlamentet har beslutat följande:
Europeiska atomenergigemenskapen,
med beaktande av rådets godkännande och
med beaktande av följande:
Föreskrifterna och de allmänna villkoren för ombudsmannens ämbetsutövning bör fastställas i enlighet med bestämmelserna i fördragen om upprättandet av Europeiska gemenskaperna.
Därför måste gemenskapens institutioner och organ på ombudsmannens begäran tillhandahålla all information som begärs och utan att det påverkar ombudsmannens skyldighet att inte avslöja sådan information.
Tillgången till sekretessbelagd information eller sekretessbelagda dokument, särskilt känsliga handlingar i den mening som avses i artikel 9 i förordning (EG) nr 1049/2001
Europaparlamentets och rådets förordning (EG) nr 1049/2001 av den 30 maj 2001 om allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar (EGT L 145, 31.5.2001, s.
43).
, bör vara förenlig med säkerhetsbestämmelserna för gemenskapsinstitutionen eller gemenskapsorganet i fråga.
Institutioner och organ som tillhandahåller sekretessbelagda uppgifter eller handlingar enligt artikel 3.2 första stycket bör underrätta ombudsmannen om att de är sekretessbelagda.
Det bör även läggas fast att ombudsmannen vid slutet av varje årlig session överlämnar en uttömmande rapport till Europaparlamentet.
Ombudsmannen och personalen måste behandla den information som de har fått under sin ämbetsutövning förtroligt; ombudsmannen måste dock underrätta de behöriga myndigheterna om förhållanden som troligen kan omfattas av straffrättslig lagstiftning och som kommit till ombudsmannens kännedom genom undersökningar.
Bestämmelser bör fastställas för ett eventuellt samarbete mellan ombudsmannen och samma slags myndigheter i vissa medlemsstater i överensstämmelse med tillämplig nationell lagstiftning.
I början av varje mandatperiod och för hela dess längd bör Europaparlamentet till ombudsman utse en person som är medborgare i unionen och som uppvisar alla erforderliga bevis för oavhängighet och kompetens.
Det bör fastställas under vilka villkor som ombudsmannens ämbetsutövning skall upphöra.
HÄRIGENOM FÖRESKRIVS FÖLJANDE
Artikel
1
1.
2.
Ombudsmannen skall utöva sitt ämbete i enlighet med de befogenheter som fördragen ger gemenskapens institutioner och organ.
3.
Ombudsmannen får inte ingripa i mål som är anhängiga vid domstol eller ifrågasätta domstolsavgöranden.
Artikel
2
1.
Inom ramarna för de ovan nämnda fördragen och de villkor som slås fast i dem skall ombudsmannen bidra till upptäckten av fel och försummelser i samband med verksamheten inom gemenskapens institutioner och organ med undantag av domstolen och förstainstansrätten i deras rättsliga funktion och föreslå åtgärder för att avhjälpa dessa fel och försummelser.
Handlingar som företas av någon annan myndighet eller person kan inte vara föremål för klagan hos ombudsmannen.
2.
Varje unionsmedborgare eller varje fysisk eller juridisk person som har sitt hemvist eller säte i en av unionens medlemsstater kan antingen direkt eller genom en ledamot av Europaparlamentet inge ett klagomål till ombudsmannen gällande fel eller försummelser i samband med verksamheten inom gemenskapens institutioner och organ med undantag av domstolen och förstainstansrätten i deras rättsliga funktion.
Ombudsmannen skall underrätta institutionen eller organet i fråga så snart ett klagomål inges.
3.
Klagomålet skall innehålla uppgifter om klagomålets innehåll och vem som framför klagomålet; denne kan begära att klagomålet behandlas förtroligt.
4.
Ett klagomål skall göras inom två år från den dag då omständigheterna på vilka klagomålet grundar sig blev kända av den person som framför klagomålet och måste föregås av lämpliga hänvändelser till de berörda institutionerna och organen.
5.
Ombudsmannen kan råda den person som framför klagomålet att vända sig till en annan myndighet.
6.
Klagomål som inges till ombudsmannen skall inte påverka tidsfrister för överklaganden i administrativa förfaranden eller domstolsförfaranden.
7.
När ombudsmannen måste avvisa ett klagomål eller avbryta sin undersökning på grund av pågående eller avslutade rättsliga åtgärder rörande omständigheter som tagits upp i ett klagomål skall resultatet av de undersökningar som redan är gjorda arkiveras utan ytterligare åtgärder.
8.
9.
Ombudsmannen skall snarast möjligt underrätta den person som har framfört klagomålet om vilka åtgärder som vidtagits.
Artikel
3
1.
Ombudsmannen skall på eget initiativ eller på grund av ett klagomål genomföra alla undersökningar som finnes vara berättigade för att reda ut misstänkta fel eller försummelser i samband med verksamheten inom gemenskapens institutioner och organ.
Ombudsmannen skall underrätta den berörda institutionen eller det berörda organet om detta och de kan ge alla relevanta upplysningar.
2.
Gemenskapens institutioner och organ ska förse ombudsmannen med all information som begärs av dem och ge ombudsmannen tillgång till relevanta dokument.
Tillgången till sekretessbelagd information eller sekretessbelagda dokument, särskilt känsliga handlingar i den mening som avses i artikel 9 i förordning (EG) nr 1049/2001, ska vara förenlig med säkerhetsbestämmelserna för gemenskapsinstitutionen eller gemenskapsorganet i fråga.
Institutioner och organ som tillhandahåller sekretessbelagda uppgifter eller handlingar enligt stycket ovan ska underrätta ombudsmannen om att de är sekretessbelagda.
Vid tillämpningen av bestämmelserna i första stycket ska ombudsmannen i förväg ha kommit överens med institutionen eller organet i fråga om villkoren för hantering av sekretessbelagd information eller sekretessbelagda dokument och annan information som omfattas av tystnadsplikt.
Institutionerna eller organen i fråga ska ge ombudsmannen tillgång till dokument som härrör från en medlemsstat och som är hemliga enligt lag eller andra författningar endast om den medlemsstaten på förhand har givit sitt samtycke.
De ska ge tillgång till andra dokument som härrör från en medlemsstat efter att ha informerat medlemsstaten i fråga.
I båda fallen får ombudsmannen i enlighet med artikel 4 inte avslöja innehållet i sådana dokument.
Tjänstemän och andra anställda inom gemenskapens institutioner och organ ska avlägga vittnesmål på begäran av ombudsmannen; de ska fortfarande vara bundna av de relevanta reglerna i tjänsteföreskrifterna, i synnerhet ska de ha fortsatt tystnadsplikt.
3.
På begäran av ombudsmannen måste medlemsstaternas myndigheter via medlemsstaternas beskickningar vid Europeiska gemenskaperna tillhandahålla all information som kan bidra till att reda ut misstänkta fel eller försummelser i samband med verksamheten inom gemenskapens institutioner och organ utom när sådan information omfattas av lagar och andra författningar om sekretess eller av bestämmelser som hindrar dess spridning.
I det senare fallet kan dock den berörda medlemsstaten tillåta ombudsmannen att ta del av informationen under förutsättning att han förbinder sig att inte avslöja den.
4.
5.
Ombudsmannen skall så långt det är möjligt försöka att tillsammans med institutionen eller organet i fråga nå en lösning som rättar till felet eller gottgör försummelsen och som tillfredsställer klagomålet.
6.
Om ombudsmannen upptäcker fall av fel eller försummelse skall institutionen eller organet i fråga meddelas och när så är lämpligt föreslå rekommendationer.
Institutionen eller organet skall inom tre månader sända ett detaljerat yttrande till ombudsmannen.
7.
Ombudsmannen skall sedan sända en rapport till Europaparlamentet och till institutionen eller organet i fråga.
Rapporten får innehålla rekommendationer.
Ombudsmannen skall underrätta den person som inlämnat klagomålet om undersökningens resultat om yttrandet från institutionen eller organet i fråga samt om ombudsmannens rekommendationer.
8.
Vid slutet av varje årlig session skall ombudsmannen överlämna en rapport om sina undersökningsresultat till Europaparlamentet.
Artikel
4
1.
Ombudsmannen och dennes personal, på vilka artikel 287 i fördraget om upprättandet av Europeiska gemenskapen och artikel 194 i fördraget om upprättandet av Europeiska atomenergigemenskapen ska tillämpas, får inte avslöja information eller innehåll i dokument som de får tillgång till i sina undersökningar.
Framför allt får de inte avslöja sekretessbelagd information eller innehåll i dokument som överlämnats till ombudsmannen, i synnerhet inte känsliga handlingar i den mening som avses i artikel 9 i förordning (EG) nr 1049/2001, eller dokument som omfattas av gemenskapslagstiftningen om skydd av personuppgifter liksom sådan information som kan skada den person som har lämnat in klagomålet eller någon annan inblandad person, dock utan att det påverkar tillämpningen av punkt 2.
2.
Ombudsmannen får även informera gemenskapsinstitutionen eller gemenskapsorganet i fråga om förhållanden som från disciplinär synpunkt ifrågasätter uppträdandet hos en av deras anställda.
Artikel
4 a
Artikel
5
1.
Ombudsmannen får samarbeta med myndigheter av samma typ i vissa medlemsstater under förutsättning att det sker i enlighet med gällande nationell lagstiftning, om det gör undersökningsarbetet mer effektivt och ger bättre skydd för rättigheter och intressen åt de personer som lämnar in klagomål.
Ombudsmannen får inte på dessa grunder begära att få se dokument som ombudsmannen inte skulle ha tillgång till enligt artikel 3.
2.
Inom ramen för sina befogenheter enligt artikel 195 i fördraget om upprättandet av Europeiska gemenskapen och artikel 107d i fördraget om upprättandet av Europeiska atomenergigemenskapen och i syfte att undvika dubbelarbete i förhållande till verksamheten inom andra institutioner och organ, får ombudsmannen, på samma villkor, samarbeta med de institutioner och organ i medlemsstaterna som ansvarar för främjande och skydd av grundläggande rättigheter.
Artikel
6
1.
Efter varje val till Europaparlamentet skall en ombudsman utses av Europaparlamentet för hela valperiodens längd.
Ombudsmannens mandat kan förlängas.
2.
Ombudsmannen skall utses bland personer som är unionsmedborgare som fullt ut äger medborgerliga och politiska rättigheter, som uppvisar alla erforderliga bevis för oavhängighet och som uppfyller kraven för utövandet av det högsta domarämbetet i sina länder eller besitter en sådan erkänd kompetens och erfarenhet som krävs för att utöva ombudsmannaämbetet.
Artikel
7
1.
Ombudsmannen skall upphöra att utöva sitt ämbete antingen vid slutet av sin ämbetsperiod eller vid frivillig avgång eller avskedande.
2.
Ombudsmannen skall stanna i sitt ämbete till dess att efterträdare har utsetts utom vid avskedande.
3.
Om ämbetet frånträds i förtid skall en efterträdare utses för den resterande delen av parlamentssessionen inom tre månader från den tidpunkt då ämbetet blev vakant.
Artikel
8
En ombudsman som inte längre uppfyller de krav som ställs för utförande av uppgifterna eller som gör sig skyldig till allvarlig försummelse kan avsättas av Europeiska gemenskapernas domstol på begäran av Europaparlamentet.
Artikel
9
1.
Ombudsmannen skall utöva sitt ämbete med fullständig oavhängighet i gemenskapernas och unionsmedborgarnas allmänna intresse.
I sin ämbetsutövning skall ombudsmannen varken begära eller acceptera instruktioner från någon regering eller från något annat organ.
Ombudsmannen skall avstå från alla handlingar som är oförenliga med ämbetsutövningen.
2.
När ombudsmannen tillträder sitt ämbete skall en högtidlig försäkran avges inför Europeiska gemenskapernas domstol att ombudsmannen ämnar utöva sitt ämbete med fullständig oavhängighet och opartiskhet samt under och efter sin ämbetsperiod kommer att respektera de åtaganden som följer av ämbetet särskilt plikten att efter ämbetstidens utgång uppträda med integritet och diskretion när det gäller att acceptera vissa befattningar eller förmåner.
Artikel
10
1.
Under ämbetsperioden får ombudsmannen inte åtaga sig någon annan politisk eller administrativ uppgift eller utöva någon annan verksamhet oavsett om den är avlönad eller inte.
2.
Ombudsmannen skall ha samma ställning som en domare vid Europeiska gemenskapernas domstol när det gäller lön, traktamenten och pension.
3.
Artikel 12-15 och artikel 18 i protokollet om immunitet och privilegier för Europeiska gemenskaperna skall tillämpas på ombudsmannen samt tjänstemännen och övriga anställda vid ombudsmannens kansli.
Artikel
11
1.
Ombudsmannen skall biträdas av ett kansli vars chefstjänsteman ombudsmannen skall utse.
2.
Tjänstemännen och andra anställda vid ombudsmannens kansli skall lyda under de regler och bestämmelser som gäller för tjänstemän och andra anställda inom Europeiska gemenskaperna.
Deras antal skall anpassas varje år som ett led i budgetprocessen.
3.
Anställda i Europeiska gemenskaperna och i medlemsstaterna som utses att tjänstgöra vid ombudsmannens kansli skall flyttas över i tjänstens intresse och skall garanteras återinträde i en tjänst vid sin ursprungliga arbetsplats.
4.
I personalärenden skall ombudsmannen ha samma status som institutionerna i den betydelse som avses i artikel 1 i tjänsteföreskrifterna för tjänstemännen i Europeiska gemenskaperna.
Artikel
12
(Utgår)
Artikel
13
Ombudsmannen skall ha samma säte som Europaparlamentet.
Artikel
14
Ombudsmannen skall anta bestämmelser för genomförandet av detta beslut.
Artikel
15
Den första ombudsman som utses efter ikraftträdandet av Fördraget om Europeiska unionen skall utses för den resterande delen av parlamentets valperiod.
Artikel
16
(Utgår)
Artikel
17
Detta beslut skall offenliggöras i Europeiska gemenskapernas officiella tidning.
Det träder i kraft samma dag som det offentliggörs.
B.
Europeiska ombudsmannens beslut om antagande av genomförandebestämmelser
Antaget den 8 juli 2002 och ändrat genom ombudsmannens beslut av den 5 april 2004.
Artikel
1
Definitioner
I dessa genomförandebestämmelser avses med
a)
”berörd institution”: den gemenskapsinstitution eller det gemenskapsorgan som är föremål för ett klagomål eller en undersökning på eget initiativ,
b)
”stadgan”: föreskrifterna och de allmänna villkoren för ombudsmannens ämbetsutövning.
Artikel
2
Inkommande klagomål
2.1.
Inkommande klagomål skall identifieras, registreras och numreras.
2.2.
Mottagandet skall bekräftas till den person som lämnat in klagomålet, med angivande av klagomålets registreringsnummer och namn på den juridiska handläggare som handlägger det.
2.3.
En framställning som Europaparlamentet med framställarens medgivande överför till ombudsmannen skall behandlas som ett klagomål.
2.4.
Ombudsmannen får, när så är lämpligt och med medgivande av den person som lämnat in klagomålet, överföra ett klagomål till Europaparlamentet för behandling som en framställning.
2.5.
Ombudsmannen får, när så är lämpligt och med medgivande av den person som lämnat in klagomålet, överföra ett klagomål till en annan behörig myndighet.
Artikel
3
Klagomåls tillåtlighet
3.1.
3.2.
Om klagomålet ligger utanför ombudsmannens ämbetsområde eller är otillåtligt skall han avvisa klagomålet.
Han skall informera den person som lämnat in klagomålet om sitt beslut och om skälen mot det.
Ombudsmannen kan råda den person som lämnat in klagomålet att vända sig till annan myndighet.
Artikel
4
Undersökningar av tillåtna klagomål
4.1.
Ombudsmannen skall besluta om det finns tillräckliga grunder för att inleda en undersökning av ett tillåtligt klagomål.
4.2.
Om ombudsmannen anser att det saknas tillräckliga grunder för att motivera en undersökning skall han avsluta ärendet och informera den person som lämnat in klagomålet om detta.
4.3.
Om ombudsmannen anser att det finns tillräckliga grunder för att motivera en undersökning skall han informera den person som lämnat in klagomålet och den berörda institutionen om detta.
Han skall skicka en kopia av klagomålet till den berörda institutionen med en uppmaning att avge ett yttrande inom en angiven tidsperiod på normalt högst tre månader.
Uppmaningen till den berörda institutionen får innehålla specifikationer om särskilda aspekter av klagomålet eller särskilda frågor som bör tas upp i yttrandet.
4.4
Ombudsmannen skall skicka den berörda institutionens yttrande till den person som lämnat in klagomålet.
Denne skall beredas möjlighet att avge kommentarer till ombudsmannen inom en angiven tidsperiod på normalt högst en månad.
4.5.
Efter att ha övervägt yttrandet och eventuella kommentarer från den person som lämnat in klagomålet får ombudsmannen antingen avsluta ärendet med ett motiverat beslut eller fortsätta sin undersökning.
Han skall informera den person som lämnat in klagomålet och den berörda institutionen om detta.
Artikel
5
Undersökningsbefogenheter
5.1.
Ombudsmannen får i enlighet med de villkor som fastställs i stadgan begära att gemenskapens institutioner och organ och medlemsstaternas myndigheter inom rimlig tid tillhandahåller information eller handlingar för en undersökning.
5.2.
Ombudsmannen får inspektera den berörda gemenskapsinstitutionens samtliga handlingar i ett ärende för att kontrollera huruvida institutionen har lämnat ett korrekt och uttömmande svar.
Ombudsmannen får ta kopior på alla handlingar i ett ärende ärendet eller vissa handlingar i det.
Ombudsmannen skall informera den person som lämnat in klagomålet om att en inspektion har skett.
5.3.
På begäran av ombudsmannen skall tjänstemän eller andra anställda inom gemenskapens institutioner eller organ avlägga vittnesmål i enlighet med de villkor som fastställs i stadgan.
5.4.
Ombudsmannen kan begära att gemenskapens institutioner och organ vidtar åtgärder så att han kan utföra sina undersökningar på plats.
5.5.
Ombudsmannen får beställa de undersökningar och expertrapporter han anser nödvändiga för att för att på ett tillfredsställande sätt genomföra en undersökning.
Artikel
6
Uppgörelser i godo
6.1
Om ombudsmannen konstaterar administrativa missförhållanden skall han i så stor utsträckning som möjligt samarbeta med den berörda institutionen för att nå en uppgörelse i godo om att undanröja dem på ett tillfredsställande sätt för den person som lämnat in klagomålet.
6.2
Om ombudsmannen anser att detta samarbete har gett ett tillfredsställande resultat skall han avsluta ärendet med ett motiverat beslut.
Han skall informera den person som lämnat in klagomålet och den berörda institutionen om sitt beslut.
6.3
Om ombudsmannen anser att en uppgörelse i godo inte är möjlig, eller om försök till en sådan har misslyckats, skall han antingen avsluta ärendet med ett motiverat beslut som kan inbegripa en kritisk anmärkning eller utarbeta en rapport med förslag till rekommendationer.
Artikel
7
Kritiska anmärkningar
7.1
Ombudsmannen skall utfärda en kritisk anmärkning om han anser
a)
att det inte längre är möjligt för institutionen i fråga att undanröja fallet av administrativt missförhållande och
b)
fallet av administrativt missförhållande inte har några allmänna återverkningar.
7.2
När ombudsmannen avslutar ett ärende med en kritisk anmärkning skall han informera den person som lämnat in klagomålet om sitt beslut.
Artikel
8
Rapporter och rekommendationer
8.1.
Ombudsmannen skall lägga fram en rapport med förslag till rekommendationer till institutionen i fråga om han anser att det antingen
a)
är möjligt för institutionen i fråga att undanröja fallet av administrativt missförhållande, eller
b)
fallet av administrativt missförhållande har allmänna återverkningar.
8.2.
Ombudsmannen skall skicka en kopia av sin rapport och sina förslag till rekommendationer till den berörda institutionen och till den person som lämnat in klagomålet.
8.3.
Den berörda institutionen skall avge ett detaljerat yttrande till ombudsmannen inom tre månader.
Det detaljerade yttrandet kan bestå av ett godkännande av ombudsmannens beslut och en beskrivning av de åtgärder som vidtagits för att genomföra de föreslagna rekommendationerna.
8.4.
Om ombudsmannen inte anser att det detaljerade yttrandet är tillfredsställande kan han utarbeta en särskild rapport till Europaparlamentet om det administrativa missförhållandet.
Den särskilda rapporten kan innehålla rekommendationer.
Ombudsmannen skall skicka en kopia av rapporten till den berörda institutionen och till den person som lämnat in klagomålet.
Artikel
9
Undersökningar på eget initiativ
9.1.
Ombudsmannen får besluta att göra undersökningar på eget initiativ.
9.2.
Ombudsmannen skall vid undersökningar på eget initiativ ha samma undersökningsbefogenheter som vid undersökningar till följd av klagomål.
9.3.
De förfaranden som tillämpas vid undersökningar till följd av klagomål skall på motsvarande sätt tillämpas vid undersökningar på eget initiativ.
Artikel
10
Procedurfrågor
10.1.
Ombudsmannen skall behandla klagomålet konfidentiellt om den person som lämnat in klagomålet begär det.
Om ombudsmannen anser det nödvändigt att skydda den klagandes eller tredje parts intressen får han på eget initiativ klassificera ett klagomål som konfidentiellt.
10.2.
Om ombudsmannen anser det lämpligt får han vidta åtgärder för att se till att ett klagomål prioriteras.
10.3.
Om rättsliga förfaranden inleds rörande omständigheter som ombudsmannen utreder skall han avsluta ärendet.
Resultatet av de undersökningar som är gjorda skall arkiveras utan ytterligare åtgärder.
10.4.
Om ombudsmannen under en undersökning upptäcker förhållanden som omfattas av strafflagstiftning skall han underrätta de nationella behöriga myndigheterna och, i tillämpliga fall, en gemenskapsinstitution eller ett gemenskapsorgan.
Ombudsmannen får även informera en gemenskapsinstitution eller ett gemenskapsorgan om förhållanden som han anser kan motivera disciplinära åtgärder.
Artikel
11
Rapporter till Europaparlamentet
11.1.
Ombudsmannen skall till Europaparlamentet överlämna en årsrapport om hela sin verksamhet, inbegripet sina undersökningsresultat.
11.2.
11.3.
Årsrapporten och de särskilda rapporterna från ombudsmannen får innehålla sådana rekommendationer han anser lämpliga för att uppfylla sina förpliktelser enligt fördragen och stadgan.
Artikel
12
Samarbete med ombudsmän och liknande instanser i medlemsstaterna
Ombudsmannen får samarbeta med ombudsmän och liknande instanser i medlemsstaterna för att effektivisera sina egna undersökningar och de undersökningar som görs av ombudsmän och liknande instanser i medlemsstaterna, och för att garantera mer verksamma åtgärder för att bevaka de rättigheter och intressen som omfattas av Europeiska unionens och Europeiska gemenskapens lagstiftning.
Artikel
13
Den klagande personens rätt att se handlingar i ärendet
13.1.
13.2.
Den person som lämnat in klagomålet kan kräva att få se handlingarna på plats.
Han eller hon kan begära att ombudsmannen tillhandahåller kopior av alla handlingar i ärendet eller av specifika handlingar.
13.3.
Artikel
14
Allmänhetens tillgång till handlingar som innehas av ombudsmannen
14.1.
Allmänheten skall, på samma villkor och med samma gränser som fastställs i förordning (EG) 1049/2001 om allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar
Europaparlamentets och rådets förordning (EG) nr 1049/2001 av den 30 maj 2001 om allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar (EGT L 145, 31.5.2001, s.
43).
14.2.
14.3.
Ansökningar om tillgång till handlingar skall vara skriftliga (brev, fax eller e-post) och tillräckligt utförliga för att handlingarna skall kunna identifieras.
14.4.
a)
Det allmänna registret över klagomål.
b)
Klagomål och bifogade handlingar från klaganden.
c)
Yttranden och detaljerade yttranden från berörda institutioner och eventuella kommentarer till dessa från klaganden.
d)
Ombudsmannens beslut att avsluta ärenden.
e)
Rapporter och förslag till rekommendationer enligt artikel 8.
14.5.
Tillgång skall antingen ges på plats eller genom att sökanden får en kopia.
Ombudsmannen får ta ut rimliga avgifter för att tillhandahålla kopior.
Alla avgifter skall specificeras.
14.6.
Tillgång till de handlingar som anges i artikel 14.4 ovan skall beredas snarast.
14.7.
Om en ansökan om tillgång till en handling helt eller delvis avslås skall grunderna för beslutet anges.
15.1.
Klagomål som inges till ombudsmannen skall vara skrivet på ett av fördragsspråken.
Ombudsmannen behöver inte behandla klagomål som ingetts på andra språk än dessa.
15.3.
Ombudsmannen skall avgöra vilka handlingar som skall upprättas på det språk som används vid förhandlingarna.
15.4.
Skriftväxling med medlemsstaternas myndigheter skall ske på den berörda statens officiella språk.
15.5.
Årsrapporten, särskilda rapporter och, i den mån det är möjligt, övriga handlingar som ombudsmannen offentliggör skall finnas tillgängliga på samtliga officiella språk.
Artikel
16
Rapporternas offentliggörande
16.1.
Ombudsmannen skall offentliggöra meddelanden om antagna årliga och särskilda rapporter i Europeiska gemenskapernas officiella tidning och offentliggöra på vilket sätt allmänheten kan få tillgång till de fullständiga handlingarna.
16.2.
17.2.
Detta beslut skall träda i kraft den 1 januari 2003.
1.
och rådets förordning (Euratom) nr 1074/1999
8.
om utredningar som utförs av Europeiska byrån för bedrägeribekämpning innehåller bestämmelser om att byrån skall inleda och utföra administrativa utredningar inom de institutioner, organ och byråer som inrättats genom EG-fördraget och Euratomfördraget eller på grundval av dessa fördrag.
Det är viktigt att öka bedrägeribekämpningens omfattning och effektivitet med hjälp av de experter som finns inom området för administrativa utredningar.
Detta gäller vidare brister som kan skada dessa gemenskapers intressen och som kan leda till disciplinära åtgärder och, i förekommande fall, straffrättsliga åtgärder.
Dessa utredningar skall utföras på samma villkor inom alla institutioner, organ och byråer inom gemenskapen utan att överlämnandet av denna uppgift till byrån skall påverka institutionernas, organens och byråernas eget ansvar eller på något sätt minska de berörda personernas rättsliga skydd.
Artikel
I detta avseende skall de till byråns anställda lämna alla upplysningar och alla förklaringar som behövs.
Artikel
Talman, generalsekreterare, generaldirektörer och avdelningschefer skall utan dröjsmål till byrån överlämna alla uppgifter som de får kännedom om och som tyder på förekomsten av sådana oegentligheter som avses i första stycket.
En tjänsteman eller anställd vid Europaparlamentet får aldrig utsättas för en orättvis eller diskriminerande behandling på grund av ett sådant uppgiftslämnande som avses i första och andra styckena.
Ledamöter som får kännedom om uppgifter som avses i första stycket skall underrätta Europaparlamentets talman, eller om ledamöterna anser det vara lämpligt, byrån direkt.
Artikel
Artikel
Under inga omständigheter får slutsatser dras efter utredningen om en namngiven ledamot, tjänsteman eller anställd inom Europaparlamentet, utan att den berörde har givits möjlighet att yttra sig över alla uppgifter som rör honom.
Om inget av det som lagts ledamoten, tjänstemannen eller den anställde vid Europaparlamentet till last kan vidhållas efter en intern utredning, skall den interna utredningen mot honom eller henne läggas ned utan vidare åtgärder efter beslut av byråns direktör, som skriftligen skall underrätta den berörde om detta.
Artikel
1.
Europaparlamentet ska därför samtidigt som kommittémedlemmarna och på samma villkor få de förslag till dagordning för mötena och de förslag om genomförandeåtgärder som läggs fram för dessa kommittéer
Ordet "kommitté" ska i denna överenskommelse genomgående anses syfta på de kommittéer som inrättas i enlighet med beslut 1999/468/EG.
i enlighet med grundläggande rättsakter som antagits enligt förfarandet i artikel 251 i EG-fördraget, och även få information om resultat av omröstningar, sammanfattningar av möten och förteckningar över de myndigheter som medlemsstaternas företrädare tillhör.
Register
2.
Måldatum för upprättande av registret är den 31 mars 2008.
.
I överensstämmelse med de åtaganden som kommissionen har gjort i sitt uttalande om artikel 7.3 i beslut 1999/468/EG
-
ange etappen i förfarandet samt tidsplanen,
4.
Detta beslut ska fattas genom en skriftväxling mellan ordförandena för de båda institutionerna.
5.
6.
Se domen av den 19 juli 1999 från Europeiska gemenskapernas förstainstansrätt i mål T-188/97 Rothmans mot kommissionen REG 1999, s.
7.
8.
Finansiella tjänster
I enlighet med sitt uttalande om artikel 7.3 i beslut 1999/468/EG åtar sig kommissionen att när det gäller finansiella tjänster
Tidigare avtal
20.
Den överenskommelse som 2000 ingicks mellan Europaparlamentet och kommissionen om tillämpningsföreskrifter till rådets beslut 1999/468/EG
1.
.
BILAGA
XIII
Europaparlamentet
Parlamentets beslut av den 26 maj 2005.
D.
Det ramavtal som undertecknades i juli 2000
EGT C 121, 24.4.2001, s.
122.
bör uppdateras och ersättas av nedanstående text.
I. TILLÄMPNINGSOMRÅDE
1.
De två institutionerna beslutar om följande åtgärder för att öka kommissionens politiska ansvar och legitimitet, utvidga den konstruktiva dialogen och förbättra informationsflödet mellan de två institutionerna samt förbättra samordningen av förfaranden och planering.
2.
Kommissionens ordförande skall fullt ut ansvara för att avgöra om det finns någon eventuell intressekonflikt som gör det omöjligt för en kommissionsledamot att fullgöra sina uppgifter.
Ordföranden skall omedelbart skriftligen underrätta parlamentets talman om ett enskilt ärende omfördelats.
3.
Om parlamentet beslutar att inte ge en kommissionsledamot sitt förtroende skall kommissionens ordförande, efter att noga ha övervägt parlamentets beslut, antingen begära att kommissionsledamoten avgår, eller förklara sitt beslut för parlamentet.
4.
Parlamentet skall se till att dess förfaranden genomförs så snabbt som möjligt, så att kommissionens ordförande kan underrättas om parlamentets ståndpunkt i god tid innan kommissionsledamoten utnämns.
5.
Kommissionens ordförande skall omedelbart underrätta parlamentet om varje beslut som rör fördelningen av kommissionsledamöternas ansvarsområden.
Om en kommissionsledamots ansvarsområde väsentligt ändras skall kommissionsledamoten i fråga infinna sig i det ansvariga utskottet om parlamentet så begär.
6.
7.
Parlamentet skall i enlighet med artikel 99 i sin arbetsordning höra kommissionens nominerade ordförande i god tid innan förfarandet för godkännande av den nya kommissionen inleds.
8.
På alla områden där parlamentet handlar som lagstiftande organ eller som en del av budgetmyndigheten skall det hållas underrättat på samma sätt som rådet i varje skede av lagstiftningsprocessen och budgetförfarandet.
9.
När det gäller den gemensamma utrikes- och säkerhetspolitiken samt polissamarbete och straffrättsligt samarbete skall kommissionen vidta åtgärder för att förbättra parlamentets deltagande så att parlamentets åsikter i så stor utsträckning som möjligt beaktas.
10.
Kommissionens ordförande och/eller den vice ordförande som ansvarar för de interinstitutionella förbindelserna kommer var tredje månad att sammanträda med talmanskonferensen för att säkerställa en löpande dialog mellan de två institutionerna på högsta nivå.
Kommissionens ordförande kommer att närvara vid talmanskonferensens sammanträden minst två gånger per år.
11.
Alla kommissionsledamöter skall se till att det sker ett regelbundet och direkt informationsutbyte mellan dem själva och ordföranden för det ansvariga parlamentsutskottet.
12.
På grundval av kommissionens lagstiftnings- och arbetsprogram och av det fleråriga programmet skall de två institutionerna genom överenskommelse på förhand fastställa vilka förslag och initiativ som är av särskild vikt, i syfte att lägga fram dem vid ett plenarsammanträde i parlamentet.
13.
Om ett internt dokument från kommissionen – som parlamentet inte har fått information om i enlighet med punkterna 8, 9 och 12 – sprids utanför institutionerna, får parlamentets talman begära att detta dokument överlämnas till parlamentet utan dröjsmål så att det kan vidarebefordras till de ledamöter av parlamentet som så begär.
14.
15.
16.
17.
18.
Om sekretess åberopas i fråga om information som överlämnats i enlighet med detta ramavtal skall bestämmelserna i bilaga 1 tillämpas.
ii) Yttre förbindelser, utvidgning och internationella avtal
19.
Sådan information som avses i första stycket skall översändas till parlamentet i så god tid att parlamentet ges möjlighet att framföra sina eventuella synpunkter och kommissionen ges möjlighet att i största möjliga mån ta hänsyn till parlamentets synpunkter.
20.
Kommissionen skall vidta de åtgärder som krävs för att säkerställa att parlamentet omedelbart och till fullo informeras om
i)
ii)
en gemenskapsståndpunkt som antagits i ett organ som upprättats genom ett avtal.
21.
22.
23.
De två institutionerna är eniga om att samarbeta när det gäller valobservation.
24.
Kommissionen skall hålla parlamentet fullständigt underrättat om läget i anslutningsförhandlingar, särskilt om viktigare aspekter och händelser, så att parlamentet ges möjlighet att i god tid lämna synpunkter genom de tillämpliga parlamentariska förfarandena.
25.
iii) Budgetgenomförandet
26.
Om det kommer fram nya uppgifter om tidigare år för vilka ansvarsfrihet redan beviljats skall kommissionen översända all relevant information, i syfte att uppnå en lösning som är acceptabel för båda parter.
IV.
i) Kommissionens politiska program och lagstiftningsprogram samt Europeiska unionens fleråriga planering
27.
Kommissionen skall lägga fram förslag till Europeiska unionens fleråriga planering, i syfte att uppnå enighet kring den interinstitutionella planeringen mellan de berörda institutionerna.
28.
Varje ny kommission skall så tidigt som möjligt lägga fram sitt politiska program och lagstiftningsprogram.
29.
När kommissionen utarbetar sitt lagstiftnings- och arbetsprogram skall de två institutionerna samarbeta i enlighet med tidsplanen i bilaga 2.
Kommissionen skall tillhandahålla tillräckliga uppgifter om planerade åtgärder inom ramen för respektive punkt i lagstiftnings- och arbetsprogrammet.
30.
Den vice kommissionsordförande som ansvarar för de interinstitutionella förbindelserna åtar sig att var tredje månad inför utskottsordförandekonferensen redogöra för huvuddragen i det politiska genomförandet av lagstiftnings- och arbetsprogrammet för det berörda året och eventuella uppdateringar av detta program som är nödvändiga på grund av aktuella och viktiga politiska händelser.
ii) Allmänna lagstiftningsförfaranden
31.
Kommissionen åtar sig att noga beakta de ändringar av kommissionens lagförslag som parlamentet antagit, i syfte att ta hänsyn till dessa ändringar i eventuellt ändrade förslag.
Om kommissionen på grund av tungt vägande skäl och efter en behandling i kollegiet av kommissionsledamöter beslutar att inte anta eller stödja sådana ändringar skall den redogöra för sitt beslut inför parlamentet samt under alla förhållanden i det yttrande om parlamentets ändringar som kommissionen skall avge i enlighet med artikel 251.2 c tredje stycket.
32.
33.
Vid andra lagstiftningsförfaranden än medbeslutandeförfarandet gäller att kommissionen
i)
i god tid skall se till att rådets instanser erinras om att de inte bör träffa någon politisk överenskommelse om kommissionens förslag innan parlamentet antagit sitt yttrande; kommissionen skall begära att diskussionen slutförs på ministernivå efter det att rådsmedlemmarna har fått en rimlig tidsfrist för att behandla parlamentets yttrande,
ii)
iii)
åtar sig att, vid behov, dra tillbaka de lagstiftningsförslag som avvisats av parlamentet; om kommissionen av tungt vägande skäl och efter diskussion i kollegiet av kommissionsledamöter beslutar att vidhålla sitt förslag skall motivera detta beslut i ett uttalande inför parlamentet.
34.
I syfte att förbättra lagstiftningsplaneringen åtar sig Europaparlamentet å sin sida att
i)
planera de lagstiftningsrelaterade delarna av föredragningslistan så att de anpassas till gällande lagstiftningsprogram och till de resolutioner som parlamentet har antagit rörande detta program,
ii)
respektera rimliga tidsfrister, om detta är till fördel för förfarandet, när det gäller att anta sitt yttrande under första behandlingen i samarbetsförfarandet och medbeslutandeförfarandet eller under samrådsförfarandet,
iii)
i så hög grad som möjligt utnämna föredragande för kommande förslag så snart lagstiftningsprogrammet har antagits,
iv)
35.
Genomförandet av rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter
EGT L 184, 17.7.1999, s.
23.
19.
mellan Europaparlamentet och kommissionen om tillämpningsföreskrifter till detta beslut.
När det gäller genomförandeåtgärder avseende värdepappers-, bank- och försäkringssektorn bekräftar kommissionen de åtaganden som den avgav under parlamentets plenarsammanträde den 5 februari 2002 och upprepade den 31 mars 2004.
Kommissionen åtar sig särskilt att ta största möjliga hänsyn till parlamentets ståndpunkt och eventuella resolutioner avseende genomförandeåtgärder som överskrider de genomförandebefogenheter som föreskrivs i grunddokumentet.
I dessa fall skall kommissionen sträva efter att finna en balanserad lösning.
iv) Kontroll av tillämpningen av gemenskapsrätten
36.
På begäran av parlamentets ansvariga utskott skall kommissionen utöver de särskilda rapporterna och årsrapporten om tillämpningen av gemenskapsrätten muntligen informera parlamentet om hur långt förfarandet fortskridit.
Detta skall ske så snart ett motiverat yttrande översänts, eller, när det gäller förfaranden med anledning av underlåtenhet att lämna underrättelse om åtgärder för genomförande av direktiv eller underlåtenhet att rätta sig efter en dom från domstolen, så snart en formell underrättelse har översänts.
V. KOMMISSIONENS DELTAGANDE I PARLAMENTETS FÖRFARANDEN
37.
Parlamentet skall som en allmän regel se till att ärenden som ingår i en viss kommissionsledamots ansvarsområde behandlas vid ett och samma tillfälle.
38.
I syfte att säkra kommissionsledamöternas närvaro åtar sig parlamentet att göra sitt bästa för att inte ändra sina slutgiltiga förslag till föredragningslista.
När parlamentet ändrar sitt slutgiltiga förslag till föredragningslista eller flyttar om punkterna på föredragningslistan för en sammanträdesperiod skall det omedelbart informera kommissionen om detta.
Kommissionen skall å sin sida göra sitt bästa för att garantera att den ansvariga kommissionsledamoten närvarar.
39.
Kommissionen kan föreslå att punkter förs upp på föredragningslistan fram till det sammanträde under vilket talmanskonferensen fastställer ett slutgiltigt förslag till föredragningslista för en sammanträdesperiod.
40.
Kommissionsledamöter skall höras på egen begäran.
När det inte uttryckligen begärs att en kommissionsledamot skall närvara vid ett utskottssammanträde skall kommissionen se till att en behörig tjänsteman på lämplig nivå företräder den.
VI.
42.
Tillämpningsområde
1.1.
I denna bilaga regleras hur kommissionens sekretessbelagda information skall överlämnas till parlamentet och hanteras i samband med parlamentets utövande av sina befogenheter när det gäller lagstiftningsprocessen, budgetförfarandet, förfarandet för beviljande av ansvarsfrihet eller sina kontrollbefogenheter i allmänhet.
De båda institutionerna skall verka i enlighet med sina respektive skyldigheter att samarbeta lojalt i en anda av fullständigt ömsesidigt förtroende samt i strikt överensstämmelse med fördragens tillämpliga bestämmelser, särskilt artiklarna 6 och 46 i Fördraget om Europeiska unionen och artikel 276 i Fördraget om upprättandet av Europeiska gemenskapen.
1.2.
1.3.
Kommissionen skall se till att parlamentet får tillgång till information i enlighet med bestämmelserna i denna bilaga när någon av de parlamentsinstanser som anges i punkt 1.4 ger in en begäran om överlämnande av sekretessbelagd information.
1.4.
Följande instanser får inom ramen för denna bilaga begära sekretessbelagd information från kommissionen: parlamentets talman, berörda parlamentsutskotts ordförande, presidiet och talmanskonferensen.
1.5.
1.6.
EGT L 113, 19.5.1995, s.
1.
eller tillämpliga bestämmelser i kommissionens beslut 1999/352/EG, EKSG, Euratom av den 28 april 1999 om inrättande av en europeisk byrå för bedrägeribekämpning (OLAF)
.
2.
Allmänna bestämmelser
2.1.
-
skydd av affärshemligheter och handelsförbindelser,
-
skydd av unionens intressen, särskilt sådana intressen som rör den allmänna säkerheten, internationella förbindelser, valutastabilitet och ekonomiska intressen.
Om parterna är oeniga skall frågan hänskjutas till kommissionens ordförande och parlamentets talman för att de skall kunna finna en lösning.
2.2.
Om det råder tvivel om huruvida viss information är sekretessbelagd eller om formerna för att överlämna informationen behöver preciseras i enlighet med de alternativ som anges i punkt 3.2, skall det ansvariga parlamentsutskottets ordförande, vid behov tillsammans med föredraganden, utan dröjsmål samråda med kommissionens ansvariga ledamot.
Om de inte kan enas skall frågan hänskjutas till kommissionens ordförande och parlamentets talman för att de skall kunna finna en lösning.
2.3.
Om oenigheten kvarstår efter förfarandet i punkt 2.2 skall parlamentets talman på motiverad begäran av det ansvariga parlamentsutskottet uppmana kommissionen att inom en lämplig på vederbörligt sätt angiven tidsfrist, överlämna den berörda sekretessbelagda informationen samt precisera formerna för detta i enlighet med de alternativ som anges i avsnitt 3 i denna bilaga.
Kommissionen skall före utgången av denna tidsfrist skriftligen underrätta parlamentet om sin slutliga ståndpunkt beträffande vilken parlamentet förbehåller sig rätten att vid behov väcka talan.
3.
Former för tillgång till och behandling av sekretessbelagd information
3.1.
Sekretessbelagd information som överlämnats i enlighet med förfarandena i punkt 2.2 och, i förekommande fall, punkt 2.3 skall på kommissionsordförandens eller en kommissionsledamots ansvar överlämnas till den parlamentsinstans som har gjort begäran.
3.2.
Utan att det påverkar bestämmelserna i punkt 2.3 skall tillgången till informationen och formerna för skydd av informationens sekretess fastställas genom en överenskommelse mellan den berörda parlamentsinstansen, vederbörligen företrädd av sin ordförande, och den ansvarige kommissionsledamoten enligt något av följande alternativ:
-
information avsedd för ordföranden och föredraganden i det ansvariga parlamentsutskottet,
-
-
överlämnande av handlingar i vilka alla personuppgifter tagits bort,
-
information avsedd endast för parlamentets talman, i välmotiverade och exceptionella fall.
Det är förbjudet att offentliggöra informationen i fråga eller att vidarebefordra den till någon som helst annan mottagare.
3.3.
3.4.
ett säkert arkiveringssystem för sekretessbelagda handlingar,
-
3.5.
:
TIDSPLAN FÖR KOMMISSIONENS LAGSTIFTNINGS- OCH ARBETSPROGRAM
1.
Under sammanträdesperioden i februari mars skall de berörda institutionerna hålla en debatt om de politiska prioriteringarnas huvuddrag, på grundval av beslutet om den årliga politiska strategin för nästföljande år.
3.
Varje parlamentsutskott skall till utskottsordförandekonferensen regelbundet rapportera om resultaten av dessa möten.
4.
5.
I september skall utskottsordförandekonferensen lägga fram en sammanfattande rapport för talmanskonferensen, som i sin tur skall informera kommissionen om denna rapport.
Presentationen skall bland annat inbegripa en utvärdering av genomförandet av det pågående programmet.
Därefter skall parlamentet under december månads sammanträdesperiod anta en resolution.
7.
Följande skall ingå: tidsplan och, i förekommande fall, rättslig grund och återverkningar på budgeten.
.
Programmet skall överlämnas till parlamentet i god tid före den sammanträdesperiod då det skall diskuteras.
8.
Denna tidsplan skall tillämpas på varje normal programcykel, med undantag för år då val till Europaparlamentet sammanfaller med att kommissionens mandatperiod löper ut.
9.
BILAGA
1.
1.1
1.2
1.3
1.4
1.5
1.6
1.7
Handlingar från andra parlamentsorgan
Protokoll
-
2.
Handlingar med allmän information
2.1
Parlamentets bulletin
-
Verksamhet
-
Sammanträdeskalendrar
-
Särskild utgåva för Europeiska rådets möten
-
Europaparlamentets verksamhet - efter plenarsammanträdet
2.2
News Alert / Direct agenda
2.3
3.
Officiella handlingar översända av andra institutioner
3.1
3.2
Rådet
-
3.3
3.4
Europeiska investeringsbanken
-
Meddelanden
3.5
Meddelanden
4.2
,
Europaparlamentets yttrande av den 3 maj 2001 och rådets beslut av den 28 maj 2001.
1.
I artikel 1 andra stycket i Fördraget om Europeiska unionen stadfästs principen om öppenhet genom att det anges att fördraget markerar en ny fas i processen för att skapa en allt fastare sammanslutning mellan de europeiska folken, där besluten skall fattas så öppet och så nära medborgarna som möjligt.
2.
Öppenhet bidrar till att stärka de principer om demokrati och respekt för grundläggande rättigheter som avses i artikel 6 i EU-fördraget och i Europeiska unionens stadga om de grundläggande rättigheterna.
3.
I de slutsatser som antogs av Europeiska rådet vid dess möten i Birmingham, Edinburgh och Köpenhamn underströks nödvändigheten av att göra arbetet vid unionens institutioner öppnare.
Denna förordning konsoliderar de initiativ som institutionerna redan tagit för att förbättra öppenheten i beslutsförfarandet.
4.
Syftet med denna förordning är att ge allmänhetens rätt till tillgång till handlingar största möjliga effekt och att fastställa allmänna principer och gränser för denna rätt i enlighet med artikel 255.2 i EG-fördraget.
5.
Eftersom Fördraget om upprättandet av Europeiska kol- och stålgemenskapen och Fördraget om upprättandet av Europeiska atomenergigemenskapen inte innehåller några bestämmelser om tillgång till handlingar bör Europaparlamentet, rådet och kommissionen söka ledning i denna förordning, i enlighet med förklaring nr 41 som fogas till slutakten till Amsterdamfördraget, beträffande handlingar som gäller verksamhet som omfattas av dessa båda fördrag.
6.
Sådana handlingar bör göras direkt tillgängliga i så stor utsträckning som möjligt.
7.
I enlighet med artikel 28.1 och artikel 41.1 i EU-fördraget är rätten till tillgång till handlingar tillämplig också på handlingar som gäller den gemensamma utrikes- och säkerhetspolitiken samt polisiärt och straffrättsligt samarbete.
Varje institution bör respektera sina säkerhetsbestämmelser.
8.
För att säkerställa att denna förordning tillämpas fullt ut i samband med all unionens verksamhet bör alla organ som inrättas av institutionerna tillämpa de principer som fastställs i denna förordning.
9.
10.
Det skall i detta sammanhang påpekas att en medlemsstat, enligt förklaring nr 35 som fogas till slutakten till Amsterdamfördraget, kan begära att kommissionen eller rådet inte vidarebefordrar en handling som härrör från den staten till tredje part, utan att medlemsstaten dessförinnan har lämnat sitt medgivande.
11.
12.
13.
För att säkerställa att rätten till tillgång till handlingar respekteras fullt ut bör ett administrativt förfarande med två steg tillämpas, där det dessutom skall vara möjligt att begära domstolsprövning eller framföra klagomål till ombudsmannen.
14.
För att medborgarna lättare skall kunna utöva sina rättigheter bör varje institution ge tillgång till ett register över handlingar.
15.
Denna förordning har varken till syfte eller effekt att ändra nationell lagstiftning om tillgång till handlingar; på grund av den princip om lojalt samarbete som styr förbindelserna mellan institutionerna och medlemsstaterna, är det dock uppenbart att medlemsstaterna bör se till att inte hindra en korrekt tillämpning av denna förordning och respektera institutionernas säkerhetsbestämmelser.
16.
Denna förordning påverkar inte tillämpningen av den rätt till tillgång till handlingar som medlemsstaterna, rättsliga myndigheter eller utredande organ redan har.
17.
EGT L 340, 31.12.1993, s.
43.
9).
58.
45).
27.
Artikel 1 Syfte
a)
att fastställa principer, villkor och gränser, under hänsynstagande till allmänna eller enskilda intressen, för rätten till tillgång till Europaparlamentets, rådets och kommissionens (nedan kallade institutionerna) handlingar i enlighet med artikel 255 i EG-fördraget på ett sätt som garanterar största möjliga tillgång till handlingar,
b)
c)
1.
2.
3.
Denna förordning skall tillämpas på alla handlingar som finns hos en institution, det vill säga handlingar som upprättats eller mottagits och som innehas av institutionen, inom samtliga Europeiska unionens verksamhetsområden.
4.
Särskilt handlingar som upprättats eller mottagits under ett lagstiftningsförfarande skall göras direkt tillgängliga i enlighet med artikel 12.
5.
6.
Denna förordning skall inte påverka allmänhetens rätt till tillgång till handlingar som finns hos institutionerna, vilken kan följa av folkrättsliga instrument eller av rättsakter som institutionerna antagit för att genomföra dessa instrument.
Artikel 3 Definitioner
handling: allt innehåll, oberoende av medium (på papper eller lagrat i elektronisk form, ljud- och bildupptagningar samt audiovisuella upptagningar) som har samband med den policy, de åtgärder och de beslut som omfattas av institutionens ansvarsområde,
b)
Artikel 4 Undantag
1.
a)
-
allmän säkerhet,
-
försvar och militära frågor,
-
internationella förbindelser,
-
2.
-
-
3.
4.
5.
6.
7.
Artikel 6 Ansökningar
1.
2.
3.
4.
Artikel 7 Behandling av ursprungliga ansökningar
1.
En bekräftelse om mottagande skall skickas till sökanden.
2.
Om ansökningen helt eller delvis avslås får sökanden inom 15 arbetsdagar efter att ha mottagit institutionens besked ge in en bekräftande ansökan till institutionen med begäran om omprövning.
3.
I undantagsfall, t.ex. om en ansökan avser en mycket omfattande handling eller ett mycket stort antal handlingar, får den tidsfrist som anges i punkt 1 förlängas med 15 arbetsdagar, förutsatt att sökanden underrättas på förhand och att utförliga skäl anges.
4.
Artikel 8 Behandling av bekräftande ansökningar
1.
En bekräftande ansökan skall behandlas skyndsamt.
2.
3.
1.
2.
En ansökan om tillgång till en känslig handling i enlighet med de förfaranden som anges i artiklarna 7 och 8 skall behandlas enbart av personer som har rätt att befatta sig med sådana handlingar.
Utan att det påverkar tillämpningen av artikel 11.2 skall dessa personer även avgöra vilka hänvisningar till känsliga handlingar som kan göras i det offentliga registret.
3.
Känsliga handlingar skall registreras eller lämnas ut endast om den varifrån handlingen härrör givit sitt samtycke.
4.
5.
Medlemsstaterna skall vidta lämpliga åtgärder för att se till att principerna i den här artikeln och i artikel 4 respekteras vid behandling av ansökningar om tillgång till känsliga handlingar.
6.
Institutionernas bestämmelser om känsliga handlingar skall offentliggöras.
7.
1.
2.
3.
Handlingen skall ställas till förfogande i en befintlig version och i ett befintligt format (inklusive i elektroniskt eller i ett alternativt format såsom blindskrift, stor stil eller bandupptagning), med fullständigt beaktande av sökandens önskemål.
1.
Tillgång till registret bör ges i elektronisk form.
2.
Registret skall för varje handling innehålla ett referensnummer (inklusive i förekommande fall den interinstitutionella referensen), ämnet och/eller en kort beskrivning av innehållet i handlingen och det datum då handlingen mottogs eller upprättades och registrerades.
3
Institutionerna skall omedelbart vidta de åtgärder som är nödvändiga för att upprätta ett register som skall vara i bruk senast den 3 juni 2002.
Artikel 12 Direkt tillgång i elektronisk form eller via ett register
1.
Institutionerna skall i största möjliga utsträckning ge allmänheten direkt tillgång till handlingar i elektronisk form eller via ett register, i enlighet med den berörda institutionens bestämmelser.
2.
3.
4.
Om direkt tillgång inte ges via registret skall registret i största möjliga utsträckning ange var handlingen finns.
1.
Utöver de akter som avses i artikel 254.1 och 254.2 i EG-fördraget och artikel 163 första stycket i Euratomfördraget skall följande handlingar offentliggöras i Officiella tidningen, om inte annat följer av artiklarna 4 och 9 i denna förordning:
a)
b)
c)
De rambeslut och de beslut som avses i artikel 34.2 i EU-fördraget.
d)
Konventioner som har utarbetats av rådet enligt artikel 34.2 i EU-fördraget.
e)
Konventioner undertecknade mellan medlemsstater på grundval av artikel 293 i EG-fördraget.
f)
Internationella avtal som ingåtts av gemenskapen eller i enlighet med artikel 24 i EU-fördraget.
2.
I största möjliga utsträckning skall följande handlingar offentliggöras i Officiella tidningen:
a)
Initiativ som lagts fram för rådet av en medlemsstat i enlighet med artikel 67.1 i EG-fördraget eller i enlighet med artikel 34.2 i EU-fördraget.
b)
Gemensamma ståndpunkter enligt artikel 34.2 i EU-fördraget.
c)
3.
Varje institution får i sin arbetsordning fastställa vilka övriga handlingar som skall offentliggöras i Officiella tidningen.
Artikel 15 Förvaltningsrutiner inom institutionerna
Artikel 16 Mångfaldigande av handlingar
Denna förordning skall inte påverka tillämpningen av befintliga bestämmelser om upphovsrätt som kan begränsa tredje parts rätt att mångfaldiga eller utnyttja handlingar som lämnats ut.
Artikel 18 Tillämpningsåtgärder
Artikel 19 Ikraftträdande
Den skall tillämpas från och med den 3 december 2001.
BILAGA
XVI a
Riktlinjer för tolkning av ordningsreglerna för ledamöterna
1.
Åtskillnad bör göras mellan å ena sidan synliga former av uppträdande som kan godtas under förutsättning att uppträdandet inte är kränkande och/eller förolämpande, faller inom rimliga gränser och inte skapar konflikt, och å andra sidan sådana som direkt stör någon form av parlamentarisk verksamhet.
2.
a)
Parlamentet ska ta särskild hänsyn till könsfördelningen.
b)
i.
Om den nominerade kommissionsledamotens ansvarsområde omfattas av ett enda parlamentsutskotts behörighetsområde, utfrågas han eller hon enbart av detta utskott.
ii.
iii.
Om den nominerade kommissionsledamotens ansvarsområde omfattas av huvudsakligen ett parlamentsutskotts behörighetsområde och i mindre omfattning ett eller flera andra parlamentsutskotts behörighetsområden, utfrågas han eller hon av det utskott som huvudsakligen är behörigt, som ska inbjuda det eller de övriga parlamentsutskotten att närvara vid utfrågningen.
Den valda kommissionsordföranden ska utförligt höras om förfarandena.
Antalet skriftliga sakfrågor får vara högst fem per behörigt parlamentsutskott.
De nominerade kommissionsledamöterna ska uppmanas att hålla ett inledande anförande på högst 20 minuter.
Före utfrågningens slut ska den nominerade kommissionsledamoten beredas möjlighet att hålla ett kort slutanförande.
Utskotten ska efter utfrågningen utan dröjsmål sammanträda för att göra en bedömning av den enskilda nominerade kommissionsledamoten.
Dessa sammanträden ska hållas inom stängda dörrar.
Som avslutning på debatten får en politisk grupp eller minst fyrtio ledamöter lägga fram ett resolutionsförslag.
Artikel 103.3, 103.4 och 103.5 ska tillämpas.
Omröstningen får skjutas upp till det därpå följande sammanträdet.
2.
Tillämpningsområde
och utarbetats på grundval av artikel 192 i EGfördraget och artikel 39 i arbetsordningen.
(b) Strategiska betänkanden
(
Kvoter
2.
För utskott med underutskott ska denna kvot utökas med ett betänkande per underutskott.
Detta ytterligare betänkande ska utarbetas av underutskottet.
Följande betänkanden ingår inte i denna kvot:
- Initiativbetänkanden som avser rättsakter.
2.
3.
Handlingen ska översändas på Europeiska unionens samtliga officiella språk.
4.
tillstånd
3.
En begäran om tillstånd att utarbeta strategiska betänkanden ska beviljas av utskottsordförandekonferensen efter det att eventuella behörighetskonflikter har lösts.
4.
talmanskonferensen och lösning av behörighetskonflikter
5.
Talmanskonferensen ska fatta ett beslut om varje begäran om tillstånd att utarbeta initiativbetänkanden som avser rättsakter och initiativbetänkanden som inte avser rättsakter inom högst fyra arbetsveckor efter det att de vidarebefordrats till utskottsordförandekonferensen, såvida talmanskonferensen inte beslutar att förlänga denna frist på grund av särskilda omständigheter.
6.
Om ett utskotts behörighet att utarbeta ett betänkande bestrids, ska talmanskonferensen fatta ett beslut inom sex arbetsveckor på grundval av en rekommendation från utskottsordförandekonferensen eller, i avsaknad av en sådan, från ordföranden för utskottsordförandekonferensen.
Om talmanskonferensen inte har fattat ett beslut inom denna frist anses rekommendationen vara godkänd
Artikel
4
1.
Utskottsordförandekonferensen ska vid sitt månatliga sammanträde behandla varje begäran om att få utarbeta initiativbetänkanden och om tillämpning av artikel 47.
3.
Om talmanskonferensen inte har fattat ett beslut inom denna frist anses rekommendationen vara godkänd
Artikel
5
Slutbestämmelser
1.
2.
- Talmanskonferensens beslut av den 9 december 1999 om förfarandet för beviljande av tillstånd att utarbeta initiativbetänkanden i enlighet med artikel 45 i arbetsordningen och talmanskonferensens beslut av den 15 februari och 17 maj 2001 om uppdatering av bilagan till detta beslut.
- Talmanskonferensens beslut av den 15 juni 2000 om förfarandet för beviljande av tillstånd att utarbeta betänkanden om handlingar som Europeiska unionens övriga institutioner eller organ förelagt parlamentet för kännedom.
BILAGA
1
De mänskliga rättigheterna i världen och EU:s politik i detta sammanhang - (Utskottet för utrikesfrågor)
Övervakning och tillämpning av gemenskapslagstiftningen - (Utskottet för rättsliga frågor)
Arbetet i den gemensamma parlamentariska AVS-EU-församlingen - (Utskottet för utveckling)
Jämställdhet mellan kvinnor och män i EU - (Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män)
Rapport om sammanhållningen - (Utskottet för regionalpolitik)
Skydd av gemenskapens finansiella intressenkampen mot bedrägerier - (Budgetkontrollutskottet)
De offentliga finanserna i EMU - (Utskottet för ekonomi och valutafrågor)
ECB:s årsrapport - (Utskottet för ekonomi och valutafrågor)
Rapport om konkurrenspolitik - (Utskottet för ekonomi och valutafrågor)
Årsrapport om konsumentskydd - (Utskottet för den inre marknaden)
BILAGA
2
ÅRLIGA VERKSAMHETS- OCH ÖVERVAKNINGSRAPPORTER SOM OMFATTAS AV AUTOMATISKT TILLSTÅND OCH EN SÄRSKILD HÄNVISNING TILL ARBETSORDNINGEN (DESSA INGÅR INTE I KVOTEN PÅ SEX BETÄNKANDEN SOM FÅR UTARBETAS SAMTIDIGT)
Årsrapport om allmänhetens tillgång till parlamentets handlingar, artikel 97.7 i arbetsordningen - (Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor)
Politiska partier i Europa, artikel 200.6 i arbetsordningen - (Utskottet för konstitutionella frågor)
Arbetet i utskottet för framställningar, artikel 192.6 i arbetsordningen - (Utskottet för framställningar)
REGISTER
Romerska siffror hänvisar till bilagor.
Allmänhetens tillgång till handlingar
avslutning
IV.5
i kammaren
168
Anföranden
IV.1
Anhållan om yttrande
82
,
XIII.II
,
V.5
beslut
70
VI.XVIII
Arkiv
IX.2
47
,
81
AVS
VI.II
,
147
196
61
B
,
VI.V
70
kontroll över genomförandet
105
Budgetberäkning
IV.8
IV.3
,
XV
C
111
COSAC
124
D
Debatt
,
43
uppskjutande
165
,
170
,
,
VI.II
,
75
,
95
I.1
ledamöter
I
36
Ekonomiska och sociala kommittén
42
Ekonomisk politik
107
Ersättare /suppleanter
178
EU:s stadga om de grundläggande rättigheterna
96
eurogruppen
II
Europeiska centralbanken
102
frågor för skriftligt besvarande
111
utnämningar
102
103
29
172
VI.XX
,
103
,
II.a
108
19
,
II
24
,
32
,
99
,
120
98
,
32
VI.XVIII
Föredragande
57
,
59
,
61
-
64
,
80
,
134
24
,
115
,
130
-
133
48
,
53
-
54
,
60
,
65
115
131
,
II
59
168
43
80 a
brådskande
134
budget
69
-
70
,
45
förlikning
64
56
64
63
-
65
64
sammankallande av
63
Första behandlingen
34
-
37
,
40
,
49
-
56
,
66
avslutande
49
,
51
IV.4
i kammaren
51
-
53
i utskotten
35
-
37
,
42
-
50
54
-
56
190
Gemensam ståndpunkt
57
-
59
61
godkännande
67
122
ändring
62
Gemensamt resolutionsförslag
103
,
108
,
115
Gemensamt utkast
85
-
90
,
VI.I
,
VII.B
Gemenskapslagstiftning, förenkling
80
-
80 a
80
80 a
Gemenskapsrätten, tillämpning
176
,
VI.IX
,
VI.XVI
,
,
Generalsekretariatet
197
4
,
22
,
68
,
137
,
146
,
197
,
70
,
72
81
3
,
11
,
VI.XVI
9
,
VI.XVIII
34
,
75
,
VI.XVII
Grupper
29
,
31
-
32
,
177
29
30
30
178
31
H
Handlingar
140
,
203
,
VII.A
,
VII.B
,
XV
,
XVI
85
,
89
,
II
I
Immunitet
5
5
-
7
38 a
,
120
,
Internationella avtal
75
,
83
-
84
Kammaren
146
,
148
,
150
67
första behandlingen
51
ordningsföreskrifter
146
-
147
Europeiska centralbanken
102
194
-
53
112
anhållan om yttrande
40
ansvarsfrihet
70
XIV
frågor
108
-
110
52
genomförande
XII
99
98
62
,
142
tillbakadragande av förslag
54
,
61
-
99
årsrapport om tillämpningen av gemenskapsrätten
112
Kommittéförfarande
XII
62
,
154
-
155
3
,
11
,
127
79
Kontrollbefogenheter
81
XI
115
,
130
,
III
Kvestorer
9
,
I
frågor till
28
25
12
,
15
-
17
L
34
-
38
,
39
,
204 a
IX
9
99
IX
61
-
62
,
65
90
95
,
103
,
108
131
149
-
150
,
155
168
-
171
,
176
-
177
,
194
,
196
,
201
-
202
,
,
IV.3
,
V.4
4
56
144
100
Monetär politik
106
Motivering
42
,
44
,
48
,
202
Motivering, betänkande
150
Muntligt betänkande
134
Mänskliga rättigheter
75
,
91
,
95
,
115
,
III
,
123
-
177
98
12
nominerade kommissionsledamöter
99
talman
12
-
13
12
,
14
76
O
Oavslutade ärenden
203
i utskotten
89
,
92
,
183
plenarsammanträdenas
96
,
172
10
80 a
Ombudsmannen
194
-
195
X
avsättning
194
195
Omröstning
77
,
131
,
149
,
152
-
155
,
157
-
164
,
169
60
-
62
,
67
51
,
19
tredje behandlingen
65
uppskjuten
52
150
-
156
159
,
161
147
,
148
Ordning i kammaren
146
-
148
,
XVI.a
19
,
166
9
Ordningsregler
146
P
125
Parlamentets bulletin
28
Parlamentets sessioner
127
-
128
Parlamentets valperiod
126
Passerkort
9
5
32
Plenarsammanträden
IV
protokoll
-
47
,
92
-
29
,
31
-
32
,
177
-
178
17
,
182
,
28
IV.8
5
-
7
VI.XVI
172
28
28
utskott
184
148
R
118
192
9
,
,
XVI
,
94
,
113
-
114
,
59
190
från rådet
77
83
89
-
90
,
94
,
114
,
,
103
113
,
115
,
151
,
,
203
,
III
gemensamma
103
Revisionsrätten
V.1
,
V.6
,
VI.V
101
uttalanden
105
54
54
,
55
,
66
,
81
Rättslig grund
35
,
39
,
55
,
VI.IX
internationella avtal
83
Rättstatsprincipen
34
,
75
,
95
,
115
,
III
Röstförklaringar
19
,
163
158
parlamentet
183
Sammanträden
146
,
148
,
165
,
171
173
173 a
128
,
145
-
172
128
137
-
138
,
-
144
,
146
-
148
,
184
22
137
,
173
Sammanträdesperiod
126
-
40
77
89
Regionkommittén
118
-
83
Samtycke
75
83
,
95
31
politiska grupper
28
,
176
,
195
,
VII.A
VII.B
,
,
XVI
Session
126
-
116
,
142
Språk
22
,
139
,
143
,
176
,
X
92
-
94
,
148
,
XVI.a
omedelbara åtgärder
146
XVI.a
34
-
35
,
41
Suppleant/ersättare
178
86
128
141
-
145
,
147
Talarlista
143
,
169
Talartid
103
,
108
,
134
,
144
,
147
,
165
-
166
fördelning
115
,
142
,
III
145
Talmannen
151
uppgifter
19
,
22
,
109
,
115
,
119
,
141
-
147
198
-
200
22
28
sammansättning
23
uppgifter
24
,
147
,
200
upplysningsplikt
28
48
,
58
,
63
,
65
24
,
176
XV
till parlamentet
9
,
137
Tillåtlighet
109
110
19
,
62
Tilläggsbudget
IV
197
,
Tolkning
138
Traktamente
147
Tredje behandlingen
förlikning
63
-
64
65
i kammaren
65
Tredje land
82
82
,
190
associerade stater
190
190
förbindelser med
24
,
190
Tystnadsplikt
96
U
122
24
,
176
,
VIII
68
,
55
-
148
7
165
,
172
,
III
Utfrågningar
176
,
194
86
VI.I
,
VI.IX
,
VII.A
-
VI.XVI
177
,
185
,
,
81
,
182
protokoll
96
,
178
,
VI
sammansättning
24
,
177
sammanträden
22
,
43
,
59
,
96
,
101
-
102
,
106
156
,
181
-
184
suppleanter
178
174
-
175
tredje behandlingen
64
underutskott
179
,
181
,
179
3
179
168
Utskottsordförandekonferensen
22
Uttalanden
105
103
87
kommissionen
103
rådet
103
V
Val
203
99
12
,
15
-
17
12
-
13
,
16
-
17
vice talmän
12
,
14
,
16
-
17
12
,
16
-
17
Y
Yttranden
83
40
-
41
parlamentet
134
,
185
rekommendationer från rådet
77
utskotten
35
,
179
193
,
V.1
Å
137
11
33
39
-
40
112
Årsrapport om tillämpningen av gemenskapsrätten
112
Åsidosättande
95
Återförvisning till utskott
40
,
52
-
53
,
165
,
168
,
V.4
IV.3
,
IV.6
204 a
Ä
Ändringar, kommissionens förslag
80 a
Ändringar, tillåtlighet
80 a
Ändringsförslag
150
53
bortfall
150
IV
frister
150
förfarande utan
43
,
131
185
kommissionens ståndpunkt
50
,
53
-
54
,
57
,
143
,
XIII
kompromissändringsförslag
53
,
59
,
62
,
muntliga
90
,
155
språk
138
-
139
,
150
tillbakadragande
150
tillåtlighet
19
150
utdelning
150
185
,
,
-
97
19
begäranden
19
UPPLYSNINGAR
I enlighet med parlamentets beslut om användningen av könsneutralt språk i sina handlingar har arbetsordningen anpassats för att ta hänsyn till de riktlinjer beträffande denna fråga som antogs av högnivågruppen för jämställdhet mellan kvinnor och män samt mångfald den 13 februari 2008 och som godkändes av presidiet den 19 maj 2008.
Europaparlamentets arbetsordning utges regelbundet som trycksak och publiceras i Europeiska unionens officiella tidning.
Den kan införskaffas genom distributionsställen tillhörande Byrån för Europeiska gemenskapernas officiella publikationer.
Europaparlamentet kan emellertid ändra sin arbetsordning.
Den gällande versionen av arbetsordningen finns på Europaparlamentets hemsida (http://www.europarl.europa.eu).
Kursiveringar i texten betyder att det rör sig om en tolkning av arbetsordningen (enligt artikel 201).
Utskottet för ekonomi och valutafrågor
ECON(2008)1013_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Måndagen den 13 oktober 2008, kl. 15.00–18.30
Bryssel
Lokal: ASP 3E2
1.
Godkännande av föredragningslistan
2.
Meddelanden från ordföranden
3.
Bekämpning av skatteundandragande i samband med gemenskapsinterna transaktioner (gemensamt system för mervärdesskatt)
ECON/6/61256
* 2008/0058(CNS) KOM(2008)0147 [01] – C6-0154/2008
Föredragande:
José Manuel García-Margallo Y Marfil (PPE–DE)
AM – PE412.256v01-00 PR – PE411.932v01-00
Ansv. utsk.:
ECON
Rådg. utsk.:
CONT, IMCO, JURI
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 18 september 2008 kl. 12.00
4.
Bekämpning av skatteundandragande i samband med gemenskapsinterna transaktioner
ECON/6/61260
* 2008/0059(CNS) KOM(2008)0147 [02] – C6-0155/2008
Föredragande:
José Manuel García-Margallo Y Marfil (PPE–DE)
PR – PE411.933v01-00
Ansv. utsk.:
ECON
Rådg. utsk.:
CONT, IMCO, JURI
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 18 september 2008 kl. 12.00
5.
Krav på offentlighet för medelstora företag och skyldigheten att upprätta sammanställd redovisning
ECON/6/62018
***I 2008/0084(COD) KOM(2008)0195 – C6-0173/2008
Föredragande:
Kristian Vigenin (PSE)
PA – PE412.235v01-00
Ansv. utsk.:
JURI
Ieke van den Burg (PSE)
PR – PE412.044v01-00
Rådg. utsk.:
ECON
· Behandling av ändringsförslag
6.
Europeiska revisionsrättens särskilda rapport nr 8/2007 om administrativt samarbete i fråga om mervärdesskatt
ECON/6/64122
2008/2151(INI)
Föredragande:
Bilyana Ilieva Raeva (ALDE)
PA – PE411.931v01-00 AM – PE412.326v01-00
Ansv. utsk.:
CONT*
Bart Staes (Verts/ALE)
PR – PE409.375v02-00 AM – PE412.175v01-00
Rådg. utsk.:
ECON*
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 22 september 2008 kl. 12.00
7.
Ett europeiskt initiativ för mikrokrediter för att främja tillväxt och sysselsättning
ECON/6/62863
2008/2122(INI) KOM(2007)0708
Föredragande:
Zsolt László Becsey (PPE–DE)
DT – PE414.015v01-00
Ansv. utsk.:
ECON
Rådg. utsk.:
BUDG, EMPL, ITRE, IMCO, JURI, FEMM
· Inledande diskussion
8.
Handel och ekonomiska förbindelser med Kina
ECON/6/65383
2008/2171(INI)
Föredragande:
Jorgo Chatzimarkakis (ALDE)
PA – PE412.345v01-00
Ansv. utsk.:
INTA
Corien Wortmann-Kool (PPE-DE)
Rådg. utsk.:
AFET, DEVE, ECON, ITRE, IMCO
· Behandling av förslag till yttrande
*** Omröstning ***
9.
EMU@10: Framsteg och utmaningar efter 10 år av den ekonomiska och monetära unionen
ECON/6/62761
2008/2156(INI) KOM(2008)0238
Med-föredragande:
Pervenche Berès (PSE) Werner Langen (PPE–DE)
PR – PE409.636v01-00 AM – PE412.060v01-00
Ansv. utsk.:
ECON
Rådg. utsk.:
INTA, EMPL
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 2 september 2008 kl. 12.00
10.
Allmänna regler för punktskatt
ECON/6/60115
* 2008/0051(CNS) KOM(2008)0078 – C6-0099/2008
Föredragande:
Astrid Lulling (PPE–DE)
AM – PE412.070v01-00 PR – PE407.726v02-00
Ansv. utsk.:
ECON
Rådg. utsk.:
CONT, ITRE, IMCO, REGI, AGRI
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 8 september 2008 kl. 12.00
11.
Europeiska revisionsrättens särskilda rapport nr 8/2007 om administrativt samarbete i fråga om mervärdesskatt
ECON/6/64122
2008/2151(INI)
Föredragande:
Bilyana Ilieva Raeva (ALDE)
PA – PE411.931v01-00 AM – PE412.326v01-00
Ansv. utsk.:
CONT*
Bart Staes (Verts/ALE)
PR – PE409.375v02-00 AM – PE412.175v01-00
Rådg. utsk.:
ECON*
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 22 september 2008 kl. 12.00
12.
Krav på offentlighet för medelstora företag och skyldigheten att upprätta sammanställd redovisning
ECON/6/62018
***I 2008/0084(COD) KOM(2008)0195 – C6-0173/2008
Föredragande:
Kristian Vigenin (PSE)
PA – PE412.235v01-00
Ansv. utsk.:
JURI
Ieke van den Burg (PSE)
PR – PE412.044v01-00
Rådg. utsk.:
ECON
· Antagande av förslag till yttrande
*** Omröstningen avslutas***
13.
Övriga frågor
14.
Tid och plats för nästa sammanträde (Bryssel)
Tisdagen den 4 november kl. 9.00–12.30 och 15.00–18.30 Onsdagen den 5 november kl. 9.00–12.30
Bröderna Dardenne tog hem Europaparlamentets filmpris
Kultur
2008-10-22 - 11:38
Filmen "Lornas tystnad" utsågs idag till vinnare av LUX-priset 2008.
Europaparlamentets talman Hans-Gert Pöttering överräckte priset till regissören Luc Dardenne inför de samlade ledamöterna i kammaren.
LUX-priset syftar till att bryta språkbarriärer och underlätta distribution av europeisk film inom EU.
- Jag skulle vilja tacka alla som har hjälpt till att producera den här filmen.
Vi ser inte varandras filmer och jag hoppas att det här priset kommer att bidra till att vi texter fler filmer och därmed ökar förståelsen, sa Luc Dardenne när han tog emot priset.
Filmen "Vid himlens utkant" av Faith Akin tilldelades LUX-priset 2007.
Vinnarfilmen textas på EU:s officiella 23 språk och en kopia i 35mm format anpassas till varje EU-land.
Vidare förses originalversionen med en textning för döva och hörselskadade personer samt eventuellt med hjälpmedel för personer med nedsatt syn.
De tre utvalda filmerna (Delta, Lornas tystnad och Citizen Havel) har visats i Europaparlamentet mellan den 15 september och 17 oktober.
Om filmen
Regi: Jean-Pierre och Luc Dardenne
Produktion: Belgien, Tyskland, Frankrike, Italien, Storbritannien
År: 2008
Speltid: 105 minuter
Originalversion: Fransk
För att Lorna ska kunna gifta sig med ryssen planerar Fabio att mörda Claudy.
SV
1
LINK
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
Kritik mot passageraruppgifter i brottsbekämpning
Rättsliga och inrikes frågor
2008-11-20 - 14:03
Europaparlamentet antog idag en resolution med 512 röster för, 5 emot och 19 nedlagda som kritiserar kommissionens förslag att upprätta ett så kallat PNR-system.
Förslaget, som presenterades för ett år sedan, innebär att flygbolag skulle lämna ut uppgifter som rör passagerare som flyger till eller från EU.
Dessa uppgifter skulle göras tillgängliga för myndigheter som arbetar med brottsbekämpning.
Europaparlamentet anser att brottsbekämpande myndigheter ska få alla de verktyg de behöver för att utföra sina uppdrag på lämpligt sätt, inklusive tillgång till uppgifter.
Resolutionsförslag
SV
1
LINK
/activities/plenary/ta/calendar.do?language=SV
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
Europaparlamentets talman fördömer terroristattackerna i Mumbai
Institutioner
2008-11-27 - 14:49
Europaparlamentets talman fördömer terroristattackerna i Mumbai Efter gårdagens terroristattacker i Mumbai (Bombay) gör Europaparlamentets talman Hans-Gert Pöttering följande uttalande:
"Jag fördömer å det kraftfullaste de många tragiska terroristattackerna som lett till att fler än hundra människor dödats och hundratals skadats.
Detta är ett brott som inte kan tolereras under några som helst omständigheter.
Terrorism utgör en av de största farorna mot säkerhet, stabilitet och demokratiska värderingar i det internationella samfundet.
På Europapaparlamentets vägnar vill jag uttrycka solidaritet med det indiska folket och deras myndigheter.
Kampen mot terrorism måste fortsätta vara en politisk prioritet för det internationella samfundet.
Det är ett globalt problem och en utmaning för alla.
Vi måste använda de verktyg som rättsväsendet ger oss för att tillsammans bekämpa terrorism en gång för alla."
Delegationen bestod av sju ledamöter från utskottet för internationell handel.
20081127IPR43127 Utskottet för Internationell handel
SV
1
PHOTO
20081124PHT42906.jpg
SV
2
LINK
/activities/committees/homeCom.do?language=SV&body=INTA
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//TEXT TA P6-TA-2008-0572 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2008-0573 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2008-0574 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2008-0575 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2008-0576 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2008-0577 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2008-0578 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2008-0579 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2008-0580 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2008-0581 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2008-0582 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2008-0583 0 DOC XML V0//SV
TECKENFÖRKLARING
*
Samrådsförfarandet
** I
** II
***
Samtyckesförfarandet
***I
Medbeslutandeförfarandet (första behandlingen)
***II
Medbeslutandeförfarandet (andra behandlingen)
***III
FÖRKORTNINGAR FÖR UTSKOTTENS NAMN
AFET:
DEVE:
Utskottet för utveckling
INTA:
Utskottet för internationell handel
BUDG:
Budgetutskottet
CONT:
Budgetkontrollutskottet
ECON:
Utskottet för ekonomi och valutafrågor
EMPL:
Utskottet för sysselsättning och sociala frågor
ENVI:
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
ITRE:
Utskottet för industrifrågor, forskning och energi
IMCO:
Utskottet för den inre marknaden och konsumentskydd
TRAN:
Utskottet för transport och turism
REGI:
Utskottet för regional utveckling
AGRI:
PECH:
Fiskeriutskottet
CULT:
Utskottet för kultur och utbildning
JURI:
Utskottet för rättsliga frågor
LIBE:
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
AFCO:
Utskottet för konstitutionella frågor
FEMM:
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
PETI:
Utskottet för framställningar
FÖRKORTNINGAR FÖR DE POLITISKA GRUPPERNA
PPE-DE:
Gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater
PSE:
Europeiska socialdemokratiska partiets grupp
ALDE:
Gruppen Alliansen liberaler och demokrater för Europa
UEN:
Gruppen Unionen för nationernas Europa
Verts/ALE
Gruppen De gröna/Europeiska fria alliansen
GUE/NGL:
Gruppen Europeiska enade vänstern/Nordisk grön vänster
IND/DEM:
Gruppen Självständighet/Demokrati
NI:
Grupplösa
Öppnande av sammanträdet
Inkomna dokument
Presentation av programmet för det tjeckiska ordförandeskapet (debatt)
Omröstning
Säkerhetsdetaljer och biometriska kännetecken i pass och resehandlingar ***I (omröstning)
Offentlig upphandling inom områdena för försvar och säkerhet ***I (omröstning)
Farliga ämnen och preparat (diklormetan) ***I (omröstning)
Bemyndigande för att ratificera ILO:s konvention om arbete i fiskenäringen från 2007 (konvention nr 188) * (omröstning)
Situationen för de grundläggande rättigheterna i Europeiska unionen 2004-2008 (omröstning)
Arbetstidens organisation för sjömän 2006 (förfaranden beträffande den sociala dialogen) (omröstning)
Utvecklingen för FN:s råd för mänskliga rättigheter, inbegripet EU:s roll (omröstning)
Allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar (omröstning)
Röstförklaringar
Rättelser/avsiktsförklaringar till avgivna röster
Justering av protokollet från föregående sammanträde
Situationen i Mellanöstern/Gaza (debatt)
Gasleverans från Ryssland till Ukraina och EU (debatt)
Frågestund (frågor till rådet)
Utskottens och delegationernas sammansättning
Situationen i Afrikas horn (debatt)
Europeiska unionens strategi för Vitryssland (debatt)
11 juli som dag till minne av offren för massakern i Srebrenica (debatt)
Föredragningslista för nästa sammanträde
Avslutande av sammanträdet
NÄRVAROLISTA
PROTOKOLL
ORDFÖRANDESKAP: Hans-Gert PÖTTERING Talman
1 Öppnande av sammanträdet
Sammanträdet öppnades kl. 09.05.
2 Inkomna dokument
Talmannen hade mottagit följande förslag till resolution från ledamöterna (artikel 113 i arbetsordningen):
- Philip Claeys, Koenraad Dillen och Frank Vanhecke.
Förslag till resolution om att anordna en folkomröstning om Europeiska unionens invandrings- och asylpolitik ( B6-0035/2009 ) hänvisat till ansvarigt utskott: LIBE
3
Presentation av programmet för det tjeckiska ordförandeskapet (debatt)
Uttalande av rådet:
Presentation av programmet för det tjeckiska ordförandeskapet
Mirek Topolánek (rådets tjänstgörande ordförande) gjorde ett uttalande.
Talare:
José Manuel Barroso (kommissionens ordförande) .
Talare:
Joseph Daul för PPE-DE-gruppen,
Martin Schulz för PSE-gruppen,
Graham Watson för ALDE-gruppen,
Brian Crowley för UEN-gruppen,
Monica Frassoni för Verts/ALE-gruppen,
Miloslav Ransdorf för GUE/NGL-gruppen,
Vladimír Železný för IND/DEM-gruppen,
Jana Bobošíková , grupplös, och
Mirek Topolánek .
ORDFÖRANDESKAP: Rodi KRATSA-TSAGAROPOULOU Vice talman
Talare:
Jan Zahradil ,
Libor Rouček ,
Silvana Koch-Mehrin ,
Konrad Szymański ,
Claude Turmes ,
Jiří Maštálka ,
Philippe de Villiers ,
Frank Vanhecke ,
Timothy Kirkhope ,
Kristian Vigenin ,
Adina-Ioana Vălean ,
Mario Borghezio ,
Milan Horáček ,
Adamos Adamou ,
Kathy Sinnott ,
Hartmut Nassauer ,
Enrique Barón Crespo ,
Lena Ek ,
Ģirts Valdis Kristovskis ,
Jacek Saryusz-Wolski ,
Jo Leinen ,
Andrew Duff ,
Bogdan Pęk ,
Stefano Zappalà ,
Bernard Poignant ,
Margarita Starkevičiūtė ,
Elmar Brok ,
Edite Estrela ,
Marco Cappato ,
Gunnar Hökmark ,
Maria Berger ,
Othmar Karas ,
Gary Titley ,
Josef Zieleniec ,
Proinsias De Rossa ,
Jerzy Buzek ,
Jan Andersson ,
Rumiana Jeleva ,
Katalin Lévai ,
Zuzana Roithová ,
Katerina Batzeli ,
John Bowis ,
Józef Pinior ,
Mihael Brejc ,
Richard Falbr ,
Zita Pleštinská ,
Miloš Koterec .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Tunne Kelam ,
Silvia-Adriana Ţicău ,
Marios Matsakis ,
Mirosław Mariusz Piotrowski ,
Dimitar Stoyanov .
Talare:
Mirek Topolánek och
José Manuel Barroso .
Talmannen förklarade debatten avslutad.
ORDFÖRANDESKAP: Luigi COCILOVO Vice talman
4 Omröstning
Omröstningsresultaten (ändringsförslag, särskilda omröstningar, delade omröstningar etc.) återfinns i bilagan ”Omröstningsresultat” som bifogas protokollet.
Bilagan med resultaten av omröstningarna med namnupprop finns endast i elektronisk form på Europarl.
4.1
Säkerhetsdetaljer och biometriska kännetecken i pass och resehandlingar ***I (omröstning)
Betänkande om förslaget till Europaparlamentets och rådets förordning om ändring av rådets förordning (EG) nr 2252/2004 om standarder för säkerhetsdetaljer och biometriska kännetecken i pass och resehandlingar som utfärdas av medlemsstaterna [ KOM(2007)0619 - C6-0359/2007 - 2007/0216(COD) ] - Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor.
Föredragande: Carlos Coelho ( A6-0500/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 1)
KOMMISSIONENS FÖRSLAG
Godkändes såsom ändrat av parlamentet
(
P6_TA(2009)0015
)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs
(
P6_TA(2009)0015
)
Inlägg
Före omröstningen meddelade talmannen att den franska sammanslutningen för politiska journalister Association des journalistes parlementaires hade uttryckt önskemål om att sammanträdesordföranden alltid skulle läsa upp resultaten av omröstningen.
Efter omröstningen protesterade
Francesco Enrico Speroni och
Edward McMillan-Scott
4.2
Offentlig upphandling inom områdena för försvar och säkerhet ***I (omröstning)
Betänkande om förslaget till Europaparlamentets och rådets direktiv om samordning av förfarandena vid tilldelning av vissa offentliga kontrakt för bygg- och anläggningsarbeten, varor och tjänster på försvars- och säkerhetsområdet [ KOM(2007)0766 - C6-0467/2007 - 2007/0280(COD) ] - Utskottet för den inre marknaden och konsumentskydd.
Föredragande: Alexander Graf Lambsdorff ( A6-0415/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 2)
KOMMISSIONENS FÖRSLAG
Godkändes såsom ändrat av parlamentet
(
P6_TA(2009)0016
)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs
(
P6_TA(2009)0016
)
4.3
Farliga ämnen och preparat (diklormetan) ***I (omröstning)
Betänkande om förslaget till Europaparlamentets och rådets beslut om ändring av rådets direktiv 76/769/EEG med avseende på begränsningar för utsläppande på marknaden och användning av vissa farliga ämnen och preparat (diklormetan) [ KOM(2008)0080 - C6-0068/2008 - 2008/0033(COD) ] - Utskottet för miljö, folkhälsa och livsmedelssäkerhet.
Föredragande: Carl Schlyter ( A6-0341/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 3)
KOMMISSIONENS FÖRSLAG
Godkändes såsom ändrat av parlamentet
(
P6_TA(2009)0017
)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs
(
P6_TA(2009)0017
)
4.4
Bemyndigande för att ratificera ILO:s konvention om arbete i fiskenäringen från 2007 (konvention nr 188) * (omröstning)
Betänkande om förslaget till rådets beslut om bemyndigande för medlemsstaterna att i Europeiska gemenskapens intresse ratificera ILO:s konvention om arbete i fiskenäringen från 2007 (konvention nr 188) [ KOM(2008)0320 - C6-0218/2008 - 2008/0107(CNS) ] - Utskottet för sysselsättning och sociala frågor.
Föredragande: Ilda Figueiredo ( A6-0423/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 4)
FÖRSLAG TILL LAGSTIFTNINGSRESOLUTION
Antogs
(
P6_TA(2009)0018
)
4.5
Situationen för de grundläggande rättigheterna i Europeiska unionen 2004-2008 (omröstning)
Betänkande om situationen för de grundläggande rättigheterna i Europeiska unionen 2004-2008 [ 2007/2145(INI) ] - Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor.
Föredragande: Giusto Catania ( A6-0479/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 5)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2009)0019
)
Inlägg
Under omröstningen lade
Mogens Camre fram ett muntligt ändringsförslag till punkt 32 (beaktades);
Syed Kamall yttrade sig om omröstningslistan och
Marco Cappato meddelade att det var den engelska versionen av punkt 166 som gällde.
4.6
Arbetstidens organisation för sjömän 2006 (förfaranden beträffande den sociala dialogen) (omröstning)
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 6)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2009)0020
)
4.7
Utvecklingen för FN:s råd för mänskliga rättigheter, inbegripet EU:s roll (omröstning)
Betänkande om utvecklingen för FN:s råd för mänskliga rättigheter, inbegripet EU:s roll [ 2008/2201(INI) ] - Utskottet för utrikesfrågor.
Föredragande: Laima Liucija Andrikienė ( A6-0498/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 7)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2009)0021
)
4.8
Allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar (omröstning)
Betänkande om allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar (genomförande av förordning (EG) nr 1049/2001) [ 2007/2154(INI) ] - Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor.
Föredragande: Marco Cappato ( A6-0459/2008 )
(Enkel majoritet erfordrades)
(Omröstningsresultat: bilagan "Omröstningsresultat", punkt 8)
RESOLUTIONSFÖRSLAG
Antogs
(
P6_TA(2009)0022
)
5 Röstförklaringar
Skriftliga röstförklaringar:
Muntliga röstförklaringar:
Betänkande Carlos Coelho - A6-0500/2008
Hubert Pirker ,
Zuzana Roithová ,
Frank Vanhecke ,
Dimitar Stoyanov
Betänkande Alexander Graf Lambsdorff - A6-0415/2008
Zuzana Roithová ,
Jim Allister ,
Carlo Fatuzzo
Betänkande Carl Schlyter - A6-0341/2008
Zuzana Roithová ,
Kathy Sinnott
Betänkande Ilda Figueiredo - A6-0423/2008
Zuzana Roithová
Betänkande Giusto Catania - A6-0479/2008
Irena Belohorská ,
Hubert Pirker ,
Peter Baco ,
Zuzana Roithová ,
Simon Busuttil ,
Péter Olajos ,
Jim Allister ,
Frank Vanhecke ,
Philip Claeys ,
Carlo Fatuzzo ,
Kathy Sinnott ,
Mairead McGuinness ,
Miroslav Mikolášik ,
Michl Ebner ,
Koenraad Dillen ,
Martin Callanan ,
Daniel Hannan ,
Ewa Tomaszewska ,
Gerard Batten ,
Christopher Heaton-Harris ,
Kinga Gál ,
László Tőkés ,
Georgs Andrejevs ,
John Attard-Montalto
Betänkande Marco Cappato - A6-0459/2008
Gay Mitchell ,
Zuzana Roithová ,
Syed Kamall
6 Rättelser/avsiktsförklaringar till avgivna röster
Den elektroniska versionen på Europarl uppdateras regelbundet under högst två veckor efter den aktuella omröstningsdagen.
Därefter slutförs förteckningen över rättelserna till de avgivna rösterna för att översättas och offentliggöras i Europeiska unionens officiella tidning.
° ° ° °
Alexander Graf Lambsdorff -
A6-0415/2008 .
Patrizia Toia hade låtit meddela att hennes omröstningsapparat inte hade fungerat vid omröstningen om betänkandet av
Marco Cappato -
A6-0459/2008 .
ORDFÖRANDESKAP: Hans-Gert PÖTTERING Talman
7 Justering av protokollet från föregående sammanträde
Protokollet från föregående sammanträde justerades.
8
Situationen i Mellanöstern/Gaza (debatt)
Uttalanden av rådet och kommissionen:
Situationen i Mellanöstern/Gaza
Karel Schwarzenberg (rådets tjänstgörande ordförande) och
Benita Ferrero-Waldner (ledamot av kommissionen) gjorde uttalanden.
Talare:
José Ignacio Salafranca Sánchez-Neyra för PPE-DE-gruppen,
Martin Schulz för PSE-gruppen,
Annemie Neyts-Uyttebroeck för ALDE-gruppen,
Cristiana Muscardini för UEN-gruppen,
Daniel Cohn-Bendit för Verts/ALE-gruppen,
Luisa Morgantini för GUE/NGL-gruppen,
Bastiaan Belder för IND/DEM-gruppen,
Luca Romagnoli , grupplös,
Elmar Brok ,
Pasqualina Napoletano ,
Marielle De Sarnez ,
Roberta Angelilli ,
Hélène Flautre ,
Kyriacos Triantaphyllides ,
Patrick Louis ,
Jim Allister ,
Rodi Kratsa-Tsagaropoulou ,
Hannes Swoboda ,
Chris Davies ,
Seán Ó Neachtain ,
David Hammerstein ,
Miguel Portas ,
Kathy Sinnott ,
Tokia Saïfi ,
Véronique De Keyser ,
Frédérique Ries ,
Feleknas Uca ,
Vladimír Železný ,
Gunnar Hökmark ,
Marek Siwiec ,
Philippe Morillon ,
Zbigniew Zaleski ,
Jelko Kacin ,
Jana Hybášková ,
Libor Rouček ,
Ioannis Kasoulides ,
Giulietto Chiesa ,
Stefano Zappalà ,
Maria Eleni Koppa ,
Struan Stevenson ,
Richard Howitt ,
Michael Gahler ,
Miguel Angel Martínez Martínez och
Geoffrey Van Orden .
ORDFÖRANDESKAP: Alejo VIDAL-QUADRAS Vice talman
Talare:
Proinsias De Rossa ,
Kinga Gál ,
Gay Mitchell och
Karel Schwarzenberg .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Sajjad Karim ,
Colm Burke ,
Nickolay Mladenov ,
Neena Gill ,
Marios Matsakis ,
Christopher Beazley ,
Antonio Masip Hidalgo ,
Margrete Auken ,
Peter Šťastný ,
Marian-Jean Marinescu ,
Bairbre de Brún ,
Czesław Adam Siekierski ,
Hannes Swoboda , vilken yttrade sig om organisationen av arbetet, och
Aurelio Juri .
Talare:
Benita Ferrero-Waldner .
-
Pasqualina Napoletano och
Hannes Swoboda för PSE-gruppen ,
om situationen i Mellanöstern/Gazaremsan ( B6-0051/2009 ) ,
-
Adamos Adamou ,
Daniel Cohn-Bendit ,
Monica Frassoni ,
David Hammerstein ,
Hélène Flautre ,
Caroline Lucas ,
Margrete Auken ,
Jill Evans ,
Angelika Beer och
Cem Özdemir för Verts/ALE-gruppen ,
om konflikten i Gazaremsan ( B6-0054/2009 ) ,
-
Joseph Daul ,
José Ignacio Salafranca Sánchez-Neyra ,
Elmar Brok ,
Jana Hybášková ,
Ioannis Kasoulides och
Gunnar Hökmark för PPE-DE-gruppen ,
om situationen i Mellanöstern och Gaza ( B6-0056/2009 ) ,
-
Francis Wurtz ,
Luisa Morgantini ,
Kyriacos Triantaphyllides ,
Miguel Portas och
Feleknas Uca för GUE/NGL-gruppen ,
om situationen i Mellanöstern/Gazaremsan ( B6-0057/2009 ) ,
-
Annemie Neyts-Uyttebroeck för ALDE-gruppen ,
om situationen i Gaza ( B6-0058/2009 ) ,
-
Cristiana Muscardini ,
Adam Bielan ,
Hanna Foltyn-Kubicka ,
Konrad Szymański ,
Eugenijus Maldeikis ,
Ryszard Czarnecki och
Marcin Libicki för UEN-gruppen ,
om situationen i Gaza ( B6-0059/2009 ) .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 6.3 i protokollet av den 15.01.2009
.
9
Gasleverans från Ryssland till Ukraina och EU (debatt)
Uttalanden av rådet och kommissionen:
Gasleverans från Ryssland till Ukraina och EU
Alexandr Vondra (rådets tjänstgörande ordförande) och
Andris Piebalgs (ledamot av kommissionen) gjorde uttalanden.
ORDFÖRANDESKAP: Gérard ONESTA Vice talman
Talare:
Jacek Saryusz-Wolski för PPE-DE-gruppen,
Hannes Swoboda för PSE-gruppen,
István Szent-Iványi för ALDE-gruppen,
Hanna Foltyn-Kubicka för UEN-gruppen,
Rebecca Harms för Verts/ALE-gruppen,
Esko Seppänen för GUE/NGL-gruppen,
Gerard Batten för IND/DEM-gruppen,
Jana Bobošíková , grupplös,
Giles Chichester ,
Jan Marinus Wiersma ,
Janusz Onyszkiewicz ,
Marcin Libicki ,
Bernard Wojciechowski ,
Irena Belohorská ,
Herbert Reul ,
Reino Paasilinna ,
Henrik Lax ,
Inese Vaidere ,
Dimitar Stoyanov ,
Charles Tannock ,
Adrian Severin ,
Toine Manders ,
Dariusz Maciej Grabowski ,
Nickolay Mladenov ,
Atanas Paparizov ,
Metin Kazak ,
Eugenijus Maldeikis ,
John Purvis ,
Dariusz Rosati och
Bilyana Ilieva Raeva .
ORDFÖRANDESKAP: Diana WALLIS Vice talman
Talare:
Romana Jordan Cizelj ,
Szabolcs Fazakas ,
Ivo Belet och
Zbigniew Zaleski .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Zita Pleštinská ,
Evgeni Kirilov ,
Fiona Hall ,
András Gyürk och
Eluned Morgan .
Talare:
Alexandr Vondra ,
Benita Ferrero-Waldner (ledamot av kommissionen) och
Andris Piebalgs .
Talmannen förklarade debatten avslutad.
10
Frågestund (frågor till rådet)
B6-0001/2009 ).
Fråga 1 (Milan Horáček): Rättssystemet i Ryssland
H-0968/08 .
H-0999/08 .
H-1008/08 .
Talare:
Daniel Hannan .
Fråga 4 (Marian Harkin): Liberalisering av världshandeln
H-0969/08 .
Fråga 5 (Seán Ó Neachtain): Framtiden för jordbrukspolitiken 2013-2020
H-0971/08 .
Seán Ó Neachtain ,
Avril Doyle och
se bilagan till det fullständiga förhandlingsreferatet
) .
ORDFÖRANDESKAP: Marek SIWIEC Vice talman
11 Utskottens och delegationernas sammansättning
Grupperna PPE-DE och PSE hade begärt att följande utnämningar skulle godkännas:
utskottet JURI:
Eva-Riitta Siitonen
utskottet FEMM:
Eva-Riitta Siitonen
delegationen för förbindelserna med Folkrepubliken Kina:
Eva-Riitta Siitonen
delegationen till den gemensamma parlamentarikerkommittén EU-Kroatien:
Hannes Swoboda i stället för
Aurelio Juri
delegationen för förbindelserna med Japan:
Aurelio Juri
Dessa utnämningar skulle betraktas som godkända om det inte framställdes några invändningar mot detta före justeringen av detta protokoll.
12
Situationen i Afrikas horn (debatt)
Uttalanden av rådet och kommissionen:
Situationen i Afrikas horn
Alexandr Vondra (rådets tjänstgörande ordförande) och
Benita Ferrero-Waldner (ledamot av kommissionen) gjorde uttalanden.
Talare:
Filip Kaczmarek för PPE-DE-gruppen,
Ana Maria Gomes för PSE-gruppen,
Johan Van Hecke för ALDE-gruppen,
Mikel Irujo Amezaga för Verts/ALE-gruppen,
Tobias Pflüger för GUE/NGL-gruppen ,
Karl von Wogau ,
Corina Creţu ,
Olle Schmidt ,
Eva-Britt Svensson och
Charles Tannock .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Rareş-Lucian Niculescu och
Alexandru Nazare .
Talare:
Alexandr Vondra och
Benita Ferrero-Waldner .
Karl von Wogau ,
Filip Kaczmarek och
Charles Tannock för PPE-DE-gruppen ,
Alain Hutchinson ,
Ana Maria Gomes ,
Glenys Kinnock ,
Marie-Arlette Carlotti och
Thijs Berman för PSE-gruppen ,
Renate Weber ,
Marco Cappato ,
Olle Schmidt ,
Johan Van Hecke och
Thierry Cornillet för ALDE-gruppen ,
Mikel Irujo Amezaga för Verts/ALE-gruppen ,
Cristiana Muscardini ,
Adam Bielan ,
Ryszard Czarnecki och
Konrad Szymański för UEN-gruppen ,
Luisa Morgantini och
Eva-Britt Svensson för GUE/NGL-gruppen ,
om situationen på Afrikas horn ( B6-0033/2009 ) .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 6.4 i protokollet av den 15.01.2009
.
13
Europeiska unionens strategi för Vitryssland (debatt)
Uttalanden av rådet och kommissionen:
Europeiska unionens strategi för Vitryssland
Alexandr Vondra (rådets tjänstgörande ordförande) och
Benita Ferrero-Waldner (ledamot av kommissionen) gjorde uttalanden.
Talare:
Jacek Protasiewicz för PPE-DE-gruppen,
Justas Vincas Paleckis för PSE-gruppen,
Janusz Onyszkiewicz för ALDE-gruppen,
Ryszard Czarnecki för UEN-gruppen,
Milan Horáček för Verts/ALE-gruppen,
Věra Flasarová för GUE/NGL-gruppen,
Bastiaan Belder för IND/DEM-gruppen,
Roberto Fiore , grupplös ,
Árpád Duka-Zólyomi ,
Józef Pinior ,
Zdzisław Zbigniew Podkański ,
Esther De Lange ,
Marianne Mikko ,
Ewa Tomaszewska ,
Colm Burke och
Sylwester Chruszcz .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Zita Pleštinská ,
Alessandro Battilocchio ,
Călin Cătălin Chiriţă ,
Czesław Adam Siekierski och
Flaviu Călin Rus .
Talare:
Alexandr Vondra och
Benita Ferrero-Waldner .
-
Annemie Neyts-Uyttebroeck ,
Jeanine Hennis-Plasschaert och
Janusz Onyszkiewicz för ALDE-gruppen ,
om EU:s strategi för Vitryssland ( B6-0028/2009 ) ,
-
Jan Marinus Wiersma för PSE-gruppen ,
om EU:s strategi för Vitryssland ( B6-0029/2009 ) ,
-
Elisabeth Schroedter ,
Hélène Flautre och
Milan Horáček för Verts/ALE-gruppen ,
om EU:s strategi för Vitryssland ( B6-0030/2009 ) ,
-
Konrad Szymański ,
Adam Bielan ,
Hanna Foltyn-Kubicka ,
Wojciech Roszkowski ,
Ryszard Czarnecki ,
Inese Vaidere och
Ģirts Valdis Kristovskis för UEN-gruppen ,
om EU:s strategi för Vitryssland ( B6-0031/2009 ) ,
-
Jacek Protasiewicz ,
José Ignacio Salafranca Sánchez-Neyra ,
Charles Tannock ,
Jacek Saryusz-Wolski ,
Elmar Brok ,
Colm Burke ,
Esther De Lange och
Vytautas Landsbergis för PPE-DE-gruppen ,
om Vitryssland ( B6-0032/2009 ) .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 6.5 i protokollet av den 15.01.2009
.
14
11 juli som dag till minne av offren för massakern i Srebrenica (debatt)
Uttalanden av rådet och kommissionen:
11 juli som dag till minne av offren för massakern i Srebrenica
Alexandr Vondra (rådets tjänstgörande ordförande) och
Benita Ferrero-Waldner (ledamot av kommissionen) gjorde uttalanden.
Talare:
Doris Pack för PPE-DE-gruppen,
Richard Howitt för PSE-gruppen,
Jelko Kacin för ALDE-gruppen,
Milan Horáček för Verts/ALE-gruppen,
Erik Meijer för GUE/NGL-gruppen,
Bastiaan Belder för IND/DEM-gruppen,
Dimitar Stoyanov , grupplös ,
Anna Ibrisagic och
Diana Wallis .
Följande talare yttrade sig i enlighet med förfarandet "catch the eye":
Zita Pleštinská ,
Pierre Pribetich ,
Jelko Kacin och
Călin Cătălin Chiriţă .
Talare:
Alexandr Vondra och
Benita Ferrero-Waldner .
-
Doris Pack för PPE-DE-gruppen ,
om utropandet av den 11 juli till europeisk minnesdag för offren för folkmordet i Srebrenica den 11 juli 1995 ( B6-0022/2009 ) ,
-
Hannes Swoboda och
Jan Marinus Wiersma för PSE-gruppen ,
om utropandet av den 11 juli till europeisk minnesdag för offren för folkmordet i Srebrenica den 11 juli 1995 ( B6-0023/2009 ) ,
-
Diana Wallis och
Jelko Kacin för ALDE-gruppen ,
om utropandet av den 11 juli till europeisk minnesdag för offren för folkmordet i Srebrenica den 11 juli 1995 ( B6-0024/2009 ) ,
-
Salvatore Tatarella ,
Ryszard Czarnecki ,
Konrad Szymański ,
Hanna Foltyn-Kubicka och
Adam Bielan för UEN-gruppen ,
om att införa den 11 juli som minnesdag för dem som föll offer för massakern i Srebrenica ( B6-0025/2009 ) ,
-
Erik Meijer och
André Brie för GUE/NGL-gruppen ,
om utropandet av den 11 juli till europeisk minnesdag för offren för folkmordet i Srebrenica den 11 juli 1995 ( B6-0026/2009 ) ,
-
Daniel Cohn-Bendit ,
Gisela Kallenbach ,
Angelika Beer ,
Raül Romeva i Rueda ,
Cem Özdemir ,
Sepp Kusstatscher och
Joost Lagendijk för Verts/ALE-gruppen ,
om utropandet av den 11 juli till europeisk minnesdag för offren för folkmordet i Srebrenica den 11 juli 1995 ( B6-0027/2009 ) .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 6.6 i protokollet av den 15.01.2009
.
15 Föredragningslista för nästa sammanträde
Föredragningslistan för nästa sammanträde fastställdes ("Föredragningslista" PE 418.510/OJJE).
16 Avslutande av sammanträdet
Sammanträdet avslutades kl. 23.35.
Harald R
ømer
Gérard Onesta
Generalsekreterare
Vice talman
NÄRVAROLISTA
Följande skrev på:
Adamou
Agnoletto
Aita
Albertini
Allister
Alvaro
Andersson
Andrejevs
Andrikienė
Angelakas
Angelilli
Antinucci
Arif
Arnaoutakis
Ashworth
Assis
Atkins
Attard-Montalto
Attwooll
Aubert
Audy
Auken
Ayala Sender
Aylward
Ayuso
Baco
Badia i Cutchet
Baeva
Barón Crespo
Barsi-Pataky
Bartolozzi
Basile
Batten
Battilocchio
Batzeli
Bauer
Beaupuy
Beazley
Becsey
Bedingfield
Beer
Belder
Belet
Belohorská
Bennahmias
Berend
Berès
Berger
Berlato
Berlinguer
Berman
Blokland
Bloom
Bobošíková
Bodu
Böge
Bösch
Bono
Borghezio
Borrell Fontelles
Boso
Boştinaru
Botopoulos
Boursier
Bowis
Bowles
Bozkurt
Bradbourn
Braghetto
Brejc
Brepoels
Breyer
Březina
Brie
Brok
van Buitenen
Bulfon
Bullmann
Bulzesc
Burke
Bushill-Matthews
Busk
Buşoi
Busquin
Busuttil
Buzek
Cabrnoch
Calia
Callanan
Camre
Capoulas Santos
Cappato
Carlotti
Carnero González
Carollo
Casa
Casaca
Cashman
Caspary
Castex
del Castillo Vera
Catania
Cavada
Cederschiöld
Cercas
Chatzimarkakis
Chichester
Chiesa
Chiriţă
Chmielewski
Christensen
Chruszcz
Chukolov
Ciani
Claeys
Clark
Cocilovo
Coelho
Cohn-Bendit
Colman
Corbett
Corda
Cornillet
Paolo Costa
Cottigny
Coûteaux
Cramer
Cremers
Corina Creţu
Gabriela Creţu
Crowley
Csibi
Marek Aleksander Czarnecki
Ryszard Czarnecki
Dăianu
Daul
David
Davies
De Blasio
de Brún
Degutis
Dehaene
De Keyser
Demetriou
De Michelis
Denanot
Deprez
De Rossa
De Sarnez
Descamps
Désir
Deß
Deva
De Veyrac
De Vits
Díaz de Mera García Consuegra
Dičkutė
Didžiokas
Dillen
Dimitrakopoulos
Dobolyi
Dombrovskis
Doorn
Douay
Dover
Doyle
Drčar Murko
Droutsas
Duchoň
Dührkop Dührkop
Duff
Duka-Zólyomi
Dumitriu
Ebner
Ehler
Ek
El Khadraoui
Esteves
Estrela
Ettl
Jill Evans
Jonathan Evans
Robert Evans
Färm
Fajmon
Falbr
Farage
Fatuzzo
Fava
Fazakas
Fernandes
Fernández Martín
Ferrari
Anne Ferreira
Elisa Ferreira
Figueiredo
Fiore
Fjellner
Flasarová
Flautre
Florenz
Foglietta
Foltyn-Kubicka
Fontaine
Ford
Fouré
Fourtou
Fraga Estévez
Fraile Cantón
França
Frassoni
Freitas
Friedrich
Funeriu
Gacek
Gahler
Gál
Gaľa
Galeote
Garcés Ramón
García-Margallo y Marfil
García Pérez
Gardini
Gargani
Garriga Polledo
Gaubert
Gauzès
Gawronski
Gebhardt
Gentvilas
Geringer de Oedenberg
Gewalt
Gibault
Gierek
Giertych
Gill
Giuntini
Gklavakis
Glante
Glattfelder
Goebbels
Goepel
Golik
Gollnisch
Gomes
Gomolka
Gottardi
Grabowska
Grabowski
Graça Moura
Gräßle
de Grandes Pascual
Grau i Segú
Grech
Griesbeck
Gröner
de Groen-Kouwenhoven
Grosch
Grossetête
Guardans Cambó
Guellec
Guerreiro
Guidoni
Gurmai
Gutiérrez-Cortines
Guy-Quint
Gyürk
Hänsch
Hall
Hammerstein
Hamon
Handzlik
Hannan
Harangozó
Harbour
Harkin
Harms
Hasse Ferreira
Heaton-Harris
Hedh
Helmer
Hénin
Hennicot-Schoepges
Hennis-Plasschaert
Herrero-Tejedor
Hieronymi
Higgins
Hökmark
Holm
Honeyball
Hoppenstedt
Horáček
Howitt
Hudacký
Hudghton
Hughes
Hutchinson
Hybášková
Ibrisagic
in 't Veld
Irujo Amezaga
Isler Béguin
Itälä
Iturgaiz Angulo
Jacobs
Jałowiecki
Janowski
Járóka
Jarzembowski
Jeggle
Jeleva
Jensen
Jöns
Jørgensen
Jonckheer
Jordan Cizelj
Jouye de Grandmaison
Juknevičienė
Juri
Kacin
Kaczmarek
Kallenbach
Kamall
Karas
Karim
Kasoulides
Kastler
Kaufmann
Kazak
Tunne Kelam
Kilroy-Silk
Kindermann
Kinnock
Kirilov
Kirkhope
Klaß
Klinz
Knapman
Koch
Koch-Mehrin
Konrad
Koppa
Korhola
Kósáné Kovács
Koterec
Kozlík
Krahmer
Krasts
Kratsa-Tsagaropoulou
Krehl
Kreissl-Dörfler
Kristovskis
Krupa
Kuc
Kuhne
Kušķis
Kusstatscher
Kuźmiuk
Lagendijk
Laignel
Lamassoure
Lambert
Lambrinidis
Landsbergis
Lang
De Lange
Langen
Langendries
Laperrouze
Lauk
Lavarra
Lax
Lebech
Lechner
Le Foll
Lefrançois
Lehideux
Lehne
Lehtinen
Leichtfried
Leinen
Jean-Marie Le Pen
Marine Le Pen
Le Rachinel
Lévai
Lewandowski
Liberadzki
Libicki
Lienemann
Liese
Lipietz
Locatelli
Lo Curto
López-Istúriz White
Losco
Louis
Lucas
Lulling
Lundgren
Luque Aguilar
Lynne
Lyubcheva
Maaten
McAvan
McCarthy
McDonald
McGuinness
McMillan-Scott
Madeira
Maldeikis
Manders
Mănescu
Maňka
Erika Mann
Thomas Mann
Marinescu
Marini
Markov
Marques
Martens
David Martin
Hans-Peter Martin
Martinez
Martínez Martínez
Masiel
Masip Hidalgo
Maštálka
Mathieu
Matsakis
Matsis
Matula
Mauro
Mavrommatis
Mayer
Mayor Oreja
Medina Ortega
Meijer
Méndez de Vigo
Menéndez del Valle
Meyer Pleite
Miguélez Ramos
Mikko
Mikolášik
Millán Mon
Mitchell
Mladenov
Mölzer
Moraes
Moreno Sánchez
Morgan
Morgantini
Morillon
Elisabeth Morin
Mote
Mulder
Musacchio
Muscardini
Mussa
Musumeci
Napoletano
Naranjo Escobar
Nassauer
Nattrass
Nazare
Neris
Newton Dunn
Neyts-Uyttebroeck
Nicholson
Nicholson of Winterbourne
Niculescu
Niebler
van Nistelrooij
Novak
Öger
Özdemir
Olajos
Olbrycht
Ó Neachtain
Onesta
Onyszkiewicz
Ortuondo Larrea
Őry
Ouzký
Oviir
Paasilinna
Pack
Pafilis
Paleckis
Panayotopoulos-Cassiotou
Panayotov
Pannella
Panzeri
Papadimoulis
Paparizov
Papastamkos
Parish
Paşcu
Patriciello
Pęk
Petre
Pflüger
Pieper
Pietikäinen
Pīks
Pinior
Piotrowski
Pirker
Pittella
Pleguezuelos Aguilar
Pleštinská
Podestà
Podkański
Pöttering
Pohjamo
Poignant
Polfer
Pomés Ruiz
Popa
Portas
Posdorf
Posselt
Prets
Pribetich
Protasiewicz
Purvis
Queiró
Quisthoudt-Rowohl
Rack
Raeva
Ransdorf
Rapkay
Rasmussen
Remek
Resetarits
Reul
Ribeiro e Castro
Riera Madurell
Ries
Rivera
Rizzo
Robsahm
Robusti
Rocard
Rodust
Rogalski
Roithová
Romagnoli
Rosati
Roszkowski
Rothe
Rouček
Roure
Rovsing
Rübig
Rühle
Rus
Rutowicz
Ryan
Sacconi
Saïfi
Sakalas
Saks
Salafranca Sánchez-Neyra
Salinas García
Sánchez Presedo
dos Santos
Sanzarello
Sanz Palacio
Sârbu
Sartori
Saryusz-Wolski
Savary
Savi
Schaldemose
Schapira
Schenardi
Schierhuber
Schinas
Schlyter
Frithjof Schmidt
Olle Schmidt
Schmitt
Schnellhardt
Schöpflin
Jürgen Schröder
Schroedter
Schulz
Schuth
Schwab
Seeber
Segelström
Seppänen
Severin
Siekierski
Siitonen
Silva Peneda
Simpson
Sinnott
Siwiec
Skinner
Škottová
Smith
Sógor
Sommer
Søndergaard
Sonik
Sornosa Martínez
Sousa Pinto
Spautz
Speroni
Staes
Staniszewska
Starkevičiūtė
Šťastný
Stauner
Stavreva
Sterckx
Stevenson
Stihler
Stockmann
Stolojan
Stoyanov
Strejček
Strož
Sturdy
Sudre
Sumberg
Surján
Susta
Svensson
Swoboda
Szájer
Szejna
Szent-Iványi
Szymański
Takkula
Tannock
Tarand
Tatarella
Teychenné
Thomsen
Ţicău
Titley
Toia
Tőkés
Tomaszewska
Tomczak
Toubon
Trakatellis
Trautmann
Triantaphyllides
Trüpel
Turmes
Tzampazi
Uca
Ulmer
Urutchev
Vaidere
Vakalis
Vălean
Vanhecke
Van Hecke
Van Lancker
Van Orden
Varela Suanzes-Carpegna
Varvitsiotis
Vatanen
Vaugrenard
Veneto
Ventre
Veraldi
Vergnaud
Vernola
Vidal-Quadras
Vigenin
de Villiers
Virrankoski
Visser
Vlasák
Vlasto
Wagenknecht
Wallis
Walter
Watson
Henri Weber
Manfred Weber
Weiler
Weisgerber
Westlund
Wieland
Wielowieyski
Wiersma
Wijkman
Willmott
Iuliu Winkler
Wise
von Wogau
Wohlin
Bernard Wojciechowski
Janusz Wojciechowski
Wortmann-Kool
Wurtz
Zahradil
Zaleski
Zapałowski
Zappalà
Zatloukal
Ždanoka
Zdravkova
Železný
Zieleniec
Zīle
Zimmer
Zlotea
Zvěřina
Zwiefka
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
FEMM(2009)0210_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Tisdagen den 10 februari 2009, kl. 9.00–12.30 och kl. 15.00–18.30
Bryssel
Lokal: PHS1A02
10 februari 2009 kl. 9.00–11.00
1.
Godkännande av föredragningslistan
2.
Justering av protokollen från sammanträdena den
· 12 januari 2009 PV – PE418.215v01-00
· 19–20 januari 2009 PV – PE418.295v01-00
3.
Meddelanden från ordföranden
4.
Åtgärder för att förbättra säkerhet och hälsa på arbetsplatsen för arbetstagare som är gravida, nyligen har fött barn eller ammar
FEMM/6/68375
***I 2008/0193(COD) KOM(2008)0637 – C6-0340/2008
Föredragande:
Edite Estrela (PSE)
DT – PE418.214v01-00
Ansv. utsk.:
FEMM*
Rådg. utsk.:
EMPL
Jamila Madeira (PSE)
PA – PE418.277v01-00
ITRE – Beslut: inget yttrande
· Behandling av arbetsdokument
5.
Integrering av ett jämställdhetsperspektiv i utskottens och delegationernas verksamheter
FEMM/6/66822
2008/2245(INI)
Föredragande:
Anna Záborská (PPE-DE)
PR – PE418.282v01-00
Ansv. utsk.:
FEMM
· Behandling av förslag till betänkande
· Fastställande av tidsfrist för ingivande av ändringsförslag
10 februari 2009 kl. 11.00–12.30
6.
Anonyma förlossningar – Offentlig utfrågning
10 februari 2009 kl. 15.00–16.00
***Omröstning (elektronisk omröstning)***
7.
Kampen mot kvinnlig könsstympning inom EU
FEMM/6/60405
2008/2071(INI)
Föredragande:
Cristiana Muscardini (UEN)
AM – PE416.657v01-00 PR – PE414.287v02-00 DT – PE412.171v02-00
Ansv. utsk.:
FEMM
· Antagande
· Tidsfrist för ingivande av ändringsförslag: 16 december 2008 kl. 12.00
8.
Patienträttigheter vid gränsöverskridande hälso- och sjukvård
FEMM/6/66116
***I 2008/0142(COD) KOM(2008)0414 – C6-0257/2008
Föredragande för yttrande:
Anna Záborská (PPE-DE)
PA – PE415.154v01-00 AM – PE418.322v01-00
Ansv. utsk.:
ENVI*
John Bowis (PPE–DE)
AM – PE418.320v01-00 AM – PE418.256v01-00 AM – PE418.304v01-00 PR – PE415.355v01-00 AM – PE418.293v01-00 AM – PE418.360v01-00 AM – PE418.342v01-00
· Antagande
· Tidsfrist för ingivande av ändringsförslag: 21 januari 2009 kl. 17.00
9.
Genomförande av principen om likabehandling av personer oavsett religion eller övertygelse, funktionshinder, ålder eller sexuell läggning
FEMM/6/65318
* 2008/0140(CNS) KOM(2008)0426 – C6-0291/2008
Föredragande för yttrande:
Donata Gottardi (PSE)
Ansv. utsk.:
LIBE*
Kathalijne Maria Buitenweg (Verts/ALE)
PR – PE418.014v02-00
· Antagande
· Tidsfrist för ingivande av ändringsförslag: 22 januari 2009 kl. 12.00
10.
Ansvarsfrihet 2007: EU:s allmänna budget, avsnitt III, kommissionen
FEMM/6/65819
2008/2186(DEC) SEK(2008)2359 [01] – C6-0415/2008
Föredragande för yttrande:
Lissy Gröner (PSE)
AM – PE418.359v01-00 PA – PE418.106v01-00
Ansv. utsk.:
CONT
Jean-Pierre Audy (PPE-DE)
· Antagande
· Tidsfrist för ingivande av ändringsförslag: 22 januari 2009 kl. 17.00
11.
En gemensam invandringspolitik för Europa: principer, åtgärder och verktyg
FEMM/6/71175
2008/2331(INI) KOM(2008)0359
Föredragande för yttrande:
Iratxe García Pérez (PSE)
AM – PE418.431v01-00 PA – PE418.283v01-00
Ansv. utsk.:
LIBE
Simon Busuttil (EPP–ED)
· Antagande
12.
En förnyad social agenda
FEMM/6/71168
2008/2330(INI) KOM(2008)0412
Föredragande för yttrande:
Marie Panayotopoulos-Cassiotou (PPE–DE)
AM – PE418.424v02-00 PA – PE418.261v02-00
Ansv. utsk.:
EMPL
José Albino Silva Peneda (PPE-DE)
PR – PE418.024v01-00
· Antagande
· Tidsfrist för ingivande av ändringsförslag: 26 januari 2009 kl. 17.00
13.
Jämställdhetsperspektivet i EU:s yttre förbindelser samt freds- och nationsuppbyggnad
FEMM/6/66838
2008/2198(INI)
Föredragande för yttrande:
Rodi Kratsa-Tsagaropoulou (PPE–DE)
PA – PE416.633v01-00 AM – PE418.358v01-00
Ansv. utsk.:
AFET
Libor Rouček (PSE)
· Antagande
· Tidsfrist för ingivande av ändringsförslag: 22 januari 2009 kl. 12.00
14.
Förenta nationernas konvention om rättigheter för personer med funktionsnedsättning
FEMM/6/66576
* 2008/0170(CNS) KOM(2008)0530 [01]
Föredragande för yttrande:
Hiltrud Breyer (Verts/ALE)
AM – PE418.363v01-00 PA – PE418.117v01-00
Ansv. utsk.:
EMPL
Rumiana Jeleva (PPE–DE)
PR – PE415.258v01-00 AM – PE418.419v01-00
· Antagande
· Tidsfrist för ingivande av ändringsförslag: 22 januari 2009 kl. 17.00
15.
Förenta nationernas konvention om rättigheter för personer med funktionsnedsättning (frivilligt protokoll)
FEMM/6/66578
* 2008/0171(CNS) KOM(2008)0530 [02]
Föredragande för yttrande:
Hiltrud Breyer (Verts/ALE)
PA – PE418.159v01-00
Ansv. utsk.:
EMPL
Rumiana Jeleva (PPE–DE)
AM – PE418.418v01-00 PR – PE415.259v01-00
· Antagande
*** Slut på omröstningen***
10 februari 2009 kl. 16.00–17.30
16.
Likabehandling av kvinnor och män som är egenföretagare
FEMM/6/68377
***I 2008/0192(COD) KOM(2008)0636 – C6-0341/2008
Föredragande:
Astrid Lulling (PPE-DE)
DT – PE419.918v01-00
Ansv. utsk.:
FEMM
Rådg. utsk.:
EMPL
Luigi Cocilovo (ALDE)
AM – PE418.266v01-00 PA – PE415.010v01-00
ITRE – Beslut: inget yttrande
JURI –
Lidia Joanna Geringer de Oedenberg (PSE)
PA – PE418.396v01-00
LIBE
· Behandling av arbetsdokument
17.
Övriga frågor
18.
Datum för nästa sammanträde
10 februari 2009 kl. 17.30–18.30
Europaparlamentet arbetar för jämställdhet
Kvinnors rättigheter/Lika möjligheter
2009-02-25 - 18:10
Lagstiftning, förslag, projektstöd och egna kampanjer är några viktiga verktyg för att skapa förbättringar.
Redan i grunden för EU-samarbetet som undertecknades 1957 slås principen om lika lön för lika arbete fast.
På mitten av 1970-talet kom de första direktiven om jämställdhet på arbetsplatsen.
Ökat inflytande
Europeiska kvinnor tjänar i genomsnitt 17 procent mindre än sina manliga kollegor.
Kamp mot kvinnovåld
1997 startade EU-stödprogrammet Daphne som nu är inne på sin tredje etapp (2007-2013).
Offentliga eller privata organisationer och institutioner kan söka stöd genom Daphne för verksamhet som förebygger våld mot kvinnor, barn och ungdomar samt skyddar våldsoffer och riskgrupper.
Rött kort till tvångsprostitution
Inför fotbolls-VM i Tyskland 2006 uppmärksammade kvinnoutskottet problemet med tvångsprostitution i samband med större idrottsevenemang.
- Kampanjen under namnet ”Rött kort till tvångsprostitution” var en stor framgång eftersom den i hög grad positivt bidrog till att minska människohandeln och tvångsprostitutionen under mästerskapet, säger utskottets ordförande Anna Záborská (EPP-ED*) från Slovakien.
Nytt jämställdhetsinstitut
2006 enades parlamentet och rådet om att inrätta ett jämställdhetsinstitut i Vilnius (Litauen).
SV
1
PHOTO
-//EP//TEXT IM-PRESS 20081117BRI42139 ITEM-006-SV NOT XML V0//SV
-//EP//TEXT IM-PRESS 20090119IPR46558 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
EU måste ge samlad hjälp till bilindustrin
Valet 2009
Industri
2009-03-25 - 14:22
EU måste bidra till vidareutbildning och omskolning Jobben i den europeiska bilindustrin är hotade och Europaparlamentet efterlyser ett ökat ekonomiskt stöd från EU och en bättre samordning mellan medlemsländerna.
Parlamentet antog idag en resolution om bilindustrins framtid med 413 röster för, 44 emot och 29 nedlagda.
Ledamöterna betonar att det handlar om en europeisk kris och efterlyser en verklig europeisk handlingsram med förslag på hur både EU och medlemsländerna kan vidta de åtgärder som krävs.
Parlamentet vill även se en strategi för förnyelse av fordonsparken, genom till exempel skrotningssystem, samt åtgärder för att stimulera billeasingmarknaden.
Ledamöterna uppmanar kommissionen att använda EU-fonder för arbetsmarknadsstöd för att bidra till vidareutbildning och omskolning av anställda som har förlorat eller riskerar att förlora sina jobb.
Moderaten Gunnar Hökmark (EPP-ED) framhöll att statsstöd måste syfta till att "garantera överlevnad" under den finansiella krisen, men inte "snedvrida konkurrensen mellan medlemsstater eller mellan biltillverkare".
Hökmark uppmanade kommissionen att säkerställa att inga övertramp sker av de regler som är uppställda.
Omröstning: 25.3.2009 20090324IPR52481 Antagna texter (preliminär utgåva, välj datum 25 mars) Kommissionens hemsida om bilindustrin
SV
1
PHOTO
SV
3
LINK
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
Utskottet för transport och turism
TRAN(2009)0330_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Måndagen den 30 mars 2009 kl. 15.00–18.30
Tisdagen den 31 mars 2009 kl. 9.00–12.30, kl. 15.00–16.00 (samordnarnas sammanträde) samt kl. 16.00–17.00
Bryssel
Lokal: PHS 4B001
30 mars 2009 kl. 15.00–18.30
1.
Godkännande av föredragningslistan
2.
Justering av protokollet från sammanträdet den
· 16 mars 2009 PV – PE421.399v01-00
3.
Europeiskt järnvägsnät för konkurrenskraftig godstrafik (text av intresse för EES)
TRAN/6/71395
***I 2008/0247(COD) KOM(2008)0852 – C6-0509/2008
Föredragande:
Petr Duchoň (PPE-DE)
AM – PE420.117v01-00 PR – PE418.273v01-00
Ansv. utsk.:
TRAN –
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 3 mars 2009 kl. 12.00
4.
Passagerares rättigheter vid resor till sjöss och på inre vattenvägar
TRAN/6/71099
***I 2008/0246(COD) KOM(2008)0816 – C6-0476/2008
Föredragande:
Michel Teychenné (PSE)
PR – PE418.200v01-00 AM – PE420.079v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
IMCO – Beslut: inget yttrande
JURI –
Georgios Papastamkos (PPE‑DE)
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 5 mars 2009 kl. 12.00
5.
Passagerares rättigheter vid busstransport
TRAN/6/71096
***I 2008/0237(COD) KOM(2008)0817 – C6-0469/2008
Föredragande:
Gabriele Albertini (PPE-DE)
AM – PE420.158v01-00 PR – PE418.207v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
IMCO – Beslut: inget yttrande
JURI – Beslut: inget yttrande
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 5 mars 2009 kl. 12.00
6.
Andra Marco Polo-programmet (Marco Polo II)
TRAN/6/71297
***I 2008/0239(COD) KOM(2008)0847 – C6-0482/2008
Föredragande:
Ulrich Stockmann (PSE)
AM – PE420.162v01-00 PR – PE418.255v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
BUDG –
AD – PE419.939v02-00
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 3 mars 2009 kl. 12.00
7.
Intelligenta transportsystem på vägtransportområdet och gränssnitt mot andra transportsätt
TRAN/6/71416
***I 2008/0263(COD) KOM(2008)0887 – C6-0512/2008
Föredragande:
AM – PE421.218v01-00 PR – PE418.288v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
ITRE – Beslut: inget yttrande
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 2 mars 2009 kl. 12.00
8.
Handlingsplanen för intelligenta transportsystem
TRAN/6/66695
2008/2216(INI)
Föredragande:
PR – PE418.162v02-00 AM – PE421.220v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
REGI –
Giovanni Robusti (UEN)
AD – PE416.672v02-00 AM – PE418.364v01-00
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 2 mars 2009 kl. 12.00
9.
Handlingsplanen för rörlighet i städerna
TRAN/6/66698
2008/2217(INI)
Föredragande:
Gilles Savary (PSE)
AM – PE419.860v01-00 PR – PE416.379v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
REGI –
Jean Marie Beaupuy (ALDE)
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 18 februari 2009 kl. 12.00
31 mars 2009, kl. 9.00–12.30
*** Elektronisk omröstning ***
10.
Tillträde till den internationella marknaden för godstransporter på väg (omarbetning)
TRAN/6/71863
***II 2007/0099(COD) 11788/1/2008 – C6-0014/2009 T6-0218/2008
Föredragande:
Mathieu Grosch (PPE-DE)
PR – PE418.415v01-00 AM – PE420.083v01-00
Ansv. utsk.:
TRAN –
· Antagande av förslag till andrabehandlingsrekommendation
· Tidsfrist för ingivande av ändringsförslag: 25 februari 2009 kl. 12.00
11.
Tillträde till marknaden för busstransporter (omarbetning)
TRAN/6/71865
***II 2007/0097(COD) 11786/1/2008 – C6-0016/2009 T6-0249/2008
Föredragande:
Mathieu Grosch (PPE-DE)
PR – PE418.416v01-00 AM – PE420.081v01-00
Ansv. utsk.:
TRAN –
· Antagande av förslag till andrabehandlingsrekommendation
· Tidsfrist för ingivande av ändringsförslag: 25 februari 2009 kl. 12.00
12.
Villkor som ska uppfyllas av personer som yrkesmässigt bedriver transporter på väg
TRAN/6/71864
***II 2007/0098(COD) 11783/1/2008 – C6-0015/2009 T6-0217/2008
Föredragande:
Silvia-Adriana Ţicău (PSE)
PR – PE418.445v01-00 AM – PE420.161v02-00
Ansv. utsk.:
TRAN –
· Antagande av förslag till andrabehandlingsrekommendation
· Tidsfrist för ingivande av ändringsförslag: 25 februari 2009 kl. 12.00
13.
Europeiskt järnvägsnät för konkurrenskraftig godstrafik (text av intresse för EES)
TRAN/6/71395
***I 2008/0247(COD) KOM(2008)0852 – C6-0509/2008
Föredragande:
Petr Duchoň (PPE-DE)
AM – PE420.117v01-00 PR – PE418.273v01-00
Ansv. utsk.:
TRAN –
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 3 mars 2009 kl. 12.00
14.
Passagerares rättigheter vid resor till sjöss och på inre vattenvägar
TRAN/6/71099
***I 2008/0246(COD) KOM(2008)0816 – C6-0476/2008
Föredragande:
Michel Teychenné (PSE)
PR – PE418.200v01-00 AM – PE420.079v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
IMCO – Beslut: inget yttrande
JURI –
Georgios Papastamkos (PPE‑DE)
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 5 mars 2009 kl. 12.00
15.
Passagerares rättigheter vid busstransport
TRAN/6/71096
***I 2008/0237(COD) KOM(2008)0817 – C6-0469/2008
Föredragande:
Gabriele Albertini (PPE-DE)
AM – PE420.158v01-00 PR – PE418.207v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
IMCO – Beslut: inget yttrande
JURI – Beslut: inget yttrande
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 5 mars 2009 kl. 12.00
16.
Andra Marco Polo-programmet (Marco Polo II)
TRAN/6/71297
***I 2008/0239(COD) KOM(2008)0847 – C6-0482/2008
Föredragande:
Ulrich Stockmann (PSE)
AM – PE420.162v01-00 PR – PE418.255v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
BUDG –
AD – PE419.939v02-00
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 3 mars 2009 kl. 12.00
17.
Intelligenta transportsystem på vägtransportområdet och gränssnitt mot andra transportsätt
TRAN/6/71416
***I 2008/0263(COD) KOM(2008)0887 – C6-0512/2008
Föredragande:
AM – PE421.218v01-00 PR – PE418.288v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
ITRE – Beslut: inget yttrande
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 2 mars 2009 kl. 12.00
18.
Handlingsplanen för intelligenta transportsystem
TRAN/6/66695
2008/2216(INI)
Föredragande:
PR – PE418.162v02-00 AM – PE421.220v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
REGI –
Giovanni Robusti (UEN)
AD – PE416.672v02-00 AM – PE418.364v01-00
19.
Avtal mellan Europeiska gemenskapen och Islamiska republiken Pakistan om vissa luftfartsaspekter
TRAN/6/59549
* 2008/0036(CNS) KOM(2008)0081 – C6-0080/2009
Föredragande:
Paolo Costa (ALDE)
PR – PE404.650v01-00
Ansv. utsk.:
TRAN –
· Antagande av förslag till betänkande
20.
Protokollet för tillämpning av Alpkonventionen på transportområdet (Transportprotokollet)
TRAN/6/71756
* 2008/0262(CNS) KOM(2008)0895 – C6-0073/2009
Föredragande:
Reinhard Rack (PPE-DE)
PR – PE421.126v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
ENVI – Beslut: inget yttrande
· Antagande av förslag till betänkande
21.
Grönboken om TEN-T-politikens framtid
TRAN/6/66700
2008/2218(INI)
Föredragande:
Eva Lichtenberger (Verts/ALE)
AM – PE420.159v01-00 PR – PE418.088v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
CONT – Beslut: inget yttrande
REGI –
Iratxe García Pérez (PSE)
AM – PE418.316v01-00 AD – PE418.034v02-00
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 18 februari 2009 kl. 12.00
22.
Handlingsplanen för rörlighet i städerna
TRAN/6/66698
2008/2217(INI)
Föredragande:
Gilles Savary (PSE)
AM – PE419.860v01-00 PR – PE416.379v01-00
Ansv. utsk.:
TRAN –
Rådg. utsk.:
REGI –
Jean Marie Beaupuy (ALDE)
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 18 februari 2009 kl. 12.00
*** Den elektroniska omröstningen avslutas ***
23.
Gemensamma regler för fördelning av ankomst- och avgångstider vid gemenskapens flygplatser
TRAN/6/74278
***I 2009/0042(COD) KOM(2009)0121 – C6-0097/2009
Föredragande:
Paolo Costa (ALDE)
Ansv. utsk.:
TRAN –
· Diskussion
31 mars 2009 kl. 15.00–16.00
24.
Samordnarnas sammanträde
Inom stängda dörrar
31 mars 2009 kl. 16.00–17.00
25.
Meddelanden från ordföranden
26.
Diskussion med
Europeiska miljöbyrån
27.
Övriga frågor
Parlamentet ställer sig bakom rätt till likabehandling
Valet 2009
Rättsliga och inrikes frågor
2009-04-02 - 13:14
Diskriminering förekommer på många håll i samhället, inte bara när det gäller jobb utan även i samband med banktjänster, transport, hälsa och utbildning.
Europaparlamentet ställde sig idag bakom direktivet om bättre likabehandling.
Kommissionens lagförslag tar upp diskriminering på grund av religion, funktionshinder, ålder och sexuell läggning.
Direktivet ska ses som ett komplement till tre andra direktiv mot diskriminering.
Europaparlamentet godkände kommissionens förslag, med några ändringar, med 363 röster för och 226 emot.
I den här frågan samråder rådet med parlamentet.
Parlamentet betonar vikten av tillgänglighet för funktionshindrade i allmänna transporter och byggnader.
Vid omröstningen antogs ändringsförslag om ett särskilt skydd för mikroföretag i likhet med den amerikanska medborgarrättslagen.
Ett annat ändringsförslag om att undanta reklam och medier från direktivets tillämpningsområde godkändes också.
Svenska inlägg i debatten
Socialdemokraten Inger SEGELSTRÖM (PES) uttrycket stöd för direktivet och sa sig vara "chockad" över förslag från kollegor att helt förkasta det.
Beslutsförfarande: Samråd (*)
LINK
/activities/plenary/ta/calendar.do?language=SV
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
Utskottet för regional utveckling
REGI(2009)0416_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Torsdagen den 16 april 2009, kl. 15.00–18.30
Bryssel
Lokal: PHS P1A2
1.
Godkännande av föredragningslistan
2.
Justering av protokollen från sammanträdena den
· 30–31 mars 2009 PV – PE423.725v01-00
3.
Meddelanden från ordföranden
I närvaro av rådet och kommissionen
4.
Diskussion med
Danuta Hübner, kommissionsledmot med ansvar för regionalpolitiken, och Luc Van den Brande, Regionkommitténs ordförande, om uppnått resultat på området för sammanhållningspolitiken under denna valperiod. (från kl. 15.15)
5.
Övriga frågor
6.
Datum för nästa sammanträde Det nya utskottets konstituerande sammanträde kommer troligtvis att hålla mellan den 16 och den 21 juli 2009.
-//EP//TEXT TA P6-TA-2009-0218 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0219 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0220 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0221 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0222 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0223 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0224 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0225 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0226 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0227 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0228 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0229 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0230 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0231 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0232 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0233 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0234 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0235 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0236 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0237 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0238 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0239 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0240 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0241 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0242 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0243 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0244 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0245 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0246 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0247 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0248 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0249 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0250 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0251 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0252 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0253 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0254 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0255 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0256 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0257 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0258 0 DOC XML V0//SV -//EP//TEXT TA P6-TA-2009-0259 0 DOC XML V0//SV
Fler produkter ska energimärkas
Energi
2009-05-05 - 11:03
Dels att märka alla energirelaterade produkter inom hushålls-, handels- och industrisektorerna, dels att utvidga tillämpningen till alla produkter som förbrukar energi direkt eller som orsaker energiförbrukning (t.ex. fönster).
Industriutskottet betonar i sin behandling av förslaget att reklam ska ge information om produktens energiförbrukning.
Vidare föreslår det skattelättnader för konsumenter och industri samt påpekar att myndigheter ska köpa energieffektiva produkter.
Ny gradering av energiklasser
Föredragande Anni Podimata (PES*, Grekland) menar att märkningssystemet måste bygga på den kunskap som konsumenterna redan har om A-G-skalan.
I takt med att energieffektiva produkter har ökat har allt fler produkter hamnat i A-kategorin.
Därför lade kommissionen i mars 2009 fram ett förslag som lägger till fler A-klasser (A-20%, A-40%, A-60% etc).
Industriutskottet är emot det nya formatet, och menar att det kan leda till förvirring över om 'A' står för mer eller mindre effektiva produkter.
20090504STO54874 EP Live - direktsändning Agenda Artikel: Liberalisering av energimarknaden Industriutskottet Betänkande Anni Podimata
SV
1
PHOTO
20080130PHT20001.jpg
SV
2
LINK
//eplive/public/livebroadcast_sv.htm
SV
3
LINK
/activities/plenary/home.do?language=SV
SV
5
LINK
/activities/committees/homeCom.do?language=SV&body=ITRE
SV
7
LINK
/members/public/yourMep/view.do?language=SV&partNumber=1&name=PODIMATA&id=39317
-//EP//TEXT IM-PRESS 20090420STO53928 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Valkvällen på Facebook
Valet 2009
Institutioner
2009-06-10 - 18:31
Europaparlamentets Facebooksida besöktes flitigt på valkvällen Europaparlamentets sida på Facebook har nu över 50 000 "fans".
Hundratals uppmanade andra att rösta innan de sista röstlokalerna stängde och kommentarsfälten fylldes under kvällen och natten av reaktioner, analyser och tankar om resultatet och valdeltagandet.
Exempelvis Xavier: "Snälla rösta, detta Europaval är viktigare än vad folk inser".
Valdeltagandet
Tania var nöjd att "min lilla, lilla stad i Italien nära havet har 65 %".
Bas däremot ifrågasatte EU: "Varför stoppar vi inte hela Europa-grejen.
Folk verkar inte bry sig överhuvudtaget."
Enligt Simone handlade "(...) nästan hela valkampanjen om nationella frågor.
Jag önskar att jag hade möjlighet att rösta på någon från andra europeiska länder.
Elisabeth skrev: "Huvudorsaken här i Österrike att inte rösta var att folk inte gillade kandidaterna ..."
Luca menade att "det har varit en stor brist på kommunikation - och ingen av de europeiska institutionerna har de senaste åren gjort tillräckligt för att informera folk".
Anne-Sophie tog upp att folk inte känner till vad Europaparlamentet gör: "Det är fortfarande alldeles för många människor som inte vet vad EU gör ... det är så sorgligt."
Platsfördelningen
Saerah: "Jag hade hoppats på ett lite rödare reslutat ... ledsen för PES, ja ..."
Marta: "Jag förstår inte varför mot bakgrund av den ekonomiska nedgången det är fler som röstar på högerpartier".
Frank: "Så bra att vara tysk nu.
Liberalerna (Alde) vann! ;-)).
Bryan: "Frankrike är grönt ♥ stolt att vara fransk".
Robert: "Vilken skamfylld dag för hela Europa ... först resultaten och sen valdeltagandet? vad är det för fel med Europa???
20090608STO56951 Europaparlamentet på Facebook Europaparlamentet på YouTube Preliminära valresultat och valdeltagande i hela EU och på nationell nivå (sidan uppdateras)
SV
1
PHOTO
20090608PHT56962.jpg
SV
2
LINK
http://www.facebook.com/europeanparliament
SV
3
LINK
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Informationskampanjen på nätet i siffror
Valet 2009
Institutioner
2009-06-11 - 16:50
EP Online Election campaign Inför valet har det varit ett stort intresse för Europaparlamentets 22-språkiga webbplats.
Under själva valveckan hade den nästan 2 miljoner besökare.
Som en del av informationskampanjen har parlamentet också varit på olika plattformar på nätet, exempelvis YouTube, Flickr, Facebook, MySpace och Twitter.
Den uppdaterades allteftersom resultaten kom in har haft 120 miljoner sidvisningar .
50 000 fans har diskuterat valet och hittat information på parlamentets sida på Facebook .
Tre "viral videos" lades ut på YouTube , tillsammans har de visats ungefär 440 000 gånger.
2 189 tweets på Twitter (22 språk).
Den 7 juni var Europavalet den tredje mest debatterade frågan på Twitter ("trending topic").
SV
1
PHOTO
20090611PHT57046.jpg
SV
2
LINK
http://www.elections2009-results.eu/en/new_parliament_sv.html
SV
3
LINK
/elections2009/default.htm?language=SV
SV
4
LINK
http://www.europarltv.eu/
SV
5
LINK
http://www.facebook.com/europeanparliament
SV
6
LINK
http://www.myspace.com/europeanparliament
SV
7
LINK
http://www.youtube.com/europeanparliament
SV
8
LINK
http://twitter.com/EU_Elections_en
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Videoporträtt av Jerzy Buzek
Utfrågningar
Institutioner
2009-07-15 - 15:52
Video: porträtt av Jerzy Buzek När Jerzy Buzek var ung drömde han om att bli parlamentsledamot i ett fritt Polen.
Han kom att fullfölja sin ambition och blev senare Polens premiärminister från 1997 till 2001.
Tisdag den 14 juli 2009 blev den 69-årige vetenskapsmannen Europaparlamentets talman efter att ha valts med 555 röster.
20090710STO58041 Första presskonferensen med nye talmannen - artikel 15/7 Jerzy Buzek vald till talman - pressmeddelande 14/7 Talmannens webbplats
SV
1
EUROPARL-TV
-//EP//TEXT IM-PRESS 20090710STO58042 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Föredragningslista
Torsdagen den 16 juli 2009
09:00 Omröstning
Meddelanden om talmanskonferensens förslag
Utnämningar i utskotten
--ooOOOoo--
fr.o.m kl. 10:30 Konstituerande sammanträden i utskotten
Tidsfrister
Meddelanden om talmanskonferensens förslag
Utnämningar i utskotten
Ändringsförslag
Onsdagen den 15 juli, 19:00
De svenska ledamöternas platser i Europaparlamentets utskott
Institutioner
Sverige
2009-07-20 - 17:04
Utskottet för utrikesfrågor
Ledamot:
Suppleant:
Utskottet för utveckling
Ledamot:
- Isabella Lövin (De gröna/EFA)
- Åsa Westlund (S-D)
Utskottet för internationell handel
Ledamot:
Suppleant:
- Carl Schlyter (De gröna/EFA)
- Göran FÄRM (S-D)
Budgetkontrollutskottet
Utskottet för ekonomi och valutafrågor
Ledamot:
Suppleant:
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Ledamot:
- Åsa Westlund (S-D)
- Lena Ek (ALDE)
- Marita Ulvskog (S-D)
Suppleant:
- Gunnar Hökmark (EPP)
Utskottet för den inre marknaden och konsumentskydd
Ledamot:
- Anna Hedh (S-D)
Utskottet för rättsliga frågor
Suppleant:
Vice ordförande:
- Lena Ek (ALDE) Utskottet för fiskeri
Ledamot:
- Isabella Lövin (De gröna/EFA)
Utskottet för kultur och utbildning
Inga svenska ledamöter
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Suppleant:
- Anna Maria CORAZZA BILDT (EPP, SE)
- Cecilia Wikström (ALDE)
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
Ordförande:
- Eva-Britt Svensson (GUE/NGL)
Utskottet för framställningar
Inga svenska ledamöter
Underutskottet för säkerhet och försvar
Suppleant:
- Anna Ibrisagic (EPP)
Ledamot:
- Eva-Britt Svensson (GUE/NGL)
SV
1
LINK
/members/expert/groupAndCountry/search.do?language=SV&country=IE
-//EP//DTD IM-PRESS 20050901 AVI DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 AVI DOC XML V0//EN
NÄRVAROLISTA
Följande skrev på:
Abad Damien
Áder János
Agnew John Stuart
Albertini
Albrecht Jan Philipp
Alfano Sonia
Alfonsi François
Allam Magdi Cristiano
Alvarez Magdalena
Alvaro
Alves Luís Paulo
Andreasen Marta
Andrikienė
Angelilli
Antinoro Antonello
Antonescu Elena Oana
Antoniozzi
Arif
Arlacchi Pino
Arsenis Kriton
Ashworth
Atkins
Attard-Montalto
Audy
Auken
Ayala Sender
Aylward
van Baalen Johannes Cornelis
Bach Georges
Badia i Cutchet
Balčytis Zigmantas
Balczó Zoltán
Baldassarre Raffaele
Balz Burkhard
Balzani Francesca
Barnier Michel
Bartolozzi
Băsescu Elena
Olejniczak
Batten
Baudis Dominique
Bauer
Becali George
Béchu Christophe
Belder
Belet
Bélier Sandrine
Benarab-Attou Malika
Bendtsen Bendt
Bennahmias
Berès
Berlato
Berlinguer Luigi
Besset Jean-Paul
Bielan
Bilbao Barandica Izaskun
Binev Slavi
Bisky Lothar
Bizzotto Mara
Blinkevičiūtė Vilija
Bloom
Böge
Bokros Lajos
Bonsignore
Bontes Louis
Borsellino Rita
Borys Piotr
Boştinaru Victor
Bové José
Bowles
Bozkurt
Myller
Brantner Franziska Katharina
Brepoels
Březina
Briard Auconie Sophie
Brok
Brons Andrew Henry William
Brzobohatá Zuzana
Bufton John
Bullmann
Buşoi
Busuttil
Bütikofer Reinhard
Buzek
Cadec Alain
Callanan
van de Camp Wim
Campbell Bannerman David
Cancian Antonio
Canfin Pascal
Capoulas Santos
Caronna Salvatore
Carvalho Maria Da Graça
Casa
Caspary
Castex
del Castillo Vera
Cavada
Cercas
Češková Andrea
Chatzimarkakis
Chichester
Childers Nessa
Chountis
Christensen
Philip Claeys
Clark
Coelho
Cofferati Sergio Gaetano
Cohn-Bendit
Colman Trevor
Comi Lara
Corazza Bildt Anna Maria
Cornelissen Marije
Correia De Campos António Fernando
Cortés Lastra Ricardo
Costa Silvia
Cozzolino Andrea
Cramer
Corina Creţu
Creutzmann Jürgen
Crocetta Rosario
Crowley
Cutaş George Sabin
Cymański Tadeusz
Ryszard Czarnecki
Daerden Frederic
Dăncilă Vasilica Viorica
Danjean Arnaud
Dantin Michel
Daul
David Mário
Davies
de Brún
Dehaene
De Keyser
Delli Karima
Delvaux Anne
de Magistris Luigi
De Mita
De Sarnez
Désir
Deß
Deutsch Tamás
Deva
De Veyrac
Díaz de Mera García Consuegra
Dodds Diane
Domenici Leonardo
Donskis Leonidas
Dorfmann Herbert
Duff
Durant Isabelle
Dušek Robert
Ehler
Ehrenhauser Martin
Eickhout Bas
Ek
El Khadraoui
Elles
Enciu Ioan
Engel Frank
Engström Christian
Eppink Derk Jan
Ernst Cornelia
Ertug Ismail
Essayah Sari
Estaras Ferragut Rosa
Estrela
Väyrynen
Fajmon
Fajon Tanja
Falbr
Farage
Färm
Feio Diogo
Ferber
Fernandes José Manuel
Ferreira João
Fidanza Carlo
Figueiredo
Fisas Ayxela Santiago
Fjellner
Beňová
Flautre
Fleckenstein Knut
Florenz
Fontana Lorenzo
Ford Vicky
Andersson
Fox Ashley
Fraga Estévez
Franco Gaston
Gahler
Gál
Gallagher
Gallo Marielle
García-Margallo y Marfil
García Pérez
Gardini Elisabetta
Garriga Polledo
Gauzès
Gebhardt
Geier Jens
Geringer de Oedenberg
Giegold Sven
Gierek
Girling Julie
Glante
Glattfelder
Godmanis Ivars
Konrad
Goerens Charles
Gollnisch
Gomes
Göncz Kinga
Goulard Sylvie
de Grandes Pascual
Gräßle
Grech
Grelier Estelle
Greze Catherine
Griesbeck
Griffin Nick
Gróbarczyk Marek Józef
Groote
Grosch
Grossetête
Gruny Pascale
Grzyb
Gualtieri Roberto
Guerrero Salom Enrique
Guillaume Sylvie
Gutiérrez-Cortines
Győri Enikő
Gyürk
Hadjigeorgiou Takis
Häfner Gerald
Haglund Carl
Hall
Händel Thomas
Handzlik
Hankiss Ágnes
Cederschiöld
Harbour
Harkin
Harms
Hassi
Haug
Häusling Martin
Hautala
Havel Jiří
Hedh
Helmer
Henin
Hennis-Plasschaert
Herczog
Herranz García
Hibner Jolanta Emilia
Higgins
Hirsch Nadja
Hoang Ngoc Liem
Hoarau Elie
Hohlmeier Monika
Hökmark
Poupakis
Howitt
Hübner Danuta Maria
Hudghton
Hughes
Husmenova
Iacolino Salvatore
Ibrisagic
Ilchev
Imbrasas Juozas
in 't Veld
Iotova Iliana Malinova
Itälä
Iturgaiz Angulo
Ivan Cătălin Sorin
Ivanova Iliana
Jaakonsaari Liisa
Jäätteenmäki
Jadot Yannick
Jahr Peter
Jauregui Atondo Ramon
Jazłowiecka Danuta
Jędrzejewska Sidonia Elżbieta
Jeggle
Jensen
Jimenez-Becerril Barrio Teresa
Joly Eva
de Jong Cornelis
Junqueras Vies Oriol
Juvin Philippe
Kacin
Kaczmarek
Kadenbach Karin
Kalfin Ivaylo
Kalinowski Jarosław
Kalniete Sandra
Kamall
Kamiński
Kammerevert Petra
Karas
Karim
Kariņš Arturs Krišjānis
Kasoulides
Kastler
Kazak Metin
Tunne Kelam
Keller Franziska
Kelly Alan
Kelly Seán
Kiil-Nielsen Nicole
Kirilov
Kirkhope
Klaß
Klinz
Klute Jürgen
Koch
Koch-Mehrin
Kohlíček
Kolarska-Bobińska Lena Barbara
Koppa Maria Eleni
Korhola
Kósa Ádám
Köstinger Elisabeth
Kovatchev Andrey
Kowal Paweł Robert
Kozlík
Kožušník Edvard
Krahmer
Kratsa-Tsagaropoulou Rodi
Krehl
Kreissl-Dörfler
Kuhn Werner
Kukan Eduard
Lamassoure
Lamberts Philippe
Lambrinidis
Lambsdorff
Landsbergis
Lange
De Lange
Langen
La Via Giovanni
Lechner
Le Foll
Legutko Ryszard Antoni
Lehne
Le Hyaric Patrick
Leichtfried
Lepage Corinne
Jean-Marie Le Pen
Marine Le Pen
Lewandowski
Lichtenberger
Liese
Liotard
Lisek Krzysztof
Lochbihler Barbara
Lövin Isabella
Lope Fontagné Veronica
López Aguilar Juan Fernando
López-Istúriz White
Lösing Sabine
Ludford
Ludvigsson Olle
Luhan Petru Constantin
Łukacijewska Elżbieta Katarzyna
Lulling
Lunacek Ulrike
Lynne
McAvan
McCarthy
Mcclarkin Emma
McGuinness
McMillan-Scott
Macovei Monica Luisa
Madlener Barry
Manders
Mănescu Ramona Nicole
Maňka
Thomas Mann
Manner Riikka
Marcinkiewicz Bogdan Kazimierz
Marinescu
David Martin
Hans-Peter Martin
Martínez Martínez
Masip Hidalgo
Maštálka
Mastella
Matera Barbara
Mathieu
Matias Marisa
Mato Adrover Gabriel
Matula Iosif
Mauro
Mavronikolas Kyriakos
Mayer
Mayor Oreja
Mazzoni Erminia
Meissner Gesine
Mélenchon Jean-Luc
Melo Nuno
Méndez de Vigo
Merkies Judith A.
Messerschmidt Morten
Meyer Pleite
Michel Louis
Migalski Marek Henryk
Mihaylova Nadezhda
Mikolášik
Milana Guido
Millán Mon
Mirskis Aleksandrs
Mölzer
Moraes
Moreira Vital
Morin
Morkūnaitė Radvilė
Morvai Krisztina
Motti Tiziano
Muñiz De Urquiza María Paloma
Muscardini
Nattrass
Nedelcheva Mariya
Neuser Norbert
Newton Dunn
Annemie Neyts-Uyttebroeck
Nicholson
Nicolai Norica
Niculescu Rareş-Lucian
Niebler
van Nistelrooij
Nitras Sławomir Witold
Obermayr Franz
Olbrycht
Olejniczak Wojciech Michał
Ford
Őry
Ouzký
Oviir
Pack
Padar Ivari
Paksas Rolandas
Paleckis
Pallone Alfredo
Panayotov Vladko Todorov
Panzeri
Papadopoulou Antigoni
Papastamkos
Pargneaux Gilles
Parvanova
Paşcu
Paška Jaroslav
Patriciello
Paulsen
Peillon
Perello Rodriguez Andres
Alojz Peterle
Pieper
Piotrowski
Pirillo Mario
Pittella
Plumb
Poc Pavel
Podimata Anni
Ponga Maurice
Poręba Tomasz Piotr
Portas
Posselt
Pöttering
Poupakis Konstantinos
Preda Cristian Dan
Vittorio Prodi
Protasiewicz
Provera Fiorello
Quisthoudt-Rowohl
Rangel Paulo
Ranner Hella
Rapkay
Rapti Sylvana
Reimers Britta
Remek
Repo Mitro
Reul
Riera Madurell
Ries
Rinaldi Niccolò
Riquet Dominique
Rivasi Michèle
Rivellini Crescenzio
Rochefort Robert
Rodust Ulrike
Roithová
Romero López Carmen
Romeva i Rueda
Ronzulli Licia
Rosbach Anna
Rossi Oreste
Roth-Behrendt
Rouček
Rübig
Rubiks Alfreds
Rühle
Saïfi
Salafranca Sánchez-Neyra
Salatto Potito
Salvini
Sanchez-Schmid Marie-Thérèse
Sánchez Presedo
Sârbu
Sargentini Judith
Sartori
Saryusz-Wolski
Saudargas Algirdas
Schaake Marietje
Schaldemose
Schlyter
Olle Schmidt
Schmitt
Schnellhardt
Schnieber-Jastram Birgit
Scholz Helmut
Schöpflin
Schroedter
Schulz
Schulz Werner
Schwab
Scicluna Edward
Scotta" Giancarlo
Scurria Marco
Seeber
Sehnalová Olga
Senyszyn Joanna
Serracchiani Debora
Severin
Siekierski
Silvestris Sergio Paolo Francesco
Simon Peter
Simpson
Sinclaire Nicole
Sippel Birgit
Siwiec
Skinner
Skrzydlewska Joanna Katarzyna
Skylakakis Theodoros
Smith
Smolková Monika
Sógor Csaba
Soini Timo
Sommer
Søndergaard
Sonik
Sosa Wagner Francisco
Soullie Catherine
Speroni
Obiols
Stassen Laurence J.A.J.
Šťastný
Stavrakakis Georgios
Steinruck Jutta
Sterckx
Stevenson
Stihler
van der Stoep Daniël
Stolojan Theodor Dumitru
Stoyanov
Stoyanov Emil
Strasser Ernst
Strejček
Striffler Michèle
Sturdy
Surján
Susta
Svensson Alf
Svensson
Swinburne Kay
Swoboda
Szymański
Tabajdi
Takkula
Tănăsescu Claudiu Ciprian
Tannock
Marc Tarabella
Tarand Indrek
Tatarella
Tavares Rui
Teixeira Nuno
Thaler Zoran
Thein Alexandra
Theocharous Eleni
Theurer Michael
Thomsen
Thun Und Hohenstein Róża, Gräfin von
Thyssen
Tirolien Patrice
Tőkés László
Tomaševski Valdemar
Tošenovský Evžen
Toussas
Trautmann
Tremopoulos Michail
Tremosa I Balcells Ramon
Triantaphyllides
Trüpel
Trzaskowski Rafał Kazimierz
Tsoukalas Ioannis
Turunen Emilie
Tzavela Niki
Uggias Giommaria
Ulmer
Ulvskog Marita
Ungureanu Traian
Urutchev Vladimir
Uspaskich Viktor
Vadim Tudor Corneliu
Vaidere
Vajgl Ivo
Vălean
Buşoi
Vanhecke
Bösch
Vattimo
Vaughan Derek
Vergiat Marie-Christine
Vergnaud
Verheyen Sabine
Verhofstadt Guy
McCarthy
Vigenin
de Villiers
Vlasák
Zdravkova
Wałęsa Jarosław Leszek
Wallis
Henri Weber
Weber Renate
Weiler
Werthmann Angelika
Westlund
Westphal Kerstin
Wieland
Wikström Cecilia
Willmott
Wils Sabine
Winkler Hermann
Winkler Iuliu
Włosowicz Jacek
Janusz Wojciechowski
Wortmann-Kool
Yannakoudakis Marina
Záborská
Zahradil
Zala Boris
Zalba Bidegain Pablo
Zalewski Paweł Ksawery
Zasada Artur
Ždanoka
Zeller Joachim
Zemke Janusz Władysław
Zīle
Zimmer
Ziobro Zbigniew
Zver Milan
Zwiefka
EU:s utrikesfrågor - många ämnen på agendan för nya Europaparlamentariker
Institutioner
2009-09-22 - 17:17
Dessa är några av de ämnen som de nya Europaparlamentarikerna kommer att ta itu med under hösten.
Här kan du läsa vad dessa utskott kommer att ha på agendan i höst.
Under slutet av året kommer alla utskott att genomföra intervjuer med de tilltänkta kommissionärerna inom deras expertområde.
När det gäller dessa fem utskott så kommer de att hålla utfrågningar med de tilltänkta kommissionärerna för Utrikesfrågor, Utveckling samt Handel.
Utrikesfrågor: Afghanistan och utvecklingsrapporter om kandidatländerna
Kommissionär Olli Rehn kommer att presentera årets utvecklingsrapporter den 15 oktober i utskottet för Utrikesfrågor.
Island ansökte om medlemskap den 23 juli.
Under de kommande månaderna kommer utskottet för Utveckling att se över Cotonouavtalet, vars mål är att minska och på sikt utrota fattigdomen samt att gradvis integrera staterna i Afrika, Västindien och Stillahavsområdet i världsekonomin.
Utskottet kommer också att förbereda en rapport som granskar finanskrisens effekt på utvecklingsländerna.
Dessutom kommer utskottet att delta i FN:s klimatkonferens i Köpenhamn i mitten av december.
Internationell handel: sociala och miljömässiga frågor på agendan
Utskottet för Internationell handel har bokat in två utfrågningar i november och december.
Den andra utfrågningen kommer att handla om hur sociala och miljömässiga frågor kan inkluderas i de internationella handelsavtalen.
Utskottet för säkerhet och försvar: utvärderar EU:s åtgärder mot pirater
Utskottet kommer att skicka en delegation till Djibouti i slutet av oktober för att utvärdera EU:s åtgärder för att förhindra piratattacker i Adenviken utanför Somalia.
Underutskottet mänskliga rättigheter: Sacharovpriset
Den 30 september kommer Europaparlamentarikerna att presentera de kandidater som de har utnämnt.
Den 6 oktober efter en omröstning i Strasbourg kommer en lista med tre kandidater att presenteras.
Den första resan för de nya Europaparlamentarikerna kommer att gå till Mozambique där det kommer att hållas val den 28 oktober.
Andra potentiella uppdrag är valet den 28 november i republiken Elfenbenskusten och den 6 december i Bolivia.
20090921STO60931 Lista över ständiga utskott The EU’s external relations Progress reports Sacharovpriset Somaliska pirater: lösningen finns på land
SV
1
PHOTO
20090915PHT60686.jpg
SV
2
LINK
/activities/committees/committeesList.do?language=SV
SV
3
LINK
/parliament/expert/displayFtu.do?language=EN&ftuId=theme6.html&id=73
SV
4
LINK
http://ec.europa.eu/enlargement/how-does-it-work/progress_reports/index_en.htm
SV
5
LINK
/sakharov/default_sv.htm
-//EP//TEXT IM-PRESS 20081211STO44303 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
EUROPAPARLAMENTET
2009 - 2014
Utskottet för utrikesfrågor
AFET(2009)0928_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Måndagen den 28 september 2009, kl. 15.00–18.30
Tisdagen den 29 september 2009, kl. 9.00–12.30 och kl. 15.00–18.30
Onsdagen den 30 september 2009, kl. 9.00–13.00
Bryssel
Lokal: JAN 2 Q 2
1.
Godkännande av föredragningslistan
2.
Justering av protokollet från sammanträdena den
· 1–2 september 2009 PV – PE427.984v01-00
· 10 september 2009 PV – PE428.139v01-00
3.
Meddelanden från ordföranden
4.
Antagande av sammanträdeskalendern för 2010
5.
Övriga frågor
28 september 2009 kl. 15.00
INOM STÄNGDA DÖRRAR
INOM STÄNGDA DÖRRAR
7.
Det utvidgade presidiet (se separat program)
29 september 2009 kl. 10.30–12.30
8.
Inrättande av ett finansieringsinstrument för samarbete med industriländer (ändring av förordning (EG) nr 1934/2006)
AFET/7/00010
* 2009/0059(CNS) KOM(2009)0197 – C7-0101/2009
Ansv. utsk.:
INTA –
Helmut Scholz (GUE/NGL)
· Diskussion
9.
Upprättande av stabilitetsinstrumentet
AFET/7/00005
***I 2009/0058(COD) KOM(2009)0195 – C7-0042/2009
Ansv. utsk.:
AFET –
Rådg. utsk.:
DEVE –
Eva Joly (Verts/ALE)
PA – PE428.241v01-00
INTA – Beslut: inget yttrande
· Diskussion
10.
Förteckningen över tredjeländer vars medborgare omfattas av eller är undantagna från viseringskrav när de passerar medlemsstaternas yttre gränser
AFET/7/00448
* 2009/0104(CNS) KOM(2009)0366 – C7-0112/2009
Ansv. utsk.:
LIBE –
Tanja Fajon (S&D)
PR – PE428.146v01-00
· Diskussion
· Tidsfrist för ingivande av ändringsförslag: 1 oktober 2009 kl. 12.00
29 september 2009 kl. 15.00–16.30
11.
Diskussion med Benita Ferrero-Waldner, kommissionsledamot med ansvar för yttre förbindelser och den europeiska grannskapspolitiken, om resultatet av ministerveckan vid FN:s generalförsamling och om kommissionens meddelande om en ny agenda för EU:s förbindelser med Latinamerika
29 september 2009 kl. 17.00
Tillsammans med delegationen till den parlamentariska samarbetskommittén EU ‑ Moldavien
12.
Diskussion med Vlad Filat, Moldaviens premiärminister, i sällskap med Iurie Leanca, Moldaviens utrikesminister, om den nuvarande politiska situationen i Moldavien efter parlamentsvalet den 29 juli 2009
30 september 2009 kl. 9.00–10.30
Tillsammans med utvecklingsutskottet och underutskottet för mänskliga rättigheter (se särskild föredragningslista)
13.
Redogörelse för nomineringarna till Sacharovpriset 2009
30 september 2009 kl. 10.45–12.45
14.
Diskussion med Javier Solana, EU:s höge representant för den gemensamma utrikes- och säkerhetspolitiken, om prioriteringarna för den gemensamma utrikes- och säkerhetspolitiken
15.
Datum och plats för nästa sammanträde
· Måndagen den 12 oktober 2009 kl. 18.00–19.00 (i Bryssel)
· Torsdagen den 15 oktober 2009 kl. 9.00–10.30 (i Bryssel)
· Tisdagen den 6 oktober 2009 kl. 9.00–12.30 och kl. 15.00–19.00 (i Bryssel)
Föredragningslista
Onsdagen den 21 oktober 2009
9:00 - 11:50 Uttalanden av rådet och kommissionen
Föreberedelser för Europeiska rådet (29-30 oktober 2009)
12:00 - 13:00 Omröstning
Resolutionsförslag
Informationsfrihet i Italien och i andra medlemsstater i Europeiska unionen
15:00 - 18:00 Gemensam debatt
Europeisk avdelning för yttre åtgärder
Betänkande Elmar Brok 19/10
De institutionella aspekterna av inrättandet av den europeiska avdelningen för yttre åtgärder
De institutionella aspekterna av inrättandet av den europeiska avdelningen för yttre åtgärder
[ 2009/2133(INI) ]
Utskottet för konstitutionella frågor
Uttalanden av rådet och kommissionen
Inrättande av en europeisk avdelning för yttre åtgärder: Läget för förhandlingarna med medlemsstaterna
Slut på den gemensamma debatten
Gemensam debatt
Transatlantiska förbindelser
Uttalanden av rådet och kommissionen
Förberedelser för CET-mötet och toppmötet mellan EU och USA (2-3 november 2009)
Uttalanden av rådet och kommissionen
Juridiskt och polisiärt transatlantiskt samarbete
Slut på den gemensamma debatten
18:00 - 19:00 Frågestund med frågor till rådet B7-0212/2009
Talartid ( artikel 149 i arbetsordningen)
9:00 - 11:50 Rådet (inklusive repliker)
Kommissionen (inklusive repliker)
Talarlista Ledamöter
PPE
28,5
S&D
20,5
ALDE
10,5
Verts/ALE
7,5
ECR
7,5
GUE/NGL
5,5
EFD
5
NI
5
"Catch the eye"
15:00 - 18:00 Rådet (inklusive repliker)
Kommissionen (inklusive repliker)
Föredragande
Talarlistor Ledamöter
PPE
23
S&D
17
ALDE
9
Verts/ALE
6
ECR
6
GUE/NGL
5
EFD
5
NI
4
"Catch the eye"
Tidsfrister
Resolutionsförslag
Informationsfrihet i Italien och i andra medlemsstater i Europeiska unionen
Resolutionsförslag
har löpt ut
Ändringsförslag och gemensamma resolutionsförslag
Måndagen den 19 oktober, 21:00
Begäran om särskild omröstning, delad omröstning eller omröstning med namnupprop
Tisdagen den 20 oktober, 19:00
Betänkande Elmar Brok 19/10
De institutionella aspekterna av inrättandet av den europeiska avdelningen för yttre åtgärder
Ändringsförslag
Tisdagen den 20 oktober, 20:00
Begäran om särskild omröstning, delad omröstning eller omröstning med namnupprop
Onsdagen den 21 oktober, 17:00
Uttalanden av rådet och kommissionen
Förberedelser för CET-mötet och toppmötet mellan EU och USA (2-3 november 2009)
Resolutionsförslag
Måndagen den 19 oktober, 19:00
Ändringsförslag och gemensamma resolutionsförslag
Onsdagen den 21 oktober, 10:00
Begäran om särskild omröstning, delad omröstning eller omröstning med namnupprop
Onsdagen den 21 oktober, 17:00
Särskild omröstning - delad omröstning - omröstning med namnupprop Texter som kommer att gå till omröstning tisdag
har löpt ut
Texter som kommer att gå till omröstning onsdag
Måndagen den 19 oktober, 19:00
Texter som kommer att gå till omröstning torsdag
Tisdagen den 20 oktober, 19:00
Resolutionsförslag om debatter om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer ( artikel 122 i arbetsordningen)
Torsdagen den 22 oktober, 10:00
EUROPAPARLAMENTET
2009 - 2014
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
FEMM(2009)1104_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Onsdagen den 4 november 2009, kl. 9.00–12.30 och kl. 15.00–18.30
Bryssel
Lokal: ASP 3G2
4 november 2009 kl. 09.00 – 11.15
1.
Godkännande av föredragningslistan
2.
Justering av protokollen från sammanträdet den
· 29–30 september 2009 PV – PE429.566v03-00
3.
Meddelanden från ordföranden
4.
Diskussion med
Eva Uddén Sonnegård ( statssekreterare, arbetsmarknadsdepartementet), svenska ordförandeskapet
*** Elektronisk omröstning ***
5.
Jämställdhet genom att förena arbete med familjerättigheter och familjeansvar
FEMM/7/00918
AM – PE429.686v01-00 RE – PE428.244v01-00
· Behandling och antagande
· Tidsfrist för ingivande av ändringsförslag: 8 oktober 2009 kl. 12.00
*** Den elektroniska omröstningen avslutas***
6.
Förberedelser inför utfrågningen av nominerade kommissionsledamöter – Ordföranden informerar om de praktiska arrangemangen
FEMM/7/01331
· Behandling och antagande av förslag till frågor (ännu ej bekräftat)
4 november 2009 kl. 11.15 – 12.30
Inom stängda dörrar
7.
Samordnarnas sammanträde
4 november 2009 kl. 15.00 – 18.30
8.
Diskussion med
Vladimír Špidla (kommissionsledamot med ansvar för sysselsättning, sociala frågor och lika möjligheter)
*** Elektronisk omröstning ***
9.
Avskaffande av våld mot kvinnor
FEMM/7/00917
AM – PE430.297v01-00 RE – PE428.239v02-00
· Behandling och antagande
· Tidsfrist för ingivande av ändringsförslag: 12 oktober 2009 kl. 12.00
*** Den elektroniska omröstningen avslutas***
10.
Förebyggande och bekämpning av människohandel samt skydd av offren
FEMM/7/00282
* 2009/0050(CNS) KOM(2009)0136 – C7-0008/2009
Föredragande:
Edit Bauer
Ansv. utsk.:
LIBE –
Anna Hedh
· Behandling och godkännande av två muntliga frågor (ännu ej bekräftat)
· Diskussion
11.
Ordföranden informerar om samordnarnas rekommendationer
12.
Övriga frågor
13.
Datum för nästa sammanträde
· Måndagen den 30 november 2009 kl. 15.00–18.30 (Bryssel)
· Tisdagen den 1 december 2009 kl. 9.00–12.30 (Bryssel)
Föredragningslista
Torsdagen den 12 november 2009
9:00 - 10:50 Betänkande Chrysoula Paliadeli A7-0020/2009
Europeiska ombudsmannens verksamhet (2008)
om årsrapporten om Europeiska ombudsmannens verksamhet 2008
[ 2009/2088(INI) ]
Utskottet för framställningar
I närvaro av Nikiforos Diamandouros
Betänkande Alain Lamassoure A7-0045/2009
Övergångsriktlinjer för budgetförfarandet för att beakta ikraftträdandet av Lissabonfördraget
om övergångsriktlinjer för budgetförfarandet för att beakta ikraftträdandet av Lissabonfördraget
[ 2009/2168(INI) ]
Budgetutskottet
11:00 - 13:00 Omröstning
Betänkande Tanja Fajon A7-0042/2009
Förteckningen över tredjeländer vars medborgare omfattas av eller är undantagna från viseringskrav när de passerar medlemsstaternas yttre gränser
om förslaget till rådets förordning om ändring av rådets förordning (EG) nr 539/2001 om fastställande av förteckningen över tredje länder vars medborgare är skyldiga att inneha visering när de passerar de yttre gränserna och av förteckningen över de tredje länder vars medborgare är undantagna från detta krav
[ KOM(2009)0366 - C7-0112/2009 - 2009/0104(CNS) ]
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Resolutionsförslag
Progress årliga arbetsprogram för 2010 och förteckningen över verksamheter per politikavsnitt
Artikel 88 i arbetsordningen
B7-0135/2009 Resolutionsförslag
Toppmötet mellan EU och Ryssland i Stockholm den 18 november 2009
RC B7-0128/2009 , B7-0128/2009 , B7-0129/2009 , B7-0130/2009 , B7-0131/2009 , B7-0132/2009 , B7-0134/2009 Resolutionsförslag
Gemensam programplanering av forskning för att bekämpa neurodegenerativa sjukdomar
B7-0133/2009 Betänkande Chrysoula Paliadeli A7-0020/2009
Europeiska ombudsmannens verksamhet (2008)
om årsrapporten om Europeiska ombudsmannens verksamhet 2008
[ 2009/2088(INI) ]
Utskottet för framställningar
Betänkande Alain Lamassoure A7-0045/2009
Övergångsriktlinjer för budgetförfarandet för att beakta ikraftträdandet av Lissabonfördraget
om övergångsriktlinjer för budgetförfarandet för att beakta ikraftträdandet av Lissabonfördraget
[ 2009/2168(INI) ]
Budgetutskottet
Talartid ( artikel 149 i arbetsordningen)
9:00 - 10:50 Kommissionen (inklusive repliker)
Ombudsmannen
Föredragande (2 x 6')
Talarlista Ledamöter
PPE
12,5
S&D
9
ALDE
5,5
Verts/ALE
4
ECR
4
GUE/NGL
3,5
EFD
3,5
NI
3
"Catch the eye" (2 x 5')
Tidsfrister
Betänkande Chrysoula Paliadeli A7-0020/2009
Europeiska ombudsmannens verksamhet (2008)
Ändringsförslag
har löpt ut
Betänkande Alain Lamassoure A7-0045/2009
Övergångsriktlinjer för budgetförfarandet för att beakta ikraftträdandet av Lissabonfördraget
Ändringsförslag
har löpt ut
Resolutionsförslag
Progress årliga arbetsprogram för 2010 och förteckningen över verksamheter per politikavsnitt
Ändringsförslag
har löpt ut
Särskild omröstning - delad omröstning - omröstning med namnupprop Texter som kommer att gå till omröstning torsdag
har löpt ut
EUROPAPARLAMENTET
2009 - 2014
Budgetutskottet
BUDG(2009)1116_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Måndagen den 16 november 2009, kl. 15.00–18.30
Bryssel
Lokal: JAN 2Q2
SAMORDNARNAS SAMMANTRÄDE
1.
Godkännande av föredragningslistan
2.
Meddelanden från ordföranden
Punkt 3, 4 och 5 BAKOM STÄNGDA DÖRRAR
BUDGETEN FÖR 2010
3.
Budgeten för 2010: alla avsnitt
BUDG/7/01518
2009/2002(BUD) 11902/2009[01] – C7-0127/2009
Föredragande:
László Surján (PPE) Vladimír Maňka (S&D)
Ansv. utsk.:
BUDG –
· Diskussion
– Resultatet av trepartsmötet den 12 november och förberedelse inför medlingen den 19 november – Ändringsskrivelse nr 2/2009 till det preliminära förslaget till budget för 2010 – Genomförbarhetsskrivelse
4.
Ändring av det interinstitutionella avtalet av den 17 maj 2006 om budgetdisciplin och sund ekonomisk förvaltning när det gäller den fleråriga budgetramen
BUDG/7/01467
2009/2184(ACI) KOM(2009)0600 – C7-0256/2009
Föredragande:
Reimer Böge (PPE)
Ansv. utsk.:
BUDG –
· Diskussion
BUDGETEN FÖR 2009
5.
Ändringsbudget nr 10/2009: minskning av betalningsbemyndigandena, ekonomisk återhämtningsplan för Europa
BUDG/7/01456
2009/2185(BUD)
Föredragande:
Jutta Haug (S&D)
Ansv. utsk.:
BUDG –
· Diskussion
*** Omröstning ***
6.
Inrättande av ett finansieringsinstrument för samarbete med industriländer (ändring av förordning (EG) nr 1934/2006)
BUDG/7/00011
* 2009/0059(CNS) KOM(2009)0197 – C7-0101/2009
Föredragande:
Alain Lamassoure (PPE)
AM – PE430.614v01-00 PA – PE430.373v01-00
Ansv. utsk.:
INTA –
Helmut Scholz (GUE/NGL)
PR – PE428.224v01-00
· Behandling och antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 9 november 2009 kl. 12.00
7.
Europeiska året för volontärarbete (2011)
BUDG/7/00316
* 2009/0072(CNS) KOM(2009)0254 – C7-0054/2009
Föredragande:
Barbara Matera (PPE)
PA – PE430.546v02-00 AM – PE430.598v01-00
Ansv. utsk.:
CULT –
Marco Scurria (PPE)
PR – PE430.366v01-00
· Behandling och antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 6 november 2009 kl. 12.00
BUDGETEN FÖR 2009
8.
2009 års budget: Avsnitt III – Kommissionen Föredragande: Jutta Haug (S&D) – DEC 35, 40, 43, 44, 45, 48, 51 och 52 – Övriga eventuella önskemål om överföringar
9.
FASTIGHETSPOLITIKEN
10.
*** Omröstningen avslutas***
BUDGETEN FÖR 2009
11.
Utnyttjande av Europeiska fonden för justering för globaliseringseffekter: Sverige/Volvo – Österrike/Steiermark - Nederländerna/Heijmans
BUDG/7/01441
2009/2183(BUD) KOM(2009)0602 – C7-0254/2009
Föredragande:
Reimer Böge (PPE)
Ansv. utsk.:
BUDG –
· Presentation av förslaget till betänkande
12.
Budgetprognosvarningar – Diskussion
13.
Övriga frågor
14.
Datum för nästa sammanträde
Tisdagen den 1 december kl. 15.00–18.30 Onsdagen den 2 december kl. 9.00–12.30
-//EP//TEXT TA P7-TA-2009-0094 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2009-0095 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2009-0096 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2009-0097 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2009-0098 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2009-0099 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2009-0100 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2009-0101 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2009-0102 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2009-0103 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2009-0104 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2009-0105 0 DOC XML V0//SV
NÄRVAROLISTA
Följande skrev på:
Abad
Áder
Agnew
Albertini
Albrecht
Alfonsi
Allam
Alvarez
Alvaro
Alves
Andreasen
Andrés Barea
Andrikienė
Aggourakis
Antinoro
Antonescu
Antoniozzi
Arias Echeverría
Arif
Arlacchi
Ashworth
Atkins
Attard-Montalto
Audy
Ayala Sender
Aylward
Ayuso
Bach
Badia i Cutchet
Balčytis
Balczó
Baldassarre
Balz
Balzani
Barnier
Băsescu
Bastos
Baudis
Bauer
Bearder
Béchu
Belder
Belet
Benarab-Attou
Bendtsen
Bennahmias
Berès
Berlato
Berlinguer
Besset
Bielan
Bilbao Barandica
Bisky
Bizzotto
Blinkevičiūtė
Bloom
Bodu
Böge
Bokros
Bonsignore
Bontes
Borghezio
Borsellino
Borys
Boştinaru
Bowles
Bozkurt
Bradbourn
Brantner
Brepoels
Březina
Briard Auconie
Brok
Brons
Brzobohatá
Bufton
Bullmann
Buşoi
Busuttil
Bütikofer
Buzek
Cabrnoch
Cadec
Callanan
van de Camp
Cancian
Canfin
Capoulas Santos
Caronna
Casa
Cashman
Casini
Caspary
Castex
del Castillo Vera
Cavada
Cercas
Češková
Chatzimarkakis
Chichester
Chountis
Christensen
Claeys
Clark
Coelho
Cofferati
Cohn-Bendit
Collino
Colman
Comi
Corazza Bildt
Cornelissen
Correia De Campos
Cortés Lastra
Silvia Costa
Cozzolino
Cramer
Creţu
Creutzmann
Crocetta
Crowley
Cutaş
Cymański
Czarnecki
Daerden
van Dalen
Dăncilă
Danellis
Danjean
Dantin
(The Earl of) Dartmouth
Dati
Daul
David
Davies
De Angelis
Dehaene
Delli
Delvaux
de Magistris
De Mita
De Rossa
De Sarnez
Désir
Deß
Deva
De Veyrac
Díaz de Mera García Consuegra
Dodds
Domenici
Dorfmann
Duff
Durant
Dušek
Ehrenhauser
El Khadraoui
Elles
Enciu
Engel
Engström
Eppink
Ernst
Ertug
Essayah
Estaràs Ferragut
Evans
Fajmon
Fajon
Falbr
Färm
Feio
Ferber
Fernandes
Elisa Ferreira
Fidanza
Figueiredo
Fjellner
Flašíková Beňová
Flautre
Fleckenstein
Fontana
Ford
Foster
Fox
Fraga Estévez
Franco
Gahler
Gál
Gallagher
Gallo
García Pérez
Gardiazábal Rubial
Garriga Polledo
Gauzès
Gebhardt
Geier
Gerbrandy
Geringer de Oedenberg
Giannakou
Giegold
Gierek
Girling
Glattfelder
Godmanis
Goerens
Gollnisch
Gomes
Göncz
Goulard
de Grandes Pascual
Gräßle
Grech
Grelier
Greze
Griesbeck
Gróbarczyk
Grosch
Grossetête
Gruny
Grzyb
Gualtieri
Guerrero Salom
Guillaume
Gurmai
Gutiérrez-Cortines
Győri
Hadjigeorgiou
Haglund
Hall
Händel
Handzlik
Hankiss
Harbour
Harkin
Haug
Häusling
Hautala
Havel
Hedh
Hénin
Hennis-Plasschaert
Herczog
Herranz García
Hibner
Jim Higgins
Joe Higgins
Hoang Ngoc
Hohlmeier
Hökmark
Honeyball
Howitt
Danuta Maria Hübner
Hudghton
Hughes
Hyusmenova
Iacolino
Ibrisagic
Ilchev
Imbrasas
in 't Veld
Iotova
Itälä
Iturgaiz Angulo
Ivan
Ivanova
Jaakonsaari
Jahr
Járóka
Jáuregui Atondo
Jazłowiecka
Jędrzejewska
Jeggle
Jensen
Jiménez-Becerril Barrio
Joly
de Jong
Juvin
Kacin
Kaczmarek
Kadenbach
Kalfin
Kalinowski
Kalniete
Kamall
Kamiński
Kammerevert
Karas
Karim
Kariņš
Kasoulides
Kastler
Kazak
Tunne Kelam
Keller
Alan Kelly
Seán Kelly
Kiil-Nielsen
Kirilov
Klaß
Klinz
Klute
Koch
Koch-Mehrin
Kohlíček
Kolarska-Bobińska
Koppa
Korhola
Kósa
Köstinger
Koumoutsakos
Kovatchev
Kozlík
Kožušník
Krahmer
Kratsa-Tsagaropoulou
Krehl
Kreissl-Dörfler
Kuhn
Kukan
Kurski
Lamassoure
Lambert
Lamberts
Lambrinidis
Landsbergis
Lange
de Lange
Langen
La Via
Lechner
Le Foll
Legutko
Lehne
Le Hyaric
Leichtfried
Jean-Marie Le Pen
Marine Le Pen
Lewandowski
Liberadzki
Lichtenberger
Liese
Liotard
Lisek
Lochbihler
Lövin
Løkkegaard
Lope Fontagné
López Aguilar
López-Istúriz White
Lösing
Lucas
Ludford
Ludvigsson
Luhan
Łukacijewska
Lulling
Lunacek
Lynne
Lyon
McCarthy
Mcclarkin
McGuinness
McMillan-Scott
Madlener
Manders
Mănescu
Maňka
Mann
Marcinkiewicz
Marinescu
David Martin
Hans-Peter Martin
Martínez Martínez
Masip Hidalgo
Maštálka
Mastella
Mathieu
Mato Adrover
Matula
Mauro
Mavronikolas
Mayer
Mayor Oreja
Mazzoni
Meissner
Mélenchon
Melo
Méndez de Vigo
Menéndez del Valle
Messerschmidt
Mészáros
Meyer
Louis Michel
Migalski
Mikolášik
Milana
Millán Mon
Mirsky
Mitchell
Mölzer
Moraes
Moreira
Morganti
Morin-Chartier
Morkūnaitė
Motti
Muñiz De Urquiza
Muscardini
Nattrass
Nedelcheva
Neuser
Neveďalová
Newton Dunn
Mihaylova
Neyts-Uyttebroeck
Nicholson
Nicolai
Niebler
van Nistelrooij
Nuttall
Obiols
Ojuland
Olbrycht
Olejniczak
Oomen-Ruijten
Őry
Oviir
Pack
Padar
Paksas
Paleckis
Paliadeli
Pallone
Panayotov
Panzeri
Papadopoulou
Papanikolaou
Papastamkos
Parvanova
Paşcu
Paška
Patrão Neves
Patriciello
Paulsen
Peillon
Alojz Peterle
Pieper
Pietikäinen
Piotrowski
Pirillo
Pittella
Plumb
Poc
Ponga
Poręba
Portas
Posselt
Pöttering
Poupakis
Preda
Protasiewicz
Provera
Quisthoudt-Rowohl
Rangel
Ransdorf
Rapkay
Rapti
Regner
Reimers
Remek
Reul
Riera Madurell
Ries
Rinaldi
Rivasi
Rivellini
Rochefort
Rodust
Rohde
Roithová
Romero López
Romeva i Rueda
Rossi
Roth-Behrendt
Rouček
Rübig
Rubiks
Rühle
Saïfi
Salatto
Salavrakos
Salvini
Sanchez-Schmid
Sánchez Presedo
Sârbu
Sargentini
Sartori
Saryusz-Wolski
Sassoli
Saudargas
Savisaar
Schaake
Schaldemose
Schlyter
Olle Schmidt
Schmitt
Schnellhardt
Schnieber-Jastram
Scholz
Schöpflin
Schroedter
Martin Schulz
Werner Schulz
Schwab
Scicluna
Scotta'
Scurria
Seeber
Sehnalová
Senyszyn
Serracchiani
Severin
Siekierski
Silvestris
Simon
Simpson
Sinclaire
Sippel
Siwiec
Skrzydlewska
Smith
Smolková
Sógor
Soini
Sommer
Søndergaard
Sonik
Sosa Wagner
Speroni
Staes
Stassen
Šťastný
Stavrakakis
Steinruck
Sterckx
Stevenson
Stihler
van der Stoep
Stolojan
Dimitar Stoyanov
Strejček
Striffler
Sturdy
Surján
Susta
Alf Svensson
Eva-Britt Svensson
Swinburne
Swoboda
Szájer
Szegedi
Szymański
Tabajdi
Takkula
Tănăsescu
Tannock
Tarabella
Tarand
Tatarella
Tavares
Teixeira
Thaler
Thein
Theocharous
Theurer
Thomsen
Thun Und Hohenstein
Thyssen
Ţicău
Tirolien
Toia
Tomaševski
Tošenovský
Toussas
Trautmann
Tremopoulos
Tremosa I Balcells
Triantaphyllides
Trüpel
Trzaskowski
Tsoukalas
Turunen
Tzavela
Uggias
Ulmer
Uspaskich
Vaidere
Vajgl
Van Brempt
Vanhecke
Van Orden
Vattimo
Vaughan
Vergiat
Vergnaud
Verheyen
Vidal-Quadras
Vigenin
Vlasák
Vlasto
Voss
Jarosław Leszek Wałęsa
Wallis
Manfred Weber
Renate Weber
Weiler
Weisgerber
Werthmann
Westlund
Westphal
Wikström
Willmott
Wils
Hermann Winkler
Iuliu Winkler
Włosowicz
Wojciechowski
Wortmann-Kool
Yáñez-Barnuevo García
Yannakoudakis
Záborská
Zahradil
Zalba Bidegain
Zalewski
Zasada
Ždanoka
Zemke
Zīle
Zimmer
Ziobro
Milan Zver
Zwiefka
NÄRVAROLISTA
Följande skrev på:
Abad
Áder
Agnew
Albertini
Albrecht
Alfano
Alfonsi
Alvarez
Alves
Andreasen
Andrikienė
Angelilli
Angourakis
Antinoro
Antonescu
Antoniozzi
Arias Echeverría
Arif
Arsenis
Ashworth
Atkins
Audy
Auken
Ayala Sender
Aylward
Ayuso
van Baalen
Bach
Badia i Cutchet
Balčytis
Balczó
Baldassarre
Balz
Balzani
Bartolozzi
Băsescu
Bastos
Batten
Baudis
Bauer
Bearder
Becali
Béchu
Belder
Belet
Bélier
Benarab-Attou
Bendtsen
Bennahmias
Berès
Berlato
Berlinguer
Berman
Besset
Bielan
Bilbao Barandica
Binev
Bisky
Bizzotto
Blinkevičiūtė
Bloom
Bodu
Böge
Bokros
Bonsignore
Bontes
Borghezio
Borsellino
Borys
Boştinaru
Bové
Bowles
Bozkurt
Bradbourn
Brantner
Brepoels
Březina
Briard Auconie
Brok
Brons
Brzobohatá
Bufton
Bullmann
Busuttil
Bütikofer
Buzek
Cabrnoch
Cadec
Callanan
van de Camp
Campbell Bannerman
Cancian
Canfin
Capoulas Santos
Caronna
Carvalho
Casa
Cashman
Casini
Caspary
Castex
del Castillo Vera
Cavada
Cercas
Češková
Chatzimarkakis
Chichester
Childers
Chountis
Christensen
Claeys
Clark
Coelho
Cohn-Bendit
Collino
Colman
Comi
Cornelissen
Correia De Campos
Cortés Lastra
Silvia Costa
Cozzolino
Cramer
Creţu
Creutzmann
Crocetta
Cutaş
Cymański
Czarnecki
Daerden
van Dalen
Dăncilă
Danellis
Danjean
Dantin
(The Earl of) Dartmouth
Dati
Daul
David
De Angelis
de Brún
De Castro
Dehaene
De Keyser
Delli
Delvaux
de Magistris
De Mita
De Rossa
De Sarnez
Désir
Deß
Deutsch
Deva
De Veyrac
Díaz de Mera García Consuegra
Dodds
Domenici
Donskis
Dorfmann
Duff
Durant
Dušek
Ehler
Ehrenhauser
Eickhout
Ek
El Khadraoui
Elles
Enciu
Engel
Engström
Eppink
Ernst
Ertug
Essayah
Estaràs Ferragut
Estrela
Evans
Fajmon
Fajon
Falbr
Farage
Färm
Feio
Ferber
Fernandes
Elisa Ferreira
João Ferreira
Fidanza
Figueiredo
Fisas Ayxela
Fjellner
Flašíková Beňová
Flautre
Fleckenstein
Florenz
Fontana
Ford
Foster
Fox
Fraga Estévez
Franco
Gahler
Gál
Gallagher
Gallo
García-Margallo y Marfil
García Pérez
Gardiazábal Rubial
Gardini
Garriga Polledo
Gauzès
Gebhardt
Geier
Gerbrandy
Geringer de Oedenberg
Giannakou
Giegold
Gierek
Girling
Glante
Glattfelder
Godmanis
Goebbels
Goerens
Gollnisch
Gomes
Göncz
Goulard
de Grandes Pascual
Gräßle
Grech
Grelier
Greze
Griesbeck
Griffin
Gróbarczyk
Groote
Grosch
Grossetête
Gruny
Grzyb
Gualtieri
Guerrero Salom
Guillaume
Gurmai
Gutiérrez-Cortines
Győri
Gyürk
Hadjigeorgiou
Häfner
Haglund
Hall
Händel
Handzlik
Hannan
Harbour
Harkin
Hassi
Haug
Häusling
Hautala
Jiří Havel
Hedh
Helmer
Hénin
Hennis-Plasschaert
Herczog
Herranz García
Hibner
Jim Higgins
Joe Higgins
Nadja Hirsch
Hoang Ngoc
Hohlmeier
Hökmark
Honeyball
Howitt
Danuta Maria Hübner
Hudghton
Hughes
Hyusmenova
Iacolino
Ilchev
Imbrasas
in 't Veld
Iotova
Iovine
Itälä
Iturgaiz Angulo
Ivan
Ivanova
Jaakonsaari
Jäätteenmäki
Jadot
Jahr
Járóka
Jáuregui Atondo
Jazłowiecka
Jędrzejewska
Jeggle
Jensen
Jiménez-Becerril Barrio
Joly
de Jong
Jordan Cizelj
Jørgensen
Junqueras Vies
Juvin
Kacin
Kaczmarek
Kadenbach
Kalfin
Kalinowski
Kalniete
Kamall
Kammerevert
Karas
Kariņš
Kasoulides
Kastler
Kazak
Tunne Kelam
Keller
Alan Kelly
Seán Kelly
Kiil-Nielsen
Kirilov
Kirkhope
Klaß
Klinz
Klute
Koch
Koch-Mehrin
Kohlíček
Kolarska-Bobińska
Koppa
Korhola
Kósa
Köstinger
Koumoutsakos
Kovatchev
Kowal
Kozlík
Kožušník
Krahmer
Kratsa-Tsagaropoulou
Krehl
Kreissl-Dörfler
Kuhn
Kukan
Kurski
Lamassoure
Lambert
Lamberts
Lambrinidis
Lambsdorff
Landsbergis
Lange
de Lange
Langen
La Via
Lechner
Le Foll
Legutko
Lehne
Le Hyaric
Leichtfried
Leinen
Lepage
Jean-Marie Le Pen
Marine Le Pen
Lewandowski
Liberadzki
Lichtenberger
Liese
Liotard
Lisek
Lochbihler
Lövin
Løkkegaard
Lope Fontagné
López Aguilar
López-Istúriz White
Lösing
Lucas
Ludford
Ludvigsson
Luhan
Łukacijewska
Lulling
Lunacek
Lynne
Lyon
McAvan
McCarthy
McClarkin
McGuinness
McMillan-Scott
Macovei
Madlener
Manders
Mănescu
Maňka
Mann
Marcinkiewicz
Marinescu
David Martin
Hans-Peter Martin
Martínez Martínez
Masip Hidalgo
Maštálka
Mastella
Matera
Mathieu
Matias
Mato Adrover
Matula
Mauro
Mayer
Mayor Oreja
Mazzoni
Meissner
Mélenchon
Melo
Méndez de Vigo
Menéndez del Valle
Merkies
Messerschmidt
Mészáros
Meyer
Louis Michel
Migalski
Mikolášik
Milana
Millán Mon
Mirsky
Mitchell
Mölzer
Moraes
Moreira
Morganti
Morin-Chartier
Morkūnaitė-Mikulėnienė
Morvai
Muñiz De Urquiza
Muscardini
Nattrass
Nedelcheva
Neuser
Neveďalová
Newton Dunn
Neynsky
Neyts-Uyttebroeck
Nicholson
Nicolai
Niculescu
Niebler
van Nistelrooij
Nuttall
Obermayr
Obiols
Ojuland
Olbrycht
Olejniczak
Oomen-Ruijten
Őry
Ouzký
Oviir
Pack
Padar
Paksas
Paleckis
Paliadeli
Pallone
Panayotov
Panzeri
Papadopoulou
Papanikolaou
Papastamkos
Pargneaux
Parvanova
Paşcu
Paška
Patrão Neves
Patriciello
Paulsen
Peillon
Perello Rodriguez
Alojz Peterle
Pieper
Pietikäinen
Piotrowski
Pirillo
Pittella
Poc
Podimata
Ponga
Poręba
Portas
Posselt
Pöttering
Poupakis
Preda
Vittorio Prodi
Protasiewicz
Provera
Rangel
Ranner
Ransdorf
Rapkay
Rapti
Regner
Reimers
Remek
Reul
Riera Madurell
Ries
Rinaldi
Riquet
Rivasi
Rivellini
Rochefort
Rodust
Rohde
Roithová
Romero López
Romeva i Rueda
Ronzulli
Rosbach
Rossi
Roth-Behrendt
Rouček
Rübig
Rubiks
Saïfi
Salafranca Sánchez-Neyra
Salatto
Salavrakos
Salvini
Sanchez-Schmid
Sánchez Presedo
Sârbu
Sargentini
Sartori
Saryusz-Wolski
Sassoli
Saudargas
Savisaar
Schaake
Schaldemose
Schlyter
Olle Schmidt
Schnellhardt
Schnieber-Jastram
Scholz
Schöpflin
Schroedter
Martin Schulz
Werner Schulz
Schwab
Scicluna
Scotta'
Scurria
Seeber
Sehnalová
Senyszyn
Serracchiani
Severin
Siekierski
Silvestris
Simon
Simpson
Sinclaire
Sippel
Siwiec
Skinner
Skrzydlewska
Skylakakis
Smolková
Sógor
Soini
Sommer
Søndergaard
Sonik
Sosa Wagner
Soullie
Speroni
Staes
Stassen
Šťastný
Stavrakakis
Steinruck
Sterckx
Stevenson
Stihler
van der Stoep
Stolojan
Emil Stoyanov
Strasser
Strejček
Striffler
Sturdy
Surján
Susta
Alf Svensson
Eva-Britt Svensson
Swinburne
Swoboda
Szájer
Szegedi
Szymański
Tabajdi
Takkula
Tănăsescu
Tannock
Tarabella
Tarand
Tavares
Teixeira
Thaler
Thein
Theocharous
Theurer
Thomsen
Thun Und Hohenstein
Thyssen
Ţicău
Toia
Tőkés
Tomaševski
Tošenovský
Toussas
Trautmann
Tremopoulos
Tremosa i Balcells
Triantaphyllides
Trüpel
Trzaskowski
Tsoukalas
Turmes
Turunen
Tzavela
Uggias
Ulmer
Ulvskog
Ungureanu
Urutchev
Uspaskich
Vajgl
Vălean
Van Brempt
Vanhecke
Van Orden
Vattimo
Vaughan
Vergiat
Vergnaud
Verheyen
Vidal-Quadras
Vigenin
de Villiers
Vlasák
Vlasto
Voss
Jarosław Leszek Wałęsa
Wallis
Watson
Henri Weber
Manfred Weber
Renate Weber
Weiler
Weisgerber
Werthmann
Westlund
Westphal
Wieland
Wikström
Willmott
Wils
Hermann Winkler
Iuliu Winkler
Włosowicz
Wojciechowski
Wortmann-Kool
Yáñez-Barnuevo García
Yannakoudakis
Záborská
Zahradil
Zala
Zalewski
Zanicchi
Zasada
Ždanoka
Zeller
Zemke
Zīle
Zimmer
Ziobro
Milan Zver
Zwiefka
EU-korrespondenter: det går åt många skor att bevaka Bryssel
Kultur
2010-03-05 - 09:56
Europaparlamentets journalistpris finns i fyra kategorier: press, radio, TV och Internet Den 31 mars är sista datum för tävlingsbidrag till Europaparlamentets journalistpris.
Men hur är det att jobba som journalist i den stora apparat som stavas parlamentet?
Vi frågade några av de fler än tusen ackrediterade reportrar som har satts att bevaka Bryssel.
"Mängden information från de olika institutionerna är överväldigande", säger Maria Laura Franciosi, före detta byråchef på nyhetsbyrån Ansa.
"Att jobba här handlar om att röra sig mellan många olika institutioner, slita ut många skor, ha örat mot otaliga informationskällor - och att sedan i slutändan sitta ner och försöka gör allt begripligt för läsaren."
"Vi har ett på många sätt privilegierat jobb", säger Ann Cahill, korrespondent för Irish Examiner.
"Vi får möjlighet att följa en idé från att den föds och se hur den jobbar sig upp genom regering, näringsliv, samhälle och EU-institutionerna."
"EU-nyheter säljer ju inte direkt som smör i solsken", säger Mikael Stabenow på en av Tysklands ledande dagstidningar, Frankfurter Allgemeine Zeitung.
"Det svåra är att förmedla nyheterna till allmänheten så att de förstår att det som händer är relevant även för dem - även om de inte kan någonting om EU", säger Anna Cahill.
"Man knyter an för dåligt till vanligt folk: det är det som saknas i Europa", säger Maria Laura Franciosi.
"Det spelar ingen roll hur väl man bevakar aktiviteterna i EU-institutionerna om du inte kan förklara för folk hur besluten här påverkar även deras liv."
20100226STO69653 Europaparlamentets journalistpris
SV
1
PHOTO
20100303PHT69895.jpg
SV
2
LINK
http://www.eppj.eu/view/sv/introduction.html
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
EUROPAPARLAMENTET
2009 - 2014
Utskottet för rättsliga frågor
JURI(2010)0308_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Extra sammanträde
Måndagen den 8 mars 2010 kl. 19.00–20.30
Strasbourg
Lokal: SDM S5
I närvaro av rådet och kommissionen
8 mars 2010 kl. 19.00–20.30
1.
Godkännande av föredragningslistan
2.
Meddelanden från ordföranden
3.
Justering av protokollen från sammanträdena den
· 18 januari 2010 PV – PE439.080v01-00
· 27–28 januari 2010 PV – PE438.502v01-00
4.
Europeiska avdelningen för yttre åtgärder: förordning om ändring av anställningsvillkoren för övriga anställda i Europeiska gemenskaperna
JURI/7/02214
Föredragande:
Bernhard Rapkay (S&D)
· Diskussion
5.
Befogenhet att delegera lagstiftning
JURI/7/02156
2010/2021(INI)
Föredragande:
József Szájer (PPE)
PR – PE439.171v01-00
Ansv. utsk.:
JURI –
Rådg. utsk.:
ENVI –
Jo Leinen (S&D)
PA – PE439.162v01-00 AM – PE439.269v01-00
· Behandling av förslag till betänkande
6.
Förvaltning av alternativa investeringsfonder
JURI/7/00301
***I 2009/0064(COD) KOM(2009)0207 – C7-0040/2009
Föredragande:
Evelyn Regner (S&D)
PA – PE438.149v01-00 AM – PE439.261v01-00
Ansv. utsk.:
ECON* –
Jean-Paul Gauzès (PPE)
PR – PE430.709v01-00 AM – PE439.111v02-00 AM – PE438.497v01-00 AM – PE439.125v01-00 AM – PE439.132v01-00 AM – PE439.135v01-00 AM – PE439.134v01-00 AM – PE439.133v01-00 DT – PE428.292v01-00
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 23 februari 2010 kl. 12.00
*** Omröstning ***
7.
Gemensamt system för mervärdesskatt, när det gäller regler om fakturering
JURI/7/00235
* 2009/0009(CNS) KOM(2009)0021 – C6-0078/2009
Föredragande:
Alexandra Thein (ALDE)
PA – PE438.143v01-00 AM – PE438.508v01-00
Ansv. utsk.:
ECON –
David Casa (PPE)
PR – PE430.975v01-00 AM – PE438.381v01-00
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 5 februari 2010 kl. 12.00
8.
Värdepapper som erbjuds till allmänheten och harmonisering av insynskraven (ändring av direktiven 2003/71/EG och 2004/109/EG)
JURI/7/01051
***I 2009/0132(COD) KOM(2009)0491 – C7-0170/2009
Föredragande:
Sebastian Valentin Bodu (PPE)
PA – PE438.405v01-00
Ansv. utsk.:
ECON –
Wolf Klinz (ALDE)
PR – PE431.183v01-00
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 19 februari 2010 kl. 12.00
9.
Betänkande om kommissionens vitbok ”Anpassning till klimatförändring: en europeisk handlingsram”
JURI/7/01305
2009/2152(INI) KOM(2009)0147
Föredragande:
Eva Lichtenberger (Verts/ALE)
PA – PE438.387v01-00 AM – PE439.160v01-00
Ansv. utsk.:
ENVI –
Vittorio Prodi (S&D)
PR – PE430.965v01-00 AM – PE439.124v01-00 AM – PE439.169v01-00
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 17 februari 2010 kl. 12.00
RÄTTSLIG GRUND
10.
Rörlighet för personer med visering för längre vistelse
JURI/7/02241
***I 2009/0028(COD) KOM(2009)0091 – C6-0076/2009
Föredragande:
Kurt Lechner (PPE)
Ansv. utsk.:
LIBE –
Carlos Coelho (PPE)
RR – PE430.461v03-00
· Prövning av den rättsliga grunden
+ Viseringar för längre vistelse och registrering på spärrlista i Schengens informationssystem – 2009/0025(CNS)
*** Omröstningen avslutas ***
Gemensam debatt (punkterna 11 till 15)
11.
Europeiska bankmyndigheten
JURI/7/01058
***I 2009/0142(COD) KOM(2009)0501 – C7-0169/2009
Föredragande:
Klaus-Heiner Lehne (PPE)
PA – PE438.267v01-00
Ansv. utsk.:
ECON –
José Manuel García-Margallo Y Marfil (PPE)
PR – PE438.408v01-00 DT – PE430.734v03-00
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 1 mars 2010 kl. 12.00
12.
Makroprudentiell tillsyn över det finansiella systemet på gemenskapsnivå och inrättande av ett europeiskt systemriskråd
JURI/7/01064
***I 2009/0140(COD) KOM(2009)0499 – C7-0166/2009
Föredragande:
Evelyn Regner (S&D)
PA – PE438.153v01-00
Ansv. utsk.:
ECON –
Sylvie Goulard (ALDE)
PR – PE438.496v01-00
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 1 mars 2010 kl. 12.00
13.
En europeisk värdepappers- och marknadsmyndighet
JURI/7/01069
***I 2009/0144(COD) KOM(2009)0503 – C7-0167/2009
Föredragande:
Raffaele Baldassarre (PPE)
PA – PE430.969v01-00
Ansv. utsk.:
ECON –
Sven Giegold (Verts/ALE)
PR – PE438.409v01-00
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 1 mars 2010 kl. 12.00
14.
En europeisk försäkrings- och tjänstepensionsmyndighet
JURI/7/01074
***I 2009/0143(COD) KOM(2009)0502 – C7-0168/2009
Föredragande:
Françoise Castex (S&D)
PA – PE438.266v02-00
Ansv. utsk.:
ECON –
Peter Skinner (S&D)
PR – PE438.410v01-00
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 1 mars 2010 kl. 12.00
15.
Befogenheterna för Europeiska bankmyndigheten, Europeiska försäkrings- och tjänstepensionsmyndigheten och Europeiska värdepappers- och marknadsmyndigheten (ändring av direktiv 1998/26/EG, 2002/87/EG, 2003/6/EG, 2003/41/EG, 2003/71/EG, 2004/39/EG, 2004/109/EG, 2005/60/EG, 2006/48/EG, 2006/49/EG och 2009/65/EG)
JURI/7/01475
***I 2009/0161(COD) KOM(2009)0576 – C7-0251/2009
Föredragande:
Sajjad Karim (ECR)
PA – PE438.379v01-00
Ansv. utsk.:
ECON –
Antolín Sánchez Presedo (S&D)
PR – PE439.086v02-00
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 1 mars 2010 kl. 12.00
Inom stängda dörrar
16.
Mål som berör parlamentet
17.
Valprövning
18.
Övriga frågor
19.
Datum för nästa sammanträde
· 22 mars 2010 kl. 15.00–18.30 (Bryssel)
· 23 mars 2010 kl. 9.00–18.30 (Bryssel)
Samordnarnas sammanträde
EUROPAPARLAMENTET
2009 - 2014
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
FEMM(2010)0419
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Måndagen den 19 april 2010, kl. 21.00–22.30
Strasbourg
Lokal: SDM-S1
1.
Godkännande av föredragningslistan
2.
Meddelanden från ordföranden
3.
Diskussion
Viviane Reding (kommissionens vice ordförande)
4.
Övriga frågor
5.
Datum för nästa sammanträde
• 3 maj 2010 kl. 15.00–18.30
• 4 maj 2010 kl. 9.00–12.30
EUROPAPARLAMENTET
2009 - 2014
Budgetutskottet
BUDG(2010)0421_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Extra sammanträde
Onsdagen den 21 april 2010 kl. 14.00–15.30
Strasbourg
Lokal: LOW N1.3
1.
Godkännande av föredragningslistan
2.
Meddelanden från ordföranden
BUDGETEN FÖR 2010
3.
Ändringsbudget nr 1/2010: Avsnitt I – Parlamentet
BUDG/7/02585
2010/2045(BUD)
Föredragande:
Vladimír Maňka (S&D)
Ansv. utsk.:
BUDG –
· Diskussion
4.
Ändringsbudget nr 2/2010: Avsnitt III – Kommissionen, Avsnitt VI - Europeiska ekonomiska och sociala kommittén, Avsnitt VII – Regionkommittén
BUDG/7/02584
2010/2046(BUD)
Ansv. utsk.:
BUDG –
· Diskussion
5.
Ändringsbudget nr 3/2010: Avsnitt III – Kommissionen – Kompletterande åtgärder för banansektorn
BUDG/7/02663
2010/2048(BUD)
Föredragande:
László Surján (PPE)
Ansv. utsk.:
BUDG –
· Diskussion
6.
Ändringsbudget nr 4/2010 – Överskottet för 2009 Föredragande: László Surján (PPE) Ansv. utsk.: BUDG – – Diskussion
7.
Den fleråriga budgetramen – det interinstitutionella avtalet: Muntlig fråga och resolutionsförslag – Föredragande: Reimer Böge Antagande (eventuellt)
8.
Beräkningen av inkomster och utgifter för 2011 – Avsnitt I – Parlamentet
BUDG/7/01997
2010/2005(BUD)
Föredragande:
Helga Trüpel (Verts/ALE)
PR – PE439.956v01-00
Ansv. utsk.:
BUDG –
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 15 april 2010 kl. 15.00
9.
Övriga frågor
10.
Datum för nästa sammanträde
· 27 april 2010 kl. 9.00 – 12.30 (Bryssel)
· 27 april 2010 kl. 9.00 – 12.30 och 12.30 – 13.30 (Bryssel)
· 28 april 2010 kl. 9.00 – 12.30 (Bryssel)
Folkhälsoutskottet tar upp kampen mot förfalskade läkemedel
Folkhälsa
2010-05-03 - 19:26
Ledamöterna i parlamentets hälsoutskott har röstat om nya regler för handeln med läkemedel.
Syftet är att ta itu med problemet med förfalskade läkemedel - även på internet.
I november och december 2008 beslagtog tulltjänstemän runtom i EU över 34 miljoner illegala piller.
Förfalskade läkemedel är en lukrativ handel: höga vinstmarginaler, låg risk och dessutom saknas tillräcklig reglering på EU-nivå.
Kontrollera internetförsäljningen
Den 27 april röstade utskottet för folkhälsa om kommissionens förslag till regler för handeln med läkemedel.
En stor del av läkemedelsförsäljningen sker på internet.
En försäljning som är legaliserad i en del medlemsländer.
Jag tror att förfalskare idag uppmuntras av att det saknas regler.
Förfalskade läkemedel är "tysta mördare" eftersom de allvarligt kan skada patienterna.
Tillräckligt ambitiöst?
Franska ledamoten Françoise Grossetête från EPP-gruppen var osäker på om resultaten är så utomordentliga:
– Jag beklagar att reglerna inte är lika hårda för läkemedel som för livsmedel.
Exempelvis tillåter vi ompaketering av läkemedel, men det går inte att paketera om ett pastapaket.
Tyska socialdemokratiska ledamoten Dagmar Roth-Behrendt (S&D) varnar för att stora mängder förfalskade produkter kan komma till EU:
- Det är ett bra resultat men det är inte tillräckligt ambitiöst.
Jag tror att den största delen handlar om kontroll på internet ...
Är vi verkligen villiga att tillämpa reglerna gentemot länder som vi har handelsavtal med, exempelvis Kina?
Betänkandet är en del av kommissionens läkemedelspaketet ("Pharmacy Package").
20100430STO73837 Artikel: Tydligare läkemedelsinformation Utskottet för miljö, folkhälsa och livsmedelssäkerhet Pressemeddelande: Fake medicines: MEPs want to target online sales Följ ärendet
SV
1
EUROPARL-TV
-//EP//TEXT IM-PRESS 20100305STO70032 0 NOT XML V0//SV
-//EP//TEXT IM-PRESS 20100426IPR73469 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Utskottet för utrikesfrågor
AFET(2010)0622_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Tisdagen den 22 juni 2010 kl. 9.00–12.30 och kl. 15.00–18.30
Onsdagen den 23 juni 2010 kl. 9.00–12.30
Bryssel
Lokal: PHS 3 C 50
22 juni 2010 kl. 9.00–10.45
1.
Godkännande av föredragningslistan
2.
Justering av sammanträdesprotokollen från den
· 27–28 april 2010 PV – PE441.046v01-00
· 17 maj 2010 PV – PE441.219v01-00
3.
Meddelanden från ordföranden
4.
Diskussion med Pieter Feith, EU:s särskilde representant i Kosovo
5.
Förslag till resolution om den europeiska integrationsprocessen för Kosovo
AFET/7/02446
Föredragande:
Ulrike Lunacek (Verts/ALE)
AM – PE441.194v02-00 RE – PE440.996v01-00
· Behandling av utkast till resolutionsförslag
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 18 maj 2010 kl. 18.00
22 juni 2010 kl. 10.45–12.30
6.
Förslag till resolution om Islands ansökan om medlemskap i Europeiska unionen
AFET/7/02372
Föredragande:
Cristian Dan Preda (PPE)
AM – PE441.321v01-00 RE – PE439.374v01-00
· Behandling av utkast till resolutionsförslag
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 3 juni 2010 kl. 18.00
7.
Halvtidsöversikt över de europeiska programmen för satellitnavigering: bedömning av genomförandet, framtida utmaningar och finansieringsutsikter
AFET/7/01771
2009/2226(INI)
Föredragande:
Maria Eleni Koppa (S&D)
PA – PE440.114v01-00 AM – PE441.280v01-00
Ansv. utsk.:
ITRE –
Vladimír Remek (GUE/NGL)
DT – PE439.881v01-00
· Behandling av förslag till yttrande
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 11 maj 2010 kl. 12.00
8.
Partnerskaps- och samarbetsavtal: förhandling och slutande av avtal med Turkmenistan
AFET/7/00040
1998/0031(NLE) 05606/1998 – C4-0371/1998
Föredragande:
Norica Nicolai (ALDE)
Ansv. utsk.:
AFET –
Rådg. utsk.:
INTA – Beslut: inget yttrande
BUDG – Beslut: inget yttrande
· Diskussion
9.
Redogörelse för den gemensamma AFET/DEVE/BUDG-delegationen till Mellanöstern (den 24–28 maj 2010)
22 juni 2010 kl. 15.00–17.00
*** Elektronisk omröstning ***
10.
Medlemsstaternas kontroll av kommissionens utövande av sina genomförandebefogenheter
AFET/7/02481
***I 2010/0051(COD) KOM(2010)0083 – C7-0073/2010
Föredragande:
Gabriele Albertini (PPE)
PA – PE441.196v01-00 AM – PE442.872v01-00
Ansv. utsk.:
JURI –
József Szájer (PPE)
PR – PE441.207v02-00 AM – PE442.936v01-00
· Behandling av förslag till yttrande och ändringsförslag
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 3 juni 2010 kl. 12.00
*** Den elektroniska omröstningen avslutas ***
Tillsammans med underutskottet för säkerhet och försvar
11.
Offentlig utfrågning om “En ny transatlantisk säkerhetsarkitektur?" (se separat program)
22 juni 2010 kl. 17.00–18.30
12.
Europeiska avdelningen för yttre åtgärder
AFET/7/02461
2010/0816(NLE) 08029/2010 – C7-0090/2010
Föredragande:
Elmar Brok (PPE)
Ansv. utsk.:
AFET* –
Rådg. utsk.:
DEVE –
Filip Kaczmarek (PPE)
INTA –
Jan Zahradil (ECR)
AD – PE440.219v03-00 AM – PE441.195v01-00
BUDG –
Roberto Gualtieri (S&D)
CONT –
Ivailo Kalfin (S&D)
PA – PE441.269v01-00 DT – PE441.318v01-00
ENVI – Beslut: inget yttrande
JURI – Beslut: inget yttrande
LIBE –
AFCO* –
Guy Verhofstadt (ALDE)
FEMM –
Franziska Katharina Brantner (Verts/ALE)
PA – PE441.063v01-00 AM – PE442.788v01-00
· Diskussion
23 juni 2010 kl. 9.00–10.00
*** Elektronisk omröstning ***
13.
Förslag till resolution om den europeiska integrationsprocessen för Albanien
AFET/7/02452
Föredragande:
Nikolaos Chountis (GUE/NGL)
AM – PE441.221v01-00 RE – PE440.129v02-00
· Antagande av ett utkast till resolutionsförslag
· Tidsfrist för ingivande av ändringsförslag: 5 maj 2010 kl. 12.00
14.
Förslag till resolution om den europeiska integrationsprocessen för Kosovo
AFET/7/02446
Föredragande:
Ulrike Lunacek (Verts/ALE)
AM – PE441.194v02-00 RE – PE440.996v01-00
· Antagande av ett utkast till resolutionsförslag
· Tidsfrist för ingivande av ändringsförslag: 18 maj 2010 kl. 18.00
15.
Förslag till resolution om Islands ansökan om medlemskap i Europeiska unionen
AFET/7/02372
Föredragande:
Cristian Dan Preda (PPE)
AM – PE441.321v01-00 RE – PE439.374v01-00
· Antagande av ett utkast till resolutionsförslag
· Tidsfrist för ingivande av ändringsförslag: 3 juni 2010 kl. 18.00
16.
Halvtidsöversikt över de europeiska programmen för satellitnavigering: bedömning av genomförandet, framtida utmaningar och finansieringsutsikter
AFET/7/01771
2009/2226(INI)
Föredragande:
Maria Eleni Koppa (S&D)
PA – PE440.114v01-00 AM – PE441.280v01-00
Ansv. utsk.:
ITRE –
Vladimír Remek (GUE/NGL)
DT – PE439.881v01-00
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 11 maj 2010 kl. 12.00
*** Den elektroniska omröstningen avslutas ***
23 juni 2010 kl. 10.00–11.00
Tillsammans med delegationen för förbindelserna med Maghrebländerna och Arabiska Maghrebunionen
17.
Diskussion med kommissionen om ramavtalet mellan EU och Libyen
23 juni 2010 kl. 11.00–12.00
18.
Diskussion om läget i Kirgizistan
23 juni 2010 kl. 12.00–12.30
Inom stängda dörrar
19.
Utvidgat presidium (se separat program)
20.
Övriga frågor
21.
Datum för nästa sammanträde
· 13 juli 2010 kl. 15.00–18.30 (Bryssel)
· 14 juli 2010 kl. 9.00–12.30 och 15.00–18.30 (Bryssel)
Fler rättigheter för båtpassagerare men ännu oklart för bussresenärer
Transporter
Plenarsammanträde
2010-07-06 - 14:47
Båtpassagerare kommer att få fler rättigheter från och med 2012, tack vare en förordning som godkändes av Europaparlamentet på tisdagen.
De nya reglerna möjliggör för stöd och ersättning vid förseningar, samt fri assistans till personer med funktionshinder.
Enligt de nya reglerna får resenärerna rätt till ombokning eller pengarna tillbaka när en passagerarbåt ställs in eller blir försenad med 90 minuter eller mer.
Undantag gäller när förseningen beror på vädret eller andra förhållanden utom operatörens kontroll.
Passagerarna måste också ges mellanmål eller måltider, om det möjligt.
Ersättningen kommer att betalas kontant om resenären kräver det.
Rättigheter för personer med funktionshinder eller nedsatt rörlighet
Av förordningen framgår att funktionshinder inte får användas som ett skäl att neka en passagerare rätt att gå ombord.
Gratis stöd måste ges till funktionshindrade personer i hamnar, under förutsättning att transportören eller hamnoperatören meddelas när bokningen görs eller minst 48 timmar innan avgång.
Detta kommer också att gälla för kryssningspassagerare.
Dessa regler träder i kraft år 2012 och gäller för passagerarfartyg som medför fler än 12 passagerare, med vissa undantag, t.ex. för utflykter och rundturer.
Båtpassagerare kommer därmed att få fler rättigheter än de som nu föreskrivs i EU: s lagstiftning för flygpassagerare, som inte garanteras ersättning för förseningar (endast för inställda flyg).
Bussresor: förhandlingar pågår
Parlamentet har också antagit ändringar av ett förordningsförslag som fastställer busspassagerares rättigheter, som återbetalning av biljettkostnaderna eller ombokning vid förseningar på mer än två timmar samt ersättning på upp till 1800 € för förlorat eller skadat bagage .
I händelse av en passagerares död i en bussolycka bör ersättningsbeloppet inte begränsas alls, tycker ledamöterna.
De krävde också gratis hjälp eller ersättning om ett fel på bussen orsaker försenad ankomst.
Gratis hjälp till passagerare med funktionshinder måste också finnas, säger de.
Parlamentet vill att förordningen gäller inte bara för långa sträckor utan även för regionala bussar.
Eftersom förhandlingarna med rådet inte har lett till någon överenskommelse kommer ärendet sannolikt att gå till förlikning.
20100705IPR77798 Antagna texter (klicka på 6 juli 2010)
SV
1
LINK
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
Polens president besöker Europaparlamentet
Institutioner
2010-09-02 - 10:09
Polens president Bronisław Komorowski och Europaparlamentets talman Jerzy Buzek Polens president Bronislaw Komorowski besökte igår, den 1 september, Europaparlamentet.
Den nyvalde presidenten valde att göra sin första officiella resa till Bryssel - en symbolisk gest för att visa hur viktigt Europa är för Polen.
Han mötte bland andra talmannen, Jerzy Buzek, och diskuterade det polska EU-ordförandeskapet 2011.
Den polske presidenten fick ett varmt och personligt mottagande av Jerzy Buzek, som Komorowski skämtsamt kallade "min gamla chef".
2000-2001 var Komorowski nämligen försvarsminister i Buzeks polska regering.
I mötet kom bland annat prioriteringar för Polens EU-ordförandeskap 2011, Polens strategiska roll i europeisk försvars- och utrikespolitik och den framtida EU-diplomattjänsten upp.
- Jag är glad att den fransk-polsk-tyska stridsgruppen kommer att vara operativ 2013 som ett konkret exempel på europeisk samarbete mellan våra tre länder, sa Bronislaw Komorowski.
Jerzy Buzek sa att han såg fram emot "nya impulser" från 2011 års ordförandeländer Ungern och Polen.
20100831STO80669 Europaparlamentets talman Polens president
SV
1
PHOTO
20100901PHT80866.jpg
SV
2
LINK
/president/view/en/the_president/latest_news.html
SV
3
LINK
http://www.president.pl/en/
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Underutskottet för säkerhet och försvar
SEDE(2010)0927_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Måndagen den 27 september 2010, kl. 16.45–19.00
Bryssel
Lokal: ASP - 1G-2
27 september 2010 kl. 16.45–19.00
1.
Godkännande av föredragningslistan
2.
Meddelanden från ordföranden
3.
Civilt och militärt samarbete, och utvecklingen av civila och militära resurser
AFET/7/02857
2010/2071(INI)
Föredragande:
Christian Ehler (PPE)
PR – PE448.660v01-00
Ansv. utsk.:
AFET –
· Behandling av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 30 september 2010 kl. 12.00
4.
SEDE:s delegation till EU:s övervakningsuppdrag i Georgien (13–16 juli 2010) – Diskussion
5.
Övriga frågor
6.
Datum för nästa sammanträde
· 28 september 2010 kl. 9.00–12.30 och 14.30–18.00 (Bryssel)
(AFET/SEDE interparlamentariskt utskottssammanträde)
* * *
Inom stängda dörrar Det utvidgade presidiet (se separat dagordning)
* * *
Utskottet för kultur och utbildning
CULT(2010)0927_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Måndagen den 27 september 2010, kl. 15.00–17.30 och kl. 17.30–18.30
Tisdagen den 28 september 2010, kl. 9.00–12.30
Bryssel
Lokal: PHS - 5B001
27 september 2010 kl. 15.00–17.30
1.
Godkännande av föredragningslistan
2.
Justering av protokollen från sammanträdena den
· 13–14 juli 2010 PV – PE445.693v01-00
· 2 september 2010 PV – PE445.956v01-00
3.
Meddelanden från ordföranden
I närvaro av rådet och kommissionen
4.
Medborgarinitiativ
CULT/7/02759
***I 2010/0074(COD) KOM(2010)0119 – C7-0089/2010
Föredragande:
Róża Gräfin Von Thun Und Hohenstein (PPE)
PA – PE445.900v01-00
Ansv. utsk.:
AFCO* –
Alain Lamassoure (PPE) Zita Gurmai (S&D)
DT – PE443.095v01-00
· Behandling av förslag till yttrande
· Beslut om tidsfrist för ingivande av ändringsförslag
5.
6.
Diskussion med Gian Francesco Lupattelli (ordförande i ACES Europe)
27 september 2010 kl. 17.30–18.30
Inom stängda dörrar
7.
Samordnarnas sammanträde
* * *
28 september 2010 kl. 9.00–12.30
I närvaro av rådet och kommissionen
*** Omröstning ***
8.
Offentligägd radio och TV i den digitala tidsåldern: framtiden för det dubbla systemet
CULT/7/02205
2010/2028(INI)
Föredragande:
Ivo Belet (PPE)
PR – PE442.905v01-00 AM – PE442.961v01-00 DT – PE441.270v01-00
Ansv. utsk.:
CULT –
· Antagande av förslag till betänkande
9.
Bekämpande av sexuella övergrepp mot barn, sexuell exploatering av barn och barnpornografi (upphävande av rambeslut 2004/68/RIF)
CULT/7/02675
***I 2010/0064(COD) KOM(2010)0094 – C7-0088/2010
Föredragande:
Petra Kammerevert (S&D)
PA – PE442.976v01-00 AM – PE442.977v01-00
Ansv. utsk.:
LIBE –
Roberta Angelilli (PPE)
· Antagande av förslag till yttrande
*** Omröstningen avslutas ***
10.
– Inledande diskussion
11.
Europa, världens främsta resmål – en ny politisk ram för europeisk turism
CULT/7/03813
2010/2206(INI) KOM(2010)0352
Föredragande:
Hella Ranner (PPE)
Ansv. utsk.:
TRAN –
· Inledande diskussion
12.
Redogörelse för en studie om Lissabonfördraget och EU: s idrottspolitik (”The Lisbon Treaty and EU Sports Policy”) av Richard Parrish (professor vid Edge Hill University i Storbritannien) och Borja Garcia (doktor vid University of Loughborough i Storbritannien)
13.
Godkännande av samordnarnas beslut
14.
Övriga frågor
15.
Datum för nästa sammanträde
· 26 oktober 2010 kl. 15.00–17.45 och kl. 17.45–18.30 i Bryssel
· 27 oktober 2010 kl. 9.00–12.30 i Bryssel
Utskottet för jordbruk och landsbygdens utveckling
AGRI(2010)1117_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Onsdagen den 17 november 2010 kl. 13.00–15.00
Bryssel
1.
Godkännande av föredragningslistan
2.
Meddelanden från ordföranden
3.
Kommissionsledamot Dacian Ciolos redogör för meddelandet ”CAP towards 2020: meeting the food, natural resource and territorial challenges of the future”
4.
Övriga frågor
5.
Datum för nästa sammanträde
· 30 november 2010 kl. 15.00–18.30 (Bryssel)
· 1 december 2010 kl. 9.00–18.30 (Bryssel)
PETI Välkomstord
Här finns information om arbetet och aktiviteterna i utskottet, som jag har varit ordförande för sedan 2009.
Att göra framställningar är ett viktigt och ofta effektivt sätt för människor att direkt engagera sig i parlamentets verksamhet och påverka utskottets ledamöter att särskilt koncentrera sig på deras intressefrågor, förslag eller klagomål.
Vårt utskott besvarar ofta framställningar från EU-medborgare genom att försöka lösa kränkningar av medborgarnas rättigheter enligt fördraget, och genom att samarbeta med nationella, regionala och lokala myndigheter i frågor som rör tillämpningen av EU:s lagar inom områden som miljö, sociala frågor, fri rörlighet och så vidare.
Vårt utskott kan även anordna informationsbesök och lägga fram betänkanden i kammaren.
Vi spelar alltså en viktig roll för förbindelserna med EU-medborgarna och för underbyggandet av den demokratiska legitimiteten och ansvarsskyldigheten inom EU:s beslutsprocess.
Erminia Mazzoni
Presentation och befogenheter Utskottet har ansvar för frågor som rör följande områden:
Utskottet för ekonomi och valutafrågor
ECON(2011)0316_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Onsdagen den 16 mars 2011 kl. 9.00–12.30 och kl. 15.00–18.30
Bryssel
Lokal: PHS - 3C050
1.
Godkännande av föredragningslistan
2.
Justering av protokollet från sammanträdena den
· 6 september 2010 PV – PE456.657v01-00
· 13 september 2010 PV – PE452.668v01-00
· 27–28 september 2010 PV – PE456.871v01-00
· 18 oktober 2010 PV – PE456.692v01-00
· 30 november 2010–1 december 2010 PV – PE456.658v01-00
· 13 januari 2011 PV – PE456.993v01-00
· 17 januari 2011 PV – PE458.619v01-00
· 24–25 januari 2011 PV – PE456.994v01-00
· 1 februari 2011 PV – PE456.986v01-00
· 7 februari 2011 PV – PE458.670v01-00
3.
Meddelanden från ordföranden
16 mars 2011 kl. 9.00–10.00
4.
Diskussion med Johnny Åkerholm, ordförande för Europeiska rådgivande organet för statistikstyrning
ECON/7/02197
16 mars 2011 kl. 10.30–12.00
5.
Utnämning av en ledamot av Europeiska centralbankens direktion: Peter Praet (BE)
ECON/7/05430
2011/0802(NLE) 00003/2011 – C7-0058/2011
Föredragande:
Sharon Bowles (ALDE)
PR – PE460.742v01-00
Ansv. utsk.:
ECON –
· Diskussion med Peter Praet, kandidat till posten
16 mars 2011 kl. 12.00–12.20
Inom stängda dörrar
6.
Utnämning av en ledamot av Europeiska centralbankens direktion: Peter Praet (BE)
ECON/7/05430
2011/0802(NLE) 00003/2011 – C7-0058/2011
Föredragande:
Sharon Bowles (ALDE)
PR – PE460.742v01-00
Ansv. utsk.:
ECON –
· Diskussion
16 mars 2011 kl. 12.20–12.30
7.
Yrkesmässiga gränsöverskridande vägtransporter av eurokontanter mellan medlemsstaterna i euroområdet
ECON/7/03539
***I 2010/0204(COD) KOM(2010)0377 – C7-0186/2010
Föredragande:
Sophie Auconie (PPE)
PR – PE454.357v01-00 AM – PE456.920v01-00
Ansv. utsk.:
ECON –
Rådg. utsk.:
EMPL, TRAN
· Behandling av ändringsförslag
16 mars 2011 kl. 15.00–15.15
8.
Politiska alternativ för främjande av en europeisk avtalsrätt för konsumenter och företag
ECON/7/05011
2011/2013(INI) KOM(2010)0348
Föredragande av yttrande:
Sirpa Pietikäinen (PPE)
PA – PE456.822v01-00 AM – PE458.830v01-00
Ansv. utsk.:
JURI* –
Diana Wallis (ALDE)
PR – PE456.886v01-00 AM – PE460.697v01-00
Rådg. utsk.:
ECON, IMCO*
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 18 februari 2011 kl. 12.00
16 mars 2011 kl. 15.15–16.20
9.
System för garanti av insättningar (omarbetning)
ECON/7/03448
***I 2010/0207(COD) KOM(2010)0368 – C7-0177/2010
Föredragande:
Peter Simon (S&D)
PR – PE460.614v01-00
Ansv. utsk.:
ECON –
Rådg. utsk.:
IMCO, JURI, JURI(AL)
· Behandling av förslag till betänkande
16 mars 2011 kl. 16.20–17.10
*** Omröstning ***
10.
Kreditvärderingsinstitut: framtidsperspektiv
ECON/7/04338
2010/2302(INI)
Föredragande:
Wolf Klinz (ALDE)
PR – PE454.361v01-00 AM – PE454.677v01-00
Ansv. utsk.:
ECON –
Rådg. utsk.:
JURI
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 17 januari 2011 kl. 17.00
11.
Företagsstyrning i finansiella institut
ECON/7/04549
2010/2303(INI) KOM(2010)0284
Föredragande:
Ashley Fox (ECR)
PR – PE454.525v03-00 AM – PE456.724v01-00
Ansv. utsk.:
ECON* –
Rådg. utsk.:
DEVE, EMPL, IMCO, JURI*
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 17 januari 2011 kl. 17.00
12.
Utnämning av en ledamot av Europeiska centralbankens direktion: Peter Praet (BE)
ECON/7/05430
2011/0802(NLE) 00003/2011 – C7-0058/2011
Föredragande:
Sharon Bowles (ALDE)
PR – PE460.742v01-00
Ansv. utsk.:
ECON –
· Antagande av förslag till betänkande
13.
EIB:s årsrapport för 2009
ECON/7/04197
2010/2248(INI)
Föredragande:
George Sabin Cutaş (S&D)
PR – PE454.577v01-00 AM – PE458.499v01-00
Ansv. utsk.:
ECON –
Rådg. utsk.:
CONT
· Antagande av förslag till betänkande
14.
Yrkesmässiga gränsöverskridande vägtransporter av eurokontanter mellan medlemsstaterna i euroområdet
ECON/7/03539
***I 2010/0204(COD) KOM(2010)0377 – C7-0186/2010
Föredragande:
Sophie Auconie (PPE)
PR – PE454.357v01-00 AM – PE456.920v01-00
Ansv. utsk.:
ECON –
Rådg. utsk.:
EMPL, TRAN
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 27 januari 2011 kl. 12.00
15.
Utvidgning av tillämpningsområdet för Europaparlamentets och rådets förordning (EU) om yrkesmässiga gränsöverskridande vägtransporter av eurokontanter mellan medlemsstaterna i euroområdet
ECON/7/03542
2010/0206(APP) 17787/2010 – C7-0025/2011
Föredragande:
Sophie Auconie (PPE)
PR – PE454.641v01-00
Ansv. utsk.:
ECON –
Rådg. utsk.:
EMPL, TRAN
· Antagande av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 27 januari 2011 kl. 12.00
16.
Framtiden för sociala tjänster av allmänt intresse
ECON/7/01752
2009/2222(INI)
Föredragande av yttrande:
Sophie Auconie (PPE)
PA – PE452.520v01-00 AM – PE452.844v01-00
Ansv. utsk.:
EMPL –
Proinsias De Rossa (S&D)
PR – PE438.251v02-00
Rådg. utsk.:
ECON, IMCO, REGI, FEMM
· Antagande av förslag till yttrande
*** Omröstningen avslutas ***
16 mars 2011 kl. 17.10–17.55
17.
Försäkringsgarantisystem
ECON/7/04779
2011/2010(INI) KOM(2010)0370
Föredragande:
Peter Skinner (S&D)
PR – PE456.981v01-00
Ansv. utsk.:
ECON –
Rådg. utsk.:
IMCO, JURI
· Behandling av förslag till betänkande
16 mars 2011 kl. 17.55–18.30
18.
Global ekonomisk styrning
ECON/7/04780
2011/2011(INI)
Föredragande:
Gunnar Hökmark (PPE)
Ansv. utsk.:
ECON –
Rådg. utsk.:
INTA, EMPL
· Inledande diskussion
19.
Övriga frågor
20.
Datum för nästa sammanträde
Måndagen den 21 mars 2011 kl. 15.00–18.30 Tisdagen den 22 mars 2011 kl. 9.00–12.30 och kl. 15.00–18.30
Michelle Bachelet: Demokrati är också integration, pluralism och mångfald
Kvinnors rättigheter/Lika möjligheter
2011-03-30 - 17:19
Demokrati handlar inte bara om att rösta, det är också om integration, pluralism och mångfald sa Bachelet när vi pratade med henne om hinder för jämställdhet, kvinnors roll i politiken och om hennes egen erfarenhet.
Vilka är de största hindren för jämställdhet?
Michelle Bachelet : Kvinnors brist på makt.
Därför är den viktigaste uppgiften att stärka kvinnorna.
När kvinnor har makt, när deras röstar blir hörda det är då de deltar i politiken, när de aktivt deltar i sina länders ekonomiska och sociala utveckling - då kan vi stärka deras potential som arbetare med rättigheter, som entreprenörer i små- och medelstora företag med tillgång till kredit eller mark, när det gäller jordbrukare, eller med fler kvinnor på beslutsfattande poster i den privata sektorn.
Med fler kvinnor på direktörsposter kommer jämställdhetsfrågor att få en särskild dimension.
Med fler kvinnor i politiken ändras dessutom politiken.
Kvaliteten ändras och blir bättre.
Därför är det så viktigt att ha både män och kvinnor.
Våld mot kvinnor är ett annat hinder för jämställdhet.
Slutligen är en viktig aspekt garanti för att hänsyn tas till kvinnors oro och problem i konflikter eller i länder som är på väg ut ur konflikter.
Hur ser du på kvinnornas roll i revolutionerna i arabvärlden?
M.B .: Jag har precis varit i Egypten.
Jag tror att det är väldigt viktigt att se till att kvinnornas närvaro på Tahrirtorget, där unga män och kvinnor kämpade för ett mer demokratiskt land, inte går förlorad.
Låt inte deras närvaro, delaktighet och syn försvinna.
Kvinnor är också med i utformningen och uppbyggnaden av ett mer demokratiskt samhälle.
Har du i ditt yrkesliv stött på hinder bara för att du är kvinna?
Jag fick inte uppfattningen att världen var begränsad för kvinnor.
Tvärtom, den som jobbar hårt och lägger ner all sin intelligens, kunskap och passion i värderingar och saker den tror på kan uppnå sina drömmar.
Detta är ett viktigt budskap: ofta syns inte kvinnor i områden med makt, utan i tjänster, och den symboliska bilden av kvinnor med makt går förlorad.
Michelle Bachelet
Född: 1951
Chef för UN Women sedan september 2010
SV
1
PHOTO
20110329PHT16601.jpg
SV
2
LINK
/wps-europarl-internet/frd/vod/player?eventCode=20110324-0900-COMMITTEE&language=EN&byLeftMenu=researchcommittee&category=COMMITTEE&format=wmv#anchor1
SV
3
LINK
http://www.unwomen.org/2011/03/executive-director-michelle-bachelet-addresses-european-parliament/
SV
4
LINK
/sv/headlines/content/20110223FCS14178/html/Internationella-kvinnodagen-2011-Dags-f%C3%B6r-handling!
SV
5
LINK
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Ledamöterna oense om kärnkraftens framtid i Europa
Energi
Plenarsammanträde
2011-04-07 - 14:06
Europaparlamentet avslog på torsdagen en resolution om kärnkraftssäkerhet i Europa med 264 ja-röster mot 300 nej-röster och 61 nedlagda röster.
Parlamentets politiska grupper var oeniga på flera frågor, vilket ledde till att sluttexten, så som den ändrats av de antagna ändringsförslagen, avslogs.
Debatten om kärnkraft hölls på onsdagen den 6 april.
20110407IPR17186 Se på debatten igen (klicka på 6 april 2011) Sammanfattning av debatten
SV
1
LINK
/wps-europarl-internet/frd/vod/research-by-date?language=sv
SV
2
LINK
/sv/headlines/content/20110324FCS16438/9/html/Debatt-om-k%C3%A4rnkraften-i-Europa-k%C3%A4rnkraftverken-ska-stresstestas
-//EP//DTD IM-PRESS 20050901 IPR DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 IPR DOC XML V0//EN
Utskottet för kultur och utbildning
CULT(2011)0411_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Måndagen den 11 april 2011 kl. 15.00–18.30
Tisdagen den 12 april 2011 kl. 9.00–12.30
Lokal: ASP 3G-2
11 april 2011 kl. 15.00–18.30
1.
Godkännande av föredragningslistan
2.
Justering av protokollen från sammanträdena den
· 3 mars 2011 PV – PE458.863v01-00
· 16–17 mars 2011 PV – PE460.793v01-00
3.
Meddelanden från ordföranden
I närvaro av rådet och kommissionen
4.
Diskussion med Neelie Kroes (kommissionens vice ordförande och kommissionsledamot med ansvar för den digitala agendan)
5.
Meddelande från kommissionen till Europaparlamentet, rådet, Europeiska ekonomiska och sociala kommittén och Regionkommittén: En agenda för ny kompetens och arbetstillfällen – EU:s bidrag till full sysselsättning
KOM(2010)0682
Föredragande av yttrande: Katarína Nevedalová (S&D) Ansv. utsk.: EMPL – Diskussion
6.
Den europeiska plattformen mot fattigdom och social utestängning
CULT/7/05571
2011/2052(INI) KOM(2010)0758
Föredragande av yttrande:
Silvia Costa (S&D)
Ansv. utsk.:
EMPL –
Frédéric Daerden (S&D)
· Diskussion
7.
Den europeiska terminen för samordning av den ekonomiska politiken KOM(2011)0011 Föredragande av yttrande: Hannu Takkula (ALDE) Diskussion
Inom stängda dörrar
8.
Samordnarnas sammanträde
* * *
12 april 2011 kl. 9.00–12.30
I närvaro av rådet och kommissionen
*** Omröstning ***
9.
Unga på väg – En ram för att förbättra de europeiska utbildningssystemen
CULT/7/04823
2010/2307(INI) KOM(2010)0477
Föredragande:
Milan Zver (PPE)
PR – PE454.698v01-00 AM – PE460.798v01-00
Ansv. utsk.:
CULT* –
Rådg. utsk.:
EMPL* –
Jutta Steinruck (S&D)
AD – PE456.784v03-00 AM – PE458.607v01-00
· Antagande av förslag till betänkande
10.
Investering i framtiden: en ny flerårig budgetram för ett konkurrenskraftigt och hållbart Europa för alla
CULT/7/04980
2010/2211(INI)
Föredragande av yttrande:
Cătălin Sorin Ivan (S&D)
PA – PE456.926v01-00 AM – PE460.772v01-00 DT – PE456.827v01-00 DT – PE456.968v02-00
Ansv. utsk.:
SURE –
Salvador Garriga Polledo (PPE)
PR – PE458.649v02-00 DT – PE454.599v01-00 DT – PE454.604v02-00 DT – PE454.602v01-00
· Antagande av förslag till yttrande
11.
Ett samlat grepp på skyddet av personuppgifter i Europeiska unionen
CULT/7/05178
2011/2025(INI) KOM(2010)0609
Föredragande av yttrande:
Seán Kelly (PPE)
PA – PE458.791v01-00 AM – PE460.957v01-00
Ansv. utsk.:
LIBE –
Axel Voss (PPE)
PR – PE460.636v01-00 DT – PE460.638v01-00 DT – PE460.637v01-00
· Antagande av förslag till yttrande
*** Omröstningen avslutas ***
12.
Diskussion med Androulla Vassiliou (kommissionsledamot för utbildning, kultur, flerspråkighet och ungdom)
13.
Utveckling av idrottens europeiska dimension KOM(2011)0012 Föredragande: Santiago Fisas Ayxela (PPE) – Inledande diskussion
14.
Insatser för att minska antalet elever som lämnar skolan i förtid KOM(2011)0019 Föredragande: Mary Honeyball (S&D) – Inledande diskussion
15.
Godkännande av samordnarnas beslut
16.
Övriga frågor
17.
Nästa sammanträde
· 25 maj 2011 kl. 15.00–18.30
· 26 maj 2011 kl. 9.00–12.30
Budgetutskottet
BUDG(2011)0502_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Måndagen den 2 maj 2011 kl. 15.00–18.30
Bryssel
Lokal: PHS 1A002
1.
Godkännande av föredragningslistan
2.
Meddelanden från ordföranden
3.
Justering av protokollet från sammanträdet den
· 31 mars 2011 PV – PE462.740v01-00
Lissabonpaketet: den fleråriga budgetramen och det interinstitutionella avtalet
4.
Den fleråriga budgetramen för 2007–2013
BUDG/7/04291
2010/0048(APP) 16973/2010 – C7-0024/2011
Föredragande:
Reimer Böge (PPE)
Ansv. utsk.:
BUDG –
· Diskussion
5.
Det interinstitutionella avtalet om samarbete i budgetfrågor
BUDG/7/02927
2010/2073(INI)
Föredragande:
Reimer Böge (PPE)
Ansv. utsk.:
BUDG –
· Diskussion
* * *
6.
Finansiella bestämmelser för unionens årliga budget
BUDG/7/04994
***I 2010/0395(COD) KOM(2010)0815 – C7-0016/2011
Medföredragande:
Crescenzio Rivellini (PPE) Ingeborg Gräßle (PPE)
DT – PE458.811v01-00
Ansv. utsk.:
BUDG –
· Diskussion
7.
Utnyttjande av Europeiska fonden för justering för globaliseringseffekter: General Motors Belgien
BUDG/7/05844
2011/2074(BUD) KOM(2011)0212 – C7-0096/2011
Föredragande:
Barbara Matera (PPE)
Ansv. utsk.:
BUDG –
· Diskussion
*** Omröstning ***
8.
EU:s tecknande av nya kapitalandelar i Europeiska banken för återuppbyggnad och utveckling (EBRD)
BUDG/7/05290
***I 2011/0014(COD) KOM(2011)0034 – C7-0038/2011
Föredragande av yttrande:
Ivailo Kalfin (S&D)
PA – PE460.940v01-00 AM – PE462.763v01-00
Ansv. utsk.:
ECON –
Sharon Bowles (ALDE)
PR – PE462.517v01-00
· Behandling och antagande
9.
Nytt protokoll om fastställande av de fiskemöjligheter och den ekonomiska ersättning som föreskrivs i partnerskapsavtalet om fiske mellan Europeiska unionen och Republiken Seychellerna
BUDG/7/04742
2010/0335(NLE) 17238/2010 – C7-0031/2011
Föredragande av yttrande:
François Alfonsi (Verts/ALE)
PA – PE458.616v01-00
Ansv. utsk.:
PECH –
Alain Cadec (PPE)
PR – PE460.600v01-00
· Behandling och antagande
10.
Nytt protokoll om fastställande av de fiskemöjligheter och den ekonomiska ersättning som föreskrivs i partnerskapsavtalet om fiske mellan Demokratiska Republiken São Tomé e Príncipe och EG
BUDG/7/04877
2010/0355(NLE) KOM(2010)0735
Föredragande av yttrande:
François Alfonsi (Verts/ALE)
PA – PE458.615v01-00
Ansv. utsk.:
PECH –
Luis Manuel Capoulas Santos (S&D)
PR – PE458.638v01-00
· Behandling och antagande
11.
2011 års budget: avsnitt III – kommissionen Föredragande: Sidonia Elżbieta Jędrzejewska (PPE) – DEC 07/2011 – Eventuellt andra önskemål om överföringar
12.
2011 års budget: övriga avsnitt Föredragande: Helga Trüpel (Verts/ALE) – ReK EST 1/2011 – Eventuellt andra önskemål om överföringar
13.
Fastighetspolitik
BUDG/7/04688
Föredragande:
Monika Hohlmeier (PPE)
DT – PE456.906v02-00 DT – PE445.867v02-00
· Diskussion
*** Omröstningen avslutas ***
Studier
Studie om Europeiska investeringsbanken
14.
Övriga frågor
15.
Datum för nästa sammanträde
· 5 maj 2011 kl. 9.00–12.30 och kl. 12.30–13.30 (samordnarnas sammanträde) (i Bryssel)
Karlspriset för ungdomar 2011 till "Europe & Me"
Ungdom
2011-05-31 - 16:38
Jerzy Buzek delar ut Europeiska Karlspriset för ungdomar 2011 Det brittiska webbmagasinet "Europe & Me" fick på tisdagen, 31 maj, årets europeiska Karlspris för ungdomar vid en ceremoni i tyska Aachen.
Talman Jerzy Buzek sa vid prisceremonin att Europe & Me fick priset eftersom det är "extremt originellt".
- Jag tror att projektets huvudbudskap är att Europa är, kan och bör vara cool.
"Europe & Me" är ett livsstilsmagasin på nätet, det skapades 2007 av unga européer för unga européer.
Mottot är att göra "Europa mer personligt" och skapa en plats för initiativ där det också går att finna likasinnade.
Andrapriset gick till det grekiska kortfilmsprojektet "Balkans Beyond Borders" och tredjepriset till det spanska kulturella utbytesprogrammet "Escena Erasmus Project".
tjänar som förebild för ungdomar i Europa och ger praktiska exempel på européer som lever i samhörighet med varandra.
20110526STO20295 Pressmeddelande Europeiska Karlspriset för ungdomar Pressmeddelande: Svensk nyhetssajt tävlar för att vinna ungdomspris Webbmagasin vann Karlspriset för ungdomar Video
SV
1
PHOTO
20110527PHT20386.jpg
SV
2
LINK
/en/pressroom/content/20110530IPR20497/html/Europe-Me-wins-European-Charlemagne-Youth-Prize-2011
SV
3
LINK
http://www.charlemagneyouthprize.eu/view/sv/introduction.html
SV
4
LINK
/sv/pressroom/content/20110322IPR16119/html/Svensk-nyhetssajt-t%C3%A4vlar-f%C3%B6r-att-vinna-ungdomspris
SV
5
MULTIMEDIA
20110530MLT20487.mp4
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
TECKENFÖRKLARING
*
Samrådsförfarande
***
Godkännandeförfarande
***I
Ordinarie lagstiftningsförfarande (första behandlingen)
***II
Ordinarie lagstiftningsförfarande (andra behandlingen)
***III
FÖRKORTNINGAR FÖR UTSKOTTENS NAMN
AFET:
DEVE:
Utskottet för utveckling
INTA:
Utskottet för internationell handel
BUDG:
Budgetutskottet
CONT:
Budgetkontrollutskottet
ECON:
Utskottet för ekonomi och valutafrågor
EMPL:
Utskottet för sysselsättning och sociala frågor
ENVI:
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
ITRE:
Utskottet för industrifrågor, forskning och energi
IMCO:
Utskottet för den inre marknaden och konsumentskydd
TRAN:
Utskottet för transport och turism
REGI:
Utskottet för regional utveckling
AGRI:
PECH:
Fiskeriutskottet
CULT:
Utskottet för kultur och utbildning
JURI:
Utskottet för rättsliga frågor
LIBE:
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
AFCO:
Utskottet för konstitutionella frågor
FEMM:
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
PETI:
Utskottet för framställningar
DROI:
Underutskottet för mänskliga rättigheter
SEDE:
Underutskottet för säkerhet och försvar
FÖRKORTNINGAR FÖR DE POLITISKA GRUPPERNA
PPE:
Europeiska folkpartiets grupp (kristdemokrater)
S&D:
Gruppen Progressiva förbundet av socialdemokrater och demokrater i Europaparlamentet
ALDE:
Gruppen Alliansen liberaler och demokrater för Europa
Verts/ALE:
Gruppen De gröna/Europeiska fria alliansen
ECR:
Gruppen Europeiska konservativa och reformister
GUE/NGL:
Gruppen Europeiska enade vänstern/Nordisk grön vänster
EFD:
Gruppen Frihet och demokrati i Europa
NI:
Grupplösa
Återupptagande av sessionen
Uttalanden av talmannen
Justering av protokollet från föregående sammanträde
Tolkning av arbetsordningen
Parlamentets sammansättning
Begäran om fastställelse av parlamentarisk immunitet
Valprövning
Utskottens och delegationernas sammansättning
Undertecknande av rättsakter som antagits i enlighet med det ordinarie lagstiftningsförfarandet
Rättelser (artikel 216 i arbetsordningen)
Inkomna dokument
Bortfallna skriftliga förklaringar
Muntliga frågor och skriftliga förklaringar (ingivande)
Avtalstexter översända av rådet
Kommissionens åtgärder till följd av parlamentets resolutioner
Framställningar
Anslagsöverföringar
Arbetsplan
Högtidlighållande av 10-årsdagen av den 11 september 2001 (uttalande av talmannen)
Pågående Doha-förhandlingar (debatt)
En effektiv råvarustrategi för Europa (debatt)
Anföranden på en minut om frågor av politisk vikt
EU:s strategi för terrorismbekämpning: viktiga framsteg och kommande utmaningar (kortfattad redogörelse)
Revisionspolitik: lärdomar av krisen (kortfattad redogörelse)
Fiske i Svarta havet (kortfattad redogörelse)
En säker olje- och gasverksamhet till havs (kortfattad redogörelse)
Kvinnors företagande i små och medelstora företag (kortfattad redogörelse)
Situationen för kvinnor som närmar sig pensionsåldern (kortfattad redogörelse)
Föredragningslista för nästa sammanträde
Avslutande av sammanträdet
NÄRVAROLISTA
EUROPAPARLAMENTET
SESSIONEN 2011
− 2012
Sammanträdena den 12
− 15 september 2011
1 Återupptagande av sessionen
Sammanträdet öppnades kl. 17.05.
2 Uttalanden av talmannen
Talmannen gjorde ett uttalande om de initiativ som EU nyligen tagit för att bekämpa den ekonomiska krisen och ett uttalande om resultatet av konflikten i Libyen.
Talare:
Talmannen meddelade att parlamentet skulle delta i FN:s internationella demokratidag den 15 september 2011.
Talmannen fördömde det våld som ledamoten Sajjad Karim hade utsatts för den 2 juli 2011 och uttryckte sitt stöd.
Talare:
Niccolò Rinaldi och
Mario Mauro yttrade sig om den italienske premiärministerns besök.
3 Justering av protokollet från föregående sammanträde
Protokollet från föregående sammanträde justerades.
° ° ° °
Danuta Maria Hübner hade meddelat att hon hade avsett att rösta för punkt 16 led b (originaltexten) i betänkandet
A7-0210/2011 vid omröstningen den 6 juli 2011.
4 Tolkning av arbetsordningen
Tolkning av artikel 51 i arbetsordningen:
"
"
Tolkning av artikel 192 i arbetsordningen:
"
De grupplösa ledamöterna utgör inte en politisk grupp i den mening som avses i artikel 30 och får därför inte utse samordnare, vilka är de enda som har rätt att delta i samordnarnas möten.
Syftet med samordnarnas möten är att förbereda utskottens beslut, och de får inte ersätta utskottsmötena utan uttrycklig delegering.
Därför måste behörigheten att fatta beslut vid samordnarnas möten delegeras på förhand.
I avsaknad av en sådan delegering får samordnarna endast anta rekommendationer, som måste godkännas formellt av utskottet i efterhand.
Under alla omständigheter måste de grupplösa ledamöternas tillgång till information garanteras i enlighet med principen om icke-diskriminering genom överlämnande av information och genom att en person från de grupplösas sekretariat närvarar vid samordnarnas möten.
"
Om så är fallet ska frågan gå till omröstning i parlamentet.
5 Parlamentets sammansättning
° ° ° °
De belgiska myndigheterna hade meddelat att Philippe De Backer hade valts till ledamot av Europaparlamentet i stället för
Dirk Sterckx .
Parlamentet noterade att detta skulle gälla från och med den 7 september 2011.
° ° ° °
De behöriga italienska myndigheterna hade den 19 juli 2011 meddelat att
Luigi de Magistris plats var vakant med verkan från och med den 19 juli 2011 och noterade valet av Andrea Zanoni med verkan från samma datum.
° ° ° °
6 Begäran om fastställelse av parlamentarisk immunitet
Den före detta ledamoten av Europaparlamentet
7 Valprövning
På förslag från utskottet JURI beslutade parlamentet att godkänna mandaten för
Tarja Cronberg och
Dimitrios Droutsas med verkan från och med den 22 juni 2011 samt för Franck Proust med verkan från och med den 23 juni 2011.
8 Utskottens och delegationernas sammansättning
Grupperna ALDE, Verts/ALE och GUE/NGL hade begärt att följande utnämningar skulle godkännas:
utskottet AFET:
Tarja Cronberg
utskottet CONT:
Giommaria Uggias
utskottet IMCO:
Cornelis de Jong i stället för
Kyriacos Triantaphyllides
utskottet TRAN: Andrea Zanoni i stället för
Giommaria Uggias , Philippe De Backer
utskottet PECH:
Jorgo Chatzimarkakis i stället för
Britta Reimers
utskottet LIBE:
Kyriacos Triantaphyllides i stället för
Cornelis de Jong
delegationen för förbindelserna med Mashrekländerna: Andrea Zanoni
delegationen till den gemensamma parlamentarikerkommittén EU-Mexiko: Philippe De Backer
delegationen till den parlamentariska församlingen EU-Latinamerika: Philippe De Backer
Dessa utnämningar skulle betraktas som godkända om det inte framställdes några invändningar mot detta före justeringen av detta protokoll.
9 Undertecknande av rättsakter som antagits i enlighet med det ordinarie lagstiftningsförfarandet
Talmannen meddelade att han tillsammans med rådets ordförande på onsdagen skulle underteckna följande antagna rättsakter, i enlighet med det ordinarie lagstiftningsförfarandet (artikel 74 i arbetsordningen):
- Europaparlamentets och rådets förordning om ändring av förordning (EG) nr 2006/2004 om samarbete mellan de nationella tillsynsmyndigheter som ansvarar för konsumentskyddslagstiftningen (00023/2011/LEX - C7-0240/2011 - 2011/0001(COD) )
- Europaparlamentets och rådets förordning om upphävande av rådets förordning (EG) nr 1541/98 om ursprungsbevis för vissa textilprodukter enligt avdelning XI i Kombinerade nomenklaturen som övergått till fri omsättning i gemenskapen och om villkoren för godkännande av dessa ursprungsbevis, och om ändring av rådets förordning (EEG) nr 3030/93 om gemensamma regler för import av vissa textilprodukter från tredje land (00025/2011/LEX - C7-0239/2011 - 2010/0272(COD) )
- Europaparlamentets och rådets beslut om Europaåret för aktivt åldrande och solidaritet mellan generationerna (2012) (00020/2011/LEX - C7-0238/2011 - 2010/0242(COD) )
- Europaparlamentets och rådets direktiv om ändring av direktiv 2000/25/EG vad gäller bestämmelser om traktorer som släpps ut på marknaden enligt flexibilitetssystemet (00019/2011/LEX - C7-0237/2011 - 2010/0301(COD) )
10 Rättelser
(artikel 216 i arbetsordningen)
Rättelse (
P7_TA-PROV(2011)0313(COR01)
)
till Europaparlamentets ståndpunkt fastställd vid första behandlingen den 5 juli 2011 inför antagandet av Europaparlamentets och rådets direktiv 2011/.../EU om ändring av Europaparlamentets och rådets direktiv 97/9/EG om system för ersättning till investerare
P7_TA-PROV(2011)0313 - ( KOM(2010)0371 – C7-0174/201 0 – 2010/0199(COD) - ECON
- Rättelse (
P7_TA-PROV(2011)0218(COR01)
)
till Europaparlamentets ståndpunkt fastställd vid andra behandlingen den 11 maj 2011 inför antagandet av Europaparlamentets och rådets förordning (EU) nr .../2011 om benämningar på textilfibrer och etikettering och märkning av fibersammansättningen i textilprodukter och om upphävande av rådets direktiv 73/44/EEG, Europaparlamentets och rådets direktiv 96/73/EG och Europaparlamentets och rådets direktiv2008/121/EG
I enlighet med artikel 216.4 i arbetsordningen ska dessa rättelser anses ha godkänts om det inte senast 48 timmar efter tillkännagivandet inkommit en begäran från en politisk grupp eller minst 40 ledamöter om att de ska bli föremål för omröstning.
Rättelserna finns tillgängliga på webbplatsen Séance en direct.
11 Inkomna dokument
Talmannen hade mottagit följande dokument:
1) från parlamentets utskott, betänkanden:
- ***I Betänkande om förslaget till Europaparlamentets och rådets beslut om Europeiska unionens tecknande av nya kapitalandelar i Europeiska banken för återuppbyggnad och utveckling (EBRD) till följd av beslutet att utöka detta kapital ( KOM(2011)0034 - C7-0038/2011 - 2011/0014(COD) ) - utskottet ECON - Föredragande: Sharon Bowles ( A7-0227/2011 )
- Betänkande om nuvarande och framtida förvaltning av fisket i Svarta havet ( 2010/2113(INI) ) - utskottet PECH - Föredragande: Iliana Malinova Iotova ( A7-0236/2011 )
- Betänkande om försäkringsgarantisystem ( 2011/2010(INI) ) - utskottet ECON - Föredragande: Peter Skinner ( A7-0243/2011 )
- *** Rekommendation om förslaget till rådets beslut om ingående av avtalet mellan Europeiska unionen, Schweiziska edsförbundet och Furstendömet Liechtenstein om ändring av tilläggsavtalet mellan Europeiska gemenskapen, Schweiziska edsförbundet och Furstendömet Liechtenstein om utvidgning av tillämpningsområdet för avtalet mellan Europeiska gemenskapen och Schweiziska edsförbundet om handel med jordbruksprodukter till att även omfatta Furstendömet Liechtenstein (16209/2010 - C7-0125/2011 - 2010/0313(NLE) ) - utskottet INTA - Föredragande: Béla Glattfelder ( A7-0248/2011 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets förordning om upphävande av förordning (EEG) nr 429/73 om särskilda bestämmelser om import till gemenskapen av vissa varor som omfattas av förordning (EEG) nr 1059/69 och med ursprung i Turkiet samt förordning (EG) nr 215/2000 om förlängning under 2000 av åtgärder som avses i förordning (EG) nr 1416/95 om införande av vissa koncessioner i form av gemenskapstullkvoter under 1995 för vissa bearbetade jordbruksprodukter ( KOM(2010)0756 - C7-0004/2011 - 2010/0367(COD) ) - utskottet INTA - Föredragande: Vital Moreira ( A7-0250/2011 )
- Betänkande om bättre lagstiftning, subsidiaritet och proportionalitet samt smart lagstiftning ( 2011/2029(INI) ) - utskottet JURI - Föredragande: Sajjad Karim ( A7-0251/2011 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets förordning om upphävande av vissa obsoleta rådsrättsakter inom området för den gemensamma jordbrukspolitiken ( KOM(2010)0764 - C7-0006/2011 - 2010/0368(COD) ) - utskottet AGRI - Föredragande: Paolo De Castro ( A7-0252/2011 )
- Betänkande om en ny handelspolitik för Europa i samband med Europa 2020-strategin ( 2010/2152(INI) ) - utskottet INTA - Föredragande: Daniel Caspary ( A7-0255/2011 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets förordning om ändring av förordning (EG) nr 428/2009 om upprättande av en gemenskapsordning för kontroll av export, överföring, förmedling och transitering av produkter med dubbla användningsområden ( KOM(2010)0509 - C7-0289/2010 - 2010/0262(COD) ) - utskottet INTA - Föredragande: Vital Moreira ( A7-0256/2011 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets förordning om upphävande av vissa obsoleta rådsrättsakter ( KOM(2010)0765 - C7-0009/2011 - 2010/0369(COD) ) - utskottet INTA - Föredragande: Vital Moreira ( A7-0257/2011 )
- Betänkande om att främja arbetskraftens rörlighet inom Europeiska unionen ( 2010/2273(INI) ) - utskottet EMPL - Föredragande: Traian Ungureanu ( A7-0258/2011 )
- *** Rekommendation om utkastet till rådets beslut om ingående av ett avtal mellan Europeiska unionen och Förbundsrepubliken Brasiliens regering om civil luftfartssäkerhet (13989/1/2010 - C7-0336/2010 - 2010/0143(NLE) ) - utskottet TRAN - Föredragande: Silvia-Adriana Ţicău ( A7-0259/2011 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets beslut om närmare föreskrifter för den offentliga reglerade tjänst (PRS) som erbjuds via det globala satellitnavigeringssystem via satellit som upprättats genom Galileoprogrammet ( KOM(2010)0550 - C7-0318/2010 - 2010/0282(COD) ) - utskottet ITRE - Föredragande: Norbert Glante ( A7-0260/2011 )
- * Betänkande om utkastet till rådets förordning om ändring av förordning (EG) nr 521/2008 om bildande av det gemensamma företaget för bränsleceller och vätgas ( KOM(2011)0224 - C7-0120/2011 - 2011/0091(NLE) ) - utskottet ITRE - Föredragande: Herbert Reul ( A7-0261/2011 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets förordning om ändring av rådets förordning (EG) nr 1234/2007 vad gäller avtalsvillkor inom sektorn för mjölk och mjölkprodukter ( KOM(2010)0728 - C7-0408/2010 - 2010/0362(COD) ) - utskottet AGRI - Föredragande: James Nicholson ( A7-0262/2011 )
- Betänkande om rörlighet och integrering av personer med funktionsnedsättning och EU:s handikappstrategi 2010–2020 ( 2010/2272(INI) ) - utskottet EMPL - Föredragande: Ádám Kósa ( A7-0263/2011 )
- Betänkande om europeisk trafiksäkerhet 2011–2020 ( 2010/2235(INI) ) - utskottet TRAN - Föredragande: Dieter-Lebrecht Koch ( A7-0264/2011 )
- Betänkande om Europa, världens främsta resmål – en ny politisk ram för europeisk turism ( 2010/2206(INI) ) - utskottet TRAN - Föredragande: Carlo Fidanza ( A7-0265/2011 )
- ***I Betänkande om förslag till Europaparlamentets och rådets förordning om kvalitetsordningar för jordbruksprodukter ( KOM(2010)0733 - C7-0423/2010 - 2010/0353(COD) ) - utskottet AGRI - Föredragande: Iratxe García Pérez ( A7-0266/2011 )
- Betänkande om begäran om upphävande av Hans-Peter Martins immunitet ( 2011/2104(IMM) ) - utskottet JURI - Föredragande: Tadeusz Zwiefka ( A7-0267/2011 )
- *** Rekommendation om utkastet till rådets beslut om ingående av avtal mellan Europeiska unionen och Republiken Island och Konungariket Norge om förfarande för överlämnande mellan Europeiska unionens medlemsstater och Island och Norge (05307/2010 - C7-0032/2010 - 2009/0192(NLE) ) - utskottet LIBE - Föredragande: Rui Tavares ( A7-0268/2011 )
- Betänkande om ensidiga förklaringar i protokoll från rådets möten ( 2011/2090(INI) ) - utskottet AFCO - Föredragande: Rafał Trzaskowski ( A7-0269/2011 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets direktiv om bedömning av inverkan på miljön av vissa offentliga och privata projekt (kodifiering) ( KOM(2011)0189 - C7-0095/2011 - 2011/0080(COD) ) - utskottet JURI - Föredragande: Sajjad Karim ( A7-0272/2011 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets förordning om integritet och öppenhet på energimarknaderna ( COM(2010)0726 - C7-0407/2010 - 2010/0363(COD) ) - utskottet ITRE - Föredragande: Jorgo Chatzimarkakis ( A7-0273/2011 )
- *** Rekommendation om utkastet till rådets beslut om ingående, på Europeiska unionens vägnar, av konventionen om bevarande och förvaltning av det fria havets fiskeresurser i södra Stilla havet (08135/2011 - C7-0098/2011 - 2011/0047(NLE) ) - utskottet PECH - Föredragande: Carmen Fraga Estévez ( A7-0274/2011 )
- Betänkande om tillämpning av direktivet om medling i medlemsstaterna, dess inverkan på medlingen och dess utnyttjande i domstolarna ( 2011/2026(INI) ) - utskottet JURI - Föredragande: Arlene Mccarthy ( A7-0275/2011 )
- *** Rekommendation om förslaget till rådets beslut om ingående av avtalet genom skriftväxling mellan Europeiska unionen och Konungariket Norge om ytterligare handelsförmåner för jordbruksprodukter, uppnådda på grundval av artikel 19 i avtalet om Europeiska ekonomiska samarbetsområdet (14206/2010 - C7-0101/2011 - 2010/0243(NLE) ) - utskottet INTA - Föredragande: Helmut Scholz ( A7-0276/2011 )
- Betänkande om förslaget till Europaparlamentets och rådets beslut om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning (ansökan EGF/2010/007 AT/Steiermark och Niederösterreich från Österrike) ( KOM(2011)0340 - C7-0159/2011 - 2011/2124(BUD) ) - utskottet BUDG - Föredragande: Barbara Matera ( A7-0277/2011 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets förordning om ändring av rådets förordning (EG) nr 2007/2004 om inrättande av en europeisk byrå för förvaltningen av det operativa samarbetet vid Europeiska unionens medlemsstaters yttre gränser (Frontex) ( KOM(2010)0061 - C7-0045/2010 - 2010/0039(COD) ) - utskottet LIBE - Föredragande: Simon Busuttil ( A7-0278/2011 )
- Betänkande om förslaget till Europaparlamentets och rådets beslut om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning (ansökan EGF/2010/008 AT/AT&S från Österrike) ( KOM(2011)0339 - C7-0160/2011 - 2011/2125(BUD) ) - utskottet BUDG - Föredragande: Barbara Matera ( A7-0279/2011 )
- *** Rekommendation om utkastet till rådets beslut om ingående på Europeiska unionens vägnar av 2006 års internationella avtal om tropiskt timmer (05812/2011 - C7-0061/2011 - 2006/0263(NLE) ) - utskottet INTA - Föredragande: Vital Moreira ( A7-0280/2011 )
- ***I Betänkande om förslaget till Europaparlamentets och rådets förordning om ändring av rådets förordning (EG) nr 1234/2007 vad gäller handelsnormer ( KOM(2010)0738 - C7-0422/2010 - 2010/0354(COD) ) - utskottet AGRI - Föredragande: Iratxe García Pérez ( A7-0281/2011 )
- Betänkande om EU:s policyram för att hjälpa utvecklingsländer att stärka livsmedelsförsörjningen ( 2010/2100(INI) ) - utskottet DEVE - Föredragande: Gabriele Zimmer ( A7-0284/2011 )
- Betänkande om EU:s strategi för terrorismbekämpning: viktiga framsteg och kommande utmaningar ( 2010/2311(INI) ) - utskottet LIBE - Föredragande: Sophia In 't Veld ( A7-0286/2011 )
- Betänkande om en effektiv råvarustrategi för Europa ( 2011/2056(INI) ) - utskottet ITRE - Föredragande: Reinhard Bütikofer ( A7-0288/2011 )
- Betänkande med Europaparlamentets rekommendationer till rådet, kommissionen och Europeiska utrikestjänsten om förhandlingarna om associeringsavtalet mellan EU och Moldavien ( 2011/2079(INI) ) - utskottet AFET - Föredragande: Graham Watson ( A7-0289/2011 )
- Betänkande om utmaningen att uppnå en säker olje- och gasverksamhet till havs ( 2011/2072(INI) ) - utskottet ITRE - Föredragande: Vicky Ford ( A7-0290/2011 )
- Betänkande om situationen för kvinnor som närmar sig pensionsåldern ( 2011/2091(INI) ) - utskottet FEMM - Föredragande: Edit Bauer ( A7-0291/2011 )
2) från ledamöterna
2.2) förslag till ändring av arbetsordningen (artikel 212 i arbetsordningen)
hänvisat till
ansvarigt utskott :
AFCO
12 Bortfallna skriftliga förklaringar
13 Muntliga frågor och skriftliga förklaringar
(ingivande)
Talmannen hade mottagit följande dokument från ledamöterna:
1) muntliga frågor (artikel 115 i arbetsordningen):
- (
O-000135/2011 ) från
Jo Leinen ,
Richard Seeber och
Theodoros Skylakakis , för utskottet ENVI, till kommissionen:
Ett helhetsbetonat grepp på frågan om antropogena utsläpp av annat slag än koldioxid och av relevans för klimatet ( B7-0418/2011 ) ;
- (
O-000148/2011 ) från
Monica Luisa Macovei ,
Mariya Nedelcheva ,
Simon Busuttil och
Manfred Weber för PPE-gruppen , till rådet:
Åtgärder för att minska klyftan mellan korruptionslagstiftningen och verkligheten ( B7-0419/2011 ) ;
- (
O-000149/2011 ) från
Monica Luisa Macovei ,
Mariya Nedelcheva ,
Simon Busuttil och
Manfred Weber för PPE-gruppen , till kommissionen:
Åtgärder för att minska klyftan mellan korruptionslagstiftningen och verkligheten ( B7-0420/2011 ) ;
- (
O-000153/2011 ) från
Pervenche Berès och
Karima Delli , för utskottet EMPL, till kommissionen:
EU:s strategi mot hemlöshet ( B7-0421/2011 ) ;
- (
O-000154/2011 ) från
Cornelis de Jong ,
Cornelia Ernst ,
Nikolaos Chountis ,
Søren Bo Søndergaard och
Alfreds Rubiks för GUE/NGL-gruppen , till rådet:
Skärpta åtgärder mot korruption ( B7-0422/2011 ) ;
- (
O-000155/2011 ) från
Cornelis de Jong ,
Cornelia Ernst ,
Nikolaos Chountis ,
Søren Bo Søndergaard och
Alfreds Rubiks för GUE/NGL-gruppen , till kommissionen:
Skärpta åtgärder mot korruption ( B7-0423/2011 ) ;
- (
O-000172/2011 ) från
Jan Philipp Albrecht och
Judith Sargentini för Verts/ALE-gruppen , till rådet:
Åtgärder för att minska klyftan mellan korruptionslagstiftningen och verkligheten ( B7-0424/2011 ) ;
- (
O-000173/2011 ) från
Jan Philipp Albrecht och
Judith Sargentini för Verts/ALE-gruppen , till kommissionen
Åtgärder för att minska klyftan mellan korruptionslagstiftningen och verkligheten ( B7-0425/2011 ) ;
- (
O-000178/2011 ) från
Ana Gomes ,
Claude Moraes ,
Rita Borsellino och
Rosario Crocetta för S&D-gruppen , till rådet:
Genomförande av EU:s åtgärdspaket för korruptionsbekämpning ( B7-0427/2011 ) ;
- (
O-000179/2011 ) från
Ana Gomes ,
Claude Moraes ,
Rita Borsellino och
Rosario Crocetta för S&D-gruppen , till kommissionen:
Genomförande av EU:s åtgärdspaket för korruptionsbekämpning ( B7-0428/2011 ) ;
- (
O-000180/2011 ) från
Herbert Reul , för utskottet ITRE, till kommissionen:
EU:s politiska strategi för ITU:s världskonferens om radiokommunikationer (WRC-12) ( B7-0429/2011 ) ;
- (
O-000185/2011 ) från
Michael Theurer ,
Niccolò Rinaldi ,
Catherine Bearder ,
Marielle De Sarnez och
Jürgen Creutzmann för ALDE-gruppen ,
Godelieve Quisthoudt-Rowohl ,
Othmar Karas ,
Daniel Caspary och
Cristiana Muscardini för PPE-gruppen ,
Robert Sturdy för ECR-gruppen , till kommissionen:
Internationalisering av europeiska små och medelstora företag ( B7-0430/2011 ) ;
- (
O-000190/2011 ) från
Timothy Kirkhope för ECR-gruppen , till rådet:
Åtgärder för att bekämpa korruption ( B7-0431/2011 ) ;
- (
O-000191/2011 ) från
Timothy Kirkhope för ECR-gruppen , till kommissionen:
Åtgärder för att bekämpa korruption ( B7-0432/2011 ) ;
- (
O-000193/2011 ) från
Sonia Alfano ,
Renate Weber ,
Sarah Ludford ,
Jan Mulder ,
Louis Michel ,
Nathalie Griesbeck ,
Ramon Tremosa i Balcells ,
Nadja Hirsch ,
Stanimir Ilchev och
Jens Rohde för ALDE-gruppen , till rådet:
Åtgärder för att minska klyftan mellan korruptionslagstiftningen och verkligheten ( B7-0433/2011 ) ;
- (
O-000194/2011 ) från
Sonia Alfano ,
Renate Weber ,
Sarah Ludford ,
Jan Mulder ,
Louis Michel ,
Nathalie Griesbeck ,
Ramon Tremosa i Balcells ,
Nadja Hirsch ,
Stanimir Ilchev och
Jens Rohde för ALDE-gruppen , till kommissionen:
Åtgärder för att minska klyftan mellan korruptionslagstiftningen och verkligheten ( B7-0434/2011 ) .
2) skriftliga förklaringar införda i registret (artikel 123 i arbetsordningen)
-
Patrick Le Hyaric ,
Robert Atkins ,
Margrete Auken ,
Véronique De Keyser och
Niccolò Rinaldi ,
om Europeiska unionens erkännande av den palestinska staten (0027/2011);
-
Marian-Jean Marinescu ,
Ádám Kósa ,
Eva Lichtenberger ,
Gesine Meissner och
Gianni Pittella ,
om behovet av allmänt tillgängliga 112-larmtjänster (0035/2011);
-
Valdemar Tomaševski ,
om stärkande av kärnsäkerheten i EU och i angränsande länder (0036/2011);
-
Spyros Danellis ,
Maria Da Graça Carvalho ,
Kyriakos Mavronikolas ,
Alyn Smith och
Giommaria Uggias ,
om inrättandet av pakten mellan öar som ett officiellt europeiskt initiativ (0037/2011);
-
Harlem Désir ,
Cornelis de Jong ,
Corinne Lepage ,
Ulrike Lunacek och
Mariya Nedelcheva ,
om att erkänna diskrimineringstester, där de ger positiva resultat, som rättsliga bevisa på rasdiskriminering
(0038/2011).
14 Avtalstexter översända av rådet
Rådet hade översänt vidimerade kopior av följande dokument:
– a
–
–
–
avtal mellan Europeiska unionen och Republiken Indonesiens regering om vissa luftfartsaspekter,
–
samarbetsmemorandum mellan Europeiska unionen och internationella civila luftfartsorganisationen om en ram för utökat samarbete,
–
–
protokoll mellan Europeiska unionen och Republiken Kap Verde om fastställande av de fiskemöjligheter och den ekonomiska ersättning som föreskrivs i det gällande partnerskapsavtalet om fiske mellan de två parterna.
16 Framställningar
Den 26 juli 2011
Joachim Ledwoch (nr 0707/2011); Widla Renata Michalska (Stowarzyszenie Przyjazna Rokietnica) (nr 0708/2011); (namnet konfidentiellt) (nr 0709/2011); Jozef Adamski (nr 0710/2011); T S Ostrowski (4 underskrifter) (nr 0711/2011); Helmut Geuking (Partei Soziale Gerechtigkeit) (nr 0712/2011); Dieter Schädlich (nr 0713/2011); Jadwiga Szczodra (nr 0714/2011); Rita Kasumu (11 underskrifter) (nr 0715/2011); Adolf Śmieszek (nr 0716/2011); Dietrich Bechstein (Flugtouristik Deitzsch e.V.) (nr 0717/2011); Robert Wilk (nr 0718/2011); Daniela Theiss (nr 0719/2011); Siegfried Schäfer (nr 0720/2011); Vincent Grünberg (nr 0721/2011); Ingeborg Flandergan (nr 0722/2011); Simon Jakob (Jakob & Kollegen) (nr 0723/2011); Kazimierz Gała (nr 0724/2011); Bernhard Kempen (Universität zu Köln) (nr 0725/2011); Enrico Venezia (nr 0726/2011); Mihai Dulgheru (nr 0727/2011); Kosyo Kosev (KOSKO LTD) (nr 0728/2011); Fiona Munro (nr 0729/2011); Agostino Furfaro (nr 0730/2011); Kevin Forbes (nr 0731/2011); Clive Smith (nr 0732/2011); Christian Nekvedavicius (Lithuanian association for the protection of human rights) (nr 0733/2011); Patrick Pearse Heffernan (nr 0734/2011); (namnet konfidentiellt) (nr 0735/2011); Mario Marocco (Associazione nazionale operatori elettrici indipendenti) (nr 0736/2011); Hugo Wolff (nr 0737/2011); Carina Diana Lintia (nr 0738/2011); Desislava Rayanovo (nr 0739/2011); Antonio Luis García Martínez (nr 0740/2011); Francisco Bernal Alfonso (nr 0741/2011); (namnet konfidentiellt) (nr 0742/2011); Jaime Sanfelix Palau (Laserood 2007, S.L.) (nr 0743/2011); María Antonia Busto Ortiz (nr 0744/2011); Alberto de la Pe
ña Guillén (nr 0745/2011); Cristina Díaz Espiñeira (nr 0746/2011); Asunción Cremades Campos (nr 0747/2011); José Ramón Gil Benito (nr 0748/2011).
Den 3 augusti 2011
Ritva Suortti (nr 0749/2011); (namnet konfidentiellt) (nr 0750/2011); Jean-Louis Posté (Président de Mauves Vivantes) (nr 0751/2011); (namnet konfidentiellt) (nr 0752/2011); Dries Emmen (O.O.B.T.) (nr 0753/2011); Salvador Peiró Gómez (Centro de Acuicultura Experimental) (nr 0754/2011); Adorjáni István (nr 0755/2011); (namnet konfidentiellt) (nr 0756/2011); Zacharias Tsirtos (nr 0757/2011); Victor Alexandru Kovacs (nr 0758/2011); Elise Michaud (nr 0759/2011); Rodulfo Galido Torres (nr 0760/2011); Silvia Beltrán Pallarés (Plataforma Europea de los Consumidores y del Medio Ambiente) (nr 0761/2011); André Goretti (Président de la Fédération Autonome des Sapeurs-pompiers professionnels) (nr 0762/2011); Judit Szima (Tettrekész Magyar Rend
ő rség Szakszervezete) (nr 0763/2011).
Den 12 augusti 2011
Ewa Rydzyńska (nr 0764/2011); Symanski Botho (nr 0765/2011); Heinz Greiner Walter (nr 0766/2011); Aartur Hirschmann (nr 0767/2011); Józef Suszczewicz (nr 0768/2011); Helga Hung (nr 0769/2011); Wolfgang Panthel (nr 0770/2011); Algimantas Jonas Petraitis (nr 0771/2011); Tsvetan Georgiev Rangelov (nr 0772/2011); Marek Iwanowski (nr 0773/2011); Jerzy Aplej (nr 0774/2011); Wilfried Gesing (nr 0775/2011); Martin Wagner (2 underskrifter) (nr 0776/2011); Agata Szczęśniak-Sevastiadi (nr 0777/2011); Krzysztof Tokarz (nr 0778/2011); Georg Schömer (nr 0779/2011); Igor Herzog (nr 0780/2011); Manfred Tröger (nr 0781/2011); Krzysztof Tomasik (nr 0782/2011); Ehrhardt Bekeschus (nr 0783/2011); Stefanija Groh (nr 0784/2011); Jolanta Smagłowska (nr 0785/2011); (namnet konfidentiellt) (nr 0786/2011); Edelmiro Cuadrado Alba (nr 0787/2011); (namnet konfidentiellt) (nr 0788/2011); Alejandro Pastor (nr 0789/2011); Pepe Montes Guillén (Agrupación de Labradores del Pozuelo S.A) (nr 0790/2011); Mikel Basabe Kortabarria (Aralar) (nr 0791/2011); Sebastiano Licciardello (Studio Legale Prof.
Avv.
Sebastiano Licciardello) (90 underskrifter) (nr 0792/2011); José Ignacio Francés Sánchez (IFS ABOGADOS) (74 underskrifter) (nr 0793/2011); Joaquim Boadas De Quintana (FECASARM ) (nr 0794/2011); Antonio Luis García Martínez (nr 0795/2011); (namnet konfidentiellt) (nr 0796/2011); (namnet konfidentiellt) (nr 0797/2011); Giorgio Gurrieri (nr 0798/2011); Giuseppe Sorrentino (Federconsumatori) (nr 0799/2011); Henryk Nowakowski (nr 0800/2011); Vladimirs Strazdi
ņš (Austrumu Medic
īn a Co., Ltd.) (nr 0801/2011); European Policy Office WWF (WWF European Policy Office) (nr 0802/2011); Vladimir Dimitrov (BAR - Association Bulgare de Recyclage) (nr 0803/2011); Sergio López (nr 0804/2011); Sándor Polgár (nr 0805/2011); Diego Zunino (3 973 underskrifter) (nr 0806/2011); Milcho Georgiev Stanoev (nr 0807/2011); Helene Lopes (nr 0808/2011); María Inés Barcia (Asociación AAPV) (nr 0809/2011); (namnet konfidentiellt) (nr 0810/2011); Garbis Vincentiu Kehaiyan (nr 0811/2011); Silvia Beltrán Pallarés (Plataforma Europea de los Consumidores y del Medio Ambiente) (nr 0812/2011); Catherine Abéguilé-Petit (nr 0813/2011); Sara Consuegra (nr 0814/2011); Anna Poulsen (nr 0815/2011); Pavlos Arvanitopoulos (nr 0816/2011); Jean-Antoine Enrile (nr 0817/2011); Samir Bekenniche (nr 0818/2011); (namnet konfidentiellt) (nr 0819/2011); Jan a.a.
Huijsman (nr 0820/2011); Εmmanuel Perrakis (nr 0821/2011); Juan Carlos Uriarte Amarica (Agaden Association) (nr 0822/2011); (namnet konfidentiellt) (nr 0823/2011); (namnet konfidentiellt) (nr 0824/2011); (namnet konfidentiellt) (2 underskrifter) (nr 0825/2011); Andrea Cocco (nr 0826/2011); Anita Brandt (ART OPUS GmbH) (2 underskrifter) (nr 0827/2011); Patrick Anazonwu (nr 0828/2011); John Hadman (nr 0829/2011); Polykarpos Markaras (nr 0830/2011); Leszek Janczyk (nr 0831/2011); (namnet konfidentiellt) (nr 0832/2011); Markus Knops (nr 0833/2011);
Ö mer Cakmak (nr 0834/2011); Peter Spyrka (nr 0835/2011); Noelia Ferrer Martínez (Ebame & Associats) (nr 0836/2011); Gianfranco Concetti (nr 0837/2011); Hans Lennros (Upadek AB) (nr 0838/2011); (namnet konfidentiellt) (nr 0839/2011); Arabadzhieva Neli Petrova (3 underskrifter) (nr 0840/2011); Magdalena Zdravkova Slavova (4 underskrifter) (nr 0841/2011); Finn Skovgaard (nr 0842/2011); Alessandro Michelucci (nr 0843/2011); Remo Pulcini (Progetto Mezzogiorno) (nr 0844/2011); Mark Borda (nr 0845/2011); Giuseppe Giacomini (Conte & Giacomini) (nr 0846/2011); Mohammad Reza Fardoom (Solidarity, Independence, Democracy (SID)) (nr 0847/2011); Antonio Luis García Martínez (nr 0848/2011); (namnet konfidentiellt) (nr 0849/2011); Basem Kasem (för 156 syriska studenter) (156 underskrifter) (nr 0850/2011).
Den 8 september 2011
Kurt Bilogan (nr 0851/2011); Wolfgard Christine Ruckershauer (nr 0852/2011); P Kuecklich-Scheer (115 underskrifter) (nr 0853/2011); Wilhelm Hök (nr 0854/2011); Ralf Schneeweiss (nr 0855/2011); Edward Zytka (nr 0856/2011); (namnet konfidentiellt) (nr 0857/2011); Ryszard Kopera (nr 0858/2011); Schmid Peter (nr 0859/2011); Kind Paul (nr 0860/2011); Christel Krombolz (2 underskrifter) (nr 0861/2011); Maria Klein (nr 0862/2011); Michał Combik (nr 0863/2011); Mehl Ulrich (nr 0864/2011); Günter Dillikrath (nr 0865/2011); Peter Mohr (nr 0866/2011); Appel c/o Schmidt Manfred (nr 0867/2011); Michael Stoltenberg (nr 0868/2011); Safet Alimehaj (www.klage-gegen-ljubljanska-banka.de) (nr 0869/2011); Reinhold Leckert (nr 0870/2011); K. T. Baranowska (nr 0871/2011); Georg Geisenfelder (nr 0872/2011); (namnet konfidentiellt) (nr 0873/2011); Michael Witfer (Sportboot Gemeinschaft Saale-Elster e.V.) (nr 0874/2011); Ursula Lehmann (nr 0875/2011); Prof.
Dr.
ří H
ů lka (Union of Municipalities of the Sumava national park) (nr 0904/2011); Michele Bertucco (Associazione Legambiente Veneto) (6 underskrifter) (nr 0905/2011); Alessandro Lanci (Nuovo Senso Civico) (2 underskrifter) (nr 0906/2011); Ljubima Jordanova Dimitrova (nr 0907/2011); (namnet konfidentiellt) (nr 0908/2011); Maria Teresa Motas de Oliveira (nr 0909/2011).
17 Anslagsöverföringar
18 Arbetsplan
Nästa punkt på föredragningslistan var fastställandet av arbetsplanen.
Det slutgiltiga förslaget till föredragningslista för sammanträdesperioden september I 2011 (PE 470.595/PDOJ) hade delats ut.
Följande ändringar hade föreslagits i enlighet med artikel 140 i arbetsordningen:
Måndag, tisdag, onsdag
Inga ändringar hade föreslagits.
Torsdag
PPE-gruppen begärde att man redan under innevarande sammanträdesperiod skulle rösta om resolutionsförslag framlagda som avslutning på debatten om situationen i Libyen
(punkt 180 i PDOJ)
.
Talare:
Cristian Dan Preda för PPE-gruppen motiverade begäran;
Niccolò Rinaldi för ALDE-gruppen uttalade sig för denna begäran och
Rebecca Harms för Verts/ALE-gruppen emot.
Följande tidsfrister hade fastställts:
resolutionsförslag: tisdagen den 13 september kl. 10.00
ändringsförslag och gemensamma förslag till resolution: onsdagen den 14 september kl. 10.00
ändringsförslag till gemensamma förslag till resolution: onsdagen den 14 september kl. 11.00
Omröstningen skulle äga rum på torsdagen.
° ° ° °
Arbetsplanen var därmed fastställd.
19 Högtidlighållande av 10-årsdagen av den 11 september 2001
(uttalande av talmannen)
Talmannen gjorde ett uttalande med anledning av 10-årsdagen av den 11 september 2001.
Parlamentet höll en tyst minut.
20
Pågående Doha-förhandlingar
(debatt)
Uttalande av kommissionen:
Pågående Doha-förhandlingar
Karel De Gucht (ledamot av kommissionen) gjorde ett uttalande.
Talare:
Godelieve Quisthoudt-Rowohl för PPE-gruppen,
Vital Moreira för S&D-gruppen,
Niccolò Rinaldi för ALDE-gruppen,
Keith Taylor för Verts/ALE-gruppen, och
Helmut Scholz för GUE/NGL-gruppen .
Talare:
William (The Earl of) Dartmouth för EFD-gruppen,
Nicole Sinclaire , grupplös,
Daniel Caspary ,
George Sabin Cutaş , som även besvarade en fråga ("blått kort") från
Hans-Peter Martin ,
Yannick Jadot ,
João Ferreira ,
Bastiaan Belder ,
Hans-Peter Martin ,
Georgios Papastamkos ,
Corina Creţu ,
Judith Sargentini ,
Christofer Fjellner ,
Béla Glattfelder och
Elisabeth Köstinger .
Talare:
Antonio Tajani (vice ordförande för kommissionen) .
-
Vital Moreira , för utskottet INTA,
om läget i förhandlingarna om utvecklingsagendan från Doha ( B7-0478/2011 ) .
Talmannen förklarade debatten avslutad.
Omröstning:
punkt 5.12 i protokollet av den 14.9.2011
.
21
En effektiv råvarustrategi för Europa
(debatt)
Betänkande om en effektiv råvarustrategi för Europa [ 2011/2056(INI) ] - Utskottet för industrifrågor, forskning och energi.
Föredragande: Reinhard Bütikofer ( A7-0288/2011 )
Reinhard Bütikofer redogjorde för sitt betänkande.
Talare:
Antonio Tajani (vice ordförande för kommissionen) .
Talare:
Birgit Schnieber-Jastram (föredragande av yttrande från utskottet DEVE) ,
Bernd Lange (föredragande av yttrande från utskottet INTA),
Daciana Octavia Sârbu (föredragande av yttrande från utskottet AGRI),
Pilar del Castillo Vera för PPE-gruppen,
Marita Ulvskog för S&D-gruppen,
Lena Ek för ALDE-gruppen,
Bas Eickhout för Verts/ALE-gruppen,
Julie Girling för ECR-gruppen,
Marisa Matias för GUE/NGL-gruppen,
Jaroslav Paška för EFD-gruppen,
Adam Gierek ,
Michael Theurer ,
Ilda Figueiredo ,
Bastiaan Belder ,
Jolanta Emilia Hibner ,
Riikka Manner ,
Esther de Lange ,
Silvia-Adriana Ţicău ,
Karl-Heinz Florenz ,
Csaba Sándor Tabajdi ,
Theodor Dumitru Stolojan ,
Herbert Reul och
Marian-Jean Marinescu .
Följande talare yttrade sig i enlighet med ögonkontaktsförfarandet:
Mairead McGuinness ,
Monika Smolková ,
Andreas Mölzer ,
Seán Kelly ,
Vasilica Viorica Dăncilă ,
Oreste Rossi ,
Elena Băsescu och
Talare:
Antonio Tajani och
Reinhard Bütikofer .
ORDFÖRANDESKAP: Rainer WIELAND Vice talman
Omröstning:
punkt 5.22 i protokollet av den 13.9.2011
.
22 Anföranden på en minut om frågor av politisk vikt
Följande ledamöter höll, i enlighet med artikel 150 i arbetsordningen, ett anförande på en minut för att uppmärksamma parlamentet på frågor av politisk vikt:
Rosa Estaràs Ferragut ,
Vasilica Viorica Dăncilă ,
Chris Davies ,
Rui Tavares ,
Marek Henryk Migalski ,
Kyriacos Triantaphyllides ,
Oreste Rossi ,
Slavi Binev ,
László Tőkés ,
Cătălin Sorin Ivan ,
Georgios Toussas ,
Gerard Batten ,
Andrew Henry William Brons ,
Jim Higgins ,
Silvia-Adriana Ţicău ,
Ilda Figueiredo ,
Alajos Mészáros ,
Maria Eleni Koppa ,
Willy Meyer ,
Georgios Papanikolaou ,
Antigoni Papadopoulou ,
Eleni Theocharous ,
George Sabin Cutaş ,
Jarosław Kalinowski ,
Boris Zala ,
Mairead McGuinness ,
Luís Paulo Alves ,
Seán Kelly och
Nuno Melo .
23
EU:s strategi för terrorismbekämpning: viktiga framsteg och kommande utmaningar
(kortfattad redogörelse)
Betänkande om EU:s strategi för terrorismbekämpning: viktiga framsteg och kommande utmaningar [ 2010/2311(INI) ] - Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor.
Föredragande: Sophia in 't Veld ( A7-0286/2011 )
Sophia in 't Veld redogjorde för betänkandet.
Följande talare yttrade sig i enlighet med ögonkontaktsförfarandet:
Agustín Díaz de Mera García Consuegra ,
Juan Fernando López Aguilar ,
Izaskun Bilbao Barandica ,
Jan Philipp Albrecht ,
Jaroslav Paška ,
Martin Ehrenhauser ,
Teresa Jiménez-Becerril Barrio ,
Anna Hedh ,
Elena Băsescu och
Monika Flašíková Beňová .
Talare:
Antonio Tajani (vice ordförande för kommissionen) .
ORDFÖRANDESKAP: Roberta ANGELILLI Vice talman
Omröstning:
punkt 5.23 i protokollet av den 13.9.2011
.
24
Revisionspolitik: lärdomar av krisen
(kortfattad redogörelse)
Betänkande om revisionspolitik: lärdomar av krisen [ 2011/2037(INI) ] - Utskottet för rättsliga frågor.
Föredragande: Antonio Masip Hidalgo ( A7-0200/2011 )
Antonio Masip Hidalgo redogjorde för betänkandet.
Följande talare yttrade sig i enlighet med ögonkontaktsförfarandet:
Monika Flašíková Beňová ,
Evelyn Regner ,
Rui Tavares ,
Kay Swinburne och
Jaroslav Paška .
Talare:
Michel Barnier (ledamot av kommissionen) .
Talmannen förklarade punkten avslutad.
Omröstning:
punkt 5.17 i protokollet av den 13.9.2011
.
25
Fiske i Svarta havet
(kortfattad redogörelse)
Betänkande om nuvarande och framtida förvaltning av fiske i Svarta havet [ 2010/2113(INI) ] - Fiskeriutskottet.
Föredragande: Iliana Malinova Iotova ( A7-0236/2011 )
Iliana Malinova Iotova redogjorde för betänkandet.
Följande talare yttrade sig i enlighet med ögonkontaktsförfarandet:
Guido Milana ,
Vasilica Viorica Dăncilă ,
Josefa Andrés Barea ,
Silvia-Adriana Ţicău ,
Evgeni Kirilov och
João Ferreira .
Talare:
Antonio Tajani (vice ordförande för kommissionen) .
Talmannen förklarade punkten avslutad.
Omröstning:
punkt 5.24 i protokollet av den 13.9.2011
.
26
En säker olje- och gasverksamhet till havs
(kortfattad redogörelse)
Betänkande om utmaningen att uppnå en säker olje- och gasverksamhet till havs [ 2011/2072(INI) ] - Utskottet för industrifrågor, forskning och energi.
Föredragande: Vicky Ford ( A7-0290/2011 )
Vicky Ford redogjorde för betänkandet.
Följande talare yttrade sig i enlighet med ögonkontaktsförfarandet:
Alajos Mészáros ,
Monika Flašíková Beňová ,
Silvia-Adriana Ţicău ,
Ilda Figueiredo och
Michèle Rivasi .
Talare:
Antonio Tajani (vice ordförande för kommissionen) .
Talmannen förklarade punkten avslutad.
Omröstning:
punkt 5.25 i protokollet av den 13.9.2011
.
27
Kvinnors företagande i små och medelstora företag
(kortfattad redogörelse)
Betänkande om kvinnors företagande i små och medelstora företag [ 2010/2275(INI) ] - Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män.
Föredragande: Marina Yannakoudakis ( A7-0207/2011 )
Marina Yannakoudakis redogjorde för betänkandet.
Följande talare yttrade sig i enlighet med ögonkontaktsförfarandet:
Regina Bastos ,
Miroslav Mikolášik ,
Vasilica Viorica Dăncilă ,
Monika Flašíková Beňová ,
Silvia-Adriana Ţicău ,
Ilda Figueiredo ,
Elena Băsescu ,
Jaroslav Paška ,
Alajos Mészáros ,
Katarína Neveďalová ,
Antigoni Papadopoulou och
Angelika Werthmann .
Talare:
Antonio Tajani (vice ordförande för kommissionen) .
Talmannen förklarade punkten avslutad.
Omröstning:
punkt 5.26 i protokollet av den 13.9.2011
.
28
Situationen för kvinnor som närmar sig pensionsåldern
(kortfattad redogörelse)
Betänkande om situationen för kvinnor som närmar sig pensionsåldern [ 2011/2091(INI) ] - Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män.
Föredragande: Edit Bauer ( A7-0291/2011 )
Edit Bauer redogjorde för betänkandet.
Följande talare yttrade sig i enlighet med ögonkontaktsförfarandet:
Christa Klaß ,
Miroslav Mikolášik ,
Vasilica Viorica Dăncilă ,
Ilda Figueiredo ,
Monika Flašíková Beňová ,
Katarína Neveďalová och
Antigoni Papadopoulou .
Talare:
Antonio Tajani (vice ordförande för kommissionen) .
Talmannen förklarade punkten avslutad.
Omröstning:
punkt 5.18 i protokollet av den 13.9.2011
.
29 Föredragningslista för nästa sammanträde
Föredragningslistan för nästa sammanträde fastställdes ("Föredragningslista" PE 470.595/OJMA).
30 Avslutande av sammanträdet
Sammanträdet avslutades kl. 22.50.
Klaus Welle
Miguel Angel Martínez Martínez
Generalsekreterare
Vice talman
NÄRVAROLISTA
Följande skrev på:
Abad
Áder
Albrecht
Alfano
Alvaro
Alves
Andreasen
Andrés Barea
Andrikienė
Angourakis
Antinoro
Antonescu
Antoniozzi
Arias Echeverría
Arif
Arlacchi
Arsenis
Ashworth
Atkins
Attard-Montalto
Auconie
Audy
Auken
Aylward
Ayuso
Bach
Badia i Cutchet
Bagó
Balčytis
Baldassarre
Bartolozzi
Băsescu
Bastos
Batten
Bauer
Bearder
Belder
Belet
Bélier
Benarab-Attou
Bendtsen
Bennahmias
Berès
Berlato
Berlinguer
Berman
Bielan
Bilbao Barandica
Binev
Bisky
Bizzotto
Blinkevičiūtė
Bodu
Bokros
Bonsignore
Borghezio
Borsellino
Boştinaru
Boulland
Bové
Bozkurt
Bradbourn
Brantner
Březina
Brons
Brzobohatá
Bufton
Bullmann
Buşoi
Busuttil
Bütikofer
Buzek
Cabrnoch
Callanan
van de Camp
Campbell Bannerman
Cancian
Capoulas Santos
Caronna
Carvalho
Casa
Cashman
Casini
Caspary
Castex
del Castillo Vera
Cavada
Cercas
Češková
Chatzimarkakis
Chichester
Childers
Chountis
Claeys
Clark
Coelho
Cofferati
Colman
Comi
Corazza Bildt
Silvia Costa
Cozzolino
Cramer
Creţu
Creutzmann
Crocetta
Cutaş
Cymański
Czarnecki
Frédéric Daerden
van Dalen
Dăncilă
Danellis
Danjean
Dantin
(The Earl of) Dartmouth
Daul
David
Davies
De Angelis
De Backer
de Brún
Dehaene
De Keyser
Delvaux
De Mita
De Rossa
De Sarnez
Deß
De Veyrac
Díaz de Mera García Consuegra
Dodds
Domenici
Donskis
Dorfmann
Droutsas
Duff
Durant
Dušek
Ehler
Ehrenhauser
Eickhout
Ek
El Khadraoui
Elles
Enciu
Engström
Eppink
Ernst
Ertug
Essayah
Estaràs Ferragut
Estrela
Evans
Fajmon
Fajon
Falbr
Farage
Färm
Feio
Ferber
Fernandes
Elisa Ferreira
João Ferreira
Fidanza
Figueiredo
Fisas Ayxela
Fjellner
Flašíková Beňová
Flautre
Fleckenstein
Florenz
Fontana
Ford
Foster
Fox
Fraga Estévez
Franco
Gahler
Gál
Gallagher
Gallo
Gáll-Pelcz
García-Margallo y Marfil
García Pérez
Gardini
Gargani
Garriga Polledo
Gauzès
Gebhardt
Geier
Geringer de Oedenberg
Giannakou
Giegold
Gierek
Glante
Glattfelder
Godmanis
Goebbels
Goerens
Gollnisch
Gomes
Göncz
Goulard
de Grandes Pascual
Gräßle
Grech
Grelier
Grèze
Griesbeck
Griffin
Gróbarczyk
Groote
Grosch
Grossetête
Grzyb
Gualtieri
Guerrero Salom
Guillaume
Gurmai
Gutiérrez-Cortines
Gutiérrez Prieto
Gyürk
Haglund
Fiona Hall
Händel
Handzlik
Hannan
Harbour
Harkin
Hartong
Hassi
Haug
Häusling
Hedh
Helmer
Hénin
Herczog
Herranz García
Hibner
Higgins
Nadja Hirsch
Hoang Ngoc
Hohlmeier
Hökmark
Honeyball
Hortefeux
Danuta Maria Hübner
Hughes
Hyusmenova
Iacolino
Ibrisagic
Ilchev
Imbrasas
in 't Veld
Iotova
Iovine
Itälä
Iturgaiz Angulo
Ivan
Ivanova
Jaakonsaari
Jäätteenmäki
Jadot
Jahr
Jazłowiecka
Jędrzejewska
Jeggle
Jensen
Jiménez-Becerril Barrio
Joly
de Jong
Jordan Cizelj
Junqueras Vies
Juvin
Kacin
Kaczmarek
Kadenbach
Kalinowski
Kalniete
Kamall
Kamiński
Karas
Karim
Kasoulides
Kastler
Kazak
Kelam
Kelly
Kiil-Nielsen
Kirilov
Kirkhope
Klaß
Klinz
Klute
Koch
Koch-Mehrin
Kohlíček
Kolarska-Bobińska
Koppa
Korhola
Kósa
Köstinger
Koumoutsakos
Kovatchev
Kowal
Kozlík
Kozłowski
Kožušník
Krahmer
Kratsa-Tsagaropoulou
Krehl
Kreissl-Dörfler
Kuhn
Kukan
Lamassoure
Lambert
Lamberts
Landsbergis
Lange
de Lange
Langen
La Via
Lechner
Le Grip
Legutko
Lehne
Leinen
Lepage
Jean-Marie Le Pen
Liberadzki
Lichtenberger
Liese
Lisek
Lochbihler
Løkkegaard
López Aguilar
Lösing
Ludford
Ludvigsson
Luhan
Łukacijewska
Lulling
Lunacek
Lynne
Lyon
McAvan
McCarthy
McClarkin
McGuinness
McMillan-Scott
Macovei
Madlener
Manders
Mănescu
Mann
Manner
Marcinkiewicz
Marinescu
David Martin
Hans-Peter Martin
Martínez Martínez
Masip Hidalgo
Mastella
Mathieu
Matias
Mato Adrover
Matula
Mauro
Mavronikolas
Mayer
Mazzoni
Meissner
Melo
Méndez de Vigo
Menéndez del Valle
Merkies
Mészáros
Meyer
Migalski
Mikolášik
Milana
Millán Mon
Mirsky
Mölzer
Moraes
Moreira
Morin-Chartier
Mulder
Murphy
Muscardini
Nattrass
Nedelcheva
Neuser
Neveďalová
Newton Dunn
Neynsky
Nicholson
Nicolai
Niculescu
Niebler
van Nistelrooij
Nitras
Nuttall
Obermayr
Ojuland
Olbrycht
Olejniczak
Oomen-Ruijten
Őry
Ouzký
Oviir
Pack
Padar
Paksas
Paleckis
Paliadeli
Pallone
Panayotov
Panzeri
Papadopoulou
Papanikolaou
Papastamkos
Pargneaux
Paška
Patrão Neves
Patriciello
Paulsen
Peillon
Perello Rodriguez
Peterle
Pieper
Pietikäinen
Piotrowski
Pirillo
Pirker
Pittella
Plumb
Poc
Podimata
Ponga
Portas
Posselt
Pöttering
Poupakis
Preda
Provera
Quisthoudt-Rowohl
Rangel
Ransdorf
Rapkay
Rapti
Regner
Reimers
Remek
Repo
Reul
Riera Madurell
Ries
Rinaldi
Riquet
Rivasi
Rivellini
Rochefort
Rodust
Rohde
Roithová
Romero López
Romeva i Rueda
Ronzulli
Rosbach
Rossi
Roth-Behrendt
Rouček
Rübig
Rubiks
Rühle
Saïfi
Sánchez Presedo
Sanchez-Schmid
Sârbu
Sargentini
Sartori
Saryusz-Wolski
Sassoli
Saudargas
Schaake
Schaldemose
Schlyter
Olle Schmidt
Schnellhardt
Schnieber-Jastram
Scholz
Schöpflin
Schroedter
Martin Schulz
Schwab
Scottà
Scurria
Seeber
Sehnalová
Senyszyn
Serracchiani
Siekierski
Silvestris
Simon
Simpson
Sinclaire
Sippel
Siwiec
Skinner
Skrzydlewska
Skylakakis
Smith
Smolková
Sógor
Sommer
Søndergaard
Sonik
Sosa Wagner
Speroni
Staes
Stassen
Šťastný
Stavrakakis
Steinruck
Stevenson
Stihler
Stolojan
Emil Stoyanov
Strejček
Striffler
Sturdy
Surján
Susta
Svensson
Swinburne
Szájer
Tabajdi
Takkula
Tănăsescu
Tannock
Tarabella
Tarand
Tatarella
Tavares
Taylor
Teixeira
Terho
Thein
Theocharous
Theurer
Thyssen
Ţicău
Toia
Tőkés
Tomaševski
Tošenovský
Toussas
Trautmann
Tremopoulos
Tremosa i Balcells
Triantaphyllides
Trüpel
Tsoukalas
Turmes
Uggias
Ulmer
Ulvskog
Ungureanu
Urutchev
Uspaskich
Vadim Tudor
Vaidere
Vajgl
Vălean
Van Brempt
Vanhecke
Van Orden
Vattimo
Vaughan
Vergnaud
Verheyen
Vidal-Quadras
Vigenin
de Villiers
Vlasák
Vlasto
Voss
Wallis
Watson
Manfred Weber
Renate Weber
Weiler
Weisgerber
Werthmann
Westphal
Wieland
Wikström
Wils
Hermann Winkler
Iuliu Winkler
Wortmann-Kool
Yáñez-Barnuevo García
Yannakoudakis
Záborská
Zala
Zalba Bidegain
Zalewski
Zanicchi
Zanoni
Zasada
Ždanoka
Zeller
Zemke
Zimmer
Zver
Zwiefka
Lewandowski: parlamentet är mer mänskligt
Institutioner
2011-09-20 - 17:27
Janusz Lewandowski Parlamentets ledamöter har olika bakgrund och skilda erfarenheter.
I dag berättar Janusz Lewandowski om sina erfarenheter av att ta steget åt andra hållet - och gå från ledamot till att bli kommissionär.
Vad har flytten från parlamentet till kommissionen inneburit för dig?
Rent praktiskt var det en enorm förändring.
Men det finns också andra skillnader.
Förklara ...
I Europaparlamentet är det mer insyn i processen, öppnare, en slags politisk teater.
I kommissionen är det mer internt.
Efter att kollegiet har fattat beslut ska vi inte tala om skillnader mellan kommissionärerna.
Det handlar om enhet och att tala med en röst.
Parlamentet är också mer mänskligt, vänligare, och kommissionen är kallare, med fler koder och förfaranden.
Har du ändrat syn på parlamentet?
Min syn på parlamentet har förändrats.
Men huvudanledningen är inte min "förflyttning" utan att Europaparlamentet har fått nya befogenheter genom Lissabonfördraget.
Nu är det ett fullfjädrat lagstiftande organ med verkligt budgetansvar.
Mer fokus på lagstiftning och beslutsfattande än på resolutioner som ofta är tidskrävande och med liten praktisk nytta.
Jag tycker också om att parlamentet har bevarat en europeisk anda - trots större och mer "högröstade" euroskeptiker den här valperioden.
Har du nytta av din bakgrund i förhandlingar med Europaparlamentet?
Min insiderkunskap och förståelse för såväl Europaparlamentet som kommissionen är min stora fördel.
Jag tror dessutom att jag har mer trovärdighet [i Europaparlamentet] och jag har lyckats behålla informella och vänskapliga kontakter i parlamentet, främst i budgetutskottet.
Det är till stor nytta, särskilt i krissituationer.
Och mina erfarenheter från parlamentet bidrar också till kommissionens arbete.
20110916STO26854 Intervju Danuta Hubner Janusz Lewandowski i Europaparlamentet Kommissionär Janusz Lewandowski
SV
1
PHOTO
20110913PHT26592.jpg
SV
3
LINK
/members/expert/inOut/viewOutgoing.do?language=SV&id=23781
SV
4
LINK
http://ec.europa.eu/commission_2010-2014/lewandowski/index_en.htm
-//EP//TEXT IM-PRESS 20110902STO25898 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Budgetkontrollutskottet
CONT(2011)0919_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Utfrågning
Måndagen den 19 september 2011 kl. 15.00–18.30
Bryssel
Lokal: ASP - 3G-2
19 september 2011 kl. 15.00–18.30
1.
Godkännande av föredragningslistan
2.
Meddelanden från ordföranden
3.
Val av ordförande för CONT-utskottet
4.
Utfrågning om Europeiska revisionsrättens framtida roll: utmaningar framöver och möjliga reformer
CONT/7/06136
Föredragande:
Inés Ayala Sender (S&D)
5.
Övriga frågor
6.
Nästa sammanträde(n)
· 22 september 2011 kl. 9.00–12.30 (Bryssel)
· 22 september 2011 kl. 15.00–16.30 (Bryssel)
Håller livsmedel samma kvalitet i alla EU-länder?
Konsumenter
2011-10-10 - 15:30
©BELGA/Belpress Det kanske är ett relativt okänt fenomen i Västeuropa, men det kommer regelbundet klagomål från konsumenter i Central- och Östeuropa på skillnader mellan produkter som ska vara identiska.
I miljöutskottet tog Elena Oana Antonescu nyligen upp frågan om kvalitetsskillnader mellan olika livsmedelsprodukter som saluförs i EU.
I början av april 2011 genomförde den slovakiska konsumentorganisationen en undersökning av märkta livsmedelsprodukter i åtta EU-länder.
Bland annat testades Coca Cola-drycker, Tchibo espressokaffe och Milka-choklad.
Testet visade att olika ingredienser används i produkterna, endast Milka-chokladen var av identisk kvalitet i alla exemplar som testades.
Som svar på den muntliga frågan från Elena Oana Antonescu (EPP, Rumänien) förklarade kommissionens representant att tillverkarna ändrar ingredienser utifrån konsumenternas preferenser.
Exempelvis är det en lösare Nutella som säljs på den franska marknaden jämfört med Tyskland, helt enkelt eftersom brödet har olika konsistens.
Kommissionens representant sa att EU inte kan bestämma över receptet, men konsumenterna har rätt till information om ingredienserna.
Elena Oana Antonescu menade att konsumenterna visst är medvetna om kvalitetsskillnader och varnade för att det kan uppstå olika klassers konsumenter.
Pavel Poc (S&D, Tjeckien) sa att han dagligen får svara på frågor om detta.
En av hans väljare undrade exempelvis "vad EU tjänar till om den inte kan skydda sina konsumenter".
Antonescu beklagade att det inte finns någon "europeisk lagstiftning som straffar diskriminerande beteende" och insisterade på att kommissionen snabbt ska göra "ytterligare undersökningar och studier".
20111007STO28689 Muntlig fråga Miljöutskottet
SV
1
PHOTO
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//TEXT TA P7-TA-2011-0520 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0521 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0522 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0523 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0524 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0525 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0526 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0527 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0528 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0529 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0530 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0531 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0532 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0533 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0534 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0535 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0536 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0537 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0538 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0539 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0540 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0541 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0542 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0543 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0544 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0545 0 DOC XML V0//SV -//EP//TEXT TA P7-TA-2011-0546 0 DOC XML V0//SV
TECKENFÖRKLARING
*
Samrådsförfarande
***
Godkännandeförfarande
***I
Ordinarie lagstiftningsförfarande (första behandlingen)
***II
Ordinarie lagstiftningsförfarande (andra behandlingen)
***III
FÖRKORTNINGAR FÖR UTSKOTTENS NAMN
AFET:
DEVE:
Utskottet för utveckling
INTA:
Utskottet för internationell handel
BUDG:
Budgetutskottet
CONT:
Budgetkontrollutskottet
ECON:
Utskottet för ekonomi och valutafrågor
EMPL:
Utskottet för sysselsättning och sociala frågor
ENVI:
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
ITRE:
Utskottet för industrifrågor, forskning och energi
IMCO:
Utskottet för den inre marknaden och konsumentskydd
TRAN:
Utskottet för transport och turism
REGI:
Utskottet för regional utveckling
AGRI:
PECH:
Fiskeriutskottet
CULT:
Utskottet för kultur och utbildning
JURI:
Utskottet för rättsliga frågor
LIBE:
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
AFCO:
Utskottet för konstitutionella frågor
FEMM:
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
PETI:
Utskottet för framställningar
DROI:
Underutskottet för mänskliga rättigheter
SEDE:
Underutskottet för säkerhet och försvar
FÖRKORTNINGAR FÖR DE POLITISKA GRUPPERNA
PPE:
Europeiska folkpartiets grupp (kristdemokrater)
S&D:
Gruppen Progressiva förbundet av socialdemokrater och demokrater i Europaparlamentet
ALDE:
Gruppen Alliansen liberaler och demokrater för Europa
Verts/ALE:
Gruppen De gröna/Europeiska fria alliansen
ECR:
Gruppen Europeiska konservativa och reformister
GUE/NGL:
Gruppen Europeiska enade vänstern/Nordisk grön vänster
EFD:
Gruppen Frihet och demokrati i Europa
NI:
Grupplösa
Öppnande av sammanträdet
Inkomna dokument
Val av Europaparlamentets talman
Val av Europaparlamentets talman (fortsättning)
Val av Europaparlamentets vice talmän (tidsfrist för inlämning av nomineringar)
Val av Europaparlamentets vice talmän
Val av Europaparlamentets vice talmän (fortsättning)
Val av Europaparlamentets vice talmän (fortsättning)
Föredragningslista för nästa sammanträde
Avslutande av sammanträdet
NÄRVAROLISTA
Bilaga 1
Bilaga 2
PROTOKOLL
ORDFÖRANDESKAP: Jerzy BUZEK
Talman
1 Öppnande av sammanträdet
Sammanträdet öppnades kl. 09.00.
2 Inkomna dokument
Talmannen hade mottagit följande dokument från rådet och kommissionen:
- Förslag till Europaparlamentets och rådets förordning om programmet för europeisk statistik 2013–2017 ( COM(2011)0928 - C7-0001/2012 - 2011/0459(COD) )
hänvisat till
ansvarigt utskott :
ECON
rådgivande utskott :
FEMM, ENVI, EMPL, BUDG, REGI
- Förslag till rådets beslut om ingående av protokollet mellan Europeiska unionen och Republiken Guinea-Bissau om fastställande av de fiskemöjligheter och den ekonomiska ersättning som föreskrivs i det gällande partnerskapsavtalet om fiske mellan de två parterna (15178/2011 - C7-0003/2012 - 2011/0257(NLE) )
hänvisat till
ansvarigt utskott :
PECH
rådgivande utskott :
DEVE, BUDG
hänvisat till
ansvarigt utskott :
IMCO
rådgivande utskott :
CULT, AFET, ENVI, EMPL, ITRE, JURI, ECON, LIBE, INTA, TRAN, REGI
- Förslag till Europaparlamentets och rådets förordning om ändring av rådets förordningar (EG) nr 2008/97, (EG) nr 779/98 och (EG) nr 1506/98 på områdena import av olivolja och andra jordbruksprodukter från Turkiet när det gäller delegerade befogenheter och genomförandebefogenheter som ska ges kommissionen ( COM(2011)0918 - C7-0005/2012 - 2011/0453(COD) )
hänvisat till
ansvarigt utskott :
INTA
rådgivande utskott :
AGRI
hänvisat till
ansvarigt utskott :
IMCO
rådgivande utskott :
AFET, ENVI, EMPL, ITRE, JURI, ECON, LIBE, INTA, TRAN, REGI
- Förslag till rådets förordning om Europeiska atomenergigemenskapens forsknings- och utbildningsprogram (2014–2018) som kompletterar Horisont 2020 – ramprogrammet för forskning och innovation ( COM(2011)0812 - C7-0009/2012 - 2011/0400(NLE) )
hänvisat till
ansvarigt utskott :
ITRE
rådgivande utskott :
ENVI, BUDG, JURI
hänvisat till
ansvarigt utskott :
ENVI
rådgivande utskott :
IMCO
hänvisat till
ansvarigt utskott :
ECON
rådgivande utskott :
JURI, IMCO
hänvisat till
ansvarigt utskott :
ECON
rådgivande utskott :
ITRE, JURI, IMCO
- Förslag till Europaparlamentets och rådets förordning om inrättande av ett instrument för stöd inför anslutningen (IPA II) ( COM(2011)0838 - C7-0491/2011 - 2011/0404(COD) )
hänvisat till
ansvarigt utskott :
AFET
rådgivande utskott :
FEMM, AGRI, EMPL, BUDG, LIBE, INTA, REGI
- Förslag till Europaparlamentets och rådets förordning om inrättande av ett europeiskt grannskapsinstrument ( COM(2011)0839 - C7-0492/2011 - 2011/0405(COD) )
hänvisat till
ansvarigt utskott :
AFET
rådgivande utskott :
DEVE, CULT, ENVI, EMPL, BUDG, ITRE, LIBE, INTA, TRAN, REGI
- Förslag till Europaparlamentets och rådets förordning om inrättande av ett finansieringsinstrument för utvecklingsarbete ( COM(2011)0840 - C7-0493/2011 - 2011/0406(COD) )
hänvisat till
ansvarigt utskott :
DEVE
rådgivande utskott :
FEMM, AFET, BUDG, LIBE, INTA
- Förslag till Europaparlamentets och rådets förordning om inrättande av ett partnerskapsinstrument för samarbete med tredjeländer ( COM(2011)0843 - C7-0495/2011 - 2011/0411(COD) )
hänvisat till
ansvarigt utskott :
INTA
rådgivande utskott :
DEVE, AFET, BUDG, ITRE
- Förslag till Europaparlamentets och rådets förordning om inrättande av ett finansieringsinstrument för främjande av demokrati och mänskliga rättigheter i hela världen ( COM(2011)0844 - C7-0496/2011 - 2011/0412(COD) )
hänvisat till
ansvarigt utskott :
AFET
rådgivande utskott :
FEMM, DEVE, BUDG
- Förslag till Europaparlamentets och rådets förordning om inrättande av ett stabilitetsinstrument ( COM(2011)0845 - C7-0497/2011 - 2011/0413(COD) )
hänvisat till
ansvarigt utskott :
AFET
rådgivande utskott :
DEVE, BUDG, INTA, ITRE
hänvisat till
ansvarigt utskott :
PECH
rådgivande utskott :
DEVE, ENVI
- Förslag till rådets beslut om inrättande av det särskilda programmet för genomförande av Horisont 2020 - ramprogrammet för forskning och innovation (2014-2020) ( COM(2011)0811 - C7-0509/2011 - 2011/0402(CNS) )
hänvisat till
ansvarigt utskott :
ITRE
rådgivande utskott :
CULT, AGRI, ENVI, EMPL, BUDG, JURI, TRAN
- Förslag till rådets beslut om ingående av avtalet mellan Amerikas förenta stater och Europeiska unionen om användning och överföring av passageraruppgifter till Förenta staternas Department of Homeland Security (17433/2011 - C7-0511/2011 - 2011/0382(NLE) )
hänvisat till
ansvarigt utskott :
LIBE
rådgivande utskott :
AFET, TRAN
- Förslag till rådets förordning om unionsstöd för stödprogrammen för kärnkraftsavveckling i Bulgarien, Litauen och Slovakien ( COM(2011)0783 - C7-0514/2011 - 2011/0363(NLE) )
hänvisat till
ansvarigt utskott :
ITRE
rådgivande utskott :
BUDG
- Förslag till rådets beslut om ingående av avtalet genom skriftväxling mellan Europeiska unionen och Ryska federationen om förvaltningen av tullkvoter på export av trä från Ryska federationen till Europeiska unionen och protokollet mellan Europeiska unionen och Ryska federationens regering om tekniska förfaringssätt enligt det avtalet (16775/2011 - C7-0515/2011 - 2011/0322(NLE) )
hänvisat till
ansvarigt utskott :
INTA
rådgivande utskott :
AGRI
- Förslag till rådets direktiv om ett gemensamt system för beskattning av räntor och royaltyer som betalas mellan närstående bolag i olika medlemsstater (omarbetning) ( COM(2011)0714 - C7-0516/2011 - 2011/0314(CNS) )
hänvisat till
ansvarigt utskott :
ECON
rådgivande utskott :
JURI
- Förslag till rådets beslut om ingående av avtalet mellan Europeiska unionen och Ryska federationens regering om handel med delar och komponenter till motorfordon mellan Europeiska unionen och Ryska federationen (16806/2011 - C7-0517/2011 - 2011/0324(NLE) )
hänvisat till
ansvarigt utskott :
INTA
rådgivande utskott :
ITRE
- Förslag till Europaparlamentets och rådets förordning om europeisk befolkningsstatistik ( COM(2011)0903 - C7-0518/2011 - 2011/0440(COD) )
hänvisat till
ansvarigt utskott :
EMPL
rådgivande utskott :
FEMM, ENVI, ECON, REGI
- Förslag till rådets beslut om ingående av avtalet genom skriftväxling mellan Europeiska unionen och Ryska federationen om införande eller höjning av exporttullar på råvaror (16827/2011 - C7-0520/2011 - 2011/0332(NLE) )
hänvisat till
ansvarigt utskott :
INTA
rådgivande utskott :
AFET
- Förslag till Europaparlamentets och rådets beslut om makroekonomiskt stöd till Kirgizistan ( COM(2011)0925 - C7-0521/2011 - 2011/0458(COD) )
hänvisat till
ansvarigt utskott :
INTA
rådgivande utskott :
AFET, BUDG
- Förslag till rådets beslut om ingående av avtalet genom skriftväxling mellan Europeiska unionen och Ryska federationens regering om bibehållande av de åtaganden om handel med tjänster som ingår i det nuvarande partnerskaps- och samarbetsavtalet mellan EU och Ryssland (16815/2011 - C7-0522/2011 - 2011/0328(NLE) )
hänvisat till
ansvarigt utskott :
INTA
rådgivande utskott :
AFET
- Förslag till Europaparlamentets och rådets beslut om ändring av avtalet om upprättande av Europeiska banken för återuppbyggnad och utveckling (EBRD) i syfte att utvidga den geografiska räckvidden för EBRD:s verksamhet till södra och östra Medelhavsområdet ( COM(2011)0905 - C7-0523/2011 - 2011/0442(COD) )
hänvisat till
ansvarigt utskott :
ECON
rådgivande utskott :
AFET, INTA
- Förslag till Europaparlamentets och rådets förordning om ändring av rådets förordning (EG) nr 774/94 om öppnande och förvaltning av vissa gemenskapstullkvoter för nötkött av hög kvalitet, griskött, fjäderfäkött, vete och blandsäd samt kli och andra restprodukter ( COM(2011)0906 - C7-0524/2011 - 2011/0445(COD) )
hänvisat till
ansvarigt utskott :
INTA
rådgivande utskott :
AGRI
3 Val av Europaparlamentets talman
Han förtydligade att ogiltiga röstsedlar inte räknas.
Talmannen utsåg sedan åtta rösträknare genom slumpmässigt urval.
Följande ledamöter utsågs:
Rita Borsellino ,
Csaba Sógor ,
Vladko Todorov Panayotov ,
Pavel Poc ,
Zoltán Bagó ,
Jarosław Kalinowski ,
Ivailo Kalfin och
Andres Perello Rodriguez .
Han informerade plenarförsamlingen om valförfarandet.
Talare:
Carl Schlyter .
Valet av talman inleddes.
ORDFÖRANDESKAP: Jerzy BUZEK
Talman
4 Val av Europaparlamentets talman
(fortsättning)
- antal röstdeltagande: 699
- blanka eller ogiltiga valsedlar: 29
- avgivna röster: 670
- absolut majoritet: 336
Valresultat:
-
Nirj Deva 142 röster
-
Martin Schulz 387 röster
-
Diana Wallis 141 röster
ORDFÖRANDESKAP: Martin SCHULZ
Talman
Talare:
Joseph Daul för PPE-gruppen,
Maria Badia i Cutchet för S&D-gruppen,
Guy Verhofstadt för ALDE-gruppen,
Rebecca Harms för Verts/ALE-gruppen,
Martin Callanan för ECR-gruppen,
Kartika Tamara Liotard för GUE/NGL-gruppen,
Nigel Farage för EFD-gruppen,
Barry Madlener , grupplös, och
José Manuel Barroso (kommissionens ordförande) .
Talmannen gjorde ett kort uttalande.
Punkten avslutades.
5
Val av Europaparlamentets vice talmän
(
tidsfrist för inlämning av nomineringar
)
På förslag av talmannen fastställdes tidsfristen för inlämning av nomineringar till kl. 18.30.
Valet skulle äga rum kl. 19.30.
ORDFÖRANDESKAP: Martin SCHULZ
Talman
6 Val av Europaparlamentets vice talmän
Talmannen meddelade att följande nomineringar av kandidater till valet av vice talmän hade lämnats in:
Alexander Alvaro ,
Roberta Angelilli ,
Isabelle Durant ,
Othmar Karas ,
Miguel Angel Martínez Martínez ,
Edward McMillan-Scott ,
Georgios Papastamkos ,
Gianni Pittella ,
Anni Podimata ,
Jacek Protasiewicz ,
László Surján ,
Indrek Tarand ,
Alejo Vidal-Quadras ,
Oldřich Vlasák och
Rainer Wieland .
Valet av vice talmän inleddes.
(Sammanträdet avbröts kl. 20.05 för rösträkning och återupptogs kl. 21.15)
ORDFÖRANDESKAP: Martin SCHULZ
Talman
7 Val av Europaparlamentets vice talmän
(fortsättning)
Talmannen redogjorde för omröstningsresultatet av första valomgången:
- antal röstdeltagande: 703
- blanka eller ogiltiga valsedlar: 14
- avgivna röster: 689
- absolut majoritet: 345
Röstfördelning, med sjunkande röstetal:
-
Alejo Vidal-Quadras : 325 röster
-
Georgios Papastamkos : 324 röster
-
Roberta Angelilli : 316 röster
-
Gianni Pittella : 306 röster
-
Othmar Karas : 305 röster
-
Miguel Angel Martínez Martínez : 276 röster
-
Anni Podimata : 269 röster
-
Rainer Wieland : 268 röster
-
Jacek Protasiewicz : 267 röster
-
László Surján : 256 röster
-
Edward McMillan-Scott : 225 röster
-
Alexander Alvaro : 199 röster
-
Oldřich Vlasák : 196 röster
-
Isabelle Durant : 182 röster
-
Indrek Tarand : 104 röster
Talmannen konstaterade att ingen kandidat erhållit absolut majoritet av rösterna och att samtliga platser därmed återstod att tillsätta.
Talmannen konstaterade att ingen av kandidaterna drog tillbaka sin kandidatur och att en andra valomgång skulle bli nödvändig.
Omröstningen genomfördes.
Talare:
Sergio Paolo Francesco Silvestris .
ORDFÖRANDESKAP: Martin SCHULZ Talman
8 Val av Europaparlamentets vice talmän
(fortsättning)
Talmannen redogjorde för omröstningsresultatet av andra valomgången:
- antal röstdeltagande: 637
- blanka eller ogiltiga valsedlar: 8
- avgivna röster: 629
- absolut majoritet: 315
Omröstningsresultat, med sjunkande röstetal:
-
-
-
-
-
-
-
-
Jacek Protasiewicz
-
Rainer Wieland
-
-
-
-
-
-
Omröstningen skulle hållas följande dag.
9 Föredragningslista för nästa sammanträde
Föredragningslistan för nästa sammanträde fastställdes ("Föredragningslista" PE 477.709/PDOJ).
10 Avslutande av sammanträdet
Sammanträdet avslutades kl. 22.45.
Klaus Welle
Martin Schulz
Generalsekreterare
Talman
NÄRVAROLISTA
Följande skrev på:
Abad
Áder
Agnew
Albertini
Albrecht
Alfano
Alfonsi
Alvaro
Alves
Andersdotter
Andreasen
Andrés Barea
Andrikienė
Angelilli
Angourakis
Antinoro
Antonescu
Antoniozzi
Arias Echeverría
Arif
Arlacchi
Arsenis
Ashworth
Atkins
Attard-Montalto
Auconie
Audy
Margrete Auken
Ayala Sender
Aylward
Ayuso
van Baalen
Bach
Badia i Cutchet
Bagó
Balčytis
Baldassarre
Balz
Balzani
Bartolozzi
Băsescu
Bastos
Batten
Bauer
Bearder
Becker
Belder
Belet
Bélier
Benarab-Attou
Bendtsen
Bennahmias
Berès
Berlato
Berlinguer
Berman
Besset
Bielan
Bilbao Barandica
Bizzotto
Blinkevičiūtė
Bloom
Bodu
Böge
Bokros
Bonsignore
Borghezio
Borsellino
Borys
Boştinaru
Boulland
Bové
Bowles
Bozkurt
Bradbourn
Brantner
Bratkowski
Brepoels
Březina
Brok
Brons
Brzobohatá
Bullmann
Buşoi
Busuttil
Bütikofer
Buzek
Cabrnoch
Cadec
Callanan
van de Camp
Campbell Bannerman
Cancian
Canfin
Capoulas Santos
Caronna
Carvalho
Cashman
Casini
Caspary
Castex
del Castillo Vera
Cavada
Cercas
Češková
Chatzimarkakis
Chichester
Childers
Chountis
Christensen
Claeys
Clark
Cochet
Coelho
Cofferati
Colman
Comi
Corazza Bildt
Cornelissen
Correa Zamora
Correia De Campos
Cortés Lastra
Silvia Costa
Cozzolino
Cramer
Creţu
Creutzmann
Crocetta
Cronberg
Cuschieri
Cutaş
Cymański
Czarnecki
Frédéric Daerden
van Dalen
Dăncilă
Danellis
Danjean
Dantin
(The Earl of) Dartmouth
Dati
Daul
David
Davies
De Angelis
De Backer
De Castro
Dehaene
De Keyser
Delli
Delvaux
De Mita
De Rossa
de Sarnez
Désir
Deß
Deutsch
Deva
De Veyrac
Díaz de Mera García Consuegra
Dodds
Domenici
Donskis
Dorfmann
Droutsas
Duff
Durant
Dušek
Ehler
Ehrenhauser
Eickhout
El Khadraoui
Elles
Enciu
Engel
Eppink
Ernst
Ertug
Estaràs Ferragut
Estrela
Evans
Fajmon
Fajon
Falbr
Färm
Feio
Ferber
Fernandes
Elisa Ferreira
João Ferreira
Fidanza
Figueiredo
Fisas Ayxela
Fjellner
Flašíková Beňová
Flautre
Fleckenstein
Florenz
Fontana
Ford
Foster
Fox
Franco
Gahler
Gál
Gallagher
Gallo
Gáll-Pelcz
Garcés Ramón
García-Hierro Caraballo
García Pérez
Gardiazábal Rubial
Gardini
Gargani
Garriga Polledo
Gauzès
Gebhardt
Geier
Gerbrandy
Geringer de Oedenberg
Giannakou
Giegold
Gierek
Girling
Glante
Glattfelder
Godmanis
Goebbels
Goerens
Gollnisch
Gomes
Göncz
Goulard
de Grandes Pascual
Gräßle
Grech
Grelier
Grèze
Griesbeck
Griffin
Gróbarczyk
Groote
Grosch
Grossetête
Grzyb
Gualtieri
Guerrero Salom
Guillaume
Gurmai
Gustafsson
Gutiérrez-Cortines
Gutiérrez Prieto
Gyürk
Hadjigeorgiou
Häfner
Haglund
Fiona Hall
Händel
Handzlik
Hankiss
Hannan
Harbour
Harkin
Hartong
Hassi
Haug
Häusling
Hedh
Helmer
Hénin
Herczog
Herranz García
Hibner
Higgins
Nadja Hirsch
Hoang Ngoc
Hohlmeier
Hökmark
Honeyball
Hortefeux
Howitt
Danuta Maria Hübner
Hudghton
Hughes
Hyusmenova
Iacolino
Ibrisagic
Ilchev
Imbrasas
in 't Veld
Iotova
Iovine
Irigoyen Pérez
Itälä
Iturgaiz Angulo
Ivan
Ivanova
Jaakonsaari
Jäätteenmäki
Jadot
Jahr
Járóka
Jazłowiecka
Jędrzejewska
Jeggle
Jensen
Jiménez-Becerril Barrio
Johansson
Joly
de Jong
Jordan
Jørgensen
Juvin
Kacin
Kaczmarek
Kadenbach
Kalfin
Kalinowski
Kalniete
Kamall
Kamiński
Kammerevert
Karas
Karim
Kariņš
Kasoulides
Kastler
Kazak
Kelam
Kelly
Kiil-Nielsen
Kirilov
Kirkhope
Klaß
Kleva
Klinz
Klute
Koch
Koch-Mehrin
Kohlíček
Kolarska-Bobińska
Koppa
Korhola
Kósa
Köstinger
Koumoutsakos
Béla Kovács
Kovatchev
Kowal
Kozlík
Kozłowski
Kožušník
Krahmer
Kratsa-Tsagaropoulou
Krehl
Kreissl-Dörfler
Kuhn
Kukan
Kurski
Lamassoure
Lambert
Lamberts
Lambsdorff
Landsbergis
Lange
de Lange
Langen
La Via
Le Brun
Lechner
Le Foll
Le Grip
Legutko
Lehne
Le Hyaric
Leichtfried
Leinen
Lepage
Jean-Marie Le Pen
Marine Le Pen
Liberadzki
Lichtenberger
Liese
Liotard
Lisek
Lochbihler
Løkkegaard
Lope Fontagné
López Aguilar
López-Istúriz White
Lösing
Lövin
Ludford
Ludvigsson
Luhan
Łukacijewska
Lulling
Lunacek
Lynne
Lyon
McAvan
McCarthy
McClarkin
McGuinness
McIntyre
McMillan-Scott
Macovei
Madlener
Malinov
Manders
Mănescu
Maňka
Mann
Manner
Marcinkiewicz
Marinescu
David Martin
Hans-Peter Martin
Martínez Martínez
Masip Hidalgo
Maštálka
Mastella
Matera
Mathieu
Matias
Mato Adrover
Matula
Mauro
Mavronikolas
Mayer
Mayor Oreja
Mazej Kukovič
Mazzoni
Meissner
Mélenchon
Menéndez del Valle
Merkies
Messerschmidt
Mészáros
Meyer
Louis Michel
Migalski
Mikolášik
Milana
Millán Mon
Miranda
Mirsky
Mitchell
Mölzer
Moraes
Moreira
Morganti
Morin-Chartier
Morkūnaitė-Mikulėnienė
Morvai
Motti
Mulder
Muñiz De Urquiza
Murphy
Muscardini
Naranjo Escobar
Nattrass
Nedelcheva
Neuser
Neveďalová
Newton Dunn
Neynsky
Neyts-Uyttebroeck
Nicholson
Nicolai
Niculescu
Niebler
Nilsson
van Nistelrooij
Nitras
Nuttall
Obermayr
Obiols
Ojuland
Olbrycht
Olejniczak
Omarjee
Oomen-Ruijten
Ortiz Vilella
Őry
Ouzký
Oviir
Pack
Padar
Paksas
Paleckis
Paliadeli
Pallone
Panayotov
Panzeri
Papadopoulou
Papanikolaou
Papastamkos
Pargneaux
Parvanova
Paşcu
Paška
Patrão Neves
Patriciello
Paulsen
Peillon
Perello Rodriguez
Peterle
Pieper
Pietikäinen
Piotrowski
Pirillo
Pirker
Pittella
Plumb
Poc
Podimata
Ponga
Poręba
Portas
Posselt
Pöttering
Poupakis
Preda
Prendergast
Prodi
Protasiewicz
Proust
Provera
Quisthoudt-Rowohl
Rangel
Ransdorf
Rapkay
Rapti
Regner
Reimers
Remek
Repo
Reul
Riera Madurell
Ries
Rinaldi
Riquet
Rivasi
Rivellini
Roatta
Rochefort
Rodust
Rohde
Roithová
Romero López
Romeva i Rueda
Ronzulli
Rosbach
Rossi
Roth-Behrendt
Rouček
Rübig
Rubiks
Šadurskis
Saïfi
Salafranca Sánchez-Neyra
Salatto
Salavrakos
Salvini
Sánchez Presedo
Sanchez-Schmid
Sârbu
Sargentini
Sartori
Saryusz-Wolski
Sassoli
Saudargas
Savisaar-Toomast
Schaake
Schaldemose
Schlyter
Olle Schmidt
Schnellhardt
Schnieber-Jastram
Scholz
Schöpflin
Schroedter
Martin Schulz
Werner Schulz
Schwab
Scicluna
Scurria
Sedó i Alabart
Seeber
Sehnalová
Senyszyn
Serracchiani
Severin
Siekierski
Silvestris
Simon
Simpson
Sinclaire
Sippel
Siwiec
Skinner
Skrzydlewska
Skylakakis
Smith
Smolková
Sógor
Sommer
Søndergaard
Sonik
Sosa Wagner
Speroni
Stadler
Staes
Stassen
Šťastný
Stavrakakis
Steinruck
Stevenson
Stihler
van der Stoep
Stolojan
Strejček
Striffler
Surján
Susta
Svensson
Swinburne
Swoboda
Szájer
Szegedi
Szymański
Tabajdi
Takkula
Tănăsescu
Tannock
Tarabella
Tarand
Tatarella
Tavares
Taylor
Teixeira
Terho
Thein
Theocharous
Theurer
Thomsen
Thun und Hohenstein
Thyssen
Ţicău
Tirolien
Toia
Tőkés
Tomaševski
Tošenovský
Trautmann
Trematerra
Tremopoulos
Tremosa i Balcells
Triantaphyllides
Trüpel
Trzaskowski
Tsoukalas
Turmes
Turunen
Tzavela
Uggias
Ulmer
Ulvskog
Ungureanu
Urutchev
Uspaskich
Vadim Tudor
Vaidere
Vajgl
Vălean
Van Brempt
Vanhecke
Van Orden
Vattimo
Vaughan
Vergiat
Vergnaud
Verheyen
Vidal-Quadras
Vigenin
de Villiers
Vlasák
Vlasto
Voss
Wallis
Watson
Henri Weber
Manfred Weber
Renate Weber
Weidenholzer
Weiler
Weisgerber
Werthmann
Westlund
Westphal
Wieland
Wikström
Willmott
Wils
Hermann Winkler
Iuliu Winkler
Włosowicz
Wojciechowski
Wortmann-Kool
Yáñez-Barnuevo García
Yannakoudakis
Záborská
Zahradil
Zala
Zalba Bidegain
Zalewski
Zanicchi
Zanoni
Zasada
Ždanoka
Zeller
Zemke
Zijlstra
Zīle
Zimmer
Ziobro
Zver
Zwiefka
Bilaga 1 - Val av Europaparlamentets talman
FÖRTECKNING ÖVER LEDAMÖTER SOM DELTOG I OMRÖSTNINGEN
Áder, Agnew, Albertini, Albrecht, Alfano, Alfonsi, Alvaro, Alves, Andreasen, Andrés Barea, Andrikienė, Angelilli, Angourakis, Antinoro, Antonescu, Arif, Arlacchi, Arsenis, Ashworth, Atkins, Attard-Montalto, Auconie, Audy, Auken, Ayala Sender, Aylward, Ayuso, van Baalen, Bach, Badia i Cutchet, Bagó, Balčytis, Baldassarre, Balz, Balzani, Bartolozzi, Băsescu, Bastos, Batten, Bauer, Bearder, Becker, Belder, Belet, Bélier, Benarab-Attou, Bendtsen, Bennahmias, Berès, Berlato, Berlinguer, Berman, Besset, Bielan, Bilbao Barandica, Bizzotto, Blinkevičiūtė, Bloom, Bodu, Böge, Bokros, Bonsignore, Borghezio, Borsellino, Borys, Boştinaru, Boulland, Bové, Bowles, Bozkurt, Bradbourn, Brantner, Bratkowski, Brepoels, Březina, Brok, Brons, Brzobohatá, Bullmann, Buşoi, Busuttil, Bütikofer, Buzek, Cabrnoch, Cadec, Callanan, van de Camp, Cancian, Canfin, Capoulas Santos, Caronna, Carvalho, Cashman, Casini, Caspary, Castex, del Castillo Vera, Cavada, Cercas, Češková, Chatzimarkakis, Chichester, Childers, Chountis, Christensen, Claeys, Clark, Cochet, Coelho, Cofferati, Cohn-Bendit, Colman, Comi, Corazza Bildt, Cornelissen, Correa Zamora , Correia De Campos, Cortés Lastra, Silvia Costa, Cozzolino, Cramer, Creţu, Creutzmann, Crocetta, Cronberg, Cuschieri, Cutaş, Cymański, Czarnecki, Frédéric Daerden, van Dalen, Dăncilă, Danellis, Danjean, Dantin, Dati, Daul, David, Davies, De Angelis, De Backer, De Castro, Dehaene, De Keyser, Delli, Delvaux, De Mita, De Rossa, De Sarnez, Désir, Deß, Deutsch, Deva, De Veyrac, Díaz de Mera García Consuegra, Dodds, Domenici, Donskis, Dorfmann, Droutsas, Duff, Durant, Dušek, Ehler, Ehrenhauser, Eickhout, El Khadraoui, Elles, Enciu, Engel, Eppink, Ernst, Ertug, Estaràs Ferragut, Estrela, Evans, Fajmon, Fajon, Falbr, Farage, Färm, Feio, Ferber, Fernandes, Elisa Ferreira, João Ferreira, Fidanza, Figueiredo, Fisas Ayxela, Fjellner, Flašíková Beňová, Flautre, Fleckenstein, Florenz, Fontana, Ford, Fox, Gahler, Gál, Gallagher, Gallo, Gáll-Pelcz, Garcés Ramón, García-Hierro Caraballo, Gardiazábal Rubial, Gardini, Gargani, Garriga Polledo, Gauzès, Gebhardt, Geier, Gerbrandy, Geringer de Oedenberg, Giannakou, Giegold, Gierek, Girling, Glante, Glattfelder, Godmanis, Goebbels, Goerens, Gollnisch, Gomes, Göncz, Goulard, de Grandes Pascual, Gräßle, Grech, Grelier, Grèze, Griesbeck, Griffin, Gróbarczyk, Groote, Grosch, Grossetête, Grzyb, Gualtieri, Guerrero Salom, Guillaume, Gurmai, Gustafsson, Gutiérrez-Cortines, Gutiérrez Prieto, Gyürk, Hadjigeorgiou, Häfner, Haglund, Fiona Hall, Händel, Handzlik, Hankiss, Hannan, Harbour, Harkin, Harms, Hartong, Hassi, Haug, Häusling, Hedh, Helmer, Hénin, Herczog, Herranz García, Hibner, Higgins, Nadja Hirsch, Hoang Ngoc, Hohlmeier, Hökmark, Honeyball, Hortefeux, Danuta Maria Hübner, Hughes, Hyusmenova, Iacolino, Ibrisagic, Ilchev, Imbrasas, in 't Veld, Iotova, Iovine, Irigoyen Pérez, Itälä, Iturgaiz Angulo, Ivan, Ivanova, Jaakonsaari, Jäätteenmäki, Jadot, Jahr, Járóka, Jazłowiecka, Jeggle, Jensen, Jiménez-Becerril Barrio, Johansson, Joly, de Jong, Jordan Cizelj, Jørgensen, Juvin, Kacin, Kaczmarek, Kadenbach, Kalfin, Kalinowski, Kalniete, Kamall, Kamiński, Kammerevert, Karas, Karim, Kariņš, Kasoulides, Kastler, Kazak, Kelam, Kelly, Kiil-Nielsen, Kirilov, Kirkhope, Klaß, Kleva, Klinz, Klute, Koch, Koch-Mehrin, Kohlíček, Kolarska-Bobińska, Koppa, Korhola, Kósa, Köstinger, Koumoutsakos, Kovatchev, Kowal, Kozlík, Kozłowski, Kožušník, Krahmer, Kratsa-Tsagaropoulou, Krehl, Kreissl-Dörfler, Kuhn, Kukan, Kurski, Lamassoure , Lambert, Lamberts, Lambsdorff, Landsbergis, Lange, Langen, La Via, Lechner, Le Foll, Le Grip, Legutko, Lehne, Le Hyaric, Leichtfried, Leinen, Lepage, Jean-Marie Le Pen, Liberadzki, Lichtenberger, Liese, Liotard, Lisek, Lochbihler, Løkkegaard, Lope Fontagné, López Aguilar, López-Istúriz White, Lösing, Lövin, Ludford, Ludvigsson, Łukacijewska, Lulling, Lunacek, Lynne, Lyon, McAvan, McCarthy, McClarkin, McGuinness, McIntyre, McMillan-Scott, Macovei, Madlener, Malinov, Manders, Mănescu, Maňka, Mann, Manner, Marcinkiewicz, Marinescu, David Martin, Hans-Peter Martin, Martínez Martínez, Masip Hidalgo, Maštálka, Mastella, Matera, Mathieu, Matias, Mato Adrover, Matula, Mauro, Mavronikolas, Mayer, Mayor Oreja, Mazej Kukovič , Mazzoni, Meissner, Menéndez del Valle, Merkies, Messerschmidt, Mészáros, Louis Michel, Migalski, Mikolášik, Milana, Millán Mon, Miranda , Mirsky, Mitchell, Mölzer, Moraes, Moreira, Morin-Chartier, Morkūnaitė-Mikulėnienė, Mulder, Muñiz De Urquiza, Murphy, Muscardini, Naranjo Escobar, Nattrass, Nedelcheva, Neuser, Neveďalová, Newton Dunn, Neynsky, Neyts-Uyttebroeck, Nicholson, Nicolai, Niculescu, Niebler, Nilsson, van Nistelrooij, Nitras, Obiols, Ojuland, Olbrycht, Olejniczak, Omarjee , Oomen-Ruijten, Ortiz Vilella, Őry, Ouzký, Oviir, Pack, Padar, Paleckis, Paliadeli, Pallone, Panayotov, Panzeri, Papadopoulou, Papanikolaou, Papastamkos, Pargneaux, Parvanova, Paşcu, Paška, Patrão Neves, Patriciello, Paulsen, Peillon, Perello Rodriguez, Peterle, Pieper, Pietikäinen, Piotrowski, Pirillo, Pirker, Pittella , Plumb, Poc, Podimata, Ponga, Poręba, Portas, Posselt, Pöttering, Poupakis, Preda, Prendergast, Prodi, Protasiewicz, Proust, Provera, Quisthoudt-Rowohl, Rangel, Rapkay, Rapti, Regner, Reimers, Remek, Repo, Reul, Riera Madurell, Ries, Rinaldi, Riquet, Rivasi, Rivellini, Roatta, Rodust, Rohde, Roithová, Romero López, Romeva i Rueda, Ronzulli, Rosbach, Rossi, Roth-Behrendt, Rouček, Rübig, Rubiks, Šadurskis, Saïfi, Salafranca Sánchez-Neyra, Salatto, Salavrakos, Sánchez Presedo, Sanchez-Schmid, Sârbu, Sargentini, Sartori, Saryusz-Wolski, Sassoli, Saudargas, Savisaar-Toomast, Schaake, Schaldemose, Schlyter, Olle Schmidt, Schnellhardt, Schnieber-Jastram, Scholz, Schöpflin, Schroedter, Martin Schulz, Werner Schulz, Schwab, Scicluna, Scurria, Sedó i Alabart, Seeber, Sehnalová, Senyszyn, Serracchiani, Severin, Siekierski, Silvestris, Simon, Simpson, Sippel, Siwiec, Skinner, Skrzydlewska, Skylakakis, Smith, Smolková, Sógor, Sommer, Søndergaard, Sonik, Sosa Wagner, Speroni, Stadler, Staes, Stassen, Šťastný, Stavrakakis, Steinruck, Stevenson, Stihler, van der Stoep, Stolojan, Strejček, Striffler, Surján, Susta, Svensson, Swinburne, Swoboda, Szájer, Szegedi, Szymański, Tabajdi, Takkula, Tănăsescu, Tannock, Tarabella, Tarand, Tatarella, Tavares, Taylor, Teixeira, Terho, Thein, Theocharous, Theurer, Thomsen, Thun und Hohenstein, Thyssen, Ţicău, Tirolien, Toia, Tőkés, Tomaševski, Tošenovský, Trautmann, Trematerra, Tremosa i Balcells, Triantaphyllides, Trüpel, Trzaskowski, Tsoukalas, Turmes, Turunen, Tzavela, Uggias, Ulmer, Ulvskog, Ungureanu, Urutchev, Vadim Tudor, Vaidere, Vajgl, Vălean, Van Brempt, Vanhecke, Van Orden, Vattimo, Vaughan, Vergnaud, Verheyen, Verhofstadt, Vidal-Quadras , Vigenin, de Villiers, Vlasák, Vlasto, Voss, Wallis, Watson, Henri Weber, Manfred Weber, Renate Weber, Weidenholzer, Weiler, Weisgerber, Werthmann, Westlund, Westphal, Wieland, Wikström, Willmott, Wils, Hermann Winkler, Iuliu Winkler, Włosowicz, Wojciechowski, Wortmann-Kool, Yáñez-Barnuevo García, Yannakoudakis, Záborská, Zahradil, Zala, Zalba Bidegain, Zanicchi, Zanoni, Zasada, Ždanoka, Zeller, Zemke, Zijlstra, Zīle, Zimmer, Zver, Zwiefka
Bilaga 2 - Val av Europaparlamentets vice talmän
VAL AV EUROPAPARLAMENTETS VICE TALMÄN (första valomgången)
FÖRTECKNING ÖVER LEDAMÖTER SOM DELTOG I OMRÖSTNINGEN
Áder, Albertini, Albrecht, Alfano, Alfonsi, Alvaro, Alves, Andersdotter, Andreasen, Andrés Barea, Andrikienė, Angelilli, Angourakis, Antinoro, Antonescu, Antoniozzi, Arias Echeverría, Arif, Arlacchi, Arsenis, Ashworth, Atkins, Attard-Montalto, Auconie, Audy, Auken, Ayala Sender, Aylward, Ayuso, van Baalen, Bach, Badia i Cutchet, Bagó, Balčytis, Baldassarre, Balz, Balzani, Bartolozzi, Băsescu, Bastos, Bauer, Bearder, Becker, Belder, Belet, Bélier, Benarab-Attou, Bendtsen, Bennahmias, Berès, Berlato, Berlinguer, Berman, Besset, Bielan, Bilbao Barandica, Bizzotto, Blinkevičiūtė, Bodu, Böge, Bokros, Bonsignore, Borghezio, Borsellino, Borys, Boştinaru, Boulland, Bové, Bowles, Bozkurt, Bradbourn, Bratkowski, Brepoels, Březina, Brok, Brons, Brzobohatá, Bullmann, Busuttil, Bütikofer, Buzek, Cabrnoch, Cadec, Callanan, van de Camp, Campbell Bannerman, Cancian, Capoulas Santos, Caronna, Carvalho, Cashman, Casini, Caspary, Castex, del Castillo Vera, Cavada, Cercas, Češková, Chatzimarkakis, Chichester, Childers, Chountis, Christensen, Claeys, Cochet, Coelho, Cofferati, Cohn-Bendit, Colman, Comi, Corazza Bildt, Cornelissen, Correa Zamora , Correia De Campos, Cortés Lastra, Silvia Costa, Cozzolino, Cramer, Creţu, Creutzmann, Crocetta, Cronberg, Cuschieri, Cutaş, Cymański, Czarnecki, Frédéric Daerden, van Dalen, Dăncilă, Danellis, Dantin, Daul, David, Davies, De Angelis, De Backer, De Castro, Dehaene, De Keyser, Delli, Delvaux, De Mita, De Rossa, De Sarnez, Deß, Deutsch, Deva, De Veyrac, Díaz de Mera García Consuegra, Dodds, Domenici, Donskis, Dorfmann, Droutsas, Duff, Durant, Dušek, Ehler, Ehrenhauser, Eickhout, El Khadraoui, Elles, Enciu, Engel, Eppink, Ernst, Ertug, Estaràs Ferragut, Estrela, Evans, Fajmon, Fajon, Falbr, Farage, Färm, Feio, Ferber, Fernandes, Elisa Ferreira, João Ferreira, Fidanza, Figueiredo, Fisas Ayxela, Fjellner, Flašíková Beňová, Flautre, Fleckenstein, Fontana, Ford, Foster, Fox, Franco, Gahler, Gál, Gallagher, Gallo, Gáll-Pelcz, Garcés Ramón, García-Hierro Caraballo, García Pérez, Gardiazábal Rubial, Gardini, Gargani, Garriga Polledo, Gauzès, Gebhardt, Geier, Gerbrandy, Geringer de Oedenberg, Giannakou, Giegold, Gierek, Girling, Glante, Glattfelder, Godmanis, Goebbels, Goerens, Gomes, Göncz, Goulard, de Grandes Pascual, Grech, Grelier, Grèze, Griesbeck, Griffin, Gróbarczyk, Groote, Grosch, Grossetête, Grzyb, Gualtieri, Guerrero Salom, Guillaume, Gurmai, Gustafsson, Gutiérrez-Cortines, Gutiérrez Prieto, Gyürk, Hadjigeorgiou, Häfner, Haglund, Fiona Hall, Händel, Handzlik, Hankiss, Hannan, Harbour, Harkin, Harms, Hartong, Hassi, Haug, Häusling, Hedh, Helmer, Hénin, Herczog, Herranz García, Hibner, Higgins, Nadja Hirsch, Hoang Ngoc, Hohlmeier, Hökmark, Honeyball, Hortefeux, Howitt, Danuta Maria Hübner, Hudghton, Hughes, Hyusmenova, Iacolino, Ibrisagic, Ilchev, Imbrasas, in 't Veld, Iotova, Iovine, Irigoyen Pérez, Itälä, Iturgaiz Angulo, Ivan, Ivanova, Jaakonsaari, Jäätteenmäki, Jadot, Jahr, Járóka, Jazłowiecka, Jędrzejewska, Jeggle, Jensen, Jiménez-Becerril Barrio, Johansson, Joly, de Jong, Jordan Cizelj, Jørgensen, Juvin, Kacin, Kaczmarek, Kadenbach, Kalfin, Kalinowski, Kalniete, Kamall, Kamiński, Kammerevert, Karas, Karim, Kariņš, Kasoulides, Kastler, Kazak, Kelam, Kelly, Kiil-Nielsen, Kirilov, Kirkhope, Klaß, Kleva, Klinz, Klute, Koch, Koch-Mehrin, Kohlíček, Kolarska-Bobińska, Koppa, Korhola, Kósa, Köstinger, Koumoutsakos, Kovatchev, Kowal, Kozlík, Kozłowski, Kožušník, Krahmer, Kratsa-Tsagaropoulou, Krehl, Kreissl-Dörfler, Kuhn, Kukan, Kurski, Lamassoure , Lambert, Lamberts, Lambsdorff, Landsbergis, Lange, de Lange, Langen, La Via, Le Brun, Lechner, Legutko, Lehne, Le Hyaric, Leichtfried, Leinen, Liberadzki, Lichtenberger, Liese, Liotard, Lisek, Lochbihler, Løkkegaard, Lope Fontagné, López Aguilar, López-Istúriz White, Lösing, Lövin, Ludford, Ludvigsson, Luhan, Lulling, Lunacek, Lynne, Lyon, McAvan, McCarthy, McClarkin, McGuinness, McIntyre, McMillan-Scott, Macovei, Madlener, Malinov, Mănescu, Maňka, Mann, Manner, Marcinkiewicz, Marinescu, David Martin, Hans-Peter Martin, Martínez Martínez, Masip Hidalgo, Maštálka, Mastella, Matera, Mathieu, Matias, Mato Adrover, Matula, Mauro, Mavronikolas, Mayer, Mayor Oreja, Mazej Kukovič , Mazzoni, Meissner, Mélenchon, Menéndez del Valle, Merkies, Messerschmidt, Mészáros, Meyer, Louis Michel, Migalski, Mikolášik, Milana, Millán Mon, Miranda , Mirsky, Mitchell, Mölzer, Moraes, Moreira, Morganti, Morin-Chartier, Morkūnaitė-Mikulėnienė, Morvai, Motti, Mulder, Muñiz De Urquiza, Murphy, Muscardini, Naranjo Escobar, Nattrass, Nedelcheva, Neuser, Neveďalová, Newton Dunn, Neynsky, Neyts-Uyttebroeck, Nicholson, Nicolai, Niculescu, Niebler, Nilsson, van Nistelrooij, Nitras, Obermayr, Ojuland, Olbrycht, Olejniczak, Omarjee , Oomen-Ruijten, Ortiz Vilella, Őry, Ouzký, Oviir, Pack, Padar, Paksas, Paleckis, Paliadeli, Pallone, Panayotov, Panzeri, Papadopoulou, Papanikolaou, Papastamkos, Pargneaux, Parvanova, Paşcu, Paška, Patrão Neves, Patriciello, Paulsen, Peillon, Perello Rodriguez, Peterle, Pieper, Pietikäinen, Piotrowski, Pirillo, Pirker, Pittella , Plumb, Poc, Podimata, Ponga, Poręba, Portas, Posselt, Pöttering, Poupakis, Preda, Prendergast, Prodi, Protasiewicz, Proust, Provera, Quisthoudt-Rowohl, Rangel, Ransdorf, Rapkay, Rapti, Regner, Reimers, Remek, Repo, Reul, Riera Madurell, Ries, Rinaldi, Riquet, Rivasi, Rivellini, Roatta, Rodust, Rohde, Roithová, Romero López, Romeva i Rueda, Ronzulli, Rosbach, Rossi, Roth-Behrendt, Rouček, Rübig, Rubiks, Šadurskis, Saïfi, Salafranca Sánchez-Neyra, Salatto, Salavrakos, Salvini, Sánchez Presedo, Sanchez-Schmid, Sârbu, Sargentini, Sartori, Saryusz-Wolski, Sassoli, Saudargas, Savisaar-Toomast, Schaake, Schaldemose, Schlyter, Olle Schmidt, Schnellhardt, Schnieber-Jastram, Scholz, Schöpflin, Schroedter, Martin Schulz, Werner Schulz, Schwab, Scicluna, Scurria, Sedó i Alabart, Seeber, Sehnalová, Senyszyn, Serracchiani, Severin, Siekierski, Silvestris, Simon, Simpson, Sinclaire, Sippel, Siwiec, Skinner, Skrzydlewska, Skylakakis, Smith, Smolková, Sógor, Sommer, Søndergaard, Sonik, Sosa Wagner, Speroni, Stadler, Staes, Stassen, Šťastný, Stavrakakis, Steinruck, Stevenson, Stolojan, Strejček, Striffler, Surján, Susta, Svensson, Swinburne, Swoboda, Szájer, Szegedi, Szymański, Tabajdi, Takkula, Tănăsescu, Tannock, Tarabella, Tarand, Tatarella, Tavares, Taylor, Teixeira, Terho, Thein, Theocharous, Theurer, Thomsen, Thun und Hohenstein, Thyssen, Ţicău, Tirolien, Toia, Tőkés, Tomaševski, Tošenovský, Trautmann, Tremopoulos, Tremosa i Balcells, Triantaphyllides, Trüpel, Trzaskowski, Tsoukalas, Turmes, Turunen, Tzavela, Uggias, Ulmer, Ulvskog, Ungureanu, Urutchev, Uspaskich, Vadim Tudor, Vaidere, Vajgl, Vălean, Van Brempt, Vanhecke, Van Orden, Vattimo, Vaughan, Vergiat, Vergnaud, Verheyen, Verhofstadt, Vidal-Quadras , Vigenin, Vlasák, Vlasto, Voss, Wallis, Watson, Henri Weber, Manfred Weber, Renate Weber, Weidenholzer, Weiler, Weisgerber, Werthmann, Westlund, Westphal, Wieland, Wikström, Willmott, Wils, Hermann Winkler, Iuliu Winkler, Włosowicz, Wojciechowski, Wortmann-Kool, Yáñez-Barnuevo García, Yannakoudakis, Záborská, Zahradil, Zala, Zalba Bidegain, Zalewski, Zanicchi, Zanoni, Zasada, Ždanoka, Zeller, Zemke, Zijlstra, Zīle, Zimmer, Ziobro, Zver, Zwiefka
VAL AV EUROPAPARLAMENTETS VICE TALMÄN (andra valomgången)
FÖRTECKNING ÖVER LEDAMÖTER SOM DELTOG I OMRÖSTNINGEN
Áder, Albertini, Albrecht, Alfano, Alfonsi, Alvaro, Alves, Andersdotter, Andrés Barea, Andrikienė, Angelilli, Angourakis, Antinoro, Antonescu, Antoniozzi, Arias Echeverría, Arif, Arlacchi, Arsenis, Attard-Montalto, Auconie, Audy, Auken, Ayala Sender, Aylward, Ayuso, van Baalen, Bach, Badia i Cutchet, Bagó, Baldassarre, Balz, Balzani, Bartolozzi, Băsescu, Bastos, Bauer, Bearder, Becker, Belder, Belet, Bélier, Benarab-Attou, Bendtsen, Berlato, Berlinguer, Berman, Besset, Bielan, Bilbao Barandica, Bizzotto, Blinkevičiūtė, Bodu, Böge, Bokros, Bonsignore, Borghezio, Borsellino, Borys, Boştinaru, Boulland, Bové, Bowles, Bozkurt, Bratkowski, Brepoels, Březina, Brok, Brzobohatá, Bullmann, Buşoi, Busuttil, Bütikofer, Buzek, Cabrnoch, Cadec, Callanan, van de Camp, Campbell Bannerman, Cancian, Canfin, Capoulas Santos, Caronna, Carvalho, Cashman, Caspary, Castex, del Castillo Vera, Cavada, Cercas, Češková, Chatzimarkakis, Childers, Christensen, Cochet, Coelho, Cofferati, Cohn-Bendit, Comi, Corazza Bildt, Cornelissen, Correa Zamora , Correia De Campos, Cortés Lastra, Silvia Costa, Cozzolino, Cramer, Creţu, Creutzmann, Crocetta, Cronberg, Cuschieri, Cutaş, Cymański, Czarnecki, Frédéric Daerden, van Dalen, Dăncilă, Danellis, Dantin, Daul, David, Davies, De Angelis, De Backer, De Castro, Dehaene, De Keyser, Delli, Delvaux, De Rossa, Deß, Deutsch, De Veyrac, Díaz de Mera García Consuegra, Dodds, Domenici, Donskis, Dorfmann, Droutsas, Duff, Durant, Dušek, Ehler, Ehrenhauser, El Khadraoui, Elles, Enciu, Engel, Eppink, Ernst, Ertug, Estaràs Ferragut, Estrela, Evans, Fajmon, Fajon, Falbr, Färm, Feio, Ferber, Fernandes, João Ferreira, Fidanza, Fisas Ayxela, Fjellner, Flašíková Beňová, Fleckenstein, Fontana, Ford, Foster, Fox, Franco, Gahler, Gál, Gallagher, Gallo, Gáll-Pelcz, Garcés Ramón, García-Hierro Caraballo, García Pérez, Gardiazábal Rubial, Gardini, Gargani, Garriga Polledo, Gauzès, Gebhardt, Geier, Gerbrandy, Geringer de Oedenberg, Giannakou, Giegold, Gierek, Girling, Glante, Glattfelder, Godmanis, Goebbels, Goerens, Gomes, Göncz, Goulard, de Grandes Pascual, Grech, Grelier, Grèze, Gróbarczyk, Groote, Grossetête, Grzyb, Gualtieri, Guerrero Salom, Guillaume, Gurmai, Gustafsson, Gutiérrez-Cortines, Gutiérrez Prieto, Gyürk, Häfner, Haglund, Fiona Hall, Händel, Handzlik, Hankiss, Hannan, Harbour, Harkin, Harms, Hassi, Haug, Häusling, Hedh, Helmer, Herczog, Herranz García, Hibner, Higgins, Nadja Hirsch, Hoang Ngoc, Hohlmeier, Hökmark, Hortefeux, Howitt, Danuta Maria Hübner, Hyusmenova, Iacolino, Ilchev, in 't Veld, Iotova, Iovine, Irigoyen Pérez, Itälä, Iturgaiz Angulo, Ivan, Ivanova, Jaakonsaari, Jäätteenmäki, Jadot, Jahr, Járóka, Jazłowiecka, Jędrzejewska, Jeggle, Jensen, Jiménez-Becerril Barrio, Johansson, Joly, Jordan Cizelj, Jørgensen, Juvin, Kacin, Kaczmarek, Kadenbach, Kalfin, Kalinowski, Kamall, Kammerevert, Karas, Karim, Kariņš, Kasoulides, Kastler, Kazak, Kelam, Kelly, Kiil-Nielsen, Kirilov, Kirkhope, Klaß, Kleva, Klute, Koch, Koch-Mehrin, Kohlíček, Kolarska-Bobińska, Koppa, Korhola, Kósa, Köstinger, Koumoutsakos, Béla Kovács, Kovatchev, Kowal, Kozlík, Kozłowski, Kožušník, Krahmer, Kratsa-Tsagaropoulou, Krehl, Kreissl-Dörfler, Kuhn, Kukan, Kurski, Lamassoure , Lambert, Lamberts, Lambsdorff, Landsbergis, Lange, de Lange, Langen, La Via, Le Brun, Lechner, Le Foll, Legutko, Lehne, Leichtfried, Leinen, Liberadzki, Lichtenberger, Liese, Liotard, Lisek, Lochbihler, Løkkegaard, Lope Fontagné, López Aguilar, López-Istúriz White, Lösing, Lövin, Ludford, Ludvigsson, Luhan, Lulling, Lunacek, Lynne, Lyon, McAvan, McCarthy, McClarkin, McGuinness, McIntyre, McMillan-Scott, Macovei, Madlener, Malinov, Manders, Mănescu, Maňka, Mann, Manner, Marcinkiewicz, Marinescu, David Martin, Martínez Martínez, Maštálka, Mastella, Matera, Mathieu, Matias, Mato Adrover, Matula, Mauro, Mavronikolas, Mayer, Mayor Oreja, Mazej Kukovič , Mazzoni, Meissner, Menéndez del Valle, Merkies, Mészáros, Louis Michel, Migalski, Mikolášik, Milana, Millán Mon, Miranda , Mirsky, Mitchell, Moraes, Moreira, Morganti, Morin-Chartier, Morkūnaitė-Mikulėnienė, Motti, Mulder, Muñiz De Urquiza, Murphy, Muscardini, Naranjo Escobar, Nedelcheva, Neuser, Neveďalová, Newton Dunn, Neynsky, Neyts-Uyttebroeck, Nicholson, Nicolai, Niculescu, Niebler, van Nistelrooij, Nitras, Ojuland, Olbrycht, Olejniczak, Oomen-Ruijten, Ortiz Vilella, Őry, Ouzký, Oviir, Pack, Padar, Paleckis, Paliadeli, Pallone, Panayotov, Panzeri, Papadopoulou, Papanikolaou, Papastamkos, Pargneaux, Parvanova, Paşcu, Paška, Patrão Neves, Patriciello, Paulsen, Peillon, Perello Rodriguez, Peterle, Pieper, Pietikäinen, Pirillo, Pirker, Pittella , Plumb, Poc, Podimata, Ponga, Poręba, Posselt, Pöttering, Poupakis, Preda, Prendergast, Prodi, Protasiewicz, Proust, Quisthoudt-Rowohl, Rangel, Ransdorf, Rapkay, Rapti, Regner, Reimers, Remek, Reul, Riera Madurell, Ries, Rinaldi, Rivasi, Rivellini, Roatta, Rodust, Rohde, Roithová, Romero López, Romeva i Rueda, Ronzulli, Rosbach, Rossi, Roth-Behrendt, Rouček, Rübig, Rubiks, Šadurskis, Saïfi, Salafranca Sánchez-Neyra, Salatto, Salavrakos, Salvini, Sánchez Presedo, Sanchez-Schmid, Sârbu, Sargentini, Sartori, Saryusz-Wolski, Sassoli, Saudargas, Savisaar-Toomast, Schaake, Schaldemose, Schlyter, Olle Schmidt, Schnellhardt, Schnieber-Jastram, Scholz, Schöpflin, Schroedter, Martin Schulz, Werner Schulz, Schwab, Scicluna, Scurria, Sedó i Alabart, Seeber, Sehnalová, Senyszyn, Serracchiani, Severin, Siekierski, Silvestris, Simon, Simpson, Sinclaire, Sippel, Skinner, Skrzydlewska, Skylakakis, Smolková, Sógor, Sommer, Søndergaard, Sonik, Sosa Wagner, Speroni, Stadler, Staes, Stassen, Šťastný, Stavrakakis, Steinruck, Stolojan, Strejček, Striffler, Surján, Susta, Svensson, Swinburne, Swoboda, Szájer, Szegedi, Szymański, Tabajdi, Takkula, Tănăsescu, Tarabella, Tarand, Tatarella, Tavares, Teixeira, Thein, Theocharous, Theurer, Thomsen, Thun und Hohenstein, Thyssen, Ţicău, Tirolien, Toia, Tőkés, Tošenovský, Trautmann, Tremopoulos, Tremosa i Balcells, Trzaskowski, Tsoukalas, Turmes, Turunen, Uggias, Ulmer, Ulvskog, Ungureanu, Urutchev, Vaidere, Vajgl, Vălean, Van Brempt, Van Orden, Vattimo, Vaughan, Vergnaud, Verheyen, Verhofstadt, Vidal-Quadras , Vigenin, Vlasák, Vlasto, Voss, Wallis, Watson, Henri Weber, Manfred Weber, Renate Weber, Weidenholzer, Weiler, Weisgerber, Werthmann, Westlund, Westphal, Wieland, Wikström, Willmott, Wils, Iuliu Winkler, Włosowicz, Wojciechowski, Wortmann-Kool, Yannakoudakis, Záborská, Zahradil, Zala, Zalba Bidegain, Zalewski, Zanicchi, Zanoni, Zasada, Ždanoka, Zeller, Zemke, Zīle, Zimmer, Ziobro, Zver, Zwiefka
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
ENVI(2012)0123_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Måndagen den 23 januari 2012 kl. 15.00–18.30
Tisdagen den 24 januari 2012 kl. 9.00–12.30 och kl. 15.00–18.30
Onsdagen den 25 januari 2012 kl. 9.00–12.30
Bryssel
Lokal: József Antall (4Q2)
23 januari 2012 kl. 15.00–15.45
Konstituerande sammanträde – Val av ordförande och vice ordförande
* * *
23 januari 2012 kl. 15.45–18.30
1.
Godkännande av föredragningslistan
2.
Meddelanden från ordföranden
3.
Översynen av det sjätte miljöhandlingsprogrammet och fastställandet av prioriteringar för det sjunde miljöhandlingsprogrammet
ENVI/7/06549
2011/2194(INI)
Föredragande:
Jo Leinen (S&D)
PR – PE478.523v01-00
Ansv. utsk.:
ENVI –
Rådg. utsk.:
ITRE –
Cristina Gutiérrez-Cortines (PPE)
PA – PE476.125v01-00 AM – PE478.700v01-00
REGI –
Vasilica Viorica Dăncilă (S&D)
PA – PE480.527v01-00
· Behandling av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 26 januari 2012 kl. 12.00
4.
Vår livförsäkring, vårt naturkapital – en strategi för biologisk mångfald i EU fram till 2020
ENVI/7/06548
2011/2307(INI) COM(2011)0244
Föredragande:
Gerben-Jan Gerbrandy (ALDE)
PR – PE478.540v01-00
Ansv. utsk.:
ENVI –
Rådg. utsk.:
ITRE –
Romana Jordan Cizelj (PPE)
PA – PE478.435v01-00
REGI –
Catherine Bearder (ALDE)
PA – PE478.368v01-00
AGRI –
Vasilica Viorica Dăncilă (S&D)
PA – PE480.548v01-00
PECH –
Crescenzio Rivellini (PPE)
PA – PE476.103v01-00 AM – PE478.664v01-00
· Behandling av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 27 januari 2012 kl. 12.00
5.
Rapport från delegationen till FN:s ramkonvention om klimatförändringar (COP 17) i Durban, Sydafrika
ENVI/7/08179
· Diskussion
* * *
24 januari 2012 kl. 9.00–12.30
*** Elektronisk omröstning ***
6.
Minimikrav för arbetstagares hälsa och säkerhet vid exponering för risker som har samband med fysikaliska agens (elektromagnetiska fält)
ENVI/7/06524
***I 2011/0152(COD) COM(2011)0348 – C7-0191/2011
Föredragande av yttrande:
Philippe Juvin (PPE)
PA – PE475.801v01-00 AM – PE478.387v01-00
Ansv. utsk.:
EMPL –
Elisabeth Morin-Chartier (PPE)
PR – PE474.084v02-00 AM – PE478.400v01-00
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 5 december 2011 kl. 12.00
7.
Ansvarsfrihet 2010: EU:s allmänna budget, avsnitt III, kommissionen
ENVI/7/06938
2011/2201(DEC) COM(2011)0473 [01] – C7-0256/2011
Föredragande av yttrande:
Jutta Haug (S&D)
PA – PE476.049v01-00 AM – PE478.622v01-00
Ansv. utsk.:
CONT –
Christofer Fjellner (PPE)
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 20 december 2011 kl. 18.00
8.
Ansvarsfrihet 2010: Europeiska miljöbyrån
ENVI/7/07233
2011/2217(DEC) COM(2011)0473 [15] – C7-0278/2011
Föredragande av yttrande:
Jutta Haug (S&D)
PA – PE476.052v01-00 AM – PE478.626v01-00
Ansv. utsk.:
CONT –
Monica Luisa Macovei (PPE)
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 20 december 2011 kl. 18.00
9.
Ansvarsfrihet 2010: Europeiska läkemedelsmyndigheten
ENVI/7/07239
2011/2220(DEC) COM(2011)0473 [18] – C7-0281/2011
Föredragande av yttrande:
Jutta Haug (S&D)
PA – PE476.054v01-00 AM – PE478.634v01-00
Ansv. utsk.:
CONT –
Monica Luisa Macovei (PPE)
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 20 december 2011 kl. 18.00
10.
Ansvarsfrihet 2010: Europeiska myndigheten för livsmedelssäkerhet
ENVI/7/07249
2011/2226(DEC) COM(2011)0473 [23] – C7-0286/2011
Föredragande av yttrande:
Jutta Haug (S&D)
PA – PE476.053v01-00 AM – PE478.706v01-00 AM – PE478.631v01-00
Ansv. utsk.:
CONT –
Monica Luisa Macovei (PPE)
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 20 december 2011 kl. 18.00
11.
Ansvarsfrihet 2010: Europeiskt centrum för förebyggande och kontroll av sjukdomar
ENVI/7/07251
2011/2227(DEC) COM(2011)0473 [24] – C7-0287/2011
Föredragande av yttrande:
Jutta Haug (S&D)
PA – PE476.050v01-00
Ansv. utsk.:
CONT –
Monica Luisa Macovei (PPE)
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 20 december 2011 kl. 18.00
12.
Ansvarsfrihet 2010: Europeiska kemikaliemyndigheten
ENVI/7/07266
2011/2235(DEC) COM(2011)0473 [31] – C7-0294/2011
Föredragande av yttrande:
Jutta Haug (S&D)
PA – PE476.051v01-00 AM – PE478.635v01-00
Ansv. utsk.:
CONT –
Monica Luisa Macovei (PPE)
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 20 december 2011 kl. 18.00
13.
Europeiska investeringsbanken (EIB) – Årsrapport 2010
ENVI/7/06849
2011/2186(INI)
Föredragande av yttrande:
Crescenzio Rivellini (PPE)
PA – PE476.126v01-00 AM – PE478.621v01-00
Ansv. utsk.:
CONT –
Iliana Ivanova (PPE)
PR – PE476.140v01-00
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 20 december 2011 kl. 18.00
14.
Kvinnor och klimatförändringarna
ENVI/7/06917
2011/2197(INI)
Föredragande av yttrande:
Bairbre de Brún (GUE/NGL)
PA – PE476.068v01-00 AM – PE478.614v01-00
Ansv. utsk.:
FEMM –
Nicole Kiil-Nielsen (Verts/ALE)
PR – PE476.093v01-00 AM – PE478.628v01-00
· Antagande av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 20 december 2011 kl. 12.00
*** Den elektroniska omröstningen avslutas ***
15.
Muntlig fråga 2012/01 från Linda McAvan om bristfälliga silikonbröstinplantat tillverkade av det franska företaget PIP
ENVI/7/08488
CM – PE480.508v01-00
· Diskussion med kommissionens företrädare
16.
Rapport från delegationsbesöket i Turkiet
ENVI/7/08556
· Diskussion
17.
Diskussion med Mette Gjerskov (Danmarks minister för livsmedel, lantbruk och fiske)
ENVI/7/08076
· Redogörelse för rådsordförandeskapets program
* * *
24 januari 2012 kl. 15.00–18.30
18.
Diskussion med Martin Lidegaard (Danmarks minister för klimat-, energi- och byggnadsfrågor)
ENVI/7/08077
· Redogörelse för rådsordförandeskapets program
19.
Utfrågning av de kandidater som önskar bli Europaparlamentets representanter i styrelsen för Europeiska miljöbyrån (EEA)
ENVI/7/07665
· Utfrågning
* * *
24 januari 2012 kl. 18.30–20.00
Inom stängda dörrar
20.
Samordnarnas sammanträde
* * *
25 januari 2012 kl. 9.00–12.30
21.
Diskussion med Pia Olsen Dyhr (Danmarks tillförordnade hälsovårdsminister)
ENVI/7/08078
· Redogörelse för rådsordförandeskapets program
22.
6:e världsforumet för vatten i Marseille, 12–17 mars 2012
ENVI/7/08359
· Godkännande av fråga för muntligt besvarande
· Behandling av utkast till förslag till resolution
· Tidsfrist för ingivande av ändringsförslag: 31 januari 2012 kl. 12.00
23.
Diskussion med Ida Auken (Danmarks miljöminister)
ENVI/7/08079
· Redogörelse för rådsordförandeskapets program
24.
Kommande sammanträden
· 30 januari 2012 kl. 15.00–18.30 (Bryssel)
· 31 januari 2012 kl. 9.00–12.30 (Bryssel)
Utskottet för utrikesfrågor
AFET(2012)0131_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Tisdagen den 31 januari 2012 kl. 10.00–12.00 och kl. 15.00–18.30
Bryssel
Lokal: József Antall (2Q2)
31 januari 2012 kl. 10.00–11.00
1.
Godkännande av föredragningslistan
2.
Meddelanden från ordföranden
3.
Justering av protokollet från sammanträdet den
· 12 december 2011 PV – PE478.487v01-00
4.
Diskussion med Abdul Latif Bin Rashid Al Zayani, generalsekreterare för Gulfstaternas samarbetsråd (GCC), om förbindelserna mellan EU och GCC
31 januari 2012 kl. 11.00–12.00
Inom stängda dörrar
5.
Diskussion med Sven Kuehn von Burgsdorff, nyutnämnd chef för EU:s delegation till Sydsudan
31 januari 2012 kl. 15.00–17.15
6.
Handel för att uppnå förändring: EU:s handels- och investeringsstrategi för södra Medelhavsområdet efter vårrevolutionerna i arabländerna
AFET/7/06738
2011/2113(INI)
Föredragande av yttrande:
Godelieve Quisthoudt-Rowohl (PPE)
PA – PE473.976v01-00 AM – PE478.670v01-00
Ansv. utsk.:
INTA –
Niccolò Rinaldi (ALDE)
PR – PE478.639v02-00 DT – PE478.391v01-00
· Behandling av förslag till yttrande
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 12 januari 2012 kl. 12.00
7.
Europaparlamentets resolution om 2011 års framstegsrapport om Island
AFET/7/07419
Föredragande:
Cristian Dan Preda (PPE)
AM – PE478.707v01-00
· Behandling av utkast till förslag till resolution
· Behandling av ändringsförslag
· Tidsfrist för ingivande av ändringsförslag: 12 januari 2012 kl. 12.00
8.
Rekommendation till rådet, kommissionen och Europeiska utrikestjänsten om förhandlingarna om associeringsavtalet mellan EU och Armenien
AFET/7/08278
2011/2315(INI)
Föredragande:
Tomasz Piotr Poręba (ECR)
PR – PE478.533v01-00
Ansv. utsk.:
AFET –
Rådg. utsk.:
INTA –
· Behandling av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 2 februari 2012 kl. 12.00
9.
Rekommendation till rådet, kommissionen och Europeiska utrikestjänsten om förhandlingarna om associeringsavtalet mellan EU och Azerbajdzjan
AFET/7/08279
2011/2316(INI)
Föredragande:
Anneli Jäätteenmäki (ALDE)
PR – PE478.534v01-00
Ansv. utsk.:
AFET –
Rådg. utsk.:
INTA –
· Behandling av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 2 februari 2012 kl. 12.00
31 januari 2012 kl. 17.15–18.30
Inom stängda dörrar
10.
Diskussion med Samuel Zbogar, EU:s nyutnämnda särskilda representant och chef för kontoret i Kosovo
11.
Övriga frågor
12.
Kommande sammanträden
· 6 februari 2012 kl. 15.00–18.30 (Bryssel)
Europaparlamentet i veckan: ACTA, finansiell transaktionsskatt, tvåpacket, passagerarrättigheter
Institutioner
2012-02-27 - 16:50
EP this week 27 februari - 2 mars möts Europaparlamentets politiska grupper och utskotten.
På tisdag kl. 12.30 överlämnas en framställning med över 2,4 miljoner underteckningar mot ACTA-avtalet, som syftar till att förhindra piratkopiering och varumärkesförfalskning.
Avtalet diskuteras i industriutskottet på tisdag och i utskottet för internationell handel på onsdag.
Under torsdagen arrangeras en workshop om avtalet.
Ekonomisk styrning
På onsdag är kreditvärderingsinstitut , avgifter på finansiella transaktioner samt monetär dialog med eurogruppens ordförande Jean-Claude Juncker i fokus för ekonomiutskottet.
Flyget och utsläppshandel är uppe för diskussion i transportutskottet och miljöutskottet, som dessutom röstar om strängare regler för barnmat .
Frågan om överföring av flygresenärers uppgifter ( PNR ) mellan EU och USA är återigen på dagordningen.
Utskottet för medborgerliga fri- och rättigheter diskuterar PNR på måndag.
Utrikesutskottet tar emot ministrar från Bahrain, Jordanien och Qatar.
Delegationen kommer också att möta Aung San Suu Kyi (29 februari).
20120223STO39228 Direktsändningar Europaparlamentets informationskontor i Sverige - nyhetsbrev ACTA - veckans webbutsändningar Mer om ACTA
SV
1
EPTVPHOTO
20120124PHT36092.jpg
SV
2
EUROPARL-TV
http://europarltv.europa.eu/sv/player.aspx?pid=0979eeee-077e-43f7-b95a-a000013bf422
SV
3
LINK
/ep-live/en/schedule/
SV
4
LINK
http://www.europaparlamentet.se/view/sv/Nyhetsbrev/vecka_09_12.html
SV
5
LINK
http://events.europarl.europa.eu/
-//EP//TEXT IM-PRESS 20120220FCS38611 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Hur påverkar ACTA civila friheter och tillgång till generiska läkemedel?
Handel med tredje land
Informationssamhället
2012-03-02 - 14:50
Det fruktar motståndarna till handelsavtalet som ska hindra varumärkesförfalskning.
Medborgerliga fri- och rättigheter
För juristen Oliver Vrins anger texten att handelsavtalet för bekämpning av varumärkesförfalskning (ACTA) ska genomföras med respekt för grundläggande rättigheter, som yttrandefrihet och rätt till en rättvis rättegång.
Oliver Vrins ansåg inte att ACTA-avtalet är ett allvarligt hot mot europeiska medborgares grundläggande rättigheter.
Rupert Schlegelmilch, Europeiska kommissionen, sa att hans institution verkligen tagit till sig att människor är bekymrade över respekten för medborgerliga rättigheter, men det finns ingen anledning till oro.
- Intellektuell egendom handlar om egendom, men inte bara det.
Respekt för privatlivet och internet är lika viktigt.
Vi tror att avtalet skapar en rättvis balans.
Han förklarade att inga nya standarder införs genom ACTA.
Syftet är tillämpning av nuvarande regler.
Professor Meir Pugatch från Haifas universitet ansåg inte att ACTA varken blockerar eller underlättar tillgången till generiska läkemedel.
- Det verkliga problemet är förfalskade och dåliga läkemedel som kan äventyra hälsan.
Förfalskade och dåliga läkemedel drabbar framför allt fattiga människor, sa Pugatch och betonade att generiska läkemedel behövs.
Rupert Schlegelmilch sa att utvecklingsländerna precis som tidigare kommer att kunna köpa generiska läkemedel.
Parlamentets föredragande, brittiske ledamoten David Martin (S&D) saknade tillräcklig information.
- Vi vet inte på vilket sätt gränskontrollmyndigheterna ska definiera varumärkesförfalskade läkemedel jämfört med generiska läkemedel (...).
Hur ska det fungera?
- Ett talesätt säger att "djävulen sitter i detaljerna".
Problemet med ACTA är att djävulen sitter i bristen på detaljer.
Vi saknar tillräcklig information på många av de områden vi i slutändan ska bedöma, sa David Martin.
20120223STO39243 Läs mer om ACTA ACTA: Text Oberoende analys av ACTA (på engelska)
SV
1
PHOTO
20120302PHT39811.jpg
SV
3
LINK
http://register.consilium.europa.eu/pdf/sv/11/st12/st12196.sv11.pdf
SV
4
LINK
/committees/en/INTA/studiesdownload.html?languageDocument=EN&file=43731
-//EP//TEXT IM-PRESS 20120220FCS38611 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Obligationer designade att attrahera ny finansiering till EU:s infrastruktur
Ekonomiska och monetära frågor
2012-03-08 - 16:52
©Belga/Belpress När banker inte lånar ut pengar och regeringar inte vill spendera - försök med obligationer.
Ett förslag för att göra obligationerna attraktiva är att backa upp investerarna med garantier och lån.
Kommissionen uppskattar att det fram till år 2020 behövs 150 till 200 biljoner euro per år för att modernisera EU:s infrastruktur - det vill säga exempelvis järnvägar, gasledningar och bredband.
Samtidigt erbjuder marknaden, genom kapital och banklån, bara 60 till 80 biljoner euro årligen.
Mer kapital behövs med andra ord men det är inte lätt att komma över.
Dels för att bankerna behöver extra kapital till sig själva och därför begränsar sina lån.
Dessutom har investerare blivit mer ovilliga eftersom investeringar inom infrastruktur är riskabelt.
Det är så kallade projektobligationer som kan hjälpa privata företag att finansiera olika europeiska infrastrukturprojekt, särskilt de som är strategiskt viktiga.
Socialdemokraten Göran Färm (S&D) som ansvarar för frågan om pilotprojektet av obligationerna i budgetutskottet, ger kommissionen medhåll.
- Det behövs nya sätt att samla investeringskapital, säger han.
I praktiken innebär projektobligationerna att Europeiska investeringsbanken (EIB) erbjuder lån och garantier för olika projekt vilket är tänkt ska förskjuta risken av privata investeringar.
Detta förväntas öka kreditkvaliteten på skulder vilket gör det attraktivt för institutionella investerare, det vill säga pensionsfonder och försäkringsbolag.
- Obligationerna kommer att minska riskerna för investerare att förlora pengar.
De kommer också att få flera andra effekter.
En euro från EU:s budget kan ge 15 till 20 euro från pensionsfonder och andra investerare, säger Göran Färm (S&D).
Kritiska röster
Även om de flesta av parlamentets ledamöter är positiva till idén med projektobligationer så hörs en del varnande röster.
Ekonomiutskottets ordförande, brittiska Sharon Bowles (ALDE) är en av dem.
- Det blir i själva verket en begränsad garanti för de första förlusterna.
Det här förändrar bara gradvis de potentiella förlusterna för privata ägare av obligationerna men innebär inte att risken försvinner, säger hon.
Strejček, vars partigrupp är emot idén, menar att man uppmuntrar investeringar som behöver skattebetalarnas pengar som garanti.
Obligationerna snart verklighet?
Budgetutskottet väntas rösta i april om förslaget, och hela parlamentet i juli.
Innan projektobligationerna i så fall tas i bruk år 2014 så pågår en prövoperiod.
230 miljoner euro vill budgetutskottet att man bidrar med till Europeiska investeringsbanken för att täcka riskerna de tar för att finansiera fem till tio lämpliga projekt inom transport, energi och bredband som budgetutskottet tror kan leda till investeringar på upp till 4,6 biljoner euro.
20120302STO39869 Kommissionens förslag (på engelska) Europaparlamentets resolution 08.03.2011 Frågor och svar (på engelska) EP pressmeddelande 05.07.2011 (på engelska)
SV
1
PHOTO
20120131PHT36652.jpg
SV
2
LINK
http://ec.europa.eu/economy_finance/financial_operations/investment/europe_2020/index_en.htm
SV
4
LINK
http://europa.eu/rapid/pressReleasesAction.do?reference=MEMO/11/707&format=HTML&aged=0&language=EN&guiLanguage=en
-//EP//TEXT TA P7-TA-2011-0080 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Strasbourg Måndagen den 12 mars 2012 Torsdagen den 15 mars 2012 FÖREDRAGNINGSLISTA Onsdagen den 14 mars 2012 15:58 Särskild omröstning - delad omröstning - omröstning med namnupprop
George Lyon Utskottet för jordbruk och landsbygdens utveckling Gemensam handelspolitik Betänkande: Godelieve Quisthoudt-Rowohl ( A7-0028/2012 ) 2011/0039(COD) ***I Gemensam handelspolitik COM(2011)0082 A7-0028/2012 Utskottet för internationell handel INTA/7/05563 Godelieve Quisthoudt-Rowohl Utskottet för internationell handel Betänkande om förslaget till Europaparlamentets och rådets förordning om ändring av vissa förordningar om den gemensamma handelspolitiken vad gäller förfarandena för antagande av vissa åtgärder
Europeiska rådets ordförande (inklusive repliker) 1 15:00 Rådet (inklusive repliker) 1 05:00 Kommissionen (inklusive repliker) 1 15:00 Frågeställare 1 05:00 Ledamöter Europeiska folkpartiets grupp (kristdemokrater) 34:00 Gruppen Progressiva förbundet av Socialdemokrater i Europaparlamentet 24:30 Gruppen Alliansen liberaler och demokrater för Europa 12:00 Gruppen De gröna/Europeiska fria alliansen 09:00 Gruppen Europeiska konservativa och reformister 08:00 Gruppen Europeiska enade vänstern/Nordisk grön vänster 06:00 Gruppen Frihet och demokrati i Europa 06:00 Grupplösa 05:30 Ögonkontaktsförfarandet 2 05:00 Rådet (inklusive repliker) 1 10:00 Kommissionen (inklusive repliker) 1 10:00 Ledamöter Europeiska folkpartiets grupp (kristdemokrater) 04:00 Gruppen Progressiva förbundet av Socialdemokrater i Europaparlamentet 03:30 Gruppen Alliansen liberaler och demokrater för Europa 02:30 Gruppen De gröna/Europeiska fria alliansen 02:30 Gruppen Europeiska konservativa och reformister 02:30 Gruppen Europeiska enade vänstern/Nordisk grön vänster 02:00 Gruppen Frihet och demokrati i Europa 02:00 Grupplösa 02:00 Rådet (inklusive repliker) 1 10:00 Kommissionen (inklusive repliker) 1 25:00 Föredragande 2 06:00 Ledamöter Europeiska folkpartiets grupp (kristdemokrater) 12:30 Gruppen Progressiva förbundet av Socialdemokrater i Europaparlamentet 09:30 Gruppen Alliansen liberaler och demokrater för Europa 05:30 Gruppen De gröna/Europeiska fria alliansen 04:00 Gruppen Europeiska konservativa och reformister 04:00 Gruppen Europeiska enade vänstern/Nordisk grön vänster 03:30 Gruppen Frihet och demokrati i Europa 03:30 Grupplösa 03:00 Ögonkontaktsförfarandet 3 05:00 Kommissionen (inklusive repliker) 1 15:00 Föredragande 3 06:00 Föredragande av yttrande 1 01:00 Ledamöter Europeiska folkpartiets grupp (kristdemokrater) 12:30 Gruppen Progressiva förbundet av Socialdemokrater i Europaparlamentet 09:30 Gruppen Alliansen liberaler och demokrater för Europa 05:30 Gruppen De gröna/Europeiska fria alliansen 04:00 Gruppen Europeiska konservativa och reformister 04:00 Gruppen Europeiska enade vänstern/Nordisk grön vänster 03:30 Gruppen Frihet och demokrati i Europa 03:30 Grupplösa 03:00 Ögonkontaktsförfarandet 3 05:00 Arv och inrättandet av ett europeiskt arvsintyg A7-0045/2012 Kurt Lechner Utskottet för rättsliga frågor Ändringsförslag Onsdagen den 7 mars 2012 12:00 Jämställdheten mellan kvinnor och män i Europeiska unionen - 2011 A7-0041/2012 Sophia in 't Veld Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män Ändringsförslag Onsdagen den 7 mars 2012 12:00 Kvinnor i politiskt beslutsfattande A7-0029/2012 Sirpa Pietikäinen Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män Ändringsförslag som lagts fram av föredraganden eller minst 76 parlamentsledamöter; alternativa förslag till resolution Onsdagen den 7 mars 2012 12:00 Gemensamma alternativa förslag till resolution Måndagen den 12 mars 2012 19:00 Stadgan för europeiska kooperativa föreningar vad gäller arbetstagarinflytande A7-0432/2011 Sven Giegold Utskottet för sysselsättning och sociala frågor Ändringsförslag som lagts fram av föredraganden eller minst 76 parlamentsledamöter; alternativa förslag till resolution Onsdagen den 7 mars 2012 12:00 Gemensamma alternativa förslag till resolution Måndagen den 12 mars 2012 19:00 Bologna-processen A7-0035/2012 Luigi Berlinguer Utskottet för kultur och utbildning Ändringsförslag som lagts fram av föredraganden eller minst 76 parlamentsledamöter; alternativa förslag till resolution Onsdagen den 7 mars 2012 12:00 Gemensamma alternativa förslag till resolution Måndagen den 12 mars 2012 19:00 Kvalitetsledning för den europeiska statistiken A7-0037/2012 Edward Scicluna Utskottet för ekonomi och valutafrågor Ändringsförslag som lagts fram av föredraganden eller minst 76 parlamentsledamöter; alternativa förslag till resolution Onsdagen den 7 mars 2012 12:00 Gemensamma alternativa förslag till resolution Måndagen den 12 mars 2012 19:00 Diskriminerande internetsidor och myndigheternas reaktioner Resolutionsförslag Måndagen den 12 mars 2012 19:00 Ändringsförslag och gemensamma förslag till resolution Tisdagen den 13 mars 2012 19:00 Ändringsförslag till gemensamma förslag till resolution Tisdagen den 13 mars 2012 20:00 Begäranden om särskild omröstning, delad omröstning eller omröstning med namnupprop Onsdagen den 14 mars 2012 17:00 Allmänna riktlinjer för 2013 års budget – Avsnitt III – Kommissionen A7-0040/2012 Giovanni La Via Budgetutskottet Ändringsförslag Onsdagen den 7 mars 2012 12:00 Barnarbete i kakaosektorn Resolutionsförslag Onsdagen den 7 mars 2012 12:00 Ändringsförslag Måndagen den 12 mars 2012 19:00 Begäranden om särskild omröstning, delad omröstning eller omröstning med namnupprop Tisdagen den 13 mars 2012 19:00 Åtgärder mot diabetesepidemin i EU Resolutionsförslag Onsdagen den 7 mars 2012 12:00 Ändringsförslag och gemensamma förslag till resolution Måndagen den 12 mars 2012 19:00 Ändringsförslag till gemensamma förslag till resolution Måndagen den 12 mars 2012 20:00 Begäranden om särskild omröstning, delad omröstning eller omröstning med namnupprop Tisdagen den 13 mars 2012 19:00 Gemensam handelspolitik A7-0028/2012 Godelieve Quisthoudt-Rowohl Utskottet för internationell handel Ändringsförslag Onsdagen den 7 mars 2012 12:00 Onsdagen den 14 mars 2012 PRIORITERADE DEBATTER Utvidgningsrapport för f.d. jugoslaviska republiken Makedonien 2011/2887(RSP) Uttalanden av rådet och kommissionen Utvidgningsrapport för f.d. jugoslaviska republiken Makedonien B7-0127/2012 Utvidgningsrapport för Island 2011/2884(RSP) Uttalanden av rådet och kommissionen Utvidgningsrapport för Island B7-0125/2012 Utvidgningsrapport för Bosnien och Hercegovina 2011/2888(RSP) Uttalanden av rådet och kommissionen Utvidgningsrapport för Bosnien och Hercegovina B7-0129/2012 OMRÖSTNING följd av röstförklaringar Europeiska fiskerifonden Betänkande: João Ferreira ( A7-0447/2011 ) 2011/0212(COD) ***I Europeiska fiskerifonden COM(2011)0484 A7-0447/2011 Fiskeriutskottet PECH/7/06703 João Ferreira Fiskeriutskottet Betänkande om förslaget till Europaparlamentets och rådets förordning om ändring av rådets förordning (EG) nr 1198/2006 om Europeiska fiskerifonden vad gäller vissa bestämmelser om den ekonomiska förvaltningen för vissa medlemsstater som genomgår eller hotas av allvarliga svårigheter med avseende på deras ekonomiska stabilitet Artikel 138 i arbetsordningen Debatt: Tisdagen den 13 mars 2012 Autonom tullkvot för import av nötkött av hög kvalitet Betänkande: Godelieve Quisthoudt-Rowohl ( A7-0025/2012 ) 2011/0169(COD) ***I Autonom tullkvot för import av nötkött av hög kvalitet COM(2011)0384 A7-0025/2012 Utskottet för internationell handel INTA/7/06358 Godelieve Quisthoudt-Rowohl Utskottet för internationell handel Betänkande om förslaget till Europaparlamentets och rådets förordning om ändring av rådets förordning (EG) nr 617/2009 om öppnande av en autonom tullkvot för import av nötkött av hög kvalitet
George Lyon Utskottet för jordbruk och landsbygdens utveckling Artikel 138 i arbetsordningen Debatt: Tisdagen den 13 mars 2012 Gemensam handelspolitik Betänkande: Godelieve Quisthoudt-Rowohl ( A7-0028/2012 ) 2011/0039(COD) ***I Gemensam handelspolitik COM(2011)0082 A7-0028/2012 Utskottet för internationell handel INTA/7/05563 Godelieve Quisthoudt-Rowohl Utskottet för internationell handel Betänkande om förslaget till Europaparlamentets och rådets förordning om ändring av vissa förordningar om den gemensamma handelspolitiken vad gäller förfarandena för antagande av vissa åtgärder
Debatt: Tisdagen den 13 mars 2012 Allmänna riktlinjer för 2013 års budget – Avsnitt III – Kommissionen Betänkande: Giovanni La Via ( A7-0040/2012 ) 2012/2000(BUD) Allmänna riktlinjer för 2013 års budget – Avsnitt III – Kommissionen A7-0040/2012 Budgetutskottet BUDG/7/08444 Giovanni La Via Budgetutskottet Betänkande om de allmänna riktlinjerna för utarbetandet av 2013 års budget – Avsnitt III – Kommissionen Debatt: Tisdagen den 13 mars 2012 Mandat för det särskilda utskottet för organiserad brottslighet, korruption och penningtvätt 2012/2577(RSO) Mandat för det särskilda utskottet för organiserad brottslighet, korruption och penningtvätt B7-0151/2012 Resolutionsförslag - Rättslig utbildning 2012/2575(RSP) Rättslig utbildning B7-0150/2012 O-000059/2012 Kommissionen Utskottet för rättsliga frågor Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor Rättslig utbildning Klaus-Heiner Lehne Utskottet för rättsliga frågor Juan Fernando López Aguilar Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor Debatt: Måndagen den 12 mars 2012 Barnarbete i kakaosektorn 2011/2957(RSP) Resolutionsförslag Barnarbete i kakaosektorn B7-0126/2012 Debatt: Tisdagen den 13 mars 2012 2010 års internationella kakaoavtal Rekommendation: Vital Moreira ( A7-0024/2012 ) 2010/0343(NLE) *** 2010 års internationella kakaoavtal 09771/2011 A7-0024/2012 Utskottet för internationell handel INTA/7/04746 Vital Moreira Utskottet för internationell handel Rekommendation om utkastet till rådets beslut om ingående av 2010 års internationella kakaoavtal Artikel 138 i arbetsordningen Debatt: Tisdagen den 13 mars 2012 Åtgärder mot diabetesepidemin i EU 2011/2911(RSP) Resolutionsförslag Åtgärder mot diabetesepidemin i EU RC-B7-0145/2012 B7-0145/2012 B7-0146/2012 B7-0147/2012 B7-0148/2012 Debatt: Tisdagen den 13 mars 2012 Utvidgningsrapport för f.d. jugoslaviska republiken Makedonien 2011/2887(RSP) Resolutionsförslag Utvidgningsrapport för f.d. jugoslaviska republiken Makedonien B7-0127/2012 Debatt: Onsdagen den 14 mars 2012 Utvidgningsrapport för Island 2011/2884(RSP) Resolutionsförslag Utvidgningsrapport för Island B7-0125/2012 Debatt: Onsdagen den 14 mars 2012 Utvidgningsrapport för Bosnien och Hercegovina 2011/2888(RSP) Resolutionsförslag Utvidgningsrapport för Bosnien och Hercegovina B7-0129/2012 Debatt: Onsdagen den 14 mars 2012 Debatt Resultatet av presidentvalet i Ryssland 2012/2573(RSP) Uttalande av vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik Resultatet av presidentvalet i Ryssland B7-0177/2012 Kazakstan 2012/2553(RSP) Uttalande av vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik Kazakstan RC-B7-0135/2012 B7-0135/2012 B7-0140/2012 B7-0141/2012 B7-0142/2012 B7-0143/2012 B7-0144/2012 Situationen i Nigeria 2012/2550(RSP) Uttalande av vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik Situationen i Nigeria RC-B7-0131/2012 B7-0131/2012 B7-0133/2012 B7-0134/2012 B7-0137/2012 B7-0138/2012 B7-0139/2012 B7-0149/2012 Situationen i Vitryssland 2012/2581(RSP) Uttalande av vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik Situationen i Vitryssland RC-B7-0178/2012 B7-0178/2012 B7-0179/2012 B7-0180/2012 B7-0181/2012 B7-0182/2012 B7-0183/2012 Kapningar till sjöss 2011/2962(RSP) Uttalande av kommissionen Kapningar till sjöss Omröstningen kommer att äga rum vid en senare sammanträdesperiod.
I kristider måste EU:s budget stärka tillväxten
Budget
2012-03-23 - 14:59
Konferens om EU:s nästa långtidsbudget: EP:s talman Martin Schulz och Danmarks statsminister Helle Thorning-Schmidt Konferens om EU:s nästa långtidsbudget - 2014-2020 Långtidsbudgeten sätter ramar för olika utgiftsområden varje år "Europaparlamentet kommer inte att acceptera mindre pengar för EU:s budget."
Det sa Europaparlamentets talman Martin Schulz i konferensen om EU:s långtidsbudget för 2014-2020 den 22 mars.
Bara med en rimlig budget kan Europa investera för att öka tillväxten i en tid av sparsamhet, sa Schulz.
Han la till att EU:s budget borde vara fullt finansierad av egna medel för att undvika betungande förhandlingar om nationella bidrag mellan medlemsstaterna.
Ungefär 75 procent av EU:s budget finansieras av avgifter från medlemsländerna baserat på deras bruttonationalinkomst, BNI.
Det innebär förhandlingar om hur mycket varje medlemsstat ska bidra med och vad de får tillbaka.
Kommissionen har föreslagit nya typer av finansieringsmedel för budgeten: en EU-moms och även en skatt på finansiella transaktioner (FTT) som ska minska medlemsstaternas avgifter, och därmed alltså göra det enklare att komma överens om budgeten.
Kommissionens ordförande, José Manuel Barroso , menade att EU:s budget är en budget för investeringar och inte för rådande kostnader.
Det är inte en investering för Bryssel eller institutioner utan ska stödja projekt i EU:s olika regioner och städer.
- Vi vill ha ett enklare system utan undantag och rabatter och vi vill inte ha högre nettoskatter.
Vikten av att krympa bidragen lyfte även Andreas Mavroyiannis , ställföreträdande minister för europeiska frågor i Cypern fram.
Han menade att beroendet av nationella bidrag överskuggar de riktiga frågorna.
Eva Kjer Hansen , ordförande för Europautskottet i danska folketinget varnade för den påverkan som en skatt på finansiella transaktioner kan ha på tillväxten.
Hon menade att konkurrenskraften inte är tydlig och att skatt troligtvis inte kommer gynna det nödvändiga stödet som behövs av medlemsstaterna.
Även Milan M. Cvikl från Europeiska revisionsrätten var kritisk.
Han varnade för att intäkten genom den nya skatten sannolikt kommer att vara flyktig eftersom storleken på de finansiella transaktionerna varierar.
Samtidigt menade franska EU-ledamoten Pervenche Berès (S&D) som stödjer en skatt av finansiella transaktioner att man genom den kan få in skatt från områden som hittills har lyckats fly undan.
Budgetkommissionären Janusz Lewandowski menade att den nya skatten kan minska medlemsstaternas avgift baserat på BNI med upp till 50 procent till 2020.
Det skulle ge 54 miljarder euro och två tredjedelar av inkomsten från skatten skulle gå till EU:s budget och den sista tredjedelen till de nationella budgetarna.
På konferensen om EU:s långtidsbudget så deltog 42 ledamöter från 21 medlemsstater.
20120316STO41092 Program konferensen 22.03.2012 Fördjupning om EU:s nästa långtidsbudget EP:s resolution om en ny flerårig budgetram 08.06.2011 Kommissionen pressmeddelande om skatt på finansiella transaktioner 28.09.2011
SV
1
PHOTO
20120313PHT40600.jpg
SV
2
LINK
http://ec.europa.eu/budget/reform/conference-mff-2014-2020/files/draftprogramme_mff_22oct2012.pdf
SV
5
LINK
http://europa.eu/rapid/pressReleasesAction.do?reference=IP/11/1085&format=HTML&aged=1&language=SW&guiLanguage=en
-//EP//TEXT IM-PRESS 20110429FCS18370 0 NOT XML V0//SV
-//EP//TEXT TA P7-TA-2011-0266 0 NOT XML V0//SV
-//EP//DTD IM-PRESS 20050901 STO DOC XML V0//EN
-//EP//STYLESHEET IM-PRESS 20050901 STO DOC XML V0//EN
Utskottet för sysselsättning och sociala frågor
EMPL(2012)0326_1
FÖRSLAG TILL FÖREDRAGNINGSLISTA
Sammanträde
Måndagen den 26 mars 2012 kl. 15.00–18.30
Tisdagen den 27 mars 2012 kl. 9.00–12.30 och kl. 15.00–19.00
Bryssel
Lokal: József Antall (4Q1)
26 mars 2012 kl. 15.00–17.00
1.
Godkännande av föredragningslistan
2.
Meddelanden från ordföranden
3.
Justering av protokollet från sammanträdet den
· 25–26 januari 2012 PV – PE480.894v01-00
· 13 februari 2012 PV – PE483.507v01-00
------
4.
Skärpning av den ekonomiska övervakningen och övervakningen av de offentliga finanserna i medlemsstater som har, eller hotas av, allvarliga problem i fråga om deras finansiella stabilitet i euroområdet
EMPL/7/07963
***I 2011/0385(COD) COM(2011)0819 – C7-0449/2011
Föredragande av yttrande:
Frédéric Daerden (S&D)
PA – PE480.648v01-00 AM – PE483.682v01-00
Ansv. utsk.:
ECON –
Jean-Paul Gauzès (PPE)
PR – PE483.472v02-00 AM – PE485.871v01-00
· Behandling av kompromissändringsförslag
------
5.
Gemensamma bestämmelser för övervakning och bedömning av utkast till budgetplaner och säkerställande av korrigering av alltför stora underskott i medlemsstater i euroområdet
EMPL/7/07960
***I 2011/0386(COD) COM(2011)0821 – C7-0448/2011
Föredragande av yttrande:
Tamás Deutsch (PPE)
PA – PE480.645v01-00 AM – PE483.671v01-00
Ansv. utsk.:
ECON –
Elisa Ferreira (S&D)
PR – PE483.469v01-00 AM – PE485.870v01-00
· Behandling av kompromissändringsförslag
------
6.
Tillämpning av principen om lika lön för manliga och kvinnliga anställda för samma eller likvärdigt arbete
EMPL/7/07713
2011/2285(INI)
Föredragande av yttrande:
Gabriele Zimmer (GUE/NGL)
PA – PE478.673v01-00 AM – PE480.870v01-00
Ansv. utsk.:
FEMM –
Edit Bauer (PPE)
PR – PE480.835v01-00 AM – PE483.791v01-00
· Behandling av kompromissändringsförslag
------
7.
EU:s program för social förändring och social innovation
EMPL/7/07508
***I 2011/0270(COD) COM(2011)0609 – C7-0318/2011
Föredragande:
Jutta Steinruck (S&D)
PR – PE483.795v01-00
Ansv. utsk.:
EMPL –
Rådg. utsk.:
BUDG –
Estelle Grelier (S&D)
CONT –
Jens Geier (S&D)
ITRE –
Inês Cristina Zuber (GUE/NGL)
PA – PE483.686v01-00
REGI –
CULT – Beslut: inget yttrande
FEMM –
Barbara Matera (PPE)
· Behandling av förslag till betänkande
· Tidsfrist för ingivande av ändringsförslag: 17 april 2012 kl. 12.00
------
26 mars 2012 kl. 17.00–18.00
8.
Diskussion med Jean-François Mézières och Stamatis Paleocrassas, Europaparlamentets experter i Europeiska yrkesutbildningsstiftelsens styrelse – slutet på mandatperioden
26 mars 2012 kl. 18.00–18.30
9.
Europeiska fonden för justering för globaliseringseffekter (2014–2020)
EMPL/7/07500
***I 2011/0269(COD) COM(2011)0608 – C7-0319/2011
Föredragande:
Marian Harkin (ALDE)
Ansv. utsk.:
EMPL –
Rådg. utsk.:
INTA –
Iuliu Winkler (PPE)
PA – PE483.733v01-00
BUDG –
Miguel Portas (GUE/NGL)
CONT –
Jorgo Chatzimarkakis (ALDE)
ITRE – Beslut: inget yttrande
REGI –
Jens Geier (S&D)
AGRI –
Luís Paulo Alves (S&D)
FEMM –
Vilija Blinkevičiūtė (S&D)
PA – PE483.818v01-00
· Diskussion utan dokument
* * *
27 mars 2012 kl. 9.00–9.30
10.
De 20 viktigaste problemen på den inre marknaden för europeiska företag och medborgare
EMPL/7/08654
2012/2044(INI) SEC(2011)1003
Föredragande av yttrande:
Nadja Hirsch (ALDE)
PA – PE480.882v01-00 AM – PE483.810v01-00
Ansv. utsk.:
IMCO –
Regina Bastos (PPE)
PR – PE483.745v01-00
· Behandling av ändringsförslag
27 mars 2012 kl. 9.30–10.30
*** Elektronisk omröstning ***
11.
Skärpning av den ekonomiska övervakningen och övervakningen av de offentliga finanserna i medlemsstater som har, eller hotas av, allvarliga problem i fråga om deras finansiella stabilitet i euroområdet
EMPL/7/07963
***I 2011/0385(COD) COM(2011)0819 – C7-0449/2011
Föredragande av yttrande:
Frédéric Daerden (S&D)
PA – PE480.648v01-00 AM – PE483.682v01-00
Ansv. utsk.:
ECON –
Jean-Paul Gauzès (PPE)
PR – PE483.472v02-00 AM – PE485.871v01-00
· Antagande av förslag till yttrande
12.
Gemensamma bestämmelser för övervakning och bedömning av utkast till budgetplaner och säkerställande av korrigering av alltför stora underskott i medlemsstater i euroområdet
EMPL/7/07960
***I 2011/0386(COD) COM(2011)0821 – C7-0448/2011
Föredragande av yttrande:
Tamás Deutsch (PPE)
PA – PE480.645v01-00 AM – PE483.671v01-00
Ansv. utsk.:
ECON –
Elisa Ferreira (S&D)
PR – PE483.469v01-00 AM – PE485.870v01-00
· Antagande av förslag till yttrande
13.
Tillämpning av principen om lika lön för manliga och kvinnliga anställda för samma eller likvärdigt arbete
EMPL/7/07713
2011/2285(INI)
Föredragande av yttrande:
Gabriele Zimmer (GUE/NGL)
PA – PE478.673v01-00 AM – PE480.870v01-00
Ansv. utsk.:
FEMM –
Edit Bauer (PPE)
PR – PE480.835v01-00 AM – PE483.791v01-00
· Antagande av förslag till yttrande
*** Den elektroniska omröstningen avslutas ***
27 mars 2012 kl. 10.30–11.00
14.
Diskussion om budgetförslaget för 2013 med Giovanni La Via, föredragande för 2013 års budget
27 mars 2012 kl. 11.00–12.30
15.
Utfrågning om initiativet för ungdomars möjligheter Diskussion med – Kommissionens representant (GD Empl) – Génération Precaire, Florence Morillon – Europeiska ungdomsforumet, Giuseppe Porcaro, generalsekreterare – Europeiska fackliga samorganisationen (EFS), vice generalsekreterare – Business Europe, Maxime Cerutti, direktör för sociala frågor
* * *
27 mars 2012 kl. 15.00–16.45
16.
Ändring av Europaparlamentets och rådets direktiv 2008/106/EG om minimikrav på utbildning för sjöfolk
EMPL/7/06836
***I 2011/0239(COD) COM(2011)0555 – C7-0246/2011
Föredragande av yttrande:
Ole Christensen (S&D)
PA – PE480.883v02-00
Ansv. utsk.:
TRAN –
Brian Simpson (S&D)
PR – PE480.581v01-00
· Behandling av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 29 mars 2012 kl. 12.00
------
17.
Instrument för stöd inför anslutningen
EMPL/7/08314
***I 2011/0404(COD) COM(2011)0838 – C7-0491/2011
Föredragande av yttrande:
Marije Cornelissen (Verts/ALE)
PA – PE483.844v03-00
Ansv. utsk.:
AFET –
Kristian Vigenin (S&D)
· Behandling av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 2 april 2012 kl. 12.00
------
18.
Europeiska statistikprogrammet 2013-2017
EMPL/7/08392
***I 2011/0459(COD) COM(2011)0928 – C7-0001/2012
Föredragande av yttrande:
Ádám Kósa (PPE)
PA – PE483.792v01-00
Ansv. utsk.:
ECON –
Edward Scicluna (S&D)
· Behandling av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 4 april 2012 kl. 12.00
------
19.
Stadga för europeiska ömsesidiga bolag
EMPL/7/08937
2012/2039(INI)
Föredragande av yttrande:
Regina Bastos (PPE)
PA – PE483.860v01-00
Ansv. utsk.:
JURI* –
Luigi Berlinguer (S&D)
Rådg. utsk.:
ECON –
EMPL* –
· Behandling av förslag till yttrande
· Tidsfrist för ingivande av ändringsförslag: 3 april 2012 kl. 12.00
27 mars 2012 kl. 17.00–19.00
20.
Gemensamt sammanträde med utskottet för ekonomi och valutafrågor (lokal: JAN 2Q2): – Diskussion med trojkan om den ekonomiska och sociala krisen i Grekland (se separat program)
------
21.
Övriga frågor
22.
Kommande sammanträden
· 23 april 2012 kl. 15.00–18.30 (Bryssel)
· 24 april 2012 kl. 9.00–12.30 och kl. 15.00–18.30 (Bryssel)
* * *
SLUTLIG VERSION
A6-0028/2004
*
BETÄNKANDE
om komissionens förslag till rådets förordning om standarder för säkerhetsdetaljer och biometriska kännetecken i EU-medborgarnas pass
(KOM(2004)0116 – C5‑0101/2004 – 2004/0039(CNS))
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Föredragande:
Carlos Coelho
Teckenförklaring
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................14
ÄRENDETS GÅNG..................................................................................................................20
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om kommissionens förslag till rådets förordning om standarder för säkerhetsdetaljer och biometriska kännetecken i EU-medborgarnas pass
( KOM(2004)0116 – C5‑0101/2004 – 2004/0039(CNS) )
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag ( KOM(2004)0116 )
EUT C 98, 23.4.2004, s.
39. ,
– med beaktande av artikel 67 i EG-fördraget, i enlighet med vilken rådet har hört parlamentet ( C5–0101/2004 ),
– med beaktande av protokollet om införlivande av Schengenregelverket inom Europeiska unionens ramar, i enlighet med vilket rådet har hört parlamentet
– med beaktande av artikel 51 i arbetsordningen,
– med beaktande av betänkandet från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor ( A6‑0028/2004 ).
1.
Kommissionens förslag
Parlamentets ändringar
Ändringsförslag
1
Skäl 2
(2) Minimisäkerhetsstandarder för pass infördes genom en resolution antagen av företrädarna för medlemsstaternas regeringar, församlade i rådet, av den 17 oktober 2000.
Denna resolution bör nu ersättas och uppdateras genom en gemenskapsåtgärd i syfte att skapa mer harmoniserade säkerhetsstandarder för pass som ger ett bättre skydd mot förfalskning.
Samtidigt bör biometriska kännetecken integreras i passet för att skapa en tillförlitlig koppling mellan den egentliga innehavaren och handlingen.
(2) Minimisäkerhetsstandarder för pass infördes genom en resolution antagen av företrädarna för medlemsstaternas regeringar, församlade i rådet, av den 17 oktober 2000.
Europeiska rådet har beslutat att denna resolution nu bör ersättas och uppdateras genom en gemenskapsåtgärd i syfte att skapa mer harmoniserade säkerhetsstandarder för pass som ger ett bättre skydd mot förfalskning.
Samtidigt bör biometriska kännetecken integreras i passet för att skapa en tillförlitlig koppling mellan den egentliga innehavaren och handlingen.
Motivering
Det bör understrykas att rådet fattade ett politiskt beslut att införa biometriska kännetecken i EU-pass utan att först inhämta råd från de som skall tillämpa beslutet, och utan att skaffa sig en uppfattning om problemets omfattning, om det nu föreligger ett problem.
Under alla omständigheter räcker det i detta skede med ett kännetecken, ansiktsbilden.
Skäl 2a (nytt)
Motivering
Eftersom syftet med biometriska uppgifter i pass måste vara uttryckligt, lämpligt, proportionerligt och tydligt måste det anges i lagtexten.
Ändringsförslag 3
Skäl 3
(3) Harmoniseringen av säkerhetsdetaljer och införandet av biometriska kännetecken är ett viktigt steg i användningen av nya element mot bakgrund av utvecklingen på EU-nivå för att göra resehandlingar säkrare och skapa en mer tillförlitlig koppling mellan innehavaren och passet, och därigenom hindra att passet används i bedrägligt syfte.
Specifikationerna i Internationella civila luftfartsorganisationens (ICAO) dokument nr 9303 om maskinläsbara resehandlingar bör beaktas.
(3) Harmoniseringen av säkerhetsdetaljer och införandet av biometriska kännetecken är ett viktigt steg i användningen av nya element mot bakgrund av utvecklingen på EU-nivå för att göra resehandlingar säkrare och skapa en mer tillförlitlig koppling mellan innehavaren och passet, och därigenom hindra att passet används i bedrägligt syfte.
Motivering
Det bör inte förekomma någon hänvisning till dokument nr 9303 i en EU-förordning eftersom dokumentet ändras kontinuerligt på ett sätt som inte inbjuder till insyn och som saknar demokratisk legitimitet.
Ändringsförslag
4
Skäl 7
Det måste säkerställas att inga andra uppgifter lagras i passet om det inte föreskrivs i förordningen eller dess bilagor eller anges i den aktuella resehandlingen .
Inga andra uppgifter bör lagras i passet.
Motivering
Det måste göras helt klart exakt vilka uppgifter som skall lagras i passet, och det bör inte finnas någon bestämmelse om att andra uppgifter skall lagras.
Ändringsförslag 5
2.
Medlemsstaterna får även inkludera fingeravtryck i driftskompatibla format.
2.
Passet skall vara försett med ett väl skyddat lagringsmedium som har tillräcklig kapacitet och som kan säkra de lagrade uppgifternas integritet, tillförlitlighet och konfidentialitet.
Det skall innehålla en ansiktsbild.
Medlemsstaterna får även inkludera fingeravtryck i driftskompatibla format.
Ingen central databas för Europeiska unionens pass och resehandlingar får upprättas som innehåller biometriska och andra uppgifter om samtliga innehavare av EU ‑pass.
Motivering
De tekniska specifikationerna är av avgörande betydelse för skyddet av privatlivet.
Därför bör vissa av de kriterier som de har att uppfylla nämnas särskilt.
Upprättandet av en central databas skulle strida mot såväl ändamåls- som proportionalitetsprincipen.
Det skulle dessutom öka risken för missbruk och ”function creep”(användning av datauppgifter i andra syften än det som ligger till grund för att de samlats in), liksom risken att biometriska kännetecken används som accesskoder till olika databaser varigenom uppgifter i dessa därmed kan sammanställas.
Ändringsförslag 6
1.
1.
Kompletterande tekniska specifikationer för passet som rör följande skall fastställas i enlighet med det förfarande som anges i artikel 5 :
Motivering
Artikel 2, punkt 1, led b
(b) Tekniska specifikationer för lagringsmediet för de biometriska uppgifterna och skyddet av dessa.
(b) Tekniska specifikationer för lagringsmediet för de biometriska uppgifterna och skyddet av dessa , i synnerhet för att trygga uppgifternas integritet, tillförlitlighet och konfidentialitet och säkra att de utnyttjas i enlighet med de ändamål som fastställs i denna förordning .
Motivering
1a.
Lagringsmediet får endast användas av
a) de myndigheter i medlemsstaterna som är behöriga att ta del av, lagra, ändra och stryka uppgifter, och
b) godkända organ som enligt lag har rätt att ta del av uppgifterna, i syfte att ta del av uppgifterna.
Motivering
Det bör framgå tydligt av lagtexten vilka myndigheter som skall ha tillgång till uppgifterna.
Otillåten tillgång är inte acceptabelt med hänsyn till skyddet av privatlivet.
2a.
Varje medlemsstat skall upprätta en förteckning över behöriga myndigheter samt över organ med behörighet enligt artikel 2.1 a.
Denna skall i sin tur upprätthålla en aktuell online förteckning över uppgifterna i fråga, och årligen offentliggöra en sammanställning av de nationella förteckningarna.
Motivering
För att se till att det råder vederbörlig insyn och öppenhet och därmed skydda mot missbruk bör enligt vad som föreslås här en förteckning upprättas över de myndigheter i medlemsstaterna som har behörighet att ta del av, lagra, ändra och radera uppgifter (såsom passmyndigheter) och de organ som har behörighet att ta del av dessa uppgifter (såsom gränsskyddsmyndigheter).
Ändringsförslag
10
1.
Utan att det påverkar bestämmelserna om skydd av personuppgifter, har personer till vilka pass utfärdas rätt att kontrollera personuppgifterna i passet och begära att få uppgifter rättade eller strukna.
1.
Utan att det påverkar bestämmelserna om skydd av personuppgifter, har personer till vilka pass utfärdas rätt att kontrollera personuppgifterna i passet och begära att få uppgifter rättade eller strukna.
Varje kontroll, rättelse eller strykning av dessa uppgifter skall utföras kostnadsfritt av den utsedda nationella myndigheten.
Motivering
Passinnehavaren skall alltid ha rätt att kontrollera, rätta eller stryka felaktiga uppgifter, och alla korrigeringar skall vara kostnadsfria.
Ändringsförslag
11
2.
Uppgifter i maskinläsbar form får inte finnas i passet, om inte annat följer av förordningen eller bilagan till denna eller anges i passet.
2.
Uppgifter i maskinläsbar form får inte finnas i passet, om inte annat följer av förordningen eller bilagan till denna eller anges i passet.
Inga ytterligare uppgifter får finnas i passet.
Motivering
Det måste göras helt klart exakt vilka uppgifter som skall lagras i passet, och det bör inte finnas någon bestämmelse om att andra uppgifter skall lagras.
2a.
De biometriska uppgifterna i pass skall endast utnyttjas för att kontrollera
a) dokumentets äkthet,
b) innehavarens identitet genom direkt tillgängliga jämförbara uppgifter när pass skall framläggas enligt lag.
Motivering
Eftersom syftet med att införa biometriska uppgifter i pass måste vara uttryckligt, lämpligt, proportionerligt och tydligt måste det anges i lagtexten.
Det får inte råda minsta tvivel om att dessa uppgifter endast får användas för att bekräfta dokumentets äkthet och innehavarens identitet.
2b.
Medlemsstaterna skall regelbundet översända granskningsrapporter om genomförandet av denna förordning till kommissionen, på grundval av gemensamt överenskomna standarder, särskilt vad gäller regler som begränsar de syften för vilka uppgifterna får användas och de organ som kan få tillgång till uppgifterna.
De skall även informera kommissionen om alla problem som uppkommer vid tillämpningen av denna förordning samt utbyta goda metoder med kommissionen och med varandra.
Motivering
Det är mycket viktigt att det finns ett effektivt kontrollnät för att man skall kunna skapa förtroende för biometriska metoder.
Ändringsförslag
14
3a.
Kommittén skall bistås av experter som utses av den arbetsgrupp som instiftats genom artikel 29 i direktiv 95/46/EG.
Motivering
De tekniska specifikationerna är av största vikt eftersom det är de som avgör huruvida införandet av biometriska uppgifter i pass kommer att tjäna sitt syfte och därtill trygga det fysiska uppgiftsskyddet.
De experter som granskar de tekniska specifikationerna ur uppgiftsskyddssynpunkt bör ha möjlighet att delta i den tekniska kommitténs arbete, och således även ge råd om vilka eventuella tekniska lösningar som är bäst sett till uppgiftsskyddet.
I slutändan bör de ha möjlighet att utvärdera de tekniska specifikationerna ur denna synvinkel.
Ändringsförslag
15
3b.
Motivering
Ändringsförslag
16
3c.
Kommissionen skall översända sitt förslag till beslut till Europaparlamentet, som inom tre månader kan anta en resolution genom vilken det motsätter sig förslaget till beslut om de tekniska specifikationerna.
Motivering
Ändringsförslag
17
3d.
Kommissionen skall informera Europaparlamentet om de åtgärder som den har för avsikt att vidta med hänsyn till Europaparlamentets resolution samt om sina skäl till detta.
Motivering
Ändringsförslag
18
3e.
Specifikationernas konfidentialitet skall säkras.
Motivering
Ändringsförslag
19
2.
För att denna förordning skall kunna tillämpas måste de nationella dataskyddsmyndigheterna intyga att de har de undersökande befogenheter och de resurser som krävs för att genomföra direktiv 95/46/EG när det gäller uppgifter som inhämtats i enlighet med detta.
Medlemsstaterna skall börja tillämpa denna förordning senast 18 månader efter antagandet av de åtgärder som avses i artikel 2.
Motivering
Ett stort antal medlemsstater anser det vore bättre om förordningen tillämpades 18 till 24 månader efter det att den antas.
Valet av 18 månader är därför en godtagbar kompromiss som även Förenta staterna bör respektera genom att förlänga tidsfristen för inresa utan visumhandlingar för resande med biometriska pass till ett datum senare än den 26 oktober 2005.
MOTIVERING
Som följd av den senaste tidens terroristattentat har olika uppmaningar gjorts runt om i världen om att förbättra dokumentsäkerheten.
Händelseutvecklingen har tjänat som en impuls för att ge ytterligare en skjuts åt det arbete med att introducera användningen av biometriska uppgifter som pågår på olika håll.
Tekniska utskott vid Internationella civila luftfartsorganisationen (ICAO) godkände under 2003 rekommendationer i denna riktning (ICAO:s ”Blueprint”).
I fråga om pass föreslog ICAO bland annat att man överallt i världen bör utnyttja maskinell ansiktsigenkänning som hjälpmedel för att bekräfta resandes identitet, och att de uppgifter som krävs för detta bör lagras på en kontaktlös integrerad krets (”chips”) med kapacitet på minst 32 kbyte.
Fingeravtryck och/eller inskannade irisbilder anges som eventuellt kompletterande kännetecken.
En annan impuls som drivit denna utveckling framåt har varit vissa amerikanska beslut om, i första hand, undantag från krav på visering (visa waiver programme, VWP
Genom VWP får medborgare från vissa länder resa in i Förenta staterna utan visum.
Deltagarna i programmet består av EU:s gamla medlemsstater (med undantag för Grekland) och, bland de nya medlemsstaterna, Slovenien. ).
Förenta staterna har fastställt att länder som gör anspråk på undantag från krav på visering eller förlängning av ett sådana undantag senast den 26 oktober 2004 skall ha infört ett program för att till sina medborgare kunna utfärda maskinläsbara pass som inte kan manipuleras och som innehåller biometriska kännetecken som uppfyller Internationella civila luftfartsorganisationens (ICAO) normer.
”Enhanced Border Security and Visa Entry Reform Act” från 2002, Sec.
303(b)(3).
Då det blev uppenbart att inget land skulle hinna uppfylla dessa krav inom den fastställda tidsfristen undertecknade president Bush en lag om att förlänga fristen med ett år.
H.R 4417 av den 9 augusti 2004.
På EU nivå kom ytterligare en impuls i form av Europeiska rådets slutsatser om att kommissionen bör lägga fram förslag om införande av biometriska uppgifter.
Vid sitt möte i Thessaloniki den 19–20 juni 2003 bekräftade Europeiska rådet att det behövs ”en enhetlig strategi inom EU vad gäller biometriska igenkänningstecken eller biometriska data, vilket skulle resultera i harmoniserade lösningar i fråga om tredjelandsmedborgares resehandlingar, EU-medborgares pass och informationssystem (VIS och SIS II)”.
Europeiska rådet har upprepat betydelsen av detta vid ett flertal tillfällen, bland annat vid sitt möte i Bryssel den 16–17 oktober 2003 där det med tillfredsställelse noterar ”det arbete som pågår inom unionen och internationella organ (ICAO, G8) för att införa biometriska kännetecken i viseringar, uppehållstillstånd och pass”.
II.
Föreliggande förslag
Syftet med föreliggande förslag är att göra passen säkrare genom att införa harmoniserade och rättsligt bindande säkerhetsdetaljer i EU-pass och att införa biometriska kännetecken i passen.
Till skillnad från kommissionens förslag om visumhandlingar och uppehållstillstånd föreslås här att endast ett biometriskt kännetecken, ansiktsbilden, skall vara obligatoriskt.
Medlemsstaterna bör själva få bestämma om fingeravtryck skall tas med.
Detaljerade tekniska specifikationer skall fastställas genom kommittésystemet och på grundval av ett föreskrivande förfarande.
Enligt kommissionens förslag kommer medlemsstaterna åläggas att genomföra förordningen ett år efter det att dessa specifikationer fastställts.
I sin motivering antyder kommissionen att det på längre sikt vore möjligt att upprätta ett centralt register för EU-pass.
III.
Föredragandens ståndpunkt
Föredraganden är över lag positiv till kommissionens förslag.
Han anser att biometriska uppgifter faktiskt kan bidra till att göra våra identifieringshandlingar säkrare.
Införandet av biometriska uppgifter kommer att göra det mycket svårt att förfalska pass eftersom de biometriska uppgifterna utgör en garant för att en person som visar upp ett pass faktiskt är identisk med den som passet utfärdades till.
Eftersom pass även används i det dagliga livet och inte bara för att passera gränser utgör införandet av biometriska uppgifter dessutom en lösning på problemet med identitetsstöld.
När det gäller själva rättsakten anser han dock att innan några biometriska pass utfärdas måste ett antal villkor till skydd för medborgarnas rättigheter uppfyllas, både när det gäller de tekniska specifikationerna (som även inbegriper kostnadseffektiva och säkra lösningar på hur biometriska uppgifter skall insamlas, bearbetas, lagras och användas) och medlemsstaternas genomförande.
Ur uppgiftsskyddssynpunkt är användningen av biometriska uppgifter mycket känslig.
Alla nödvändiga skyddsåtgärder måste vidtas i enlighet direktivet om dataskydd.
Direktiv 95/46/EG.
Såsom fastställs i artikel 29-arbetsgruppens allmänna arbetsdokumentet om biometriska uppgifter
Vidare måste de uppgifter som insamlas vara adekvata och relevanta och inte får omfatta mer än vad som är nödvändigt med hänsyn till de ändamål för vilka de har samlats in och för vilka de senare behandlas”
När det gäller tillämpningen av dess två grundläggande principer anser föredraganden att syftet med införandet av biometriska uppgifter måste anges och avgränsas på ett tydligare sätt i lagtexten, och att det ännu återstå att fastställa vem som har rätt att använda dessa uppgifter.
Vad gäller syftet får det inte råda minsta tvivel om att dessa uppgifter ändats får användas i verifieringssyfte och under inga villkor i andra syften, exempelvis vid dold övervakning.
Föredraganden oroas särskilt över konsekvenserna på sikt om man i enlighet med vad kommissionen skisserar i sin motivering upprättar ett europeiskt register över utfärdade pass.
En sådan central databas behövs inte om syftet är att skapa ”en säkrare länk mellan innehavaren och passet”.
Därtill är risken för ”function creep” (användning av datauppgifter i andra syften än det som ligger till grund för att de samlats in) allt för stor.
Föredraganden uppmanar samtidigt medlemsstaterna att inte lagra dessa uppgifter i nationella databaser.
De biometriska uppgifterna bör endast lagras lokalt, i själva passet.
Som kommissionen konstaterar i sin motivering medför användningen av denna teknik dessutom en ökad arbetsbörda för de myndigheter som ansvarar för dataskyddet.
Föredraganden uppmanar medlemsstaterna att se till att dessa myndigheter tilldelas de resurser som krävs för att de skall kunna fullfölja de skyldigheter de ålagts enligt lag.
Det är utomordentligt viktigt att de tekniska lösningar man slutligen enas om, efter det att de tekniska specifikationerna utarbetats genom kommittéförfarandet, håller måttet.
Det är dessa specifikationer som avgör om användningen av biometriska uppgifter i pass lyckas eller inte, och som garanterar uppgifternas fysiska säkerhet.
Se artikel 17 i dataskyddsdirektivet.
Föredraganden föreslår därför vissa ändringar i förslaget varigenom ytterligare några kriterier för det tekniska genomförandet anges.
Dessa avser en rad olika hänsyn på åtminstone tre områden: För det första, för att medborgarnas personuppgifter skall kunna skyddas måste det finnas ett adekvat skydd mot otillbörlig tillgång.
Vissa påstår att ett chips kan läsas på relativt långt håll, andra att ett chips med kapacitet motsvarande ISO-norm 14443 endast kan läsas på ett avstånd av 10–15 cm.
För det andra måste man se till att chipset är väl skyddat mot oavsiktlig skada och att det har en ”livstid” motsvarande dagens pass (som ofta har en giltighetstid på 10 år).
För det tredje måste det finnas garantier för att det chips som ligger inbakat i passet inte skapar interferens med chips i visumhandlingar som fästs i passet.
Föredraganden vill i detta sammanhang understryka vikten av att ge de tekniska experterna tid att hitta rätta lösningar.
Den tekniska utvecklingen öppnar dörren för lösningar som till och med kan göra chipset överflödigt ur såväl säkerhets- som kostnadssynpunkt.
Ett exempel på en sådan lösning är ett system med digitaliserade passfoton och fingeravtryck i kombination med en streckkodad digitalsignatur som krypterats med öppen nyckel.
Det vore knappast till hjälp om EU i hast valde att rikta in sig på vad som i dagsläget uppfattas som en given lösning endast för att i ett senare skede upptäcka att man inte förberett sig tillräckligt, eller att lösningen i fråga i allt för hög grad är beroende av föråldrad teknik.
Ett sådant handlande skulle endast bidra till att undergräva medborgarnas förtroende.
Eftersom de tekniska specifikationerna är av avgörande för graden av dataskydd föreslår föredraganden att de experter som granskar dessa specifikationer utifrån ett dataskyddsperspektiv även bör ges tillfälle att delta i utformningen av dem.
I slutändan bör de har möjlighet att utvärdera specifikationerna utifrån detta perspektiv och, i den mån det krävs, begära att arbetet med att fina lösningar på återstående problem får fortsätta.
Utöver de noggranna förberedelser som medlemsstaterna måste göra för att fastställa dessa tekniska specifikationer uppmanar föredraganden dem att fortsätta testa de tekniska lösningarna i det verkliga livet och i bred skala, innan de utfärdar nya pass.
Detta skulle även främja förtrogenheten med denna relativt nya teknik.
Det sätt på vilket medlemsstaterna väljer att genomföra de nya bestämmelserna kommer att avgöra om införandet av biometriska uppgifter blir framgångsrikt eller ej.
Föredraganden betonar att det kommer an på medlemsstaterna att se till att i god tid ge medborgarna uttömmande information om dessa nya rutiner liksom att tillhandahålla en högkvalitativ utbildning åt alla som har att verkställa dem i dess olika steg (från inläsning till övervakning och kontroll).
Vad som i slutändan är viktigast är behovet att under alla omständigheter värna om oskyldiga medborgares integritet i en atmosfär där ”misstag inte kan förekomma”.
Det måste finnas garantier för att medborgare som utsätts för felaktiga avvisanden vid gränskontroller underrättas om skälen till att de avvisas och om hur denna situation så snabbt som möjligt kan redas ut och åtgärdas.
RESERVATION
Ole Krarup, Sylvia-Yvonne Kaufmann, Mary Lou McDonald och Giusto Catania
Av flera anledningar motsätter vi oss tanken att införa biometriska kännetecken i identitetshandlingar:
För det första är vi allvarligt oroade över de enorma risker de extremt stora databaserna kommer att innebära för uppgiftsskyddet och skyddet av privatlivets helgd.
Riskerna i samband med lagring, tillträde till och överföring av uppgifter har inte undanröjts, och faran för identitetsstöld och missbruk kvarstår även om uppgifterna endast lagras på ett mikrochip.
Frågorna kring multipla identiteter, avlyssning av dataöverföringar och proaktiv övervakning har ännu inte lösts.
Biometriska system är aldrig hundraprocentigt säkra, och för flera hundra tusen människor i EU kommer inte ens fingeravtrycken vara helt tillförlitliga.
För det andra strider förslaget mot alla vedertagna standarder för lämplighet och subsidiaritet.
Hittills har varken kommissionen eller rådet på ett fullgott sätt redogjort för behovet, funktionen eller effektiviteten av eller de sannolika bieffekterna av att införa biometriska kännetecken i identitetshandlingar.
De har inte ens lagt fram någon detaljerad beräkning över de förväntade kostnaderna eller föreslagit en tydlig budget!
Till sist, biometriska metoder ökar inte säkerheten, eftersom de inte binder en person till en verklig identitet, utan bara till en identitet som fastställts genom en identitetshandling.
Om passet är falskt kan det biometriska kännetecknet som ingår i det ändå inte ändra på detta.
Framtida brottslingar kommer därför fortfarande att kunna låta sig registreras i alla tillgängliga databaser under falsk identitet och passera de framtida kontrollerna okontrollerade, vilket kommer att leda till att världen blir osäkrare istället för säkrare.
Framtida terrorister som är beredda att kasta bort sina liv kommer att vara beredda till detta, även om de därmed anger sin verkliga identitet.
ÄRENDETS GÅNG
Titel
Komissionens förslag till rådets förordning om standarder för säkerhetsdetaljer och biometriska kännetecken i EU-medborgarnas pass
Referensnummer
Kom(2004)0116 – C5-0101/2004 – 2004/0039(CNS)
Rättslig grund
Grund i arbetsordningen
Begäran om samråd med parlamentet
LIBE
Rådgivande utskott
Tillkännagivande i kammaren
Inget yttrande avges
Beslut
Förstärkt samarbete
Tillkännagivande i kammaren
Föredragande
Carlos Coelho
Utnämning
Tidigare föredragande
Förenklat förfarande
Beslut
Bestridande av den rättsliga grunden
JURI:s yttrande
Ändrad anslagstilldelning
BUDG:s yttrande
Samråd med Europeiska ekonomiska och sociala kommittén
Beslut i kammaren
Samråd med Regionkommittén
Beslut i kammaren
Behandling i utskott
Antagande
för:
26
emot:
9
nedlagda röster:
Slutomröstning: närvarande ledamöter
Alexander Nuno Alvaro, Roberta Angelilli, Edit Bauer, Kathalijne Maria Buitenweg, Giusto Catania, Charlotte Cederschiöld, Carlos Coelho, António Costa, Agustín Díaz De Mera García Consuegra, Antoine Duquesne, Kinga Gál, Lilli Gruber, Timothy Kirkhope, Ewa Klamt, Wolfgang Kreissl-Dörfler, Barbara Kudrycka, Stavros Lambrinidis, Henrik Lax, Sarah Ludford, Edith Mastenbroek, Jaime Mayor Oreja, Claude Moraes, Athanasios Pafilis, Lapo Pistelli, Martine Roure, Michele Santoro, Luciana Sbarbati, Inger Segelström, Ioannis Varvitsiotis, Manfred Weber, Stefano Zappalà, Tatjana Ždanoka
Slutomröstning: närvarande suppleanter
Frederika M.J. Brepoels, Gérard Deprez, Luis Francisco Herrero-Tejedor, Sophia Helena In 't Veld, Jean Denise Lambert, Vincent Peillon, Antonio Tajani
Slutomröstning: närvarande suppleanter (art.
178.2)
Ingivande – A6
Anmärkningar
SLUTLIG VERSION
A6-0033/2005
***I
BETÄNKANDE
om förslaget till Europaparlamentets och rådets förordning om statistik över yrkesutbildning på företag
(KOM(2004)0095 – C5‑0083/2004 – 2004/0041(COD))
Utskottet för sysselsättning och sociala frågor
Föredragande:
Ottaviano Del Turco
PE 349.855v02-00
Teckenförklaring
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................13
ÄRENDETS GÅNG..................................................................................................................15
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till Europaparlamentets och rådets förordning om statistik över yrkesutbildning på företag
( KOM(2004)0095 – C5‑0083/2004 – 2004/0041(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2004)0095 )
EUT C 98, ,
– med beaktande av artikel 51 i arbetsordningen,
– med beaktande av betänkandet från utskottet för sysselsättning och sociala frågor ( A6‑0033/2005 ).
Kommissionens förslag
Parlamentets ändringar
Ändringsförslag
1
Skäl 5a (nytt)
(5a) Denna förordning följer den definition av ”mindre gynnade personer på arbetsmarknaden” som ges i riktlinjerna för medlemsstaternas sysselsättningspolitik.
Motivering
Enligt riktlinjerna för medlemsstaternas sysselsättningspolitik är mindre gynnade personer ”personer som har särskilda svårigheter på arbetsmarknaden, till exempel personer som tidigt avbrutit sin utbildning, lågutbildade arbetstagare, funktionshindrade personer, invandrare och etniska minoriteter”.
Ändringsförslag
2
Skäl 7
(7) Särskild vikt måste fästas vid utbildning på arbetsplatsen som en väsentlig aspekt på det livslånga lärandet.
(7) Särskild vikt måste fästas vid utbildning som sker på arbetsplatsen och under arbetstid, bägge två väsentliga aspekter på det livslånga lärandet.
Motivering
Ändringsförslag
3
Skäl 13
(13) De åtgärder som krävs för genomförandet av denna förordning bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter.
(13) De åtgärder som krävs för genomförandet av denna förordning bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter.
I dessa åtgärder bör man beakta medlemsstaternas kapacitet att samla in och behandla uppgifter.
Ändringsförslag
4
(c) den andra undersökningen om yrkesinriktad fortbildning (CVTS2): den andra europeiska undersökningen av yrkesinriktad fortbildning på företag som utfördes 2000–2001 i alla medlemsstater med 1999 som referensår.
utgår
Motivering
Detta ändringsförslag är nödvändigt med tanke på ändringsförslag 12 som gäller strykning av bilagan om bruttourval.
Ändringsförslag
5
(c) Arbetsmarknadens parters roll för tillhandahållandet av adekvat yrkesinriktad fortbildning på arbetsplatsen.
(c) Arbetsmarknadens parters roll för tillhandahållandet av yrkesinriktad fortbildning på arbetsplatsen i alla dess aspekter .
Motivering
Denna ändring i förslaget till förordning tjänar till att undanröja en rent godtycklig bedömning som är svår att kvantifiera i en statistisk analys.
Genom ändringsförslaget vill man dock säkerställa arbetsmarknadsparternas roll i tillhandahållandet av yrkesinriktad fortbildning på arbetsplatsen i alla dess aspekter.
Ändringsförslag
6
(fa) Offentliga åtgärders inverkan på yrkesinriktad fortbildning på företag.
Motivering
Genom detta tillägg inkluderas inverkan av offentliga åtgärder i analysen av yrkesinriktad fortbildning.
På så sätt kan man undersöka med vilka medel yrkesutbildningen finansieras.
Ändringsförslag
7
(g) Lika möjligheter till yrkesinriktad fortbildning på företag för alla anställda, särskilt med avseende på kön.
(g) Lika möjligheter till yrkesinriktad fortbildning på företag för alla anställda, särskilt med avseende på kön och särskilda åldersgrupper .
Ändringsförslag
8
(ha) Yrkesutbildningsåtgärder avsedda för olika former av anställningskontrakt.
Motivering
Detta tillägg syftar till att uppdatera undersökningen och ta med de olika nya formerna av anställningskontrakt i analysen av yrkesutbildning.
Ändringsförslag
9
(j) Utvärdering av yrkesinriktad fortbildning på företag .
(j) Företagens förfaranden för utvärdering och övervakning av yrkesinriktad fortbildning.
Motivering
Dessa ändringar i förslaget till förordning tjänar till att undanröja en rent godtycklig bedömning som är svår att kvantifiera i en statistisk analys.
Det är sålunda lämpligare att analysera metoderna för utvärdering och övervakning av yrkesutbildning.
Övervakningen intar dessutom en särskilt viktig roll när det gäller att undersöka utbildningens effektivitet.
Ändringsförslag
10
Medlemsstaterna får, med beaktande av den specifika nationella storleksfördelningen för företag och utvecklingen av politiska behov, utvidga definitionen av en statistisk enhet i sitt land.
Kommissionen får också besluta att utvidga denna definition i enlighet med det förfarande som anges i artikel 14, om en sådan utvidgning väsentligt skulle förbättra representativiteten hos och kvaliteten på undersökningens resultat i de berörda medlemsstaterna.
Motivering
Detta tillägg behövs för att man skall kunna inbegripa företag med mindre än 10 anställda i förordningen då de specifika ekonomiska förhållandena i landet kräver detta.
Enligt uppgifter från Eurostat utgör företag med mindre än 10 anställda i genomsnitt 90 procent av företagen i det utvidgade EU och de sysselsätter 27,49 procent av arbetskraften.
I Italien t.ex. har till och med 96,85 procent av företagen mindre än 10 anställda och de sysselsätter hela 57,65 procent av arbetskraften.
Genom ändringsförslaget vill man alltså ge medlemsstaterna möjlighet att utvidga definitionen av en statistisk enhet i sina respektive länder, om de så önskar, och ge kommissionen möjlighet att fatta beslut om att utvidga denna definition i enlighet med det förfarande som anges i artikel 14.
Ändringsförslag
11
2.
I samband med undersökningen uppmanas företagen att lämna korrekta och fullständiga uppgifter inom angiven tid.
2.
I samband med undersökningen uppfordras företagen att lämna korrekta och fullständiga uppgifter inom angiven tid.
Motivering
Ändringsförslaget syftar till att förplikta och inte enbart uppmana företagen att lämna korrekta och fullständiga uppgifter inom angiven tid.
Ändringsförslag
12
3.
Medlemsstaterna får bestämma att det skall vara obligatoriskt för företagen att besvara undersökningen.
I samband med en obligatorisk undersökning skall de undersökta företagen åläggas att lämna korrekta och fullständiga uppgifter inom angiven tid.
3.
Medlemsstaterna skall bestämma på vilket sätt företagen skall besvara undersökningen.
Motivering
Syftet med ändringsförslaget är att göra det till medlemsstaternas plikt att ålägga företagen att besvara undersökningen.
Det ger dock de enskilda länderna friheten att bestämma på vilket sätt företagen skall besvara undersökningen.
Ändringsförslag
13
1.
Undersökningen skall vara en urvalsundersökning.
Urvalens storlek skall likna dem som användes under CVTS2, vilka anges i bilagan.
1.
Undersökningen skall vara en urvalsundersökning.
Motivering
Detta ändringsförslag är nödvändigt med tanke på ändringsförslag 12 som gäller strykning av bilagan om bruttourval.
Ändringsförslag
14
3.
Krav på urval och precision samt specifikationer av NACE- och storlekskategorier på vilka resultaten skall kunna uppdelas skall bestämmas av kommissionen i enlighet med det förfarande som anges i artikel 14.
3.
Krav på urval och precision och de urvalsstorlekar som behövs för att dessa krav skall uppfyllas samt specifikationer av NACE- och storlekskategorier på vilka resultaten skall kunna uppdelas skall bestämmas av kommissionen i enlighet med det förfarande som anges i artikel 14.
Motivering
Detta tillägg är nödvändigt med tanke på ändringsförslag 12 som gäller strykning av bilagan om bruttourval.
Urvalens storlek skall bestämmas av kommissionen, som biträds av Kommittén för det statistiska programmet, i enlighet med det förfarande som fastställs i artikel 14 i detta förslag till förordning.
Ändringsförslag
15
(Berör inte den svenska versionen.)
(Berör inte den svenska versionen.)
Motivering
(Berör inte den svenska versionen.)
Ändringsförslag
17
3.
Kommissionen (Eurostat) skall bedöma de överlämnade uppgifternas kvalitet.
3.
Ändringsförslag
18
Bilaga
Bruttourval, avrundade, i CVTS2
utgår
Land
Urval, brutto (avrundat)
Motivering
Bilagan är inte uppdaterad: den inbegriper nämligen inte de nya medlemsstaterna och bruttourvalen baserar sig på den andra CVTS-undersökningen som utfördes 2000–2001.
Därför föreslås att bilagan stryks och att man överlåter åt kommissionen, som biträds av Kommittén för det statistiska programmet, att bestämma urvalens storlek i de enskilda medlemsländerna (jfr ändringsförslag 11).
MOTIVERING
Tanken om livslångt lärande är en hörnsten i den europeiska sysselsättningsstrategin (vilket bl.a. betonades redan vid Europeiska rådets möte i Lissabon 2000) och har införlivats i alla medlemsstaters nationella handlingsplaner.
Det är dock nödvändigt att man vid sidan om det allmänna politiska engagemanget för en sådan politik koncentrerar ansträngningarna på att uppnå en effektiv tillämpning och uppföljning av dessa åtaganden.
De statistiska uppgifterna ger en oroväckande bild: år 1998 deltog totalt 8 procent av de anställda i fortbildningsprojekt, medan denna andel endast ökat till 8,5 procent i slutet av 2003.
Dessa siffror, som enbart hänför sig till ett EU med 15 medlemsländer, är dessutom irrelevanta om de relateras till det utvidgade EU.
En europeisk rättslig grund för insamling av jämförbara uppgifter som kan förmedla en verklighetstrogen bild av yrkesinriktad fortbildning måste ses som en av de viktigaste faktorerna när det gäller att märkbart öka EU:s engagemang för en effektiv uppföljning av denna politik.
Därför anser föredraganden det vara nödvändigt att göra det föreliggande förslaget till förordning så precist och bindande som möjligt .
II.
Förordning om statistik över yrkesutbildning på företag
Genom denna förordning upprättas en gemensam ram för sammanställning av gemenskapsstatistik över yrkesutbildning på företag.
Den första företagsundersökningen avseende yrkesinriktad fortbildning (CVTS1) genomfördes 1994.
Undersökningen var en del av handlingsprogrammet för utveckling av yrkesinriktad fortbildning i Europeiska gemenskapen (FORCE) i enlighet med rådets beslut 90/267/EEG av den 29 maj 1990.
Den andra undersökningen (CVTS2) utfördes 2000–2001 i alla medlemsstater samt i Norge och i nio kandidatländer.
Både CVTS1 och CVTS2 genomfördes enligt ”gentlemen’s agreements” mellan Eurostat och EU:s medlemsstater.
Efter CVTS2 beslöt Eurostat och EU:s medlemsstater att införa en rättslig grund för insamlingen av uppgifter inom det europeiska statistiska systemet i form av en förordning från Europaparlamentet och rådet.
Eftersom CVTS är den enda källan till internationell statistik över yrkesinriktad fortbildning på företag syftar denna förordning till att införa regelbunden insamling av uppgifter om utbildning på företag inom ramen för det europeiska statistiksystemet.
Enligt föreliggande förslag bör man särskilt utarbeta en metod som kan sätta samarbetet med företagen i medlemsstaterna på en stabil grund och förbättra uppgifternas kvalitet och fullständighet.
III.
Kommentar till de ändringsförslag som föredraganden lagt fram
Föredraganden välkomnar medlemsstaternas och Eurostats politiska beslut att införa en rättslig grund för insamlingen av uppgifter om yrkesutbildning på företag i form av en förordning från Europaparlamentet och rådet.
Föredraganden är även medveten om vikten av att denna förordning snabbt kan träda i kraft eftersom den bidrar till att sätta samarbetet med företagen i medlemsstaterna på en stabil grund och förbättra uppgifternas kvalitet och fullständighet.
Föredraganden anser det dock vara nödvändigt att lägga fram några ändringsförslag i syfte att göra förordningen verkligt bindande för företagen i alla medlemsstater och se till att den med största möjliga precision kan återspegla den reella situationen när det gäller yrkesutbildning på företag.
Ändringsförslagen gäller huvudsakligen
ü en önskan att göra det till medlemsstaternas plikt att ålägga företagen att besvara undersökningen, samtidigt som de enskilda länderna ges friheten att bestämma på vilket sätt företagen skall besvara undersökningen,
ü en önskan att inbegripa företag med mindre än 10 anställda i förordningen då de specifika ekonomiska förhållandena i landet kräver detta; enligt uppgifter från Eurostat utgör företag med mindre än 10 anställda i genomsnitt 90 procent av företagen i det utvidgade EU och de sysselsätter 27,49 procent av arbetskraften; i vissa länder, t.ex.
Frankrike, Belgien, Finland, Portugal, Spanien, Sverige, Ungern, Polen, Tjeckien, Malta och Italien, är dock denna procentsats större; i Italien t.ex. har till och med 96,85 procent av företagen mindre än 10 anställda och de sysselsätter hela 57,65 procent av arbetskraften,
ü en önskan att uppdatera undersökningen och ta med de olika nya formerna av anställningskontrakt i analysen av yrkesutbildning,
ü en önskan att inkludera inverkan av offentliga åtgärder i analysen av yrkesinriktad fortbildning,
ü en önskan att stryka den icke uppdaterade bilagan.
Denna inbegriper nämligen inte de nya medlemsstaterna och bruttourvalen baserar sig på den andra CVTS-undersökningen som utfördes 2000–2001.
ÄRENDETS GÅNG
Titel
Förslaget till Europaparlamentets och rådets förordning om statistik över yrkesutbildning på företag
Referensnummer
KOM(2004)0095 – C5‑0083/2004 – 2004/0041(COD)
Rättslig grund
art.
251.2 och art.
Grund i arbetsordningen
Framläggande för parlamentet
Föredragande Utnämning
Tidigare föredragande
Förenklat förfarande Beslut
Bestridande av den rättsliga grunden JURI:s yttrande
Ändrad anslagstilldelning BUDG:s yttrande
Behandling i utskott
Antagande
för:
emot:
nedlagda röster:
22
1
Slutomröstning: närvarande ledamöter
Jan Andersson, Philip Bushill-Matthews, Ole Christensen, Derek Roland Clark, Ottaviano Del Turco, Harald Ettl, Richard Falbr, Ilda Figueiredo, Stephen Hughes, Jan Jerzy Kułakowski, Sepp Kusstatscher, Jean Lambert, Elizabeth Lynne, Mary Lou McDonald, Thomas Mann, Jiří Maštálka, Ana Mato Adrover, Csaba Őry, Jacek Protasiewicz, Anne Van Lancker, Gabriele Zimmer
Slutomröstning: närvarande suppleanter
Jamila Madeira, Dimitrios Papadimoulis, Leopold Józef Rutowicz, Eva-Britt Svensson, Georgios Toussas
Slutomröstning: närvarande suppleanter (art.
178.2)
Ingivande – A[6]-nummer
Anmärkningar
...
SLUTLIG VERSION
A6-0123/2005
***I
BETÄNKANDE
om förslaget till Europaparlamentets och rådets förordning om internationella tågresenärers rättigheter och skyldigheter
(KOM(2004)0143 – C6‑0003/2004 – 2004/0049(COD))
Utskottet för transport och turism
Föredragande:
Dirk Sterckx
PE 347.287v02-00
Teckenförklaring
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................57
ÄRENDETS GÅNG..................................................................................................................61
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till Europaparlamentets och rådets förordning om internationella tågresenärers rättigheter och skyldigheter
( KOM(2004)0143 – C6‑0003/2004 – 2004/0049(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
EUT C ... / Ännu ej offentliggjort i EUT. ,
– med beaktande av artikel 51 i arbetsordningen,
– med beaktande av betänkandet från utskottet för transport och turism ( A6‑0123/2005 ).
Kommissionens förslag
Parlamentets ändringar
Ändringsförslag
1
Titel
Motivering
Förordningen bör gälla även den nationella tågtrafiken.
Ändringsförslag
2
Skäl 1
(1) Inom ramen för den gemensamma transportpolitiken är det viktigt att slå vakt om tjänsternas kvalitet och de internationella tågresenärernas rättigheter, och att förbättra den internationella persontrafikens kvalitet och effektivitet för att bidra till en ökning av järnvägstrafikens andel i förhållande till andra transportsätt.
(1) Inom ramen för den gemensamma transportpolitiken är det viktigt att slå vakt om tjänsternas kvalitet och tågresenärernas rättigheter, och att förbättra persontrafikens kvalitet och effektivitet för att bidra till en ökning av järnvägstrafikens andel i förhållande till andra transportsätt.
Motivering
Dessa bestämmelser bör gälla även den nationella tågtrafiken.
Ändringsförslag
3
Skäl 2a (nytt)
(2a) Det gällande fördraget om internationell järnvägstrafik (COTIF) av den 9 maj 1980 omfattar enhetliga regler för avtal om internationell järnvägsbefordran av resande (CIV ‑bihang A i fördraget).
COTIF ‑fördraget ändrades genom Vilniusprotokollet av den 2 juni 1999.
I denna förordning bör det tas hänsyn till de bestämmelser som redan finns i CIV ‑bihang A till COTIF-fördraget.
Tillämpningsområdet bör dock utvidgas på ett sådant sätt att det inte enbart skyddar resenärer som färdas i internationell trafik, utan även resenärer i nationell trafik.
Med hänsyn till rättssäkerheten är det absolut nödvändigt att avstå ifrån att bestämmelser som redan ingår i CIV-bihangen övertas ordagrant i denna förordning.
Motivering
Förhållandet mellan CIV-bihanget och de rättigheter som föreskrivs i denna förordning preciseras inte klart genom att enbart hänvisa till detta bihang.
Ändringsförslag
4
Skäl 6
(6) Järnvägsföretag bör samarbeta för att underlätta övergången från ett nät till ett annat och från en verksamhetsutövare till en annan, och genom detta samarbete garantera att tågresenärerna får samordnade biljetter.
(6) Järnvägsföretag bör samarbeta för att underlätta övergången från ett nät till ett annat och från en verksamhetsutövare till en annan, och genom detta samarbete verka för att tågresenärerna får samordnade biljetter.
Motivering
Föredraganden föreslår att man byter ut resultatkravet mot ett krav på ansträngning.
Ändringsförslag
5
Skäl 7
(7) För att garantera att internationella tågresenärer kan dra nytta av de bestämmelser som fastställs i den här förordningen måste de järnvägsföretag som bedriver persontrafik samarbeta.
Detta samarbete bör på icke-diskriminerande basis vara öppet för alla järnvägsföretag som bedriver persontrafik.
(7) För att garantera att tågresenärer kan dra nytta av de bestämmelser som fastställs i den här förordningen måste de järnvägsföretag som bedriver persontrafik samarbeta.
Detta samarbete bör på icke-diskriminerande basis vara öppet för alla järnvägsföretag som bedriver persontrafik.
Motivering
Dessa bestämmelser bör gälla även den nationella tågtrafiken.
Ändringsförslag
6
Skäl 8
(8) Den internationella persontrafiken på järnväg bör gagna allmänheten.
Funktionshindrade personer bör därför, oavsett om deras nedsatta rörelseförmåga beror på handikapp, ålder eller andra faktorer, ha samma möjligheter som andra medborgare att resa med tåg.
(8) Den internationella persontrafiken på järnväg bör gagna allmänheten.
Samtliga resenärer, inbegripet funktionshindrade personer och andra resenärer med nedsatt rörelseförmåga, bör därför ha samma möjligheter som andra medborgare att resa med tåg utan att utsättas för diskriminering .
Motivering
[Första meningen i motiveringen berör inte den svenska versionen.]
Ändringsförslaget innebär dessutom att de rättigheter som gäller för funktionshindrade personer och andra personer med nedsatt rörelseförmåga understryks med större kraft.
Ändringsförslag
7
Skäl 8a (nytt)
(8a) Järnvägsföretag och stationsförvaltare skall alltid beakta alla tänkbara problem som kan uppstå för funktionshindrade personer, så att systematiska förbättringar kan åstadkommas i samband med inköp av ny rullande materiel, ombyggnad av stationer, inrättningar för information och assistans samt järnvägsnätets generella tillgänglighet.
Motivering
Skyldigheten att göra infrastruktur och rullande materiel mera lättillgängliga bör uttryckligen nämnas.
Vi kan visserligen inte begära att alla stationer har hiss ett år efter att denna förordning har trätt i kraft, men däremot att fullständig tillgänglighet för alla medborgare är en ledstjärna vid ombyggnationer eller inköp av nya tåg.
Ändringsförslag
8
Skäl 10
(10) Införandet av gränser för järnvägsföretagens ansvarighet vid förlust av eller skada på resgods och för skada som uppkommer på grund av försening, missad anslutning eller inställd trafik torde leda till ökad klarhet och införa incitament på den internationella persontrafikmarknaden som gagnar resenärerna.
(10) Införandet av gränser för järnvägsföretagens ansvarighet vid förlust av eller skada på resgods och för skada som uppkommer på grund av försening, missad anslutning eller inställd trafik torde leda till ökad klarhet och införa incitament på persontrafikmarknaden som gagnar resenärerna.
Motivering
Denna förordning bör gälla även den nationella tågtrafiken.
Ändringsförslag
9
Skäl 19
I enlighet med proportionalitetsprincipen i samma artikel går förordningen inte utöver vad som är nödvändigt för att uppnå dessa mål.
I enlighet med proportionalitetsprincipen i samma artikel går förordningen inte utöver vad som är nödvändigt för att uppnå dessa mål.
Motivering
Dessa bestämmelser bör gälla även den nationella tågtrafiken.
Ändringsförslag
10
-1.
Genom denna förordning genomförs vissa bestämmelser i det internationella COTIF-fördraget, och den innehåller dessutom ett antal kompletterande bestämmelser.
Motivering
Föredraganden vill i förordningen så långt som möjligt ansluta till bestämmelserna i COTIF‑fördraget, när dessa är lämpliga och i linje med kommissionens avsikter.
Att införliva dessa bestämmelser ger den fördelen att vi har en ram som genast kan tillämpas i 42 länder.
Förutom EU-länderna omfattar den också ett antal grannländer, såsom Norge och Schweiz.
När unionen har blivit medlem av COTIF kommer man att kunna påverka där.
Det är inte meningen att överta COTIF:s hela regelverk.
Denna förordning innehåller lämpliga kompletteringar på vissa punkter.
Ändringsförslag
11
1.
I denna förordning fastställs rättigheter och skyldigheter för internationella tågresenärer.
1.
I denna förordning fastställs rättigheter och skyldigheter för alla tågresenärer.
Ändringsförslag
12
Även i avtal om offentliga tjänster måste minst den miniminivå som fastställs i denna förordning garanteras.
Medlemsstater kan fastställa mera omfattande rättigheter inom ramen för nationell lagstiftning eller i avtal om offentliga tjänster.
Under en period på fem år från ikraftträdandet av denna förordning kan medlemsstaterna begära undantag från denna bestämmelse.
Ändringsförslag
13
2.
Förordningen skall vara tillämplig på internationella resor inom gemenskapen där den internationella trafiken bedrivs av ett järnvägsföretag som innehar tillstånd i enlighet med rådets direktiv 95/18/EG.
utgår
Motivering
Förordningen bör inte begränsas till att gälla endast internationella resor.
Ändringsförslag
14
3.
utgår
Motivering
Bokningssystem är ett av många teman i förordningen.
Det finns ingen anledning att explicit nämna just detta tema under rubriken Syfte och tillämpningsområde.
Ändringsförslag
15
1) järnvägsföretag: offentligt eller privat företag med tillstånd enligt gällande gemenskapslagstiftning vars huvudsakliga verksamhet består i att tillhandahålla tjänster för transport av resenärer på järnväg, med kravet att företaget måste tillhandahålla dragkraft.
1) järnvägsföretag: offentligt eller privat företag med tillstånd enligt gällande gemenskapslagstiftning vars verksamhet består i att regelbundet tillhandahålla tjänster för transport av resenärer på järnväg, med kravet att företaget måste tillhandahålla dragkraft.
Motivering
De föreslagna bestämmelserna skall tillämpas av samtliga järnvägsföretag som tillhandahåller persontrafik.
Av denna anledning är det missvisande om det kommer an på huruvida företaget ”huvudsakligen” ägnar sig åt persontrafik.
Denna definition förefaller att inrikta sig på vilket förhållande som råder mellan persontrafiken och godstrafiken.
Avgörande måste dock vara huruvida persontrafiken utförs regelbundet och inte enbart i undantagsfall eller tillfälligtvis.
Därför bör i detta sammanhang den definition användas som fastställs i direktiv 91/440.
Ändringsförslag
16
6) större järnvägsstation: en järnvägsstation med internationell trafik och/eller nationell fjärrtrafik som sträcker sig över mer än 100 kilometer .
6) större järnvägsstation: en järnvägsstation som p.g.a. trafikvolym, internationell karaktär och/eller geografiskt läge betecknas som sådan av den berörda medlemsstaten .
Motivering
Föredraganden är orolig för att de kriterier som kommissionen här anger inte alltid fungerar i praktiken.
Gemenskapens järnvägsnät kan inte skäras över en kam.
Internationella förbindelser stannar ibland vid riktigt små stationer som täcks av kommissionens definition, medan nationella stationer med stor resandevolym skulle falla utanför definitionen.
Därför föreslår föredraganden att medlemsstaterna själva får avgöra, enligt ett antal kriterier, vilka som är deras större järnvägsstationer.
Ändringsförslag
17
9a) abonnemang: ett transportavtal som ger innehavaren rätt att regelbundet resa under en viss period på en viss rutt.
Motivering
Denna definition behövs när denna förordnings tillämpningsområde utvidgas till att omfatta även den nationella tågtrafiken och rätten för innehavare av tågkort (abonnemang, o.dyl.) att få kompensation vid upprepade förseningar.
Ändringsförslag
18
10) bokning: innebär att resenären har en biljett eller annat bevis för att bokningen har accepterats och registrerats av järnvägsföretaget eller researrangören .
10) bokning: innebär ett avtal som ingås mellan en resenär och järnvägsföretag, i samband med vilket en biljett eller annat färdbevis utfärdas och tillhandahålls resenären.
Motivering
Bokningen ses i detta sammanhang som ”bevis” för att ett avtal ingåtts som är bindande för båda parter och att resenären förfogar över biljett eller annat färdbevis.
Begreppet i sig säger dock inget om avtalsingåendet.
Likaså utgör bokningen ingen garanti för att resenären redan förfogar över en biljett eller liknande färdbevis.
Man kan även tänka sig andra varianter, nämligen: Resenären bokar hos en resebyrå och erhåller vanligtvis ett bokningsbevis.
Resenären binder sig på förhand utan att avtalet omedelbart är perfekt.
En researrangör kan förbehålla sig rätten till ett godkännande vid en senare tidpunkt.
Det är heller inte säkert att det vid denna tidpunkt utfärdats en biljett.
Resenären kan även boka direkt på biljettkontoret och erhåller då biljetten omedelbart.
I detta fall kan man utgå ifrån att avtalet ingåtts omedelbart.
Ändringsförslag
19
Motivering
Förenkling av definitionen.
Ändringsförslag
20
utgår
Motivering
Skillnaden mellan vanlig tågtrafik och höghastighetstrafik är relevant endast när det handlar om att fastställa ersättning (bilaga III).
Föredraganden anser att denna skillnad i ersättning är onödig och förvirrande.
I och med detta blir även denna definition överflödig.
Ändringsförslag
21
15) försening: skillnaden mellan den avgångs- och/eller ankomsttid som anges i tjänstetidtabellen eller den offentliggjorda tidtabellen (även tidtabellshäften som ställs till resenärernas förfogande) för den internationella trafiken eller den internationella höghastighetstrafiken vid avgångs- och/eller ankomststationen och den verkliga avgångs- och/eller ankomsttiden.
15) försening: skillnaden mellan den ankomsttid som anges i tidtabellen och den verkliga ankomsttiden.
Förändringar i tidtabellen som meddelats resenärerna minst 48 timmar i förväg skall inte betecknas som förseningar.
Motivering
Definitionen av förseningar kan förenklas.
Ändringsförslag
22
16) inställd trafik: indragning av planerade internationella tåg eller internationella höghastighetståg .
16) inställd trafik: indragning av planerade tåg , med undantag av avgångar vilkas indragning meddelats resenärerna minst 48 timmar i förväg .
Motivering
Denna bestämmelse bör även gälla nationella tåg.
Ändringsförslag
23
17) följdskador: omfattande skador som uppkommer till följd av en försening, en försening som leder till en missad anslutning eller inställd trafik.
utgår
Motivering
Föredraganden anser att definitionen av och bestämmelserna avseende följdskador är för vaga och för långtgående.
Föredraganden inser att en försening eller en missad anslutning i undantagsfall kan få långtgående följder.
Därför lägger föredraganden till en punkt i artikel 15 i vilken förtydligas att denna förordning inte inverkar på en passagerares rätt att kräva ytterligare kompensation, t.ex. rätt till ersättning enligt nationell lagstiftning.
Ändringsförslag
24
18) tjänstetidtabell: uppgifter om alla planerade tågrörelser och rörelser av rullande materiel som kommer att äga rum på den berörda infrastrukturen under tidtabellens giltighetstid.
utgår
Motivering
Denna definition är överflödig.
Ändringsförslag
25
20) systemleverantör: ett företag och dess filialer som ansvarar för driften eller marknadsföringen av datoriserade informations- och bokningssystem för järnvägstrafik.
Motivering
Järnvägsföretag kan inte utan vidare betraktas som systemleverantörer, eftersom de inte kan förpliktigas att ta in andra företags obegränsade tjänster i sitt bokningssystem.
Om järnvägsföretag betraktas som systemleverantörer innebär detta att de enligt artikel 5.2 är skyldiga att tillhandahålla alla övriga järnvägsföretag tillgång till all reseinformation och alla bokningssystem.
Denna konsekvens kan inte vara önskvärd eftersom den inte ger resenären några rättigheter utan påverkar konkurrensförhållandet mellan olika företag.
Ändringsförslag
26
21) funktionshindrade personer: en person vars rörelseförmåga är nedsatt på grund av fysiskt, sensoriskt, motoriskt eller psykiskt funktionshinder, eller på grund av annat handikapp eller ålder, vid användning av transportmedel och som kräver att särskild hänsyn tas och att utbudet av de tjänster som erbjuds resenärerna anpassas till personens behov.
21) funktionshindrade personer: en person vars oberoende, orienteringsförmåga, kommunikationsförmåga eller rörelseförmåga är nedsatt på grund av fysiskt, sensoriskt, motoriskt eller psykiskt funktionshinder, eller på grund av annat handikapp eller ålder, vid användning av transportmedel och som kräver att särskild hänsyn tas och att utbudet av de tjänster som erbjuds resenärerna anpassas till personens behov.
Motivering
Begreppet funktionshinder bör utvidgas kraftigt.
Ändringsförslag
27
23a) CIV: Enhetliga regler för avtal om internationell järnvägsbefordran av resande, ändrade genom Vilniusprotokollet från 1999, bilaga A i COTIF-fördraget.
Motivering
Föredraganden vill på flera ställen hänvisa till de gällande COTIF-bestämmelserna avseende resenärer.
I samtliga dessa fall hänvisas till ovan nämnda dokument.
Ändringsförslag
28
Järnvägsföretag och/eller researrangörer skall till resenären lämna åtminstone den information som anges i bilaga I.
Järnvägsföretag och/eller researrangörer skall på begäran till resenären lämna den information som anges i bilaga I om de tjänster som företaget erbjuder .
Motivering
Den information som nämns i bilaga I är mycket detaljerad.
Järnvägsföretag kommer inte alltid att ha tillgång till all denna information, när det handlar om tjänster som erbjuds av andra företag (i utlandet).
Ändringsförslag
29
Den information som enligt bilaga I skall lämnas före resan skall även omfatta trafik som erbjuds av andra järnvägsföretag.
utgår
Motivering
Den information som nämns i bilaga I är mycket detaljerad.
Järnvägsföretag kommer inte alltid att ha tillgång till all denna information, när det handlar om tjänster som erbjuds av andra företag (i utlandet).
Ändringsförslag
30
Informationen skall lämnas i den form som är lämpligast .
Informationen skall erbjudas i en form som är tillgänglig och förståelig och den skall vara avgiftsfri.
Särskild hänsyn skall tas till personer med hörsel- och/eller synskada .
Ändringsförslag
31
Järnvägsföretag och researrangörer är ansvariga för att den tryckta eller elektroniskt erbjudna informationen om deras tjänster är korrekt.
Motivering
Felaktig information i foldrar eller på Internet måste undvikas.
Det måste fastställas var ansvaret ligger.
Ändringsförslag
32
1.
Genom transportavtalet åtar sig järnvägsföretaget eller järnvägsföretagen att transportera resenären samt dennes handresgods och resgods till bestämmelseorten.
Avtalet skall bekräftas genom att en eller flera biljetter utfärdas för resenären.
Biljetterna skall betraktas som prima facie-bevis för avtalets ingående .
1.
För transportavtal gäller bestämmelserna i artiklarna 6 och 7 i CIV .
Motivering
Föredraganden vill i förordningen så långt som möjligt ansluta till bestämmelserna i COTIF‑fördraget för att förekomma att järnvägsföretag måste införa olika eller t.o.m. motstridiga bestämmelser.
Ändringsförslag
33
2.
De biljetter som järnvägsföretagen utfärdar skall omfatta åtminstone den information som anges i bilaga II.
2.
Utan att det påverkar tillämpningen av punkt 1 skall de biljetter som järnvägsföretagen utfärdar omfatta åtminstone den information som anges i bilaga II.
Motivering
Se även föregående ändringsförslag.
Bilaga II är ett bra komplement till bestämmelserna i CIV och bör således vara kvar som tilläggsbestämmelser.
Ändringsförslag
34
3.
Om biljetterna utfärdats och bokningarna gjorts i resenärens namn skall de, på de villkor som anges när biljetterna köps, kunna överlåtas till en annan person.
utgår
Motivering
Ändringsförslag
35
4.
Biljetterna och bokningarna kan ha formen av elektronisk dataregistrering, som kan överföras till läsliga skriftsymboler.
utgår
Motivering
Ändringsförslag
36
2.
En systemleverantör som erbjuder distributionstjänster avseende regelbunden persontrafik på järnväg skall ge varje järnvägsföretag som så begär möjlighet att få del av dessa tjänster på lika och icke-diskriminerande villkor inom ramen för det berörda systemets tillgängliga kapacitet med förbehåll för tekniska begränsningar som ligger utanför systemleverantörens kontroll.
2.
En systemleverantör skall ge varje järnvägsföretag som så begär möjlighet att få del av dessa distributionstjänster på lika och icke‑diskriminerande villkor inom ramen för det berörda systemets tillgängliga kapacitet med förbehåll för tekniska begränsningar som ligger utanför systemleverantörens kontroll.
Motivering
Järnvägsföretag kan inte utan vidare ses som systemleverantörer.
Föredraganden vill inte att järnvägsföretag skall vara skyldiga att utan begränsningar även inlemma andra företags tjänster i sina reservationssystem.
Ändringsförslag
37
1.
Järnvägsföretag och/eller researrangörer skall erbjuda biljetter och/eller samordnade biljetter för internationella resor åtminstone mellan större järnvägsstationer, och till järnvägsstationer som är belägna i ett område med närmaste järnvägsstation som knutpunkt.
utgår
Motivering
I praktiken erbjuder redan många järnvägsföretag biljetter som gäller inom en zon.
Med tanke på de skiftande förhållandena inom det europeiska järnvägsnätet är det svårt att lagstiftningsvägen framtvinga dylika möjligheter.
Det är faktiskt svårt att fastställa var zongränsen går i varje enskilt fall.
Föredraganden utgår från att järnvägsföretagen kommer att tillämpa eller införa zonbiljetter där så är möjligt.
Ändringsförslag
38
3.
Biljetter för internationella resor skall distribueras till resenärer åtminstone via följande försäljningsställen:
3.
Biljetter skall distribueras till resenärer åtminstone via följande försäljningsställen:
a) biljettkontor och biljettautomater (om sådana finns) på samtliga större järnvägsstationer, eller
a) biljettkontor och tillgängliga biljettautomater (om sådana finns) på samtliga större järnvägsstationer, eller
b) telefon/ Internet eller annan allmänt tillgänglig informationsteknik utan extra avgifter för användning av denna distributionskanal.
b) telefon/ tillgängliga webbplatser eller annan allmänt tillgänglig informationsteknik utan extra avgifter för användning av denna distributionskanal.
Ändringsförslag
39
3a.
Biljetter som utfärdas inom ramen för avtal om offentliga tjänster skall åtminstone distribueras via följande försäljningsställen:
a) biljettkontor och tillgängliga biljettautomater (om sådana finns) på samtliga större järnvägsstationer, och
b) telefon/tillgängliga webbplatser eller annan allmänt tillgänglig informationsteknik utan extra avgifter för användning av denna distributionskanal.
Ändringsförslag
40
3b.
Om det inte finns något biljettkontor eller någon biljettautomat på avgångsstationen skall passagerarna på järnvägsstationen åtminstone informeras om:
– möjligheten att köpa biljett per telefon, via Internet eller på tåget samt de förfaranden som skall följas,
– den närmaste stora järnvägsstationen eller platsen där det finns tillgängliga biljettkontor och/eller biljettautomater.
Ändringsförslag
41
4.
Järnvägsföretag skall emellertid, på de villkor som anges i artikel 36, ge resenärerna möjlighet att köpa biljetter för internationella resor ombord på tåget.
4.
Om inte tillträdet till tåget eller stationsbyggnaden av säkerhetsskäl är begränsat skall järnvägsföretag ge resenärerna möjlighet att köpa biljetter ombord på tåget , i synnerhet om resenärerna inte kunnat köpa sina biljetter på avgångsstationen av något av följande skäl:
– biljettkontoren var stängda,
– biljettautomaterna var i olag,
– det fanns varken biljettkontor eller biljettautomater på avgångsstationen,
– biljettkontoren eller biljettautomaterna var inte tillgängliga för funktionshindrade resenärer.
Resenären skall omedelbart informera behörig tågpersonal.
Ändringsförslag
42
Artikel 6a (ny)
Artikel 6a
2.
3.
Ett år efter det att denna förordning antagits skall kommissionen, på förslag av Europeiska järnvägsbyrån, anta de tekniska specifikationerna för driftskompatibilitet för telematikapplikationer avsedda för persontrafik.
Med TSD skall det bli möjligt att tillhandahålla den information som avses i bilaga II.
4.
Motivering
I dagsläget är det omöjligt att kräva att järnvägsföretag skall erbjuda biljetter för hela sträckan när det gäller internationella resor genom hela Europa.
Genom att utveckla TSD kan vi hjälpa järnvägsföretagen att samarbeta.
Föredraganden hoppas att man sålunda, på samma sätt som inom flyget, skall kunna ta ett antal initiativ för att göra det möjligt att sälja heltäckande biljetter för hela Europa.
Föredraganden är övertygad om att denna utveckling kommer att gå hand i hand med den fortgående konkurrensutsättningen av den europeiska marknaden.
Ändringsförslag
43
Kapitel III, rubrik
JÄRNVÄGSFÖRETAGETS ANSVARIGHET
ANSVARIGHET OCH SKADESTÅND VID RESENÄRERS DÖDSFALL ELLER SKADA
Motivering
Föredraganden vill föra samman alla bestämmelser som rör passagerares död eller skador under en enda rubrik.
Ändringsförslag
44
1.
Järnvägsföretaget skall vara ansvarigt om en resenär dödas eller skadas (fysiskt eller psykiskt), men endast om olyckan som ledde till dödsfallet eller skadan inträffade när resenären befann sig på tåget eller i samband med på- eller avstigning .
1.
Järnvägsföretaget skall vara ansvarigt om en resenär dödas eller skadas (fysiskt eller psykiskt), om olyckan som ledde till dödsfallet eller skadan inte var följden av en naturkatastrof, en krigshandling eller av terrorism .
Motivering
Ingen begränsning av ansvaret enligt platsen där passageraren befann sig, utan i stället en begränsning av ansvaret kopplat till orsak.
Man kan inte förvänta sig att järnvägsföretag skall ta ansvar för en terroristattack, som den i Madrid.
Ändringsförslag
45
Motivering
Med tanke på den allt sämre integrering mellan järnvägsföretag som blivit resultatet av alla EU-direktiv och de allt flera aktörerna inom järnvägssektorn (järnvägsföretag, infrastrukturförvaltare, självständiga företag som ansvarar för underhåll, …) är det lämpligt att, som skydd för resenärerna, vid en olycka låta dem ha juridisk kontakt med endast en part: järnvägsföretaget som har ombesörjt resan.
Det är järnvägsföretagets sak att sedan vända sig till tredje part för att utkräva deras ansvar.
Ändringsförslag
46
Artikel 7a (ny)
Artikel 7a
Skadestånd vid resenärers dödsfall eller skada
1.
Inget begränsningsbelopp gäller för järnvägsföretagets ansvarighet vid resenärers dödsfall eller kroppsskada.
2.
Vid högre belopp skall järnvägsföretaget inte vara ansvarigt för skadan om det kan bevisa att det inte handlat försumligt eller begått något fel.
3.
Om personer för vilka resenären hade eller skulle ha haft en lagstadgad underhållsskyldighet, på grund av resenärens död berövas detta stöd, skall de ha rätt till ersättning för denna förlust.
Motivering
För att göra förordningen mera lättläst föreslår föredraganden att alla bestämmelser som rör passagerares död eller skador förs samman.
Artiklarna 12 och 13 flyttas alltså till artikel 7.
Ändringsförslag
47
Artikel 7b (ny)
Artikel 7b
Vid dödsfall uppgår detta förskott till minimum 19 000 EUR.
Detta förskott utgör inget erkännande av ersättningsansvar och dras ifrån ett eventuellt senare ersättningsbelopp som utbetalas på grund av järnvägsföretagets ersättningsansvar.
Motivering
För att förordningen skall bli mer lättbegriplig föreslås att alla bestämmelser som rör resenärers dödsfall eller skador sammanfattas.
Av denna anledning införlivas artikel 13 i artikel 7.
Vidare görs anpassningar till luftfartsbestämmelserna.
Ändringsförslag
48
Kapitel IIIa (nytt)
Kapitel IIIa
ANSVARIGHET OCH SKADESTÅND VID SKADAT ELLER FÖRKOMMET RESGODS, HANDRESGODS, DJUR OCH FORDON
Motivering
För att göra förordningen mera lättläst föreslår föredraganden att alla bestämmelser som rör skador eller förluster förs samman.
Ändringsförslag
49
Artikel 8, rubrik
Handresgods
utgår
Motivering
Föredraganden föreslår att bestämmelser rörande alla resgodstyper samlas i en enda artikel (se följande ändringsförslag).
Ändringsförslag
50
1.
Om en resenär dödas eller skadas skall järnvägsföretaget vara ansvarigt för total eller partiell förlust av eller skada på personliga tillhörigheter som resenären hade med sig som handresgods .
1.
När det gäller ansvarighet och ersättning i händelse av att handresgods, husdjur, resgods, rullstol, barnvagn, cykel eller fordon helt eller delvis förstörs, förloras eller skadas skall de bestämmelser gälla som anges i kapitel III i CIV, särskilt artiklarna 33–46 .
Motivering
Den ansvarighet som anges i CIV i händelse av skada på eller förlust av resgods är betydligt mer omfattande än vad som föreslås i föreliggande förslag till förordning.
Man bör särskilt se till att ansvarigheten omfattar resgods som gör det lättare att byta transportsätt, såsom rullstolar, barnvagnar, cyklar o.s.v.
2.
I andra fall skall järnvägsföretaget inte ha något ansvar för förlust av eller skada på personliga tillhörigheter och handresgods för vilket resenären själv har tillsynsansvaret, såvida inte järnvägsföretaget begått något fel som orsakat förlusten eller skadan .
2.
Utan att det påverkar tillämpningen av punkt 1 skall järnvägsföretaget eller den stationsförvaltare som är skadeståndsansvarig vid total eller fullständig förstörelse av, förlust av eller skada på funktionshindrade resenärers rörelsehjälpmedel/medicinska hjälpmedel betala ett skadestånd som högst motsvarar ersättningskostnaden för utrustningen.
I förekommande fall skall järnvägsföretaget även erbjuda den berörda resenären ett hjälpmedel som tillfällig ersättning .
Motivering
Skadeståndet för förlust av handresgods och djur är högst 1 400 räkneenheter (ca 1 650 euro).
Föredraganden föreslår att denna gräns höjs när det gäller förlust av eller skada på rörelsehjälpmedel för funktionshindrade.
Med tanke på att funktionshindrade är beroende av sin utrustning måste det ansvariga järnvägsföretaget eller den ansvarige stationsförvaltaren också se till att det erbjuds ett tillfälligt ersättningshjälpmedel.
Ändringsförslag
52
Artikel 9
Artikel 9
utgår
Annat resgods
Järnvägsföretaget skall vara ansvarigt för den skada som lidits om en del av eller hela resgodset förstörs, förloras eller skadas, under förutsättning att den händelse som ledde till att resgodset förstördes, försvann eller skadades inträffade när järnvägsföretaget hade ansvaret för resgodset.
Motivering
Se motivering till ändringsförslaget avseende artikel 8.
Ändringsförslag
53
Artikel 10
Artikel 10
utgår
Försening
Järnvägsföretaget är ansvarigt för förseningar, inbegripet förseningar som leder till en missad anslutning, och/eller för inställd internationell trafik som drabbar resenärer och/eller transport av resgods.
Järnvägsföretaget skall inte vara ansvarigt för försenad eller inställd internationell trafik som är en följd av extrema väderförhållanden, naturkatastrofer, krigshandlingar eller terrorism.
Motivering
Föredraganden föreslår att alla bestämmelser rörande förseningar samlas i kapitel IV.
Ändringsförslag
54
Artikel 11
Artikel 11
utgår
Följdskador
Om järnvägsföretaget är ansvarigt för en försening, en försening som leder till missad anslutning eller inställd trafik, skall järnvägsföretaget vara skadeståndsansvarigt, oberoende av de villkor för ersättning vid förseningar som anges i artikel 10.
Vid förseningar på mindre än en timme skall det inte utgå någon ersättning för följdskador; detta skall dock inte påverka tillämpningen av artikel 16.
Motivering
Föredraganden anser att bestämmelserna avseende följdskador är för vaga och för långtgående.
Föredraganden inser att en försening eller en missad anslutning i undantagsfall kan få långtgående följder.
Därför lägger föredraganden till en punkt i artikel 15 i vilken förtydligas att denna förordning inte inverkar på en passagerares rätt att kräva ytterligare kompensation, t.ex. rätt till ersättning enligt nationell lagstiftning.
Ändringsförslag
55
Kapitel IV, rubrik
SKADESTÅND OCH ERSÄTTNING
ANSVARIGHET, SKADESTÅND OCH ASSISTANS VID FÖRSENINGAR
Motivering
I likhet med bestämmelserna om dödsfall eller skada och förlust av eller skada på resgods vill föredraganden även här samla alla bestämmelser rörande förseningar i ett enda kapitel.
Ändringsförslag
56
Artikel 11a (ny)
Artikel 11a
Försening
1.
Järnvägsföretaget är ansvarigt för förseningar som leder till en missad anslutning, och/eller för inställd trafik som drabbar resenärer och/eller transport av resgods.
2.
Järnvägsföretaget skall inte vara ansvarigt för förseningar, missade anslutningar eller inställd trafik om detta beror på
– extrema väderförhållanden eller naturkatastrofer, krigshandlingar eller terrorism,
– omständigheter utanför järnvägsföretagets verksamhet som företaget inte kunnat undvika, och vilkas följder man inte kunnat förhindra trots att man visat den omsorg som situationen kräver,
– resenärens vållande, eller
3.
Järnvägsföretaget och/eller stationsförvaltaren skall också vara ansvarig(a) för försenad assistans vid järnvägsstationen eller ombord på tåget som leder till att en resenär med funktionshinder missar sitt tåg vid avfärd eller sin anslutning vid ankomst.
Ändringsförslag
57
Artikel 12
Artikel 12
utgår
Skadestånd vid resenärers dödsfall eller kroppsskada
1.
Inget begränsningsbelopp gäller för järnvägsföretagets ansvarighet vid resenärers dödsfall eller kroppsskada.
2.
Vid högre belopp skall järnvägsföretaget inte vara ansvarigt för skadan om det kan bevisa att det inte handlat försumligt eller begått något fel.
3.
Om personer för vilka resenären hade eller skulle ha haft en lagstadgad underhållsskyldighet, på grund av resenärens död berövas detta stöd, skall de ha rätt till ersättning för denna förlust.
Motivering
Föredraganden föreslår att denna artikel flyttas till kapitel III och där infogas som artikel 7a (ny).
Ändringsförslag
58
Artikel 13
Artikel 13
utgår
Förskottsutbetalningar
Om en resenär dödas eller skadas skall järnvägsföretaget göra en förskottsutbetalning för att täcka omedelbara ekonomiska behov, inom 15 dagar från det att det fastställts vem som har rätt till skadestånd.
Vid dödsfall skall denna förskottsutbetalning uppgå till minst 21 000 euro.
Motivering
Se föregående ändringsförslag.
Artikel 14
Artikel 14
utgår
Ersättning för handresgods och annat resgods
1.
När järnvägsföretaget är ansvarigt enligt artikel 8 skall det betala en ersättning på högst 1 800 euro per resenärer.
2.
När järnvägsföretaget är ansvarigt enligt artikel 9 skall det betala en ersättning på högst 1 300 euro per resenärer.
Motivering
Se föregående ändringsförslag.
Ändringsförslag
60
-1.
Järnvägsföretaget skall betala tillbaka till resenären tillägg och påslag om de tillhandahållna tjänsterna inte motsvarar de angivna kriterierna för tillägg och påslag (se bilaga II, punkt 4a).
Motivering
Det ersättningssystem som föreslagits av kommissionen bör ersättas av ett mer praktiskt system som grundar sig på reella prisstrukturer (se ändringsförslaget till bilaga II från Michael Cramer).
Ändringsförslag
61
1.
Resenärer som drabbas av förseningar får, utan att därmed avsäga sig rätten till transport, begära ersättning för dessa förseningar från järnvägsföretaget.
Minimiersättningen vid förseningar anges i bilaga III .
1.
Resenärer som drabbas av förseningar får, utan att därmed avsäga sig rätten till transport, begära ersättning för dessa förseningar från järnvägsföretaget.
Minimiersättningen vid förseningar skall uppgå till:
– 25 procent vid en försening på minst 60 minuter,
– 50 % vid en försening på minst 120 minuter,
– 75 % vid en försening på minst 180 minuter.
Ändringsförslag
62
1a.
Resenärer som har ett abonnemang och som under dess giltighetstid upprepade gånger drabbats av förseningar eller inställd trafik skall på begäran få ersättning.
Denna ersättning kan utbetalas på olika sätt: gratis resor, prisreduktioner eller en förlängning av abonnemangets giltighetstid.
Järnvägsföretagen skall på förhand fastställa, och i nära samarbete med användarnas företrädare och med ansvariga myndighet i samband med avtal om offentliga tjänster, de kriterier som ska gälla i samband med tillämpningen av denna punkt när det gäller att fastställa den berörda tjänstens punktlighet och tillförlitlighet.7
Ändringsförslag
63
2.
Ersättningen får inte erläggas i form av kuponger och/eller andra tjänster, såvida resenären inte ger sitt skriftliga medgivande .
2.
Den ersättning som avses i punkt 1 skall betalas inom en månad efter det att en begäran om ersättning framställts.
Ersättningen får erläggas i form av kuponger och/eller andra tjänster, under förutsättning att villkoren är flexibla (särskilt avseende giltighetstid och destination).
Ersättningen måste utbetalas i reda pengar om resenären begär det .
Ändringsförslag
64
3a.
Tillämpningen av denna artikel påverkar inte en passagerares rätt till ytterligare kompensation.
Kompensation som beviljas i enlighet med denna förordning får räknas av från sådan kompensation.
Motivering
Denna bestämmelse har tagits från den nyligen antagna förordningen för lufttrafik och är enligt föredraganden betydligt mer realistisk än den här förordningens bestämmelser om följdskada.
Ändringsförslag
65
-1.
Järnvägsföretagens första prioritet är att se till att hålla anslutningar och att med alla till buds stående medel undvika att trafik inställs.
Motivering
Järnvägstjänsten i sig, d.v.s. det att hålla anslutningar och undvika att trafik inställs, bör stå i första ledet bland resenärers rättigheter (”befordringsplikten”).
Ändringsförslag
66
1.
Vid förseningar som leder till missade anslutningar eller vid inställd internationell trafik skall punkt 2 tillämpas, såvida järnvägsföretaget inte kan bevisa att trafiken ställdes in enbart på grund av extrema omständigheter.
1.
Vid förseningar , inbegripet förseningar i järnvägsföretagets tillhandahållande av assistans till personer med funktionshinder, som leder till missade anslutningar eller vid inställd trafik skall punkt 2 tillämpas, såvida järnvägsföretaget inte kan bevisa att trafiken försenades eller ställdes in enbart på grund av extrema omständigheter.
Ändringsförslag
67
2.
2.
När ett järnvägsföretag drabbas av en försening som kommer att leda till en missad anslutning eller om järnvägsföretaget, före den tidtabellsenliga avgångstiden, ställer in eller har rimlig anledning att förvänta sig att det kommer att ställa in trafik, skall det vidta erforderliga åtgärder för att informera resenärerna och se till att dessa kan nå den slutliga bestämmelseorten .
Motivering
Oberoende av förseningens orsaker måste järnvägsföretagen göra allt för att informera resenärerna och se till så att de kan komma fram till den slutliga bestämmelseorten.
Om resan kan genomföras längs en annan järnvägssträckning med tåg från ett annat järnvägsföretag får detta inte räknas som ett hinder.
Ändringsförslag
68
Denna ersättning skall betalas ut på samma villkor som den ersättning som avses i artikel 15.2 eller 15.3.
a) Ersättning motsvarande hela biljettpriset, enligt samma villkor som vid köpet, för den eller de delar av resan som inte fullföljts och för den eller de delar som fullföljts, om resan inte längre har något syfte med tanke på resenärens ursprungliga resplan, med en returresa till den första avgångsorten snarast möjligt om detta är relevant.
Denna ersättning skall betalas ut på samma villkor som den ersättning som avses i artikel 15.2 eller 15.3.
Motivering
Denna bestämmelse bör gälla också för nationell tågtrafik.
Ändringsförslag
69
b) Fortsatt resa eller ombokning till den slutliga bestämmelseorten på likvärdiga transportvillkor snarast möjligt.
b) Fortsatt resa eller ombokning till den slutliga bestämmelseorten på likvärdiga transportvillkor och med samma grad av tillgänglighet snarast möjligt , eventuellt med dyrare tåg utan extra kostnader .
Motivering
”Likvärdiga transportvillkor” måste tolkas på ett sådant sätt att man säkrar samma grad av tillgänglighet.
Om exempelvis en förbindelse som är tillgänglig för rullstol ställs in och nästa tåg (det ”snarast möjliga”) inte är tillgänglig för rullstol skall en resande med funktionshinder inte vara skyldig att acceptera denna otillgängliga förbindelse som alternativ resa.
Ändringsförslag
70
c) Fortsatt resa eller ombokning till den slutliga bestämmelseorten på likvärdiga transportvillkor en senare dag som resenären finner lämplig .
c) Fortsatt resa eller ombokning till den slutliga bestämmelseorten på likvärdiga transportvillkor en senare dag.
Motivering
Force majeur-klausulen bör övervägas i samband med rätten att välja huruvida man önskar fortsätta resan eller avbryta den och erhålla ersättning i samband med försening som leder till att en anslutning missas eller i samband med att ett tåg ställs in eller att ett tåg förväntas ställas in.
För oavsett av vilken anledning kan det vara möjligt att det för resenären inte längre lönar sig att påbörja resan vid en senare tidpunkt, t.ex. om denne haft ett avtalat möte som han/hon under alla omständigheter inte längre kan hinna till.
Vidare kan det inte råda någon tvekan om att biljettpriset skall återbetalas ifall järnvägsföretaget å sin sida inte kan tillhandahålla sina tjänster.
Risken för händelser beroende på force majeur ankommer alltid i sådana fall på företaget (detta gäller även andra branscher).
Järnvägsföretag bör i dylika fall inte heller kunna åberopa force majeur i samband med dessa rättigheter som gäller resenärerna.
Ändringsförslag
71
a) måltider och förfriskningar i skälig proportion till väntetiden , och/eller
a) måltider och förfriskningar i möjlig mån , och/eller
Motivering
Ändringsförslagen till punkterna a och b i denna artikel är i enlighet med de europeiska järnvägsföretagens åtagande, enligt sin egen stadga, att under angivna omständigheter tillhandahålla sådan assistans som krävs för att möta resenärers rimliga behov.
Det bör noteras att järnvägsföretagen erkänner sin förpliktelse att säkra sina kunders säkerhet och komfort (d.v.s. genom punkterna a, b och c om problem uppstår, även om det enskilda järnvägsföretaget inte är ersättningsskyldigt i enlighet med artikel 11a.2).
Dock är formuleringen ”i möjlig mån” nödvändig eftersom situationer kan uppstå då järnvägsföretaget inte har möjlighet att uppfylla detta åtagande.
Exempelvis saknar många tåg cateringfaciliteter, och det är sällan möjligt att leverera varor till ett tåg som inte står vid station, och särskilt inte om uppehållet orsakas av dåligt väder.
Ändringsförslag
72
b) hotellrum i sådana fall då övernattning under en eller flera nätter eller ytterligare vistelse blir nödvändig, och/eller
b) inkvartering, om detta inte är omöjligt under rådande omständigheter, i sådana fall då övernattning under en eller flera nätter eller ytterligare vistelse blir nödvändig, och/eller
Motivering
Ändringsförslagen till punkterna a och b i denna artikel är i enlighet med de europeiska järnvägsföretagens åtagande, enligt sin egen stadga, att under angivna omständigheter tillhandahålla sådan assistans som krävs för att möta resenärers rimliga behov.
Det bör noteras att järnvägsföretagen erkänner sin förpliktelse att säkra sina kunders säkerhet och komfort (d.v.s. genom punkterna a, b och c om problem uppstår, även om det enskilda järnvägsföretaget inte är ersättningsskyldigt i enlighet med artikel 11a.2).
Dock är formuleringen ”om detta inte är omöjligt under rådande omständigheter” nödvändig, eftersom situationer kan uppstå då järnvägsföretaget inte har möjlighet att uppfylla detta åtagande.
Exempelvis saknar många tåg cateringfaciliteter, och det är sällan möjligt att leverera varor till ett tåg som inte står vid station, och särskilt inte om uppehållet orsakas av dåligt väder.
Ändringsförslag
73
c) transport mellan järnvägsstationen och inkvarteringsstället (hotell eller annat),
c) transport mellan järnvägsstationen och inkvarteringsstället (hotell eller annat), eller
Ändringsförslag
74
Motivering
Denna ändring av punkt d är nödvändig för att fastställa en uppsättning praktiskt tillämpbara alternativ för järnvägssektorn.
Särskilda bestämmelser om avstigning utanför stationsområdet har konsekvenser som även måste beaktas ur ett säkerhetsperspektiv och bör därför inte regleras i lagstiftning om resenärers rättigheter.
I situationer där förseningen el. dyl. skylls omständigheter som ligger utanför järnvägsföretagets kontroll vore det orimligt att de skall ha skyldighet att tillhandahålla alternativ transport.
Ändringsförslag
75
3.
3.
Järnvägsföretag skall på resenärens begäran intyga på biljetten att tågtrafiken varit försenad, att förseningen lett till en missad anslutning eller att trafiken ställts in.
Om järnvägsföretag kräver sådana intyg måste de vidta lämpliga åtgärder så att resenärerna snabbt och enkelt kan få dem.
Motivering
Det är inte klart hur ett sådant här intygande skall ske, eller vilka rutiner som skall tillämpas.
Skall varje tåganställd kunna ge intyg?
Om så inte är fallet, skall resenärerna då vara tvungna att välja mellan att antingen t.ex. ta ett senare tåg eller leta reda på en viss tjänsteman som kan ge detta intyg?
Järnvägsföretag som kräver sådana intyg måste åläggas att införa snabba och enkla intygsrutiner.
Ändringsförslag
76
Upplysningar om förseningar eller inställd trafik, hotellrum eller alternativa transportmedel, ersättningsvillkor samt möjlighet till fortsatt eller ombokad resa måste meddelas på ett tillgängligt sätt.
Järnvägsföretaget skall se till att inkvartering och alternativa transportmedel är tillgängliga för funktionshindrade resenärer och att dessa erbjuds lämplig assistans i händelse av förseningar eller inställd trafik.
Motivering
Syftet med ändringsförslaget är att förtydliga texten.
Resenärer med funktionshinder har särskilda behov som måste tillgodoses i händelse av försening.
Ändringsförslag
77
1.
Bestämmelserna om ansvarighet skall även gälla när järnvägsfordon transporteras med färja på del(ar) av den internationella resan , såvida inte de regler som gäller för sjötransporten är mer förmånliga för resenären .
1.
När järnvägsfordon transporteras med färja på del(ar) av resan eller när järnvägstrafiken tillfälligt ersätts av ett annat transportmedel gäller bestämmelserna i artikel 31 i CIV .
Motivering
Föredraganden vill så långt som möjligt ansluta till bestämmelserna i COTIF-fördraget för att förekomma att järnvägsföretag måste införa olika eller t.o.m. motstridiga bestämmelser.
Ändringsförslag
78
2.
utgår
Motivering
Detta täcks av det föregående ändringsförslaget.
Ändringsförslag
79
Artikel 19
Om den internationella transporten utförs av flera på varandra följande järnvägsföretag skall de berörda järnvägsföretagen vara solidariskt ansvariga om en resenär dödas eller skadas, om resgods förstörs eller förloras, eller i händelse av förseningar, förseningar som leder till missade anslutningar eller inställd trafik.
Om transporten utförs av flera på varandra följande järnvägsföretag skall de berörda järnvägsföretagen vara solidariskt ansvariga om en resenär dödas eller skadas, om resgods förstörs eller förloras, eller i händelse av förseningar, förseningar som leder till missade anslutningar eller inställd trafik.
Motivering
Denna bestämmelse bör gälla också för nationell tågtrafik.
Ändringsförslag
80
Artikel 20
Om ett järnvägsföretag har anförtrott åt ett annat järnvägsföretag att helt eller delvis utföra transporten, skall de ordinarie järnvägsföretaget trots det förbli ansvarigt för hela transporten.
Om ett järnvägsföretag har anförtrott åt ett annat järnvägsföretag att helt eller delvis utföra transporten, skall de ordinarie järnvägsföretaget trots det förbli ansvarigt för hela transporten enligt bestämmelserna i artikel 39 i CIV .
Motivering
Artikel 39 i CIV innehåller ett antal nyttiga kompletterande bestämmelser beträffande ställföreträdande järnvägsföretag.
Ändringsförslag
81
Järnvägsföretaget skall vara ansvarigt för sin personal och andra personer vars tjänster det utnyttjar för utförandet av transporten, när dessa agerar inom ramen för sina funktioner .
Järnvägsföretaget skall vara ansvarigt för de personer som nämns i artikel 51 i CIV .
Motivering
Artikel 21 är helt och hållet i överensstämmelse med artikel 51 i CIV.
Det räcker därför att hänvisa till detta fördrag.
Ändringsförslag
82
Infrastrukturförvaltarens personal skall betraktas som personer vars tjänster järnvägsföretaget utnyttjar för utförandet av transporten.
utgår
Motivering
Artikel 21 är helt och hållet i överensstämmelse med artikel 51 i CIV.
Det räcker därför att hänvisa till detta fördrag.
Ändringsförslag
83
Artikel 23
1.
När det gäller preskriptionstider för skadeståndstalan skall bestämmelserna i artikel 60 i CIV tillämpas .
a) För resenärer: tre år från olycksdagen.
b) För andra skadelidande personer: tre år från resenärens bortgång, dock högst fem år från olycksdagen.
2.
Motivering
Föredraganden vill så långt som möjligt ansluta till bestämmelserna i COTIF-fördraget för att förekomma att järnvägsföretag måste införa olika eller t.o.m. motstridiga bestämmelser.
Ändringsförslag
84
Järnvägsföretaget skall ha rätt att kräva ersättning från infrastrukturförvaltaren för att täcka den ersättning som järnvägsföretaget betalat ut till resenärerna.
Infrastrukturförvaltarens ansvarighet skall inte påverka tillämpningen av den verksamhetsstyrning genom kvalitetskrav på utförande som fastställs i artikel 11 i Europaparlamentets och rådets direktiv 2001/14/EG.
Järnvägsföretaget skall ha rätt att kräva ersättning från infrastrukturförvaltaren för att täcka den ersättning som järnvägsföretaget betalat ut till resenärerna.
Infrastrukturförvaltarens ansvarighet skall inte påverka tillämpningen av den verksamhetsstyrning genom kvalitetskrav på utförande som fastställs i artikel 11 i Europaparlamentets och rådets direktiv 2001/14/EG , och skall stå i proportion till priset för järnvägssträckan om det inte finns något kompensationssystem fastställt i verksamhetsstyrningen .
Motivering
De ersättningar för förseningar som ingår i denna förordning uttrycks som procent av biljettpriset.
Detta pris är inte alltid proportionellt mot den ersättning som infrastrukturförvaltaren får för utnyttjandet av järnvägen.
Vid ersättningskrav riktade mot infrastrukturförvaltaren är det önskvärt att även ta hänsyn till de inkomster som denne har haft för järnvägssträckan.
Ändringsförslag
85
Artikel 27
Ett järnvägsföretag och/eller en researrangör får inte på grund av en resenärs rörelsehinder vägra att utfärda en biljett för eller boka en internationell resa från en större järnvägsstation.
Ett järnvägsföretag och/eller en researrangör får inte på grund av en resenärs rörelsehinder vägra att utfärda en biljett för eller boka en resa från en större järnvägsstation.
Ändringsförslag
86
Artikel 27a (ny)
Artikel 27a
Särskilda faciliteter på tåg
Ifall funktionshindrade personer behöver särskilda faciliteter på tåg, vilka inte kan ställas till förfogande utan mycket stora extra insatser gäller järnvägsföretagets transportskyldighet endast inom ramen för den disponibla kapaciteten.
Järnvägsföretagen uppmanas att öka sin disponibla kapacitet i förhållande till behoven.
Motivering
Järnvägsföretagen kan endast tillhandahålla transporttjänster för funktionshindrade personer i den mån detta är möjligt med hänsyn till de på tåget för sådana personer befintliga faciliteterna.
Ifall enbart begränsade speciella faciliteter finns tillgängliga på tåget och dessa redan är reserverade kan en funktionshindrad person inte tillhandahållas erforderlig transport om dessa faciliteter endast kan tillhandahållas genom mycket stora insatser.
Järnvägsföretagen bör dock bygga ut sådana faciliteter.
Ändringsförslag
87
Artikel 27b (ny)
Artikel 27b
Förbud mot prisdiskriminering
Järnvägsföretag och/eller researrangörer skall se till att resenärer med funktionshinder kan köpa biljetter till samma pris som resenärer utan funktionshinder.
Motivering
Resenärer med funktionshinder bör inte behöva betala mer än resenärer utan funktionshinder.
Ändringsförslag
88
Artikel 27c (ny)
Stationsförvaltarna skall se till att stationer, perronger och samtliga tjänster är tillgängliga för funktionshindrade personer genom att avlägsna alla arkitektoniska hinder.
Motivering
Detta är en förutsättning för att funktionshindrade personers rätt till rörlighet skall kunna garanteras.
En förordning som i bredaste mening skall skydda resenärers rättigheter kan inte bortse från behovet att avlägsna alla hinder som begränsar tillgängligheten till stationer.
Ändringsförslag
89
Artikel 27d (ny)
Järnvägsföretag skall säkra tillgängligheten till transportmedel genom att avlägsna allt som hindrar funktionshindrade personers på- och avstigning samt deras möjlighet att vistas ombord på tåget.
Motivering
Järnvägsföretagen skall i samråd med stationsförvaltare se till att tågen helt och fullt uppfyller funktionshindrade personers behov.
System skall införas som möjliggör obehindrad på- och avstigning och som ger funktionshindrade personer möjlighet att förflytta sig i tåget under färd.
Ändringsförslag
90
1.
Stationsförvaltaren på avgångsstationen, på den station där tågbyte sker eller på ankomststationen skall ge funktionshindrade personer som befinner sig på en internationell resa assistans så att de kan stiga på avgående tåg, byta till anslutande tåg eller stiga av ett ankommande tåg för vilket det köpt biljett.
1.
Stationsförvaltaren på avgångsstationen, på den station där tågbyte sker eller på ankomststationen skall ge funktionshindrade personer som befinner sig på resa assistans så att de kan stiga på avgående tåg, byta till anslutande tåg eller stiga av ett ankommande tåg för vilket det köpt biljett.
Motivering
Denna bestämmelse bör gälla också för nationell tågtrafik.
Ändringsförslag
91
2.
Den assistans som avses i punkt 1 skall lämnas under förutsättning att järnvägsföretaget och/eller researrangören minst 24 timmar innan assistans erfordras underrättats om den funktionshindrade personens behov av sådan assistans.
2.
Den assistans som avses i punkt 1 skall lämnas under förutsättning att järnvägsföretaget och/eller researrangören minst 48 timmar innan assistans erfordras underrättats om den funktionshindrade personens behov av sådan assistans.
Motivering
Förordningen tillämpningsområde skall utvidgas till att omfatta även nationella resor.
Eftersom reglerna gällande assistans i artikel 28.1 förutsätter ett mycket omfattande assistanssystem även på nationella resor bör tidsfristen för förberedelse av sådan assistans förlängas till 48 timmar.
Ändringsförslag
92
3.
3.
Motivering
Texten kan förkortas på detta sätt.
Ändringsförslag
93
Artikel 29
Artikel 29
utgår
Assistans på järnvägsstationer
1.
Stationsförvaltaren skall ansvara för assistansen till funktionshindrade personer.
2.
Stationsförvaltaren skall fastställa särskilda platser inne i och utanför järnvägsstationen där funktionshindrade personer kan meddela sin ankomst till järnvägsstationen och vid behov begära assistans.
Motivering
Föredraganden anser att assistans på järnvägsstationer garanteras tillräckligt väl genom bestämmelserna i artikel 28.
Ändringsförslag
94
Artikel 30
Järnvägsföretaget , stationsförvaltaren och/eller researrangören skall ge funktionshindrade personer assistans ombord på tåget och vid på- och avstigning, i enlighet med vad som anges i artikel 28.2.
Assistans ombord på tåget förutsätter att tåget är planenligt bemannat.
Järnvägsbolagen uppmanas att anpassa sin personalplanering efter behoven.
Motivering
Förvaltaren av den station där tjänsten tillhandahålls bör också ansvara för att funktionshindrade personer ges assistans.
Ändringsförslag
95
1.
Järnvägsföretag och researrangörer skall vidta alla erforderliga åtgärder för att vid samtliga försäljningsställen kunna ta emot underrättelser om funktionshindrade personers behov av assistans.
1.
Järnvägsföretag och researrangörer skall se till att det finns ett system som resenärer med funktionshinder kan utnyttja för att meddela järnvägsföretaget sina behov av assistans samt informera om detta system när biljetten köps .
Motivering
Föredraganden föreslår att ersätta denna detaljerade artikel med ett enklare krav på resultat.
Det är bättre att låta järnvägsföretagen och researrangörerna själva avgöra hur de vill organisera meddelanden om behov av assistans.
De måste hur som helst ordna detta på ett väl fungerande sätt, annars uppfyller de inte kraven på assistans i artikel 28.
Ändringsförslag
96
2.
utgår
Motivering
Föredraganden föreslår att ersätta denna detaljerade artikel med ett enklare krav på resultat.
Det är bättre att låta järnvägsföretagen och researrangörerna själva avgöra hur de vill organisera meddelanden om behov av assistans.
De måste hur som helst ordna detta på ett väl fungerande sätt, annars uppfyller de inte kraven på assistans i artikel 28.
Ändringsförslag
97
3.
Omedelbart efter ett nationellt eller internationellt tågs avgång skall järnvägsföretaget underrätta stationsförvaltaren vid den järnvägsstation där tågbyte sker och ankomststationen om antalet funktionshindrade personer som behöver assistans och om vilken typ av assistans som erfordras.
utgår
Motivering
Föredraganden föreslår att ersätta denna detaljerade artikel med ett enklare krav på resultat.
Det är bättre att låta järnvägsföretagen och researrangörerna själva avgöra hur de vill organisera meddelanden om behov av assistans.
De måste hur som helst ordna detta på ett väl fungerande sätt, annars uppfyller de inte kraven på assistans i artikel 28.
Ändringsförslag
98
Kapitel VII, rubrik
SÄKERHET OCH TJÄNSTEKVALITET
RESENÄRERNAS PERSONLIGA SÄKERHET SAMT KLAGOMÅL
Motivering
Rubriken är anpassad till de ändringsförslag som föredraganden föreslår i detta kapitel.
Ändringsförslag
99
Säkerhet
Resenärernas personliga säkerhet
Motivering
”Säkerhet för järnvägsföretaget” är enligt föredraganden ett felaktigt valt begrepp.
Det rör sig här om resenärernas personliga säkerhet, skydd mot brottslighet i mindre skala, etc.
Ändringsförslag
100
1.
Järnvägsföretag skall vidta erforderliga åtgärder för att sörja för en hög säkerhetsnivå på järnvägsstationer och tåg.
De skall förebygga risker som kan hota resenärernas säkerhet och på ett effektivt sätt åtgärda sådana risker som uppkommer inom järnvägsföretagets ansvarsområde.
1.
Järnvägsföretag och stationsförvaltare skall vidta erforderliga åtgärder för att sörja för en hög nivå på den personliga säkerheten på järnvägsstationer och tåg.
De skall förebygga risker som kan hota resenärernas säkerhet och på ett effektivt sätt åtgärda sådana risker som uppkommer inom järnvägsföretagets ansvarsområde.
Motivering
Det rör sig här om resenärernas personliga säkerhet, skydd mot brottslighet i mindre skala, etc. Även stationsföreståndarna måste sörja för den personliga säkerheten, särskilt på järnvägsstationerna.
Ändringsförslag
101
Artikel 33
Artikel 33
utgår
Kvalitetsnormer
1.
Kvalitetsnormerna skall åtminstone omfatta de punkter som anges i bilaga IV.
2.
Järnvägsföretag skall kontrollera kvaliteten på sin verksamhet och detta skall avspeglas i kvalitetsnormerna.
Järnvägsföretagen skall varje år, tillsammans med sin årsrapport, offentliggöra en rapport om kvaliteten på sin verksamhet.
Resultaten skall även offentliggöras på järnvägsföretagens webbplats på Internet.
Motivering
Denna förordning reglerar resenärernas rättigheter och skyldigheter vid tågresor.
Föredraganden anser att järnvägsföretagens kvalitet i första hand är en fråga för järnvägsföretagen som är bäst skickade att känna sina kunders önskningar och att svara upp mot dessa.
Det är olämpligt att lagstiftaren intar företagarens plats.
Föredraganden ser inte heller något mervärde i en rapport som ett järnvägsföretag offentliggör om sina egna kvalitetsnormer.
Det ankommer på tredje part (journalister, konsumentorganisationer, etc.) att bedöma järnvägsföretagens kvalitet och slå larm om järnvägsföretag som inte lever upp till kvalitetskraven.
Ändringsförslag
102
Artikel 33a
Oberoende genomgång
Europeiska järnvägsbyrån skall göra en oberoende genomgång av hur effektiv sektorns självreglering är och den skall göra det lättare att jämföra järnvägsföretagen med varandra.
Motivering
Förslaget innehåller fullständig självreglering.
Järnvägsföretagens resultat måste också kunna bedömas av ett mer oberoende organ.
Europeiska järnvägsbyrån skulle kunna ta på sig denna uppgift.
Ändringsförslag
103
1.
1.
Ändringsförslag
104
2.
Resenärer får rikta klagomål avseende internationella resor till vilket som helst av de järnvägsföretag som deltagit i bedrivandet av trafiken, eller till det försäljningsställe där de köpte biljetten.
2.
Resenärer får rikta klagomål till vilket som helst av de järnvägsföretag som deltagit i bedrivandet av trafiken, eller till det försäljningsställe där de köpte biljetten.
Ändringsförslag
105
3.
Klagomålet får lämnas på det eller de språk som används i de medlemsstater där resan ägde rum, på det språk som används på den ort där biljetten köptes eller på engelska , franska eller tyska .
3.
Klagomålet får lämnas åtminstone på det eller de språk som används i de medlemsstater där resan ägde rum, eller på engelska.
Ändringsförslag
106
4.
Detta kan innebära att de besvarar klagomålet i ett ställföreträdande eller efterföljande järnvägsföretags ställe, eller på stationsförvaltarens, researrangörens och/eller infrastrukturförvaltarens vägnar.
Om det försäljningsställe som tar emot klagomålet inte är ett av de järnvägsföretag som bedrev trafiken på en del av den berörda sträckan, får försäljningsstället vidarebefordra klagomålet till rätt adress; det skall då informera resenären om detta.
utgår
Ändringsförslag
107
6.
utgår
Motivering
Denna förordning reglerar resenärernas rättigheter och skyldigheter vid tågresor.
Föredraganden anser att järnvägsföretagens kvalitet i första hand är en fråga för järnvägsföretagen som är bäst skickade att känna sina kunders önskningar och att svara upp mot dessa.
Det är olämpligt att lagstiftaren intar företagarens plats.
Föredraganden ser inte heller något mervärde i en rapport som ett järnvägsföretag offentliggör om sina egna kvalitetsnormer.
Det ankommer på tredje part (journalister, konsumentorganisationer, etc.) att bedöma järnvägsföretagens kvalitet och slå larm om järnvägsföretag som inte lever upp till kvalitetskraven.
Ändringsförslag
108
Artikel 36
1.
Resenären skall vid mottagandet av biljetten kontrollera att den har utfärdats i enlighet med hans eller hennes instruktioner.
Resenären måste ha en giltig biljett från resans början, såvida det inte var omöjligt att köpa en biljett på den större järnvägsstation från vilket tåget avgick på grund av att biljettkontoret var stängt eller på grund av att biljettautomaten var ur funktion.
I detta fall skall resenären omedelbart underrätta den ansvariga tågpersonalen om detta.
Resenären skall på begäran visa sin biljett för den ansvariga tågpersonalen .
2.
Järnvägsföretagen får kräva att
a) resenärer som inte kan uppvisa en giltig biljett, utöver transportavgiften, betalar en tilläggsavgift som uppgår till högst 100 % av transportavgiften,
Järnvägsföretagen skall kräva att resenären avbryter sin resa, utan rätt till ersättning för färd- eller platsbiljetter, om resenären
a) utgör en fara för tågpersonalens eller andra resenärers säkerhet, eller
b) utgör en fara för tågets säkerhet, eller
c) stör tågpersonalen eller andra resenärer genom ett olämpligt beteende, exempelvis genom att röka där detta är förbjudet eller genom vandalism, förolämpningar eller våld .
Motivering
När förordningen och COTIF stämmer överens anser föredraganden det lämpligt att hänvisa till COTIF-fördraget.
Det måste dock understrykas att resenärer under vissa förutsättningar kan köpa biljett ombord på tåget (se vidare ändringsförslag till artikel 6.4), en möjlighet som inte finns enligt COTIF.
Ändringsförslag
109
Artikel 37
Informationsskyldighet
Information till resenärerna om deras rättigheter
Järnvägsföretag skall på lämpligt sätt informera allmänheten om sina eventuella planer på att upphöra med internationell trafik .
Järnvägsföretag , stationsförvaltare och researrangörer skall informera resenärerna om de rättigheter och skyldigheter som de har enligt denna förordning .
Kommissionen skall för detta syfte ställa en sammanfattning av denna förordning, på ett för resenärerna begripligt språk, till förfogande för järnvägsföretag, stationsförvaltare och researrangörer.
Motivering
I direktiv 2001/14, bilaga III, återfinns strikta lagstadgade tidsfrister för att fastställa tidtabeller.
Därför är det överflödigt att ta upp en sådan informationsskyldighet i denna förordning.
Föredraganden är däremot positiv till information, t.ex. via affischer, om resenärernas rättigheter.
Kommissionen har tagit fram affischer om flygresenärernas rättigheter.
Affischerna finns nu uppsatta på flygplatserna.
Föredraganden anser att liknande information bör finnas på järnvägsstationer och perronger.
Föredraganden anser att det är mycket bättre att informera resenärerna om de rättigheter och skyldigheter som de har enligt denna förordning.
Ändringsförslag
110
1.
Varje medlemsstat skall utse ett organ som skall ansvara för att kontrollera efterlevnaden av denna förordning.
I tillämpliga fall skall detta organ vidta erforderliga åtgärder för att se till att resenärernas rättigheter tillvaratas .
b) ett organ som medlar då dispyt uppstår om dess tillämpning och som efterlever de principer som anges i kommissionens rekommendation 2001/310/EG av den 4 april 2001 om principer som skall tillämpas på extrajudiciella organ som deltar i reglering av konsumenttvister,
I lämpliga fall skall dessa organ vidta de åtgärder som krävs för att se till att resenärernas rättigheter respekteras.
I detta syfte skall järnvägsföretagen se till att resenärerna får information om hur man kontaktar relevanta tillsynsmyndigheter i de enskilda medlemsstaterna .
______
1 EGT L 109, 19.4.2001, s.
56.
Motivering
Ingen uppskattning har gjorts av kostnaderna av att upprätta och administrera en tillsynsordning.
Medling skulle kunna vara ett mer kostnadseffektivt sätt att lösa många klagomål.
Tillsynen bör vara frivillig i de fall där det finns ett medlingsförfarande som uppfyller kriterierna för kompetens och oberoende (såsom dessa fastslås i kommissionens rekommendation 2001/310/EG).
Ändringsförslag
111
2a.
Järnvägsföretag och stationsförvaltare skall se till att resenärerna på lämpligt sätt på stationerna och tågen informeras om hur man kan kontakta regleringsorganet.
Motivering
Föredraganden vill med detta garantera att resenärerna ges möjlighet att lämna in klagomål.
Ändringsförslag
112
2b.
Det organ som skall upprättas enligt punkt 1 skall regelbundet offentliggöra hur många klagomål som inkommit från resenärerna och vad dessa klagomål gäller.
Motivering
Med detta ändringsförslag vill föredraganden bidra till öppenhet och stimulera järnvägsföretagen till förbättring av sitt tjänsteutbud.
Ändringsförslag
113
Denna förordning träder i kraft 20 dagar efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning träder i kraft 1 år efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Motivering
Med tanke på att det handlar om lagstiftning som är direkt tillämpbar i medlemsstaterna och som medför många förpliktelser för de berörda är det önskvärt att ge dem mera tid innan man tillämpar dessa nya bestämmelser.
Föredraganden konstaterar dessutom att den nyligen antagna förordningen om nekad ombordstigning inom luftfarten också kommer att träda i kraft först efter 1 år.
Ändringsförslag
114
Bilaga I, rubrik 1, strecksats 5
Möjligheten att ta med cyklar samt gällande villkor.
Möjligheten att ta med cyklar och andra fordon samt gällande villkor.
Motivering
Det mesta av informationen måste ges före resans början, eftersom man efter resan så snart som möjligt beger sig till bestämmelseorten, särskilt efter en försening och därav följande möjliga klagomål.
För resenärerna är all information om transportmöjligheter vid framkomsten ett plus som kommer att locka resenärer till tåget.
Ändringsförslag
115
Bilaga I, rubrik 1, strecksatserna 8a och 8b (nya)
Information om intermodala möjligheter (buss, spårvagn, tunnelbana, pendeltåg, cykeluthyrning m.m.) vid ankomsten.
Information om rutiner och kontaktmöjligheter för inlämning av klagomål och vid förlust av resgods.
Motivering
Det mesta av informationen måste ges före resans början, eftersom man efter resan så snart som möjligt beger sig till bestämmelseorten, särskilt efter en försening och därav följande möjliga klagomål.
För resenärerna är all information om transportmöjligheter vid framkomsten ett plus som kommer att locka resenärer till tåget.
Ändringsförslag
116
Bilaga I, rubrik 3, strecksats 2
Förfaranden för inlämnande av klagomål.
Förfaranden och kontaktmöjligheter för inlämnande av klagomål.
Motivering
Det mesta av informationen måste ges före resans början, eftersom man efter resan så snart som möjligt beger sig till bestämmelseorten, särskilt efter en försening och därav följande möjliga klagomål.
För resenärerna är all information om transportmöjligheter vid framkomsten ett plus som kommer att locka resenärer till tåget.
Ändringsförslag
117
Bilaga I, rubrik 3, strecksats 2a (ny)
Denna information skall ges minst på de språk som talas i den medlemsstat där tjänsten utförs.
Ändringsförslag
118
Bilaga II, strecksats 3a (ny)
Uppgifter om huruvida och till vilket datum ersättning kan erhållas.
Motivering
Eftersom det finns skräddarsydda priserbjudanden för många målgrupper uppstår det alltid problem när resenärer begär att få ersättning för en biljett med prisreduktion som de inte använt, eftersom det finns väsentliga skillnader mellan biljetter till fullt pris och nedsatta biljetter även beroende på bokningsform.
Ändringsförslag
119
Bilaga II, strecksats 4a (ny)
Kriterier som komfort, höghastighet m.m., som bidrar till att tillägg/påslag gör biljetten och/eller den tillhandahållna tjänsten dyrare en konventionella tjänster.
Motivering
Ändringsförslag
120
Bilaga III
Denna bilaga utgår.
Motivering
De skadestånd vid förseningar som kommissionen föreslår är inte anpassade till bestämmelserna i den nyligen antagna förordningen för luftfarten (förordning (EG) nr 261/2004).
Skillnaden mellan vanliga tåg och höghastighetståg är svår att tillämpa i praktiken.
Föredraganden inser inte vitsen med denna skillnad, särskilt som skadeståndet räknas som procent av biljettpriset och detta sålunda hur som helst kommer att bli större för höghastighetsförbindelser.
Hur lång tid tågresan tar är inte heller ett relevant kriterium.
Föredraganden väljer att införa ett förenklat ersättningssystem i den relevanta artikeln.
Ändringsförslag
121
Bilaga IV
Denna bilaga utgår.
Motivering
Då artikel 33 föreslås utgå faller också bilagan bort.
MOTIVERING
Kommissionens förslag
Kommissionen konstaterar att marknadsandelen för internationella tågresor minskar, framför allt som följd av konkurrensen från billiga flygbolag.
Kommissionen anser det nödvändigt, också med tanke på kundernas klagomål, att förbättra tjänsteutbudet inom den spårbundna trafiken genom en förordning som tillerkänner resenärerna vissa rättigheter.
Dessa rättigheter går ibland längre än vad som är avtalat inom den mellanstatliga organisationen för internationell tågtrafik (OTIF)
CIV-bihang i COTIF-fördraget (enhetliga regler för avtal om internationell järnvägsbefordran av resande). .
Förslaget innehåller bl.a. bestämmelser om tillgänglighet till information, hur transportavtal ingås, järnvägsföretags ansvarighet, skadestånd till resenärer, ersättning vid förseningar, funktionshindrade personers resor, transporttjänstens kvalitet och behandlingen av klagomål.
De europeiska järnvägarna undertecknade själva 2002 en stadga med kvalitetsnormer för spårbundna persontransporttjänster.
Då detta är en frivillig överenskommelse som inte medför rättigheter som kan åberopas har kommissionen ansett att man ändå måste gå lagstiftningsvägen.
Reaktioner på kommissionens förslag
Konsumentorganisationerna välkomnar detta förslag och begär att man på vissa punkter skall gå ännu längre, t.ex. genom att ge vissa grupper (äldre, funktionshindrade) ännu bättre skydd och ytterligare assistans.
Järnvägsföretagen är däremot helt emot förordningen.
De visar på sina egna ansträngningar (bl.a. den ovannämnda stadgan) och hävdar att konkurrensen mellan företagen och med andra transportsätt redan är en tillräcklig sporre för förbättring av tjänsteutbudet.
De pekar också på de stora skillnader som finns när det gäller gränsöverskridande järnvägstjänster.
Detta borde medföra skräddarsydda tjänster i stället för en gemensam europeisk (minimi)nivå för tjänsteutbudet.
Rådet verkar ge detta förslag låg prioritet.
Medan man redan har hunnit långt vad gäller förslaget till direktiv om certifiering av tågförare har man hittills inte ägnat några överläggningar åt detta förslag.
Föredragandens ståndpunkt
Föredraganden är i princip positiv till en förordning som reglerar tågresenärernas rättigheter.
Dock anser föredraganden att vi måste ta hänsyn till vad som redan finns internationellt.
Vi får inte utan vidare börja mixtra med bra internationella överenskommelser.
Helheten måste fungera och framför allt komma resenärerna till godo.
Vi måste hålla oss till det nödvändiga och ge företagen chansen att utöver detta minimum överträffa varandra i kvalitet eller ytterligare kontraktsbundna garantier.
Att utforma lagar som reglerar resenärers rättigheter och skyldigheter i hela unionen är ingen enkel sak.
Det visar förslaget från kommissionen.
På några punkter går förslaget mycket långt, texten är ofta mycket detaljerad och innehåller ett antal bestämmelser som inte är praktiskt genomförbara.
Förordningens tillämpningsområde innebär att resenärer som sitter bredvid varandra i ett tåg kan omfattas av olika bestämmelser p.g.a. att en av dem gör en internationell resa medan den andra reser inrikes.
Föredraganden lägger därför fram en rad ändringsförslag med syftet att utvidga förordningens tillämpningsområde, förenkla innehållet i en rad bestämmelser, göra strukturen mer lättläst och göra innehållet praktiskt tillämpbart.
Tillämpningsområde: garanti även för resenärer på inrikes resor
Detta förslag ger rättigheter endast åt resenärer på internationella tågresor, vilket innebär att alla resenärer som gör en internationell resa omfattas av förordningen, även när en nationell tågförbindelse utnyttjas vid resans början eller slut.
T.ex. omfattas en resenär som reser från Bryssel till Liverpool av förordningen när han sitter på Eurostar, men också när han sitter på det nationella tåget mellan London och Liverpool.
Föredraganden finner det tillämpningsområde som kommissionen föreslår förvirrande.
Resenärer på samma tåg skulle omfattas av olika bestämmelser beroende på om de gör en inrikes eller en internationell resa.
Föredraganden vill få bort denna osäkerhet och olikhet beträffande rättigheter och föreslår att tillämpningsområdet utvidgas till att gälla alla tågresor.
I gemenskapslagstiftningen avseende luftfarten görs heller ingen skillnad mellan nationella och internationella flygningar när det gäller skyddet av resenärernas rättigheter och ansvarigheten vid olyckor.
Det finns ingen anledning att ha andra utgångspunkter för järnvägstransporter.
Sambandet mellan förordningen och internationella överenskommelser
Sedan 1980 finns det detaljerade all-europeiska överenskommelser om befordran av resenärer med spårbunden trafik.
Dessa är fastställda i ett bihang till COTIF-fördraget.
CIV-bihanget) regleras i detalj ett antal rättigheter och skyldigheter för resenärerna.
Förordningen handlar till stor del om sådant som också regleras i CIV-bihanget.
I stället för att hänvisa till CIV har kommissionen gjort om samma arbete som den mellanstatliga organisationen för internationell järnvägstrafik (OTIF) har gjort, och ställt samman en ny text, löst baserad på internationella principer och terminologi.
Detta leder till att de två regelsystemen påminner starkt om varandra men skiljer sig åt vad gäller formuleringar, struktur och indelning av materialet.
Detta medför oklarheter för dem som måste rätta sig både efter CIV-bihanget och förordningen.
Föredraganden anser att förordningen bör ansluta till CIV där så är möjligt.
I många fall räcker det med en hänvisning till den relevanta CIV-artikeln.
Detta gäller t.ex. bestämmelserna om ansvarighet och skadestånd vid förkommet eller skadat resgods.
CIV är mycket tydligare inom detta område och innehåller inte bara bestämmelser om resgods och handresgods, utan även om djur som resenärerna har med sig och om fordon (t.ex. biltåg).
Endast i de fall då CIV verkligen är otillräckligt är det önskvärt med ytterligare bestämmelser.
T.ex. föreslår föredraganden att man avviker från det maximala skadestånd som CIV anger för skadad eller förkommen rullstol eller andra medicinska hjälpmedel.
Förslagets struktur
Indelningen av förordningen är inte helt logisk.
T.ex. är bestämmelserna om ansvarighet vid död eller skada placerade i ett annat kapitel än bestämmelserna om skadestånd vid död eller skada.
Föredraganden har försökt göra texten mer logisk och lättläst genom att flytta om eller sammanföra ett antal artiklar.
Föredraganden har också försökt förenkla ett antal formuleringar och definitioner.
Att göra förslaget praktiskt genomförbart
Föredraganden anser att det måste garanteras en miniminivå för rättigheterna, men att allt inte behöver regleras i detalj.
Företagen måste kunna göra kommersiella avvägningar och stimuleras att själva komma med uppfinningsrika lösningar för att göra tågresandet attraktivare för resenärerna.
Överreglering kan dessutom leda till ökande kostnader som tjänsteleverantören måste övervältra på resenärerna och som gör att tågresorna blir dyrare och ytterligare tappar mark till bilen och andra transportmedel.
På så vis skulle dessa välmenande bestämmelser förfela sin verkan.
Föredraganden slår fast att tillämpningen av kommissionens förslag på ett antal punkter kommer att leda till tunga administrativa bördor som inte står i proportion till vad en resenär rimligtvis kan förvänta sig av järnvägsföretaget.
Det gäller t.ex. systemet för skadestånd.
I tabellen i bilaga III bestäms skadestånden efter tågtyp (höghastighetståg eller vanligt tåg) och resans varaktighet.
Föredraganden anser att det finns endast ett viktigt kriterium: hur stor förseningen är.
Detta är den enda aspekt som bör spela någon roll när skadeståndet skall bestämmas.
Dessutom förordar föredraganden en höjning av miniminivån.
Obligatoriskt skadestånd är önskvärt först fr.o.m. en timmes försening (inte 30 minuter som kommissionen föreslår).
Naturligtvis kan järnvägsföretagen sätta en lägre gräns, men det är då ett kommersiellt övervägande som företagen själva står för.
Föredraganden föreslår att byta ut bestämmelserna om följdskada mot en mer realistisk formulering från den nyligen antagna förordningen om nekad ombordstigning inom luftfarten.
Enligt denna bestämmelse är det möjligt att på basis av nationell lagstiftning kräva ytterligare skadestånd vid förseningar.
Förslaget är för detaljerat på några punkter och tappar fokus på det viktigaste.
Om vi tittar på definitionen av ”försening” förklarar det ett och annat.
Föredraganden försöker därför förenkla några saker och, om det är nödvändigt, låta dem utgå.
Kompletterande förslag
Föredraganden föreslår att förslaget om att järnvägsföretagen själva skall bestämma sina kvalitetsnormer utgår, och att man i stället inrättar oberoende organ för järnvägsresenärernas klagomål.
Hit kan resenärerna vända sig om järnvägsföretagen inte respekterar resenärernas rättigheter, såsom de beskrivs i denna förordning, och sedan struntar i kundernas klagomål.
Föredraganden föreslår, såsom redan nämnts ovan, att skadestånd skall vara obligatoriskt först fr.o.m. en timmes försening.
Däremot förordar han att det skall finnas ersättningsbestämmelser för resenärer som har abonnemang och råkar ut för upprepade (kortare) förseningar inom en viss tidsperiod.
Sådana bestämmelser finns redan i ett antal medlemsstater, bl.a. i Förenade kungariket.
ÄRENDETS GÅNG
Titel
Förslag till Europaparlamentets och rådets förordning om internationella tågresenärers rättigheter och skyldigheter
Referensnummer
KOM(2004)0143 – C6-0003/2004 – 2004/0049(COD)
Rättslig grund
art.
Grund i arbetsordningen
Framläggande för parlamentet
4.3.2004
Ansvarigt utskott Tillkännagivande i kammaren
TRAN 15.9.2004
Rådgivande utskott Tillkännagivande i kammaren
IMCO 15.9.2004
Inget yttrande avges Beslut
IMCO 31.8.2004
Förstärkt samarbete Tillkännagivande i kammaren
Föredragande Utnämning
Dirk Sterckx 1.9.2004
Tidigare föredragande
Förenklat förfarande Beslut
Bestridande av den rättsliga grunden JURI:s yttrande
Ändrad anslagstilldelning BUDG:s yttrande
Samråd med Europeiska ekonomiska och sociala kommittén Beslut i kammaren
Samråd med Regionkommittén Beslut i kammaren
Behandling i utskott
6.10.2004
23.11.2004
Antagande
19.4.2005
Slutomröstning: resultat
för:
emot:
nedlagda röster:
39
3
1
Slutomröstning: närvarande ledamöter
Margrete Auken, Inés Ayala Sender, Etelka Barsi-Pataky, Philip Bradbourn, Sylwester Chruszcz, Paolo Costa, Michael Cramer, Christine De Veyrac, Armando Dionisi, Petr Duchoň, Saïd El Khadraoui, Robert Evans, Luis de Grandes Pascual, Mathieu Grosch, Ewa Hedkvist Petersen, Jeanine Hennis-Plasschaert, Stanisław Jałowiecki, Georg Jarzembowski, Dieter-Lebrecht Koch, Jaromír Kohlíček, Jörg Leichtfried, Bogusław Liberadzki, Evelin Lichtenberger, Erik Meijer, Janusz Onyszkiewicz, Josu Ortuondo Larrea, Willi Piecyk, Luís Queiró, Reinhard Rack, Luca Romagnoli, Gilles Savary, Ingo Schmitt, Dirk Sterckx, Ulrich Stockmann, Gary Titley, Marta Vincenzi, Corien Wortmann-Kool, Roberts Zīle
Slutomröstning: närvarande suppleanter
Fausto Correia, Den Dover, Willem Schuth
Slutomröstning: närvarande suppleanter (art.
178.2)
Herbert Reul, Eoin Ryan
Ingivande – A6-nummer
28.4.2005
A6-0123/2005
Anmärkningar
SLUTLIG VERSION
A6-0167/2005
***II
ANDRABEHANDLINGS-REKOMMENDATION
om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets förordning om kontroller av kontanta medel som förs in i eller ut ur gemenskapen
(14843/1/2004 – C6‑0038/2005 – 2002/0132(COD))
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Föredragande:
Vincent Peillon
PE 355.777v02-00
Teckenförklaring
* Samrådsförfarandet majoritet av de avgivna rösterna
**I Samarbetsförfarandet (första behandlingen) majoritet av de avgivna rösterna
**II Samarbetsförfarandet (andra behandlingen) majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
*** Samtyckesförfarandet majoritet av parlamentets samtliga ledamöter utom i de fall som avses i artiklarna 105, 107, 161 och 300 i EG-fördraget och artikel 7 i EU-fördraget
***I Medbeslutandeförfarandet (första behandlingen) majoritet av de avgivna rösterna
***II Medbeslutandeförfarandet (andra behandlingen) majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
***III Medbeslutandeförfarandet (tredje behandlingen) majoritet av de avgivna rösterna för att godkänna det gemensamma utkastet
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Parlamentets ändringar markeras med fetkursiv stil.
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING............................................................................................................................8
ÄRENDETS GÅNG..................................................................................................................10
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
(14843/1/2004 – C6‑0038/2005 – 2002/0132(COD) )
(Medbeslutandeförfarandet: andra behandlingen)
Europaparlamentet utfärdar denna resolution
– med beaktande av rådets gemensamma ståndpunkt (14843/1/2004 – C6‑0038/2005 ),
EUT C 67 E, 17.3.2004, s.
259. , en behandling som avsåg kommissionens förslag till Europaparlamentet och rådet ( KOM(2002)0328 )
EGT C 227 E, 24.9.2002, s.
574. ,
– med beaktande av ändringarna i kommissionens förslag ( KOM(2003)0371 )
Ännu ej offentliggjort i EUT. ,
– med beaktande av artikel 62 i arbetsordningen,
– med beaktande av andrabehandlingsrekommendationen från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor ( A6‑0167/2005 ).
1.
Rådets gemensamma ståndpunkt
Parlamentets ändringar
Ändringsförslag från Vincent Peillon
Ändringsförslag
1
Vid tillämpningen av denna förordning bör Europaparlamentets och rådets direktiv 95/46/EG av den 24 oktober 1995 om skydd för enskilda personer med avseende på behandling av personuppgifter och om det fria flödet av sådana uppgifter 1 och Europaparlamentets och rådets förordning (EG) nr 45/2001 av den 18 december 2000 om skydd för enskilda då gemenskapsinstitutionerna och gemenskapsorganen behandlar personuppgifter och om den fria rörligheten för sådana uppgifter 2 tillämpas på den behandling av personuppgifter som utförs av de behöriga myndigheterna i medlemsstaterna.
_______________________
1 EGT L 281, 23.11.1995, s.
31.
2 EGT L 8, 12.1.2001, s.
1.
Ändringsförslag
2
Skäl 14
(14) Denna förordning respekterar de grundläggande rättigheter och iakttar de principer som erkänns framför allt i Europeiska unionens stadga om grundläggande rättigheter.
Ändringsförslag från Vincent Peillon
Ändringsförslag
3
Artikel 7a (ny)
Artikel 7a
Varje uppgift som är konfidentiell eller som lämnats konfidentiellt skall omfattas av tystnadsplikt och skall inte lämnas ut av de behöriga myndigheterna utan uttryckligt tillstånd från den person eller den myndighet som lämnat uppgiften.
Uppgifter får emellertid översändas om de behöriga myndigheterna är skyldiga att göra detta i enlighet med gällande bestämmelser, särskilt inom ramen för rättsliga förfaranden.
Utlämnande och översändande av uppgifter skall ske med strikt beaktande av gällande bestämmelser för skydd av personuppgifter, särskilt direktiv 95/46/EG och förordning (EG) nr 45/2001.
MOTIVERING
Bakgrund
Den 25 juni 2002 lade kommissionen fram ett förslag till förordning om ”kontroller av kontanta medel som förs in i eller ut ur gemenskapen” i syfte att komplettera direktiv 91/308/EEG om penningtvätt.
De två huvudpunkterna i detta förslag var följande: att införa en skyldighet att deklarera in‑ och utförsel av kontanta medel som uppgår till belopp över 15 000 euro samt att förse de behöriga myndigheterna med information om transaktioner som innebär en risk för penningtvätt.
Europaparlamentet lade fram sitt yttrande vid första behandlingen den 15 maj 2003 och antog 23 ändringar.
Merparten av dessa ändringar syftade till att ändra den föreslagna rättsakten.
Europaparlamentet hade i själva verket föredragit ett direktiv i stället för en förordning.
Parlamentet föreslog även att som rättslig grund lägga till artikel 95 i EG-fördraget om tillnärmning av medlemsstaternas lagar och andra författningar om den inre marknadens sätt att fungera.
Parlamentet önskade även att medlemsstaterna skulle få välja mellan två förfaranden: skyldighet att anmäla och skyldighet att deklarera.
Vidare utökades definitionen av begreppet kontanta medel i syfte att inbegripa ett större antal typer av checkar.
Den 1 juli 2003 lade kommissionen fram ett ändrat förslag i vilket den hade godtagit två ändringar (13 och 15) helt och hållet och tre ändringar (2, 11 och 21) till viss del.
Rådets gemensamma ståndpunkt
Den 17 februari 2005 antog rådet sin gemensamma ståndpunkt med kvalificerad majoritet.
Rådet tillbakavisade parlamentets förslag om att omvandla rättsakten till ett direktiv, men det tillstyrkte att artikel 95 i EG-fördraget skulle läggas till som rättslig grund.
När det gäller obligatorisk deklaration stöder rådet kommissionens förslag, men ställer sig inte positivt till det system med valmöjlighet som parlamentet föreslagit och som skulle ha gjort det möjligt för medlemsstaterna att välja mellan ett system med deklaration och ett system med anmälan.
Icke desto mindre har rådet infört större flexibilitet genom att tillåta tre olika typer av deklaration: muntlig, skriftlig eller elektronisk.
Rådet har sänkt tröskeln till 10 000 euro, från de 15 000 euro som ursprungligen avsågs.
Definitionen av begreppet kontanta medel har utökats i enlighet med parlamentets förslag, men även i enlighet med den särskilda rekommendationen IX från arbetsgruppen för finansiella åtgärder mot penningtvätt (FATF), i syfte att åstadkomma ökad samstämdhet mellan de bestämmelser som fastställs på gemenskapsnivå respektive internationellt.
De upplysningar som tas emot med hjälp av deklarationer och kontroller skall göras tillgängliga för finansunderrättelseenheterna.
Upplysningar kan registreras även om de medel som förs in eller ut uppgår till ett värde som är lägre än 10 000 euro, om det finns tecken på olaglig verksamhet.
Vidare har rådet förenklat bestämmelserna om påföljder.
Medlemsstaterna skall införa effektiva, avskräckande och proportionerliga påföljder för brott mot skyldigheten att deklarera in- och utförsel av kontanta medel vid passage av Europeiska unionens yttre gränser.
Föredragandens hållning
Föredraganden välkomnar rådets förslag.
Med tanke på den ökande oro som penningtvätten skapar och den roll penningtvätten spelar inom organiserad brottslighet och terrorverksamhet är det viktigt att lagstifta på detta område och att effektivt kontrollera in- och utförsel av kontanta medel vid våra gränser.
I rapporten ”Moneypenny”, som var namnet på en gemensam insats som gjordes av medlemsstaternas tullmyndigheter mellan september 1999 och februari 2000, underströks att de befintliga kontrollerna i kampen mot penningtvätt delvis blir ineffektiva till följd av skillnaderna i metoder för övervakning av flödet av kontanta medel vid gränserna.
De markanta skillnader som konstaterades i medlemsstaternas tillvägagångssätt synliggjorde att det finns stora brister i övervaknings- och skyddssystemen och att det saknas ett övergripande skydd på gemenskapsnivå.
Det är därför nödvändigt och brådskande att unionen, särskilt efter det att euron infördes, skapar en enhetlig och effektiv strategi på detta område.
Föredraganden anser att den rättsakt som föreslagits är den mest lämpliga, särskilt för att underlätta informationsutbytet mellan medlemsstaterna.
Vid en jämförelse med det ursprungliga förslaget verkar denna förordning tydligare och mer användbar.
De ändringsförslag som föredraganden föreslår syftar till att införa ändringar som leder till ett bättre skydd av personuppgifter, vilket är en fråga som parlamentet uttalat sig om vid flera tillfällen (ändringsförslagen 2, 3, 4 och 5).
Med tanke på att det är brådskande att införa en effektiv bekämpning av penningtvätt önskar föredraganden, som beklagar den redan långa fördröjningen, att samarbetet med rådet blir framgångsrikt, så att det blir möjligt att nå en överenskommelse vid andra behandlingen.
ÄRENDETS GÅNG
Titel
Rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets förordning om kontroller av kontanta medel som förs in i eller ut ur gemenskapen
Referensnummer
14843/1/2004 – C6‑0038/2005 – 2002/0132(COD)
Rättslig grund
art.
251.2 och art.
95 och 135 EG-fördraget
Grund i arbetsordningen
Parlamentets första behandling – P5-nummer
15.5.2003
T5-0214/2003
Kommissionens förslag
KOM(2002)0328 – C5‑0291/2002
Kommissionens ändrade förslag
KOM(2003)0371
Mottagande av den gemensamma ståndpunkten: tillkännagivande i kammaren
24.2.2005
Ansvarigt utskott Tillkännagivande i kammaren
LIBE 24.2.2005
Föredragande Utnämning
Tidigare föredragande
Behandling i utskott
26.4.2005
26.5.2005
Antagande
26.5.2005
Slutomröstning: resultat
för:
emot:
nedlagda röster:
29
Slutomröstning: närvarande ledamöter
Alexander Nuno Alvaro, Edit Bauer, Johannes Blokland, Mihael Brejc, Michael Cashman, Giusto Catania, Charlotte Cederschiöld, Carlos Coelho, Antoine Duquesne, Patrick Gaubert, Lilli Gruber, Magda Kósáné Kovács, Wolfgang Kreissl-Dörfler, Barbara Kudrycka, Stavros Lambrinidis, Romano Maria La Russa, Henrik Lax, Edith Mastenbroek, Claude Moraes, Martine Roure, Ioannis Varvitsiotis, Stefano Zappalà
Slutomröstning: närvarande suppleanter
Ignasi Guardans Cambó, Luis Francisco Herrero-Tejedor, Sophia in 't Veld, Jean Lambert, Siiri Oviir, Vincent Peillon, Kyriacos Triantaphyllides
Slutomröstning: närvarande suppleanter (art.
178.2)
Ingivande – A6-nummer
30.5.2005
A6‑0167/2005
Anmärkningar
...
A6-0206/2005
***I
BETÄNKANDE
om förslaget till Europaparlamentets och rådets förordning om europeiska grupperingar för gränsöverskridande samarbete (EGGS)
(KOM(2004)0496 – C6‑0091/2004 – 2004/0168(COD))
Utskottet för regional utveckling
Föredragande:
Jan Olbrycht
PE 357.502v02-00
Teckenförklaring
* Samrådsförfarandet majoritet av de avgivna rösterna
**I Samarbetsförfarandet (första behandlingen) majoritet av de avgivna rösterna
**II Samarbetsförfarandet (andra behandlingen) majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
*** Samtyckesförfarandet majoritet av parlamentets samtliga ledamöter utom i de fall som avses i artiklarna 105, 107, 161 och 300 i EG-fördraget och artikel 7 i EU-fördraget
***I Medbeslutandeförfarandet (första behandlingen) majoritet av de avgivna rösterna
***II Medbeslutandeförfarandet (andra behandlingen) majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
***III Medbeslutandeförfarandet (tredje behandlingen) majoritet av de avgivna rösterna för att godkänna det gemensamma utkastet
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Parlamentets ändringar markeras med fetkursiv stil.
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................20
ÄRENDETS GÅNG..................................................................................................................24
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till Europaparlamentets och rådets förordning om europeiska grupperingar för gränsöverskridande samarbete (EGGS)
( KOM(2004)0496 – C6‑0091/2004 – 2004/0168(COD) )
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2004)0496 )
Ännu ej offentliggjort i EUT. ,
– med beaktande av artikel 51 i arbetsordningen,
– med beaktande av betänkandet från utskottet för regional utveckling ( A6‑0206/2005 ).
Kommissionens förslag
Parlamentets ändringar
Ändringsförslag
1
Titel
Förslag Europaparlamentets och rådets förordning om europeiska grupperingar för gränsöverskridande samarbete ( EGGS )
Förslag Europaparlamentets och rådets förordning om europeiska grupperingar för territoriellt samarbete ( EGTS )
Motivering
I den allmänna förordningen om strukturfonderna fastslås att territoriellt samarbete är ett nytt mål 3 som inbegriper gränsöverskridande, transnationellt och interregionalt samarbete.
För att termerna skall bli konsekventa bör titeln och förkortningen ändras.
Ändringsförslag
2
Skäl 1
För att få en harmonisk utveckling i hela EU och en starkare ekonomisk, social och regional sammanhållning måste samarbetet över nationsgränserna intensifieras.
Därför måste det skapas bättre förutsättningar för ett sådant samarbete.
För att få en harmonisk utveckling i hela EU och en starkare ekonomisk, social och regional sammanhållning måste det territoriella samarbetet intensifieras.
Därför måste det skapas bättre förutsättningar för ett sådant samarbete.
Motivering
I alla bestämmelser i förordningen där man använder uttrycket ”gränsöverskridande samarbete” eller ”samarbete över gränserna” och åsyftar territoriellt samarbete bör man ändra dessa ord till "territoriellt".
Ändringsförslag
3
Skäl 5
(5) Resurserna för det regionala samarbetet ökas genom rådets förordning (EG) nr (…) om allmänna bestämmelser för Europeiska regionala utvecklingsfonden, Europeiska socialfonden och Sammanhållningsfonden.
(5) Resurserna för det regionala eller territoriella samarbetet ökas på tre områden: gränsöverskridande, interregionalt och transnationellt samarbete, genom rådets förordning (EG) nr (…) om allmänna bestämmelser för Europeiska regionala utvecklingsfonden, Europeiska socialfonden och Sammanhållningsfonden
Ändringsförslag
4
Skäl 6
(6) Det är nödvändigt att underlätta och främja ett gränsöverskridande samarbete även i de fall där EU inte ger något ekonomiskt stöd.
(6) Det är nödvändigt att underlätta och främja ett territoriellt samarbete även i de fall där EU inte ger något ekonomiskt stöd.
Motivering
Se motiveringen till ändringsförslag 2.
Ändringsförslag
5
Skäl 7
(7) För att undanröja hindren för ett gränsöverskridande samarbete behövs det ett nytt instrument på EU-nivå som gör det möjligt att bilda samarbetsgrupperingar som har status som juridiska personer, nedan kallade ”europeiska grupperingar för gränsöverskridande samarbete” (EGGS) , eller ”grupperingar”.
Det bör emellertid inte bli obligatoriskt att bilda sådana grupperingar.
(7) För att undanröja hindren för ett territoriellt samarbete behövs det ett nytt instrument på EU-nivå som gör det möjligt att bilda samarbetsgrupperingar som har status som juridiska personer, nedan kallade ”europeiska grupperingar för territoriellt samarbete” (EGTS) , eller ”grupperingar”.
Se motiveringen till ändringsförslag 2.
Ändringsförslag
6
Skäl 7a (nytt)
(7a) De avtal som ingåtts om gränsöverskridande, interregionalt och övernationellt samarbete mellan medlemsstater och/eller regionala och lokala instanser kan fortsätta att tillämpas.
Motivering
De rättsliga bestämmelser som ligger till grund för mellanstatliga avtal, till exempel Karlsruheavtalen, får inte begränsas i sitt tillämpningsområde till följd av att förordningen träder i kraft.
Ändringsförslag
7
Skäl 9
(9) Grupperingens uppgifter och behörighet bör anges i ett samarbetsavtal som medlemmarna själva utformar, nedan kallat ”avtal”.
(Berör inte den svenska versionen.)
Motivering
(Berör inte den svenska versionen.)
Ändringsförslag
8
Skäl 10
(10) Medlemmarna kan välja mellan att bilda en gruppering som får status som separat juridisk person eller att låta en av medlemmarna fylla den funktionen.
(10) Medlemmarna bildar en gruppering som får status som separat juridisk person och som får låta en av medlemmarna fylla den funktionen.
Ändringsförslag
9
Skäl 11
(11) En gruppering bör kunna agera för att genomföra dels gränsöverskridande samarbetsprogram som medfinansieras av EU, t.ex. via strukturfonderna i enlighet med förordning (EG) nr (…) och förordning (EG) nr (…) om Europeiska regionala utvecklingsfonden, dels transnationella och interregionala samarbetsprogram, eller för att utan stöd från EU och på medlemsstaternas, regionernas eller de lokala instansernas eget initiativ genomföra ett gränsöverskridande samarbete.
(11) En gruppering bör kunna agera för att genomföra dels gränsöverskridande samarbetsprogram som medfinansieras av EU, t.ex. via strukturfonderna i enlighet med förordning (EG) nr (…) och förordning (EG) nr (…) om Europeiska regionala utvecklingsfonden, dels transnationella och interregionala samarbetsprogram, eller för att utan stöd från EU och/eller på medlemsstaternas, regionernas eller de lokala instansernas eget initiativ genomföra ett territoriellt samarbete.
Ändringsförslag
10
Skäl 11a (nytt)
(11a) Kommissionen bör säkerställa synergieffekter mellan denna förordning och Europarådets tilläggsprotokoll* till Europeiska ramkonventionen om samarbete mellan lokala och regionala samhällsorgan avseende inrättandet av euroregionala samarbetsgrupperingar (ESG).
____________
* nr 3 i form av utkast
Motivering
EGGS-förordningen rör endast medlemsstater, medan de parter som är inblandade i gränsöverskridande, transnationellt och interregionalt samarbete däremot omfattar kandidatländer och tredje länder.
För dessa gäller endast tilläggsprotokoll nr 3 till Europeiska ramkonventionen om samarbete mellan lokala och regionala samhällsorgan och därför föreslås det att kommissionen och Europarådet skall samarbeta för att harmonisera de två utkasten.
Ändringsförslag
11
Skäl 13
(13) Ett avtal bör inte få innehålla något om en regional eller lokal instans befogenhet att utöva samhällelig makt, t.ex. polismakt eller rätten att utfärda olika former av bestämmelser.
(Berör inte den svenska versionen.)
Skäl 14
(14) Det är nödvändigt att en gruppering utformar sina egna stadgar och att den skaffar sig egna organ, samt att den har regler för sin budget och för sitt ekonomiska ansvar.
(14) Det är nödvändigt att en gruppering utformar sina egna stadgar och att den skaffar sig egna organ och fastställer beslutsförfaranden samt att den har regler för sin budget och för sitt ekonomiska ansvar.
Motivering
I ett offentligt organs stadgar redogörs alltid för det sätt på vilket beslut fattas.
Därmed undviks problem i samband med beslutsförfaranden samtidigt som större öppenhet skapas i fråga om denna process.
Ändringsförslag
13
Skäl 15
(15) I enlighet med subsidiaritetsprincipen i artikel 5 i fördraget får EU vidta åtgärder om medlemsstaterna inte på ett effektivt sätt kan skapa sådana förutsättningar för ett gränsöverskridande samarbete som anges i den här förordningen och om detta på ett bättre sätt kan åstadkommas på EU-nivå.
I enlighet med den proportionalitetsprincip som åsyftas i ovan nämnda artikel går den här förordningen inte längre än vad som är nödvändigt för att nå målen, eftersom samarbetsgrupperingarna inte blir obligatoriska och eftersom varje medlemsstats egna lagar och författningar beaktas fullt ut.
(15) Eftersom medlemsstaterna inte på ett effektivt sätt kan skapa de rättsliga förutsättningarna inom hela EU för det territoriella samarbete som anges i den här förordningen är det bättre att skapa sådana förutsättningar på EU-nivå.
EU får därmed vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget.
I enlighet med den proportionalitetsprincip som åsyftas i ovan nämnda artikel går den här förordningen inte längre än vad som är nödvändigt för att nå målen, eftersom samarbetsgrupperingarna inte blir obligatoriska och eftersom varje medlemsstats egna lagar och författningar beaktas fullt ut.
Motivering
Se motiveringen till ändringsförslag 2.
Ändringsförslag
14
Artikel 1, rubrik
Europeiska grupperingar för gränsöverskridande samarbete
Europeiska grupperingar för territoriellt samarbete
Motivering
Se motiveringen till ändringsförslag 1.
Ändringsförslag
15
1.
Inom EU kan samarbetsgrupperingar bildas i form av europeiska grupperingar för gränsöverskridande samarbete, nedan kallade ”grupperingar”, enligt de villkor och regler som föreskrivs i den här förordningen.
1.
Inom EU kan samarbetsgrupperingar bildas i form av europeiska grupperingar för territoriellt samarbete, nedan kallade ”grupperingar”, enligt de villkor och regler som föreskrivs i den här förordningen.
Motivering
Se motiveringen till ändringsförslag 2.
3.
En gruppering skall ha till uppgift att underlätta och främja medlemsstaternas och de regionala och lokala instansernas gränsöverskridande samarbete , med målet att stärka den ekonomiska, sociala och regionala sammanhållningen.
3.
En gruppering skall ha till uppgift att underlätta och främja territoriellt (gränsöverskridande, transnationellt och interregionalt) samarbete mellan regionala och lokala instanser inom EU, med målet att stärka den ekonomiska, sociala och regionala sammanhållningen.
Motivering
I förordningen används begreppet regionalt eller territoriellt samarbete.
Ändringsförslag
17
Den medlemsstat vars lagstiftning är tillämplig skall informera de andra medlemsstater som berörs av avtalet om resultatet av varje genomförd kontroll.
Motivering
Det är nödvändigt att fastställa kontrollsystemet för grupperingarnas verksamhet på ett klart och transparent sätt, med beaktande av att grupperingarna består av enheter från olika medlemsstater och att själva grupperingen agerar på grundval av en rättslig ordning från en av medlemsstaterna och står under denna medlemsstats kontroll.
För att försäkra sig om att informationen verkligen når de övriga medlemsstaterna införs en regel som syftar till att informera samtliga medlemsstater som är inblandade i en gruppering om resultaten av de kontroller som genomförts.
3b.
Om det under en längre tid pågått civila eller militära konflikter i gränsområden får grupperingen även ha till uppgift att främja försoning och bistå via fredsskapande program.
Motivering
Gränsområden är ofta skådeplatser för konflikter, vilket har skapat ytterligare och specifika hinder för det gränsöverskridande samarbetet.
Ändringsförslag
19
1.
(Berör inte den svenska versionen.)
Ändringsförslag
20
1.
1.
Ändringsförslag
21
3.
3.
Medlemmarna bildar en gruppering som får status som separat juridisk person och som får låta en av medlemmarna fylla den funktionen.
Motivering
Ändringsförslag
22
Artikel 3, rubrik
Befogenheter
Uppgifter och befogenheter
Motivering
I denna artikel beskrivs inte bara grupperingens befogenheter utan även dess uppgifter.
Ändringsförslag
23
1.
En gruppering skall utföra de uppgifter som medlemmarna ger den i enlighet med den här förordningen.
Dess befogenheter skall anges i ett avtal om gränsöverskridande europeiskt samarbete, nedan kallat ”avtal”, som medlemmarna skall ingå i enlighet med artikel 4.
1.
En gruppering skall utföra de uppgifter som medlemmarna ger den i enlighet med den här förordningen.
Dess befogenheter skall anges i ett avtal om territoriellt europeiskt samarbete, nedan kallat ”avtal”, som medlemmarna skall ingå i enlighet med artikel 4.
Motivering
Se motiveringen till ändringsförslag 2.
Ändringsförslag
24
2.
Inom gränserna för de uppgifter som delegeras till den skall en gruppering agera på medlemmarnas vägnar .
En gruppering skall därför ha den status som en juridisk person har enligt den nationella lagstiftningen .
2.
Motivering
En gruppering är en juridisk person och kan utföra sina uppgifter i eget namn, på eget ansvar och egen risk.
(Naturligtvis förutsätts att en gruppering agerar i de medlemmars intressen som bildat den, även om det inte finns någon juridisk koppling).
Grupperingen har i egenskap av juridisk person den rättskapacitet som är en av de karaktäristiska egenskaperna för en juridisk person.
En gruppering kan utföra de utgifter som delegerats till den direkt (i egenskap av gruppering) eller delegera genomförandet till en av sina medlemmar.
Ändringsförslag
25
3.
En gruppering kan få i uppgift att genomföra program för gränsöverskridande samarbete som medfinansieras av EU, t.ex. via strukturfonderna, men också andra former av sådant samarbete, med eller utan ekonomiskt stöd från EU.
3.
En gruppering kan få i uppgift att genomföra program för territoriellt samarbete som medfinansieras av EU, t.ex. via strukturfonderna, men också andra former av sådant samarbete, med eller utan ekonomiskt stöd från EU.
Motivering
Se motiveringen till ändringsförslag 2.
3a.
Medlemsstater som inte är medlemmar i grupperingen skall inte ha något ekonomiskt ansvar, även om deras regionala, lokala eller offentliga organ deltar som medlemmar.
Detta skall emellertid inte påverka medlemsstaternas finansiella ansvar när det gäller gemenskapsmedel som utnyttjas av en gruppering.
Motivering
De bästa Interreg-programmen har redan infört gränsöverskridande projekt som grundar sig på sådan goodwill som följer på gemensam förvaltning, finansiering och kontroll samt gemensamma garantier.
Syftet med denna förordning är att öka och stärka gränsernas befintliga samarbetspotential genom att koppla samman skilda rättssystem och ge de regionala och lokala organisationerna möjlighet att samarbeta tvärs över gränserna utan att först erhålla medlemsstaternas tillstånd.
Detta leder till ett ökat ansvar.
Medlemsstaterna kan bli medlemmar av grupperingen, men om de inte är medlemmar skall de inte vara ekonomiskt ansvariga för grupperingens verksamhet.
Ändringsförslag
27
Artikel 4, rubrik
Ändringsförslag
28
1.
För varje gruppering skall ett avtal ingås.
1.
För en gruppering skall ett avtal ingås av dess medlemmar .
Ändringsförslag
29
2.
Avtalet skall reglera grupperingens uppgifter, varaktighet och upplösning.
2.
Avtalet skall i synnerhet reglera principerna för verksamheten, grupperingens uppgifter, varaktighet och upplösning.
Ändringsförslag
30
3.
Avtalet skall enbart avse sådant gränsöverskridande samarbete som medlemmarna fattar beslut om.
3.
Avtalet skall enbart avse sådant territoriellt samarbete som medlemmarna fattar beslut om.
Motivering
Se motiveringen till ändringsförslag 2.
Ändringsförslag
31
4.
Avtalet skall reglera varje medlems ansvar gentemot grupperingen och gentemot tredje part.
utgår
Motivering
Ändringsförslag
32
5.
5.
Avtalet skall ange vilken lagstiftning som gäller för grupperingen.
Den tillämpliga lagstiftningen skall vara lagstiftningen i en medlemsstat som berörs av avtalet och där grupperingen har sitt säte.
Ändringsförslag
33
6.
utgår
Motivering
Beskrivningen är oklar, och därför krävs det att frågan avgörs i förordningen och inte i avtalet.
Ändringsförslag
34
6a.
Grupperingen skall vara föremål för den nationella rätt avseende associationers verksamhet som valts av medlemmarna.
Motivering
I kommissionens förslag nämns inga som helst förfaranden för registrering av grupperingar eller övervakning av denna registrering eller den bildade grupperingens förenlighet med nationell lagstiftning i den medlemsstat som valts.
Ändringsförslag
35
7.
7.
Villkoren för beviljandet av koncessioner eller delegeringar av offentliga uppgifter till en gruppering inom ramen för territoriellt samarbete skall anges i avtalet, i enlighet med den tillämpliga nationella lagstiftningen.
Ändringsförslag
36
8.
8.
Avtalet skall skickas till samtliga medlemsstater som berörs av grupperingen, till kommissionen och till Regionkommittén.
Kommissionen skall registrera avtalet i ett offentligt register för alla avtal avseende sådana grupperingar.
Det verkar också motiverat att skapa en databas med alla grupperingar som kan bildas på EU:s territorium och ge Regionkommittén i uppdrag att utföra denna uppgift.
Ändringsförslag
37
2.
Stadgarna skall innehålla följande:
2.
Stadgarna skall innehålla följande:
a) En förteckning över medlemmarna.
a) En förteckning över medlemmarna.
b) Grupperingens mål och uppgifter , samt relationerna mellan grupperingen och dess medlemmar .
b) Grupperingens mål och uppgifter.
c) Grupperingens namn och säte.
c) Grupperingens namn och säte.
d) Grupperingens olika organ, deras befogenheter och funktion, samt antalet medlemsrepresentanter i organen.
d) Grupperingens olika organ, inbegripet en församling som består av företrädare för medlemmarna och en verkställande kommitté, deras befogenheter och funktion, antalet medlemsrepresentanter i organen och ett sekretariat .
Ytterligare organ kan fastställas i stadgarna.
e) Grupperingens beslutsfattande.
e) Grupperingens beslutsfattande.
Motivering
Varje juridisk person skapar sin egen uppsättning organ i enlighet med den lagstiftning som reglerar principerna för dess verksamhet.
Det bör även ingå i grupperingens befogenheter att avgöra på vilket sätt grupperingen skall företrädas, dvs. vem som får företräda grupperingen på ett visst område och huruvida det krävs att en eller flera personer ingår i denna representation när det gäller att ingå avtal, osv.
ia) Formerna för grupperingens upplösning.
Motivering
För att garantera en demokratisk ledning som medger insyn skall varje gruppering ha en församling bestående av företrädare för samtliga dess medlemmar och en ledningsgrupp och/eller en direktör som är ansvariga inför församlingen.
Stadgan kan även innehålla bestämmelser om upplösningen av grupperingen.
Föredragandens ändringsförslag 36, enligt vilket artikel 6 stryks, kompletterar detta ändringsförslag.
Ändringsförslag
39
4.
utgår
Motivering
I ändringsförslag 31 där man inför en ny bestämmelse till artikel 6a (ny), föreslås registreringsförfaranden för grupperingar på grundval av den lagstiftning som gäller för registrering av associationer.
Därför bör man fastslå att en gruppering får status som juridisk person och därmed rättskapacitet att agera i enlighet med den lagstiftning som är tillämplig på registrering av associationer.
Ändringsförslag
40
Artikel 6
Artikel 6
Organ
1.
2.
En gruppering kan inrätta en församling som består av företrädare för medlemmarna.
3.
I stadgarna får det finnas bestämmelser om ytterligare organ.
Motivering
Ändringsförslag
41
Artikel 8, stycke 1
Från och med då skall grupperingens juridiska status erkännas i samtliga medlemsstater.
MOTIVERING
1.
Allmän bakgrund
Inom ramen för den nya målsättningen ”europeiskt territoriellt samarbete” föreslår kommissionen att under perioden 2007-2013 anslå en övergripande budget på 13,5 miljarder euro till gränsöverskridande, transnationellt och interregionalt samarbete.
Detta utgör 4 procent av medlen i strukturfonderna och Sammanhållningsfonden under denna period och innebär en ökning på 14 procent jämfört med perioden 2000–2007.
Europaparlamentet har betonat vikten av gränsöverskridande, transnationellt och interregionalt samarbete för den europeiska integrationen
Den rättsliga grunden till förslaget till Europaparlamentets och rådets förordning om europeiska grupperingar för gränsöverskridande samarbete är artikel 159 tredje stycket i fördraget.
Denna artikel utgör fördragets särskilda rättsliga grund för att vidta särskilda åtgärder utanför fonderna i syfte att uppnå målet om ekonomisk och social sammanhållning enligt artikel 158 i fördraget.
I utkastet till fördrag om upprättande av en konstitution för Europa nämns vid upprepade tillfällen territoriell sammanhållning, och inte bara ekonomisk och social sammanhållning, som ett av unionens mål och som ett område med delad befogenhet.
Artiklarna I-3.3, I-14 och II-96.
Det är i artikel III-220 i konstitutionsförslaget (nuvarande artikel 158 i EG-fördraget) som särskild uppmärksamhet fästs vid bland annat gränsöverskridande regioner.
2.
Målet med kommissionens förslag
Kommissionens förslag ingår i lagstiftningspaketet med förslag till nya förordningar om strukturfonderna för perioden 2007-2013 och innehåller en allmän förordning där gemensamma regler för alla instrument fastställs och särskilda förordningar för Europeiska regionala utvecklingsfonden (ERUF), Europeiska socialfonden (ESF) och Sammanhållningsfonden.
Förslaget ingår också i det övergripande paketet med interna och externa instrument för gränsöverskridande samarbete inom Europeiska unionen (europeiska grupperingar för gränsöverskridande samarbete) med kandidatländerna eller potentiella kandidatländer (föranslutningsinstrumentet) och med tredje länder som Europeiska unionen önskar knyta goda grannskapsförbindelser med (det europeiska grannskaps- och partnerskapsinstrumentet).
Det framkommer av motiveringen och inledningen till förslaget ( skäl 1 i kommissionens förslag ) att syftet är att uppnå fördragets mål om ekonomisk och social sammanhållning (artikel 158 i EG-fördraget), att stärka det gränsöverskridande samarbetet genom att förbättra de förutsättningar under vilka gränsöverskridande åtgärder genomförs.
Kommissionens förslag syftar på så sätt till att minska hindren och svårigheterna att administrera åtgärder kring det gränsöverskridande, transnationella och interregionala samarbetet inom ramen för olika nationella regler och rutiner, genom att inrätta ett samarbetsinstrument på gemenskapsnivå som gör att möjligt att på gemenskapens territorium skapa europeiska grupperingar som är juridiska personer för gränsöverskridande samarbete (EGGS) som det inte skall vara obligatoriskt att utnyttja ( skäl 2 och 7 och artikel 1 i kommissionens förslag ).
3.
Föredragandens utvärdering av de främsta kännetecknen för ”europeiska grupperingar för gränsöverskridande samarbete” (EGGS)
Ø Förslaget till förordning om ”europeiska grupperingar för gränsöverskridande samarbete” syftar till att erbjuda en lämplig ram för att underlätta det gränsöverskridande, transnationella och interregionala samarbetet (titel, skäl 1 och artikel 1 i kommissionens förslag).
Föredraganden anser att detta nya instrument bör benämnas ”europeiska grupperingar för territoriellt samarbete” (EGTS) som en anpassning till de tre dimensionerna i det nya målet om europeiskt territoriellt samarbete som föreslagits av kommissionen för perioden 2007‑2013: gränsöverskridande, transnationellt och interregionalt ( ändringsförslag 1, 2, 5, 6, 8, 10, 12, 13, 14, 20, 22, 24, 27 och 32) .
Föredragen anser också att ikraftträdandet av denna förordning varken får påverka giltigheten i existerande överenskommelser eller möjligheterna för de medlemsstater som så önskar att förhandla bilaterala eller multilaterala internationella avtal som syftar till gränsöverskridande samarbete (ändringsförslag 7) .
1.
Sammansättningen av grupperingarna ( artikel 2.1 i kommissionens förslag): En gruppering kan bestå av medlemsstater, regionala och lokala instanser eller andra lokala offentliga organ, nedan kallade ”medlemmar”.
Föredraganden anser att det europeiska territoriella samarbetet till sin natur gör att detta instrument underlättar samarbete mellan regionala och/eller lokala myndigheter utan inblandning från medlemsstaterna ( ändringsförslag 10 och 17) .
Ø Föredraganden skulle vilja betona att inrättandet av en gruppering innebär att de offentliga myndigheterna i den medlemsstat vars lagstiftning är tillämplig har kontrollen över detta instrument inom ramen för såväl medlemsstaternas som gemenskapens ekonomiska insatser (ändringsförslag 16).
Ø Grupperingarna får den rättskapacitet som juridiska personer har i nationell lagstiftning, på grundval av den typ av verksamhet som de bedriver och de uppgifter som delegerats till dem.
Grupperingarnas rättskapacitet är den som juridiska personer har i nationell lagstiftning (artikel 3.2 i kommissionens förslag) .
Föredraganden insisterar på att grupperingarna begränsar sig till att utföra specificerade uppgifter .
En gruppering agerar inom ramen för de uppgifter som delegerats till den och som kan tilldelas en av dess medlemmar.
En gruppering bör fungera som en juridisk enhet (oavsett om den är juridisk person eller inte) på grundval av bindande nationella rättsakter såsom associationsrätt (ändringsförslag 19, 21 och 31) .
Ø Bildande av en gruppering: I kommissionens förslag erbjuds två möjligheter (artikel 2.3 i kommissionens förslag):
- Medlemmarna i grupperingen skapar en särskild enhet av den typ de behöver och i detta fall utför grupperingen själv uppgifterna inom ramen för det gränsöverskridande samarbetet.
- Medlemmarna bildar en gruppering och grupperingen fattar beslut enligt sina egna beslutsregler att delegera grupperingens uppgifter till en regional och/eller lokal myndighet som är medlem i grupperingen, om man föredrar detta.
Denna myndighet skall utföra de uppgifter som delegerats till grupperingen.
Föredraganden anser att medlemmarna inte ”kan besluta att bilda en gruppering” på ett av dessa sätt utan de ”bildar” denna (ändringsförslag 18) .
Ø Grupperingens uppgifter och befogenheter bör fastställas av dess medlemmar i ett avtal om europeiskt gränsöverskridande samarbete (artikel 4 i kommissionens förslag).
Föredraganden anser att för en gruppering skall ett avtal om europeiskt territoriellt samarbete ingås av dess medlemmar (ändringsförslag 25).
Ø I avtalet fastställs:
- grupperingens uppgifter, varaktighet och upplösning (punkt 2)
- varje medlems ansvar gentemot grupperingen och gentemot tredje part (punkt 4).
- vilken lagstiftning som gäller för grupperingen och dess tillämpning (punkt 5).
Den tillämpliga lagstiftningen skall vara en av de berörda medlemsstaternas lagstiftning, endera på grundval av landets deltagande i grupperingen, eller på grundval av deltagande i en instans under statlig nivå eller i en offentlig organisation med säte på denna medlemsstats territorium.
Det kan röra sig om lagstiftningen i den medlemsstat där grupperingen har inrättat sitt säte.
- bestämmelser om ömsesidigt erkännande i fråga om kontroller (punkt 6)
- att avtalet skall skickas till samtliga medlemmar och till de deltagande medlemsstaterna (punkt 8).
Föredraganden anser att:
– punkt 2: Avtalet bör i synnerhet fastslå (icke uttömmande lista) regler för grupperingens funktion , grupperingens uppgifter , dess varaktighet och upplösning (ändringsförslag 26) .
– punkt 4: Frågan om varje medlems ansvar utvecklas tillräckligt i artikel 7.2 om medlemsstaternas ansvar (ändringsförslag 28) .
– punkt 6: Bestämmelser om ömsesidigt erkännande bör specificeras i själva förordningen och inte i avtalets bestämmelser.
Föredraganden föreslår därför att det läggs till en ny punkt i artikel 1.3 (se ändringsförslag 16) (ändringsförslag 30) .
– Den lagstiftning som gäller för grupperingar bör vara associationsrätten i den berörda medlemsstaten (ändringsförslag 31) .
– punkt 8: Avtalet bör också skickas till Regionkommittén (ändringsförslag 33) .
Ø Grupperingen antar sina stadgar (artikel 5 i kommissionens förslag) och inrättar sina egna organ (artikel 6 i kommissionens förslag) .
Grupperingen skall alltid ha en direktör.
Däremot är frågan om att inrätta en församling som består av företrädare för medlemmarna eller andra organ något som överlåts till medlemmarna.
– Föredraganden anser att stadgarna också bör innehålla bestämmelser om hur grupperingen skall företrädas , inbegripet en församling som består av företrädare för dess medlemmar och en verkställande kommitté (ändringsförslag 34).
Här föreslås att artikel 6 om grupperingens organ stryks och att dessa tas med i artikeln om stadgarna (ändringsförslag 36) .
Ø Grupperingen skall publiceras i Europeiska unionens officiella tidning.
Från och med denna tidpunkt är grupperingens rättsliga status erkänd i alla medlemsstaterna ( artikel 7 i kommissionens förslag) .
Föredraganden anser att när grupperingen väl blivit en juridisk person enligt tillämplig nationell lagstiftning i den berörda medlemsstaten skall stadgarna med vilka en gruppering inrättas offentliggöras i Europeiska unionens officiella tidning ( ändringsförslag 37) .
ÄRENDETS GÅNG
Titel
Europeiska grupperingar för gränsöverskridande samarbete (EGGS)
Referensnummer
KOM(2004)0496 – C6‑0091/2004 – 2004/0168(COD)
Rättslig grund
art.
251.2, och.
Grund i arbetsordningen
Framläggande för parlamentet
15.7.2004
REGI
17.11.2004
BUDG 17.11.2004
CONT 17.11.2004
CONT 23.3.2005
BUDG 31.1.2005
-
Jan Olbrycht 6.10.2004
Tidigare föredragande
Förenklat förfarande Beslut
Ändrad anslagstilldelning BUDG:s yttrande
Samråd med Europeiska ekonomiska och sociala kommittén Beslut i kammaren
Behandling i utskott
7.10.2004
20.1.2005
21.4.2005
Antagande
16.6.2005
Slutomröstning: resultat
för:
emot:
nedlagda röster:
43
1
3
Slutomröstning: närvarande ledamöter
Alfonso Andria, Stavros Arnaoutakis, Jean Marie Beaupuy, Rolf Berend, Jana Bobošíková, Graham Booth, Bairbre de Brún, Giovanni Claudio Fava, Iratxe García Pérez, Eugenijus Gentvilas, Lidia Joanna Geringer de Oedenberg, Ambroise Guellec, Zita Gurmai, Konstantinos Hatzidakis, Mieczysław Edmund Janowski, Gisela Kallenbach, Miloš Koterec, Constanze Angela Krehl, Miroslav Mikolášik, Francesco Musotto, Lambert van Nistelrooij, Jan Olbrycht, István Pálfi, Markus Pieper, Francisca Pleguezuelos Aguilar, Bernard Poignant, Elisabeth Schroedter, Alyn Smith, Grażyna Staniszewska, Catherine Stihler, Kyriacos Triantaphyllides, Vladimír Železný
Slutomröstning: närvarande suppleanter
Alfredo Antoniozzi, Inés Ayala Sender, Jan Březina, Simon Busuttil, Den Dover, Mojca Drčar Murko, Richard Falbr, Věra Flasarová, Louis Grech, Ewa Hedkvist Petersen, Mirosław Mariusz Piotrowski, Richard Seeber, Thomas Ulmer
Slutomröstning: närvarande suppleanter (art.
178.2)
Sharon Margaret Bowles, Albert Deß
Ingivande – A6-nummer
21.6.2005
A6-0206/2005
Anmärkningar
...
SLUTLIG VERSION
A6-0261/2005
***I
BETÄNKANDE
om förslaget till Europaparlamentets och rådets rekommendation om ytterligare europeiskt samarbete om kvalitetssäkring i den högre utbildningen
(KOM(2004)0642 – C6‑0142/2004 – 2004/0239(COD))
Utskottet för kultur och utbildning
Föredragande:
Ljudmila Novak
PE 359.988v03-00
Teckenförklaring
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................12
ÄRENDETS GÅNG..................................................................................................................16
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till Europaparlamentets och rådets rekommendation om ytterligare europeiskt samarbete om kvalitetssäkring i den högre utbildningen
( KOM(2004)0642 – C6‑0142/2004 – 2004/0239(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2004)0642 )
EUT C ... / Ännu ej offentliggjort i EUT. ,
– med beaktande av artikel 51 i arbetsordningen,
– med beaktande av betänkandet från utskottet för kultur och utbildning ( A6‑0261/2005 ).
Kommissionens förslag
Parlamentets ändringar
Ändringsförslag
1
Skäl 1
(1) Rådets rekommendation av den 24 september 1998 om europeiskt samarbete om kvalitetssäkring i den högre utbildningen har genomförts framgångsrikt, vilket framgår av kommissionens rapport av den 30 september 2004.
Men den högre utbildningen i Europa behöver förbättras ytterligare och bli mer öppen för insyn och tillförlitlig för medborgarna och för studenter och forskare från andra delar av världen.
Motivering
Det europeiska samarbetet om kvalitetssäkring i den högre utbildningen måste i första hand bidra till att den högre utbildningens kvalitetsnivå höjs i medlemsstaterna.
Detta bör uttryckligen påpekas redan i det första skälet.
Ändringsförslag
2
Skäl 3
(3) I rådets rekommendation framhölls det att kvalitetssäkringssystemen bör bygga på ett antal viktiga komponenter, däribland utvärdering av program och högskolor genom interna och externa bedömningar där studenterna medverkar, offentliggörande av resultat och internationellt deltagande.
(3) I rådets rekommendation framhölls det att kvalitetssäkringssystemen bör bygga på ett antal viktiga komponenter, däribland utvärdering av program och högskolor genom interna och externa bedömningar där studenterna medverkar, offentliggörande av resultat och internationellt deltagande.
Dessa resultat bör systematiskt bearbetas och användas som grund för nästa bedömningsomgång.
Motivering
Resultaten av den interna och externa kvalitetssäkringen måste utgöra grunden för en kontinuerlig förbättring av högskolorna.
De skall tjäna som utgångspunkt för en systematisk utveckling av kvalitetstänkandet och anpassningen till samhällets föränderliga behov.
Ändringsförslag
3
Skäl 6
(6) Vid sitt möte i Berlin i september 2003 uppmanade utbildningsministrarna ENQA att genom sina medlemmar samarbeta med den europeiska rektorsorganisationen EUA, högskolesammanslutningen EURASHE och studentorganisationen ESIB för att utarbeta gemensamma standarder , förfaranden och riktlinjer, undersöka hur man kan utarbeta ett adekvat system för kollegiegranskning av kvalitetssäkrings- och ackrediteringsorgan samt genom uppföljningsgruppen rapportera för ministrarna 2005.
(6) Vid sitt möte i Berlin i september 2003 uppmanade utbildningsministrarna ENQA att genom sina medlemmar samarbeta med den europeiska rektorsorganisationen EUA, högskolesammanslutningen EURASHE och studentorganisationen ESIB för att utarbeta gemensamma standarder och riktlinjer, undersöka hur man kan utarbeta ett adekvat system för kollegiegranskning av kvalitetssäkrings- och ackrediteringsorgan samt genom uppföljningsgruppen rapportera för ministrarna 2005.
Inom ramen för Bolognaprocessen antog utbildningsministrarna från 45 länder vid sitt möte i Bergen den 20 maj 2005 de standarder och riktlinjer för kvalitetssäkring i det europeiska området för högre utbildning som hade förslagits av ENQA.
De välkomnade även principen om ett europeiskt register över kvalitetssäkringsorgan grundat på nationell översyn och uppmanade ENQA att i samarbete med EUA, EURASHE och ESIB ytterligare utveckla genomförandemetoderna.
Vidare underströk ministrarna vikten av samarbete mellan nationellt erkända organ i syfte att förbättra det ömsesidiga erkännandet av beslut om ackreditering eller kvalitetssäkring.
Ändringsförslag
4
Skäl 7
(7) Man bör upprätta en förteckning eller ett register över oberoende och tillförlitliga organ för kvalitetssäkring i Europa, oavsett om de är regionala eller nationella, allmänna eller specialiserade, offentliga eller privata, vinstdrivande eller inte, för att främja öppenhet och insyn i den högre utbildningen och medverka till att examensbevis och utlandsstudier erkänns.
(7) Man bör upprätta en förteckning eller ett register över oberoende och tillförlitliga organ för kvalitetssäkring i Europa, oavsett om de är regionala eller nationella, allmänna eller specialiserade, offentliga eller privata, för att främja öppenhet och insyn i den högre utbildningen och medverka till att examensbevis och utlandsstudier erkänns.
Motivering
(Berör inte den svenska versionen.)
Ändringsförslag
5
Avsnitt I, led a
A. att ålägga alla högskolor i det egna landet att införa eller utarbeta strikta mekanismer för intern kvalitetssäkring,
A. att ålägga alla högskolor i det egna landet att införa eller utarbeta strikta mekanismer för intern kvalitetssäkring, i överensstämmelse med de standarder och riktlinjer för kvalitetssäkring i det europeiska området för högre utbildning som antogs i Bergen inom ramen för Bolognaprocessen,
Ändringsförslag
6
Avsnitt I, led b
B. att ålägga alla kvalitetssäkrings- eller ackrediteringsorgan i det egna landet att göra oberoende bedömningar, tillämpa de komponenter i kvalitetssäkringen som fastställs i rådets rekommendation från september 1998 och tillämpa gemensamma standarder , förfaranden och riktlinjer vid bedömningen,
B. att ålägga alla kvalitetssäkrings- eller ackrediteringsorgan i det egna landet att göra oberoende bedömningar, tillämpa de komponenter i kvalitetssäkringen som fastställs i rådets rekommendation från september 1998 och tillämpa de allmänna gemensamma standarder och riktlinjer vid bedömningen som antogs i Bergen.
Ändringsförslag
7
Avsnitt I, led c
C. att uppmana kvalitetssäkrings- och ackrediteringsorgan att tillsammans med organisationer som företräder den högre utbildningen upprätta ett europeiskt register över kvalitetssäkrings- och ackrediteringsorgan enligt bilagan och att fastställa villkoren för att införas i registret,
C. att uppmana företrädare för kvalitetssäkrings- och ackrediteringsorgan , sektorn för högre utbildning och nationella myndigheter att upprätta ett europeiskt register över kvalitetssäkrings- och ackrediteringsorgan , grundat på en nationell bedömning, enligt bilagan och att fastställa villkoren för att införas i registret samt reglerna för att upprätthålla registret ,
Ändringsförslag
8
Avsnitt I, led d
D. att underlätta för högskolor i det egna landet att välja det organ som bäst svarar mot deras behov och profil, när de väljer bland kvalitetssäkrings- och ackrediteringsorgan i det europeiska registret,
Ändringsförslag
9
Avsnitt I, led e
E. att godta bedömningar som gjorts av kvalitetssäkrings- och ackrediteringsorgan i det europeiska registret som underlag för beslut om examensrätt för eller finansiering av högskolor, även när det gäller de studerandes rätt till studiebidrag eller studielån.
utgår
Motivering
Syftet med ändringsförslaget är att göra texten mer samstämmig.
Den åtskillnad som görs mellan examensrätt och kompletterande bedömning/ackreditering i led d och e i deras nya lydelse medför att den ursprungliga texten blir överflödig.
Ändringsförslag
10
Avsnitt I, led ea (nytt)
Ea. att främja att högskolorna eftersträvar en kompletterande transnationell bedömning eller ackreditering som gjorts av ett organ i det europeiska registret för att stärka högskolans internationella rykte,
Motivering
Det bör uttryckligen betonas att högskolorna skall sträva efter en ytterligare ackreditering eller bedömning som görs av ett internationellt organ i det europeiska registret, och att medlemsstaterna skall främja detta.
Ändringsförslag
11
Avsnitt I, led eb (nytt)
Eb. att främja samarbetet mellan organen med målet att bygga upp ömsesidigt förtroende och erkännande mellan dessa och på detta sätt underlätta erkännandet av deras examensbevis när det gäller studier och arbete i ett annat land, inbegripet studier som leder fram till ett reglerat yrke,
Ändringsförslag
12
Avsnitt I, led ec (nytt)
Ec. att främja offentliggörande av och garantera allmän tillgång till de bedömningar som kvalitetssäkrings- eller ackrediteringsorganen i det europeiska registret utfört.
Motivering
Att offentliggöra resultaten av kvalitetssäkrings- eller ackrediteringsorganens bedömningar skulle bidra till bättre information och större öppenhet för högskolorna.
Ändringsförslag
13
Bilaga, punkt 1
1.
Förteckningen bör upprättas av företrädare för kvalitetssäkrings- och ackrediteringsorgan i medlemsstaterna, i samarbete med företrädare för den högre utbildningen (universitet och övriga högskolor, studerande, högskolelärare och forskare) och arbetsmarknadens parter.
1.
Förteckningen bör upprättas av företrädare för nationella myndigheter och kvalitetssäkrings- och ackrediteringsorgan i medlemsstaterna, i samarbete med företrädare för den högre utbildningen (universitet och övriga högskolor, studerande, högskolelärare och forskare) och arbetsmarknadens parter.
Ändringsförslag
14
Bilaga, punkt 2, strecksats 3
- Organet ska agera i enlighet med de gemensamma standarder , förfaranden och riktlinjer som avses i punkt 6 i denna rekommendation.
- Organet ska agera i enlighet med de gemensamma standarder och riktlinjer som avses i led B i denna rekommendation.
Ändringsförslag
15
Bilaga, punkt 2a (ny)
2a.
Om registreringen först inte skulle godkännas är det möjligt att göra en ny bedömning på grundval av förbättringar som gjorts.
Motivering
Det är viktigt att fastställa ett förfarande enligt vilket organen på nytt kan begära att ett införande i registret prövas om en registrering först har avslagits, efter det att nödvändiga förbättringar har gjorts.
MOTIVERING
KOMMISSIONENS FÖRSLAG
Den rekommendation som skall behandlas här bygger på den rekommendation som antogs 1998 om europeiskt samarbete om kvalitetssäkring i den högre utbildningen
Rådets rekommendation av den 24 september 1998 om europeiskt samarbete om kvalitetssäkring i den högre utbildningen (98/561/EG), EGT L 270, 7.10.1998, s.
56. .
Syftet med båda rekommendationerna är att främja det ömsesidiga erkännandet av kvalitetssäkringssystemen och kvalitetsbedömningarna i Europa.
Vid mötet i Bergen den 19–20 maj 2005 diskuterade de ansvariga ministrarna för högre utbildning från 45 europeiska länder de framsteg som gjorts i Bolognaprocessen och kom överens om riktlinjerna för den fortsatta utvecklingen i det europeiska området för högre utbildning, även med avseende på kvalitetssäkringssystemen.
Det konstaterades att flera länder redan har gjort anmärkningsvärda framsteg när det gäller inrättandet av kvalitetssäkringssystem och främjandet av samarbetet.
Trots detta måste ytterligare steg tas, i synnerhet måste högskolorna fortsätta sina ansträngningar att uppnå högre kvalitet genom att systematiskt införa interna mekanismer som har direkt samband med extern kvalitetssäkring.
I detta sammanhang föreslår kommissionen att rådet och parlamentet skall anta en ny rekommendation som definierar fem steg på vägen mot ett ömsesidigt erkännande av kvalitetssäkringssystemen och kvalitetsbedömningarna:
Syftet är att uppnå ytterligare framsteg i utvecklingen och konsolideringen av mekanismerna för intern kvalitetssäkring vid högskolorna i Europa.
Den interna kvalitetsstyrningen skall samtidigt tjäna som underlag för den externa bedömningen av de europeiska högskolorna i syfte att optimera högskolornas jämförbarhet, insyn och resultat.
Genom att utveckla och tillämpa ett gemensamt system med uppsättningar av standarder, förfaranden och riktlinjer för kvalitetssäkring skall enhetliga regler skapas som framhäver likheter och skillnader mellan studieprogram utan att dessa harmoniseras.
Syftet är att upprätta ett europeiskt register över tillförlitliga kvalitetssäkringsorgan.
D. Högskolornas fria val av organ
Högskolorna skall vara fria att välja det kvalitetssäkringsorgan som passar dem bäst, förutsatt att organet i fråga finns med i registret och erkänns som oberoende och tillförlitligt i det egna landet.
Kommissionen föreslår dessutom att medlemsstaterna i samband med beslut om examensrätt och finansiering av högskolor skall godta beslut som fattats av organ i det europeiska registret.
ANMÄRKNINGAR OCH ÄNDRINGSFÖRSLAG FRÅN FÖREDRAGANDEN
Föredraganden ställer sig bakom föreliggande förslag från kommissionen som på ett positivt sätt bidrar till det ömsesidiga erkännandet av kvalitetssäkringssystemen och kvalitetsbedömningarna i Europa.
Föredraganden välkomnar särskilt att det föreslås konkreta åtgärder för att få den högre utbildningen i Europa att ge bättre resultat och bli mer öppen för insyn och attraktivare för studenter och forskare.
Det är dessutom positivt att en hög kvalitetsnivå hos utbildningsorganen kräver större rörlighet bland studenter och arbetstagare, vilket är viktigt i Lissabonstrategin.
En annan positiv aspekt är att en systematisk användning av det gemensamma kvalitetssäkringssystemet som instrument för en kontinuerlig förbättring av högskolornas kvalitet är en viktig förutsättning för det önskvärda ömsesidiga erkännandet av examensbevis och högskoleexamina i Europa.
Endast en sådan systematisk användning av mekanismer för kvalitetssäkring kan garantera en akademisk utbildning av hög kvalitet i EU, inom vars ramar undervisningen vid högskolorna främjas och jämförbarheten mellan de nationella utbildningssystemen underlättas.
Föredraganden betonar att det är nödvändigt att de interna och externa bedömningsresultaten av program eller högskolor kontinuerligt används som grund för nästa bedömningsomgång.
B. Gemensamma standarder, förfaranden och riktlinjer
Föredraganden välkomnar utarbetandet av de gemensamma standarder, förfaranden och riktlinjer för kvalitetssäkring i enlighet med mandatet från Berlin (september 2003), inom vars ramar de europeiska utbildningsministrarna uppmanade det europeiska nätverket för kvalitetssäkring i den högre utbildningen (ENQA) att utarbeta sådana gemensamma standarder, förfaranden och riktlinjer och undersöka hur man kan utarbeta ett adekvat system för kollegiegranskning av kvalitetssäkrings- och/eller ackrediteringsorgan.
Föredraganden betonar härvid att dessa standarder, förfaranden och riktlinjer för bedömning och ackreditering av högskolorna och organen kommer att främja mångfald på högskoleområdet och ge stöd till högskolornas anpassning till det moderna samhällets krav.
Kvalitetssäkringssystem får emellertid inte påtvingas.
I stället måste de frivilligt antas av alla berörda parter.
Det är därför önskvärt att det gemensamma systemet utvecklas av både organen och företrädare för högskolorna så att en gemensam identifikation med standarderna i högskolevärlden kan uppkomma.
Föredraganden välkomnar inrättandet av registret som bidrar till att utvärderings- och ackrediteringssystem och bedömningar blir vedertagna i hela Europa, vilket i sin tur kan underlätta det ömsesidiga erkännandet av examensbevis i och utanför Europa.
Mekanismerna för förvaltningen av registret och villkoren för att tas med i registret måste utvecklas ytterligare och preciseras.
De skall garantera en kontinuerlig bedömning av organen och säkra deras kvalitet, för att ett ömsesidigt godkännande och hög standard när det gäller oberoendet och yrkesmässigheten skall kunna säkerställas.
I enlighet med principen att alla berörda parter skall involveras skall den praktiska genomföranderamen även fortsättningsvis utvecklas genom ENQA i samarbete med EUA, EURASHE och ESIB.
Föredraganden betonar också betydelsen av samarbetet mellan de nationellt erkända organen som är en grundläggande förutsättning när det gäller att öka det ömsesidiga erkännandet av ackreditering och kvalitetssäkringsbeslut.
Föredraganden betonar dessutom att det är viktigt att fastställa ett förfarande i enlighet med vilket organen kan granskas på nytt om en begäran om registrering har avslagits, efter det att nödvändiga förbättringar har gjorts.
Det är viktigt att skilja mellan två olika processer: examensrätten (punkt D) och bedömningen/ackrediteringen (se punkt E).
Examensrätt betyder rätten att utfärda examina.
Vanligtvis utfärdas examen på grundval av minimistandarder och skall även i fortsättningen skötas av medlemsstaterna i den mån som medlemsstaterna står för finansieringen.
Bedömnings- och ackrediteringsförfarandena införs för att stärka allmänhetens insyn och förtroendet för högskolorna.
Den internationella ackrediteringen/bedömningen skall därför inte ersätta de nationella processerna, utan i stället utgöra ett komplement.
Respektive nationellt ministerium skall i enlighet med subsidiaritetsprincipen i princip fungera som behörig instans när det gäller högskoleutbildningens examensrätt.
Föredraganden föredrar därför en lydelse som ger medlemsstaterna utrymme att besluta i vilken utsträckning de vill lämna dörren öppen för organ från andra europeiska länder.
Medlemsstaterna skall härvid ge de högskolor som är verksamma i det egna landet möjlighet att välja ett nationellt organ eller ett utländskt organ i det europeiska registret, i den mån detta är tillåtet i det egna landet genom bestämmelser eller en överenskommelse med det behöriga ministeriet.
Det görs en åtskillnad mellan examensrätt och kompletterande bedömning/ackreditering (se punkt D).
När det gäller den andra kategorin betonar föredraganden att en sådan kompletterande ackreditering eller bedömning genom ett internationellt organ som finns i det europeiska registret skall eftersträvas av högskolorna och främjas av medlemsstaterna.
Det europeiska mervärdet av kvalitetssäkring/ackreditering uppkommer endast på grund av ett närmare samarbete mellan medlemsstaterna och deras organ.
Föredraganden ställer sig därför bakom samarbetet om kvalitetssäkring och ackreditering, som är ett viktigt steg på vägen mot ömsesidigt erkännande av utbildningsexamina.
Föredraganden betonar samtidigt att det är nödvändigt att koppla ihop de nationella kvalitetssäkrings- och ackrediteringssystemen med motsvarande europeiska ackrediteringsmekanismer.
Målet med det ömsesidiga erkännandet av kvalitetssäkringssystem samt kvalitets- och ackrediteringsbedömningar kan endast uppnås på lång sikt om det skapas ett förtroende mellan de behöriga organen.
Samarbetsmålen för EU:s medlemsstater skall fastställas på ett lika tydligt och ambitiöst sätt som i Bolognaprocessen, inte minst när det gäller dubbla utbildningsbevis och tillgången till den europeiska arbetsmarknaden.
ÄRENDETS GÅNG
Titel
Förslag till Europaparlamentets och rådets rekommendation om ytterligare europeiskt samarbete om kvalitetssäkring i den högre utbildningen
Referensnummer
( KOM(2004)0642 – C6-0142/2004 – 2004/0239(COD)
art.
Grund i arbetsordningen
art.
51
Framläggande för parlamentet
12.10.2004
Ansvarigt utskott Tillkännagivande i kammaren
CULT 26.01.2004
Rådgivande utskott Tillkännagivande i kammaren
Inget yttrande avges Utnämning
Förstärkt samarbete Tillkännagivande i kammaren
Föredragande Utnämning
Ljudmila Novak
25.11.2004
Tidigare föredragande
Behandling utskott
31.1.2005
11.7.2005
30.8.2005
Antagande
30.8.2005
Slutomröstning: resultat
för:
emot:
nedlagda röster:
24
1
1
Slutomröstning: närvarande ledamöter
María Badía i Cutchet, Giovanni Berlinguer, Guy Bono, Marie-Hélène Descamps, Milan Gaľa, Claire Gibault, Vasco Graça Moura, Lissy Gröner, Erna Hennicot-Schoepges, , Luis Herrero-Tejedor, Ruth Hieronymi, Manolis Mavrommatis, Ljudmila Novak, Doris Pack, Zdzisław Zbigniew Podkański, Christa Prets, Karin Resetarits, Nikolaos Sifunakis, Hannu Takkula, Helga Trüpel, Thomas Wise, Tomáš Zatloukal
Slutomröstning: närvarande suppleanter
Adamos Adamou, András Gyürk, Gyula Hegyi, Jaroslav Zvěřina,
Slutomröstning: närvarande suppleanter (art.
178.2)
Ingivande – A6-nummer
1.9.2005
A6-0261/2005
SLUTLIG VERSION
A6-0031/2006
om omstruktureringar och sysselsättning
(2005/2188(INI))
Utskottet för sysselsättning och sociala frågor
Föredragande:
Jean Louis Cottigny
PE 362.704v03-00
INNEHÅLL
MOTIVERING..........................................................................................................................12
ÄRENDETS GÅNG..................................................................................................................15
EUROPAPARLAMENTETS FÖRSLAG TILL RESOLUTION
om omstruktureringar och sysselsättning
( 2005/2188(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens meddelande av den 31 mars 2005 med titeln ”Omstruktureringar och sysselsättning – Att förutse omstruktureringar och ge stöd i samband med dem i syfte att utveckla sysselsättningen: Europeiska unionens roll” ( KOM(2005)0120 ) och yttrandet från EESK av den 14 december 2005 (CESE 1495/2005),
– med beaktande av stadgan om arbetstagares grundläggande sociala rättigheter från 1989 och tillhörande åtgärdsprogram,
EGT L 254, 30.9.1994, s.
EGT L 225, 12.8.1998, s.
16. ,
– med beaktande av rådets direktiv 2001/23/EG av den 12 mars 2001 om tillnärmning av medlemsstaternas lagstiftning om skydd för arbetstagares rättigheter vid överlåtelse av företag, verksamheter eller delar av företag eller verksamheter
EGT L 82, 22.3.2001, s.
16. ,
– med beaktande av Europaparlamentets och rådets direktiv 2002/14/EG av den 11 mars 2002 om inrättande av en allmän ram för information till och samråd med arbetstagare i Europeiska gemenskapen
EGT L 80, 23.3.2002, s.
29. ,
– med beaktande av sina resolutioner av den 28 oktober 1999
EGT C 154, 5.6.2000, s.
139. , den 17 februari 2000
EGT C 339, 29.11.2000, s.
280. och den 15 februari 2001
EGT C 276, 1.10.2001, s.
160. om omstruktureringar av europeiska företag,
– med beaktande av rådets rekommendation 92/443/EEG av den 27 juli 1992 om främjande inom medlemsstaterna av arbetstagares möjlighet att ta del av företagsvinster och resultat (inklusive andelsägande genom aktieförvärv)
EGT L 245, 26.8.1992, s.
53. ,
EGT C 377, 29.12.2000, s.
164. ,
P6_TA(2005)0127 . ,
– med beaktande av kommissionens meddelande om den socialpolitiska agendan ( KOM(2005)0033 ) och sin resolution av den 26 maj 2005
P6_TA(2005)0230 . om den socialpolitiska agendan 2006–2010
P6_TA(2005)0210 . ,
– med beaktande av kommissionens meddelande till rådet och Europaparlamentet med titeln ”Gemensamma insatser för tillväxt och sysselsättning: gemenskapens Lissabonprogram” ( KOM(2005)0330 ),
– med beaktande av kommissionens initiativ att utnämna år 2006 till året för arbetstagarnas rörlighet samt genomförandet av Lissabonstrategin
MEMO/05/229. ,
P6_TA(2005)0224 . om politiska utmaningar och budgetmedel i ett utvidgat EU 2007–2013 ,
– med beaktande av Europeiska rådets gemensamma ståndpunkt den 15 och 16 december 2005 i Bryssel om budgetplanen 2007–2013,
– med beaktande av förslaget till rådets förordning om allmänna bestämmelser för Europeiska regionala utvecklingsfonden, Europeiska socialfonden och Sammanhållningsfonden ( KOM(2004)0492 ),
– med beaktande av förslaget till Europaparlamentets och rådets förordning om Europeiska socialfonden ( KOM(2004)0493 ),
– med beaktande av artikel 45 i arbetsordningen,
– med beaktande av betänkandet från utskottet för sysselsättning och sociala frågor ( A6‑0031/2006 ), och av följande skäl:
A. Den ekonomiska och sociala strategin med avseende på riskerna är den huvudsakliga beståndsdelen i den europeiska sociala modellen, och den finns även med i de olika nationella politiska strategier som syftar till att bygga ett välfärdssamhälle grundat på solidaritet och social trygghet.
B. Om dessa risker inte förutses kan de drabba och skada arbetstagarna, för vilka arbetet är en av de faktorer som är avgörande för frihet och värdighet, och även arbetsgivarna och deras produktionsmedel, som utvecklas i den konkurrenssituation som råder i en öppen ekonomi.
J. Arbetsmarknadens parter och de offentliga myndigheterna bör spela en avgörande roll i samband med omstruktureringar, både på övergripande nivå genom att skapa nya arbetstillfällen och på individuell nivå genom att ge de berörda arbetstagarna möjlighet att anpassa sig till en ny verksamhet, särskilt genom utbildningsåtgärder, men också i ett förberedande skede och i sökandet efter alternativa lösningar när detta är möjligt.
M. Europaparlamentet anser att företagen som ett sätt att ta ansvar för lämpliga förebyggande insatser bör garantera bästa möjliga villkor för fortbildning av sina anställda
– vid praktikperioder under grundutbildning och lärlingskap,
– vid erkännandet och godkännandet av yrkeserfarenhet.
O. En av orsakerna till svårigheterna för de europeiska företagen är att det inte finns tillräckliga regler på internationell nivå för att skydda immateriella rättigheter och effektivt bekämpa förfalskning.
Parlamentet anser att dessa förutsättningar inte alltid finns.
Kommissionen bör utnyttja möjligheten till medling av ett oberoende organ på europeisk nivå vid fall av omoraliska åtgärder som vidtas enbart i vinstsyfte.
4.
Europaparlamentet anser att unionen är skyldig att möta de globala utmaningarna såsom omstruktureringar genom att förbättra den europeiska ekonomins och företagens konkurrenskraft och åstadkomma bättre samordning och större samstämmighet i användningen av gemenskapens fyra befintliga styrinstrument, nämligen
– konkurrenspolitiken, särskilt frågan om statligt stöd,
– politiken för den inre marknaden, särskilt inrättandet av Societas Europea och gemenskapspatentet,
– företagspolitiken, särskilt stödet till små och medelstora företag,
– solidaritetspolitiken, särskilt genom omfördelning av medel från Europeiska regionala utvecklingsfonden och Europeiska socialfonden till regioner som drabbats av omstruktureringar eller genom planer för förberedande åtgärder.
b) Europaparlamentet begär att det beaktas om ett företag i sin företagsplan inkluderar anpassningsåtgärder, särskilt om det engagerar sig i yrkesutbildning och vidareutbildning.
Europaparlamentet föreslår att miljödimensionen bör beaktas i samband med att EU ger stöd vid omstruktureringar, bland annat genom att främja industriell omställning eller omställning av jordbruk till metoder som är mindre förorenande och därmed mindre farliga för befolkningen i området och arbetstagarna.
Bland omstruktureringarnas dolda effekter fördömer Europaparlamentet också åtgärden att förtidspensionera arbetstagare som på grund av sin ålder tillhör de minst anställningsbara, eftersom detta medför stora kostnader för samhället och leder till att deras yrkeskompetens går förlorad samt till en absurd risk för brist på arbetskraft.
Europaparlamentet bekräftar den viktiga roll som gemenskapens regelverk har på det sociala området och särskilt betydelsen av de befintliga rättsliga instrumenten, som bör tillämpas till fullo och kontrolleras bättre av medlemsstaterna, som har ansvar för att bestämmelserna införlivas i lagstiftningen och tillämpas.
Detta gäller framför allt :
– rådets direktiv 94/45/EG av den 22 september 1994 om inrättandet av ett europeiskt företagsråd,
– rådets direktiv 98/59/EG av den 20 juli 1998 om kollektiva uppsägningar,
– rådets direktiv 2001/23/EG av den 12 mars 2001 om tillnärmning av medlemsstaternas lagstiftning om skydd för arbetstagares rättigheter vid överlåtelse av företag, verksamheter eller delar av företag eller verksamheter,
Europaparlamentet beklagar att den andra samrådsfasen om det europeiska företagsrådet endast är ett litet avsnitt i ett större meddelande från kommissionen och uppmanar kommissionen att, om den har för avsikt att se över det gällande direktivet om det europeiska företagsrådet, se till att det blir en ordentlig andra samrådsfas där arbetsmarknadens parter ges möjlighet att förhandla i enlighet med artikel 138 i EG‑fördraget och där öppenhetsprincipen beaktas.
19.
Europaparlamentet delar kommissionens uppfattning att den europeiska arbetsmarknadens parter bör ha en central roll i samband med och i styrningen av omstruktureringar, för att gynna arbetstagarnas rörlighet i Europa och uppmuntra till fortbildning genom hela livet närhelst detta behövs.
20.
Europaparlamentet uppmanar kommissionen att fortsätta verka för en gemenskapsram för skyddet av arbetstagarnas rättigheter vid omstruktureringar.
Europaparlamentet stöder behovet av uppföljande analyser av genomförda omstruktureringar för att kunna få kunskap om deras konkreta inverkan på det aktuella företaget och därmed få bättre beredskap inför framtida omstruktureringar.
30 Europaparlamentet kräver att unionens handelspartner inför lagar om skydd av immateriella rättigheter och att medlemsstaterna gör allt vad som står i deras makt för att effektivt bekämpa förfalskning.
En första nivå på omstruktureringar gäller dem som sker mellan branscher: dessa omvandlingar av stora branscher, till exempel tillväxten inom tjänstesektorn, har i hög grad blivit synliga i länderna i Västeuropa och berör i dag de nya medlemsstaterna i Central‑ och Östeuropa.
En andra nivå på omstruktureringar gäller de omstruktureringar och den utveckling som sker inom branscher.
Den tredje nivån omfattar hela företag där olika typer av omstruktureringar kan ske, såsom ändrade tillverkningsprocesser, outsourcing av verksamhet, omflyttningar, stängning av anläggningar, personalnedskärningar, sammanslagningar/förvärv osv.
Generellt sett finns det två kategorier av utlösande faktorer bakom omstruktureringar: en allmän utlösande faktor som hör samman med den internationella handelsutvecklingen och den nuvarande globaliseringen samt en andra utlösande faktor som hör samman med företagets strategi.
Dessa två utlösande faktorer är inbördes sammanbundna.
Företagets strategi motsvarar i själva verket ofta behovet av anpassning till utvecklingen av marknaden och verksamheten.
Europeiska kommissionen behandlar i sitt meddelande av den 31 mars 2005, ”Omstruktureringar och sysselsättning – Att förutse omstruktureringar och ge stöd i samband med dem i syfte att utveckla sysselsättningen: Europeiska unionens roll” problemen och de negativa konsekvenserna av omstruktureringar, omflyttningar och sammanslagningar.
Konsekvenserna går ofta i motsatt riktning som Lissabonmålen, närmare bestämt de mål som gäller främjandet av full sysselsättning, arbetets kvalitet, social sammanhållning och hållbar utveckling.
Europeiska unionen har sedan länge utvecklat politiska åtgärder och instrument för omstruktureringar.
Tidigare har även unionen spelat en avgörande roll för omstruktureringen av stål‑ och varvsektorn, men den senaste krisen inom textilbranschen visade att de befintliga instrumenten inte längre var tillräckliga för att bemöta så omfattande omvälvningar.
Det åligger därför Europeiska unionen att stärka åtgärderna och utveckla resurser som kan mobiliseras vid kris, men också att se över införandet av nya verktyg som gör det lättare att förutse och därmed också hantera omstruktureringar.
Ur ett horisontellt perspektiv har för övrigt många av EU:s politiska åtgärder redan bidragit till målet att förutse och följa omstruktureringar: direktiven om information till och samråd med arbetstagare (även om man bör övervaka att de tillämpas korrekt), dialogen mellan arbetsmarknadens parter på EU‑nivå, sysselsättningspolitiken, ekonomiska stödinstrument, industri‑ och företagspolitiken, politiken för landsbygdsutvecklingen osv.
I detta hänseende är det viktigt att tänka sig ett sammanhang med delat ansvar mellan arbetsgivare, offentliga myndigheter, arbetsmarknadens parter och arbetstagare för att inleda en debatt om förberedelser, uppföljning och anpassning.
Förberedelserna, hanteringen och uppföljningen av omstruktureringsprocesser kräver aktiv medverkan av alla berörda parter och måste bygga på tydliga synergier mellan politiska, rättsliga, avtalsmässiga och finansiella instrument.
Åtgärderna bör vidtas på samtliga relevanta nivåer, däribland EU‑nivå.
Det är viktigt att genom kommissionens meddelande och detta betänkande föra upp frågan om omstruktureringar på EU:s agenda, liksom dess samband med sysselsättningen och övriga politiska åtgärder på området, dialogen mellan arbetsmarknadens parter i fråga om företagens sociala ansvar, oavsett om det gäller på EU‑nivå eller nationell nivå.
Det finns en konsekvens i att Europeiska unionen på det rättsliga planet tar på sig kostnaderna och följderna av den politik den driver och vi kan beklaga bristen på politisk vilja från medlemsstaternas sida att arbeta i denna riktning.
– Finansiella resurser måste finnas tillgängliga när debatten om budgetplanen har avslutats, både inom strukturfonderna och i genomförandet av en fond för anpassning till tillväxten.
Detta är det pris unionen måste betala för de öppna marknaderna.
Genom dessa åtgärder kan arbetstagarnas rättigheter stärkas och därmed bli mer verkningsfulla.
– De arbetstagare som först drabbas av omstruktureringar måste stå i centrum för all uppmärksamhet, vara de första som beviljas stöd, tas om hand och följs upp.
Anpassad fortbildning skall alltid kunna föreslås dem för att de skall kunna möta förändringar och få sysselsättning av hög kvalitet.
– Relevanta analysinstrument måste inrättas branschvis för att få bättre kunskap om fenomenet med omstruktureringar och därmed också kunna förutse dem och anpassa bemötandet av dem.
Den harmonisering som så småningom beräknas ske av medlemsstaternas system på skatteområdet och det sociala området kommer också att innebära en mer verkningsfull kamp mot de olika former av social dumpning inom gemenskapen som är en av orsakerna till omlokaliseringar och omstruktureringar.
Här finns några av de medel som gör att unionen på ett effektivt sätt kan ingripa för att omstruktureringar inte blir liktydigt med sociala bakslag och ekonomiska förluster.
Vi måste ständigt värna om att behålla den europeiska sociala modellen och vi måste ha modet att i varje beslut sträva mot det bästa.
ÄRENDETS GÅNG
Titel
Omstruktureringar och sysselsättning
Förfarandenummer
2005/2188(INI)
Grund i arbetsordningen
Ansvarigt utskott Tillstånd: tillkännagivande i kammaren
Rådgivande utskott Tillkännagivande i kammaren
Inget yttrande avges Beslut
Förstärkt samarbete Tillkännagivande i kammaren
nej
Resolutionsförslag som återges i betänkandet
Föredragande Utnämning
Tidigare föredragande
Behandling i utskott
5.10.2005
23.11.2005
25.1.2006
Antagande
26.1.2006
Slutomröstning: resultat
för:
emot:
nedlagda röster:
34
5
5
Slutomröstning: närvarande ledamöter
Jan Andersson, Roselyne Bachelot-Narquin, Jean-Luc Bennahmias, Emine Bozkurt, Iles Braghetto, Philip Bushill-Matthews, Milan Cabrnoch, Derek Roland Clark, Luigi Cocilovo, Jean Louis Cottigny, Harlem Désir, Harald Ettl, Richard Falbr, Carlo Fatuzzo, Joel Hasse Ferreira, Roger Helmer, Stephen Hughes, Karin Jöns, Jan Jerzy Kułakowski, Sepp Kusstatscher, Bernard Lehideux, Elizabeth Lynne, Thomas Mann, Ana Mato Adrover, Maria Matsouka, Ria Oomen-Ruijten, Csaba Őry, Marie Panayotopoulos-Cassiotou, Pier Antonio Panzeri, Jacek Protasiewicz, José Albino Silva Peneda, Kathy Sinnott, Jean Spautz, Gabriele Zimmer
Slutomröstning: närvarande suppleanter
Edit Bauer, Dieter-Lebrecht Koch, Lasse Lehtinen, Jamila Madeira, Marianne Mikko, Dimitrios Papadimoulis, Luca Romagnoli, Leopold Józef Rutowicz, Elisabeth Schroedter, Barbara Weiler, Tadeusz Zwiefka
Slutomröstning: närvarande suppleanter (art.
178.2)
Ingivande – A6-nummer
9.2.2006
A6‑0031/2006
SLUTLIG VERSION
A6-0141/2006
BETÄNKANDE
om kustfiske och problem för fiskare som idkar kustfiske
(2004/2264(INI))
Fiskeriutskottet
Föredragande:
Seán Ó Neachtain
PE 357.550v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
MOTIVERING
YTTRANDE från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
ÄRENDETS GÅNG
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om kustfiske och problem för fiskare som idkar kustfiske
( 2004/2264(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av den gemensamma fiskeripolitiken,
– med beaktande av bestämmelserna för Europeiska fiskerifonden,
– med beaktande av artikel 11 i rådets förordning (EG) nr 2792/1999 av den 17 december 1999 om föreskrifter och villkor för gemenskapens strukturstöd inom fiskerisektorn
1). ,
– med beaktande av sin resolution av den 5 april 2001 om fiskeri: säkerhet och olycksorsaker
EGT C 21 E, 24.1.2002, s.
359. ,
EGT L 358, 31.12.2002, s.
59. ,
EUT L 260, 6.8.2004, s.
1. ,
Antagna texter, P6_TA(2005)0532 . ,
– med beaktande av artikel 45 i arbetsordningen,
– med beaktande av betänkandet från fiskeriutskottet och yttrandet från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män ( A6‑0141/2006 ), och av följande skäl:
B. Den ekonomiska och sociala kris som har drabbat fiskerisektorn är särskilt kännbar för de mindre konkurrenskraftiga flottsegmenten, särskilt kustfisket.
C. För närvarande finns det en mängd olika åtgärder som rör olika aspekter av småskaligt fiske i flera olika gemenskapsförordningar.
D. Den gemensamma fiskeripolitiken och dess instrument, särskilt den framtida Europeiska fiskerifonden (EFF), måste ta hänsyn till kustfisket och anpassas till kustfiskets specifika problem, framför allt i samband med småskaligt och traditionellt fiske.
E. Det är viktigt att säkerställa kustfiskets framtid i Europeiska unionen med tanke på dess viktiga bidrag till sysselsättningen i kustområdena, samtidigt som det är nödvändigt att förhindra överkapacitet i detta flottsegment och den uttömning av resurser som detta leder till.
F. Trots att arbetslösheten är hög och kustfiskebefolkningen åldras finns det en allvarlig brist på rekrytering av unga människor i vissa kustområden.
G. Det finns ett stort beroende av fiske och därmed sammanhängande industrier i vissa kustområden, särskilt i öområden och i avlägsna kustområden.
H. I de mest avlägsna regionerna utgör gemenskapsstöden en garanti för konkurrenskraft och ekonomisk livskraft hos en stor del av beredningsindustrin.
I. Det finns en allvarlig brist på tillförlitlig statistik om kustfiskesektorn i många medlemsstater, vilket omöjliggör seriösa analyser och jämförelser.
J. Det behövs ett nytt gemenskapssynsätt som inriktas på harmonisering och undviker särbehandling av fiskare från olika medlemsstater, med tanke på de oförenliga nationella politiska åtgärderna för kustfiske.
K. Med tanke på den viktiga roll som branschorganisationer och lokala myndigheter kan spela för att utveckla sektorn på lokal nivå, bör projekt och verksamheter som dessa utvecklar till stöd för kustfisket, framför allt småskaligt och traditionellt fiske, uppmuntras och stödjas på gemenskapsnivå.
L. Det är viktigt för kustfiskarna att delta i handelsprocessen, förbättra mekanismerna för att marknadsföra sina produkter och främja en översyn av den gemensamma organisationen av marknaden för fiskeriprodukter för att garantera ett rättvisare försäljningspris vid första försäljningstillfället och främja en bättre spridning av mervärdet längs hela värdekedjan.
M. Det är oerhört viktigt att se till att kustfiskare och deras intresseorganisationer deltar i den gemensamma fiskeripolitikens beslutsprocess, skyddandet av havsmiljön och återhämtningen av fiskbestånden genom att främja tillämpningen av principen om samförvaltning och decentraliseringen av den gemensamma fiskeripolitiken.
N. Sektorn präglas av osäkra inkomster och löner, vilket beror på dess marknadspraxis och prissättningsmetoder vid första försäljningstillfället samt verksamhetens oregelbundna karaktär.
O. Att de rörliga kostnaderna ökar och bränslepriserna är mycket instabila påverkar också kustfiskesektorn.
P. Det finns tilltagande spänningar och konkurrens om resurserna mellan kustfiskare som fiskar för sitt uppehälle och fritidsfiskare, vilket är ett problem som måste lösas.
Q. Det är nödvändigt att se till att kustfiskets metoder även bidrar till bättre miljöskydd och till en hållbar utveckling av fiskesektorn.
Europaparlamentet betonar att kustfisket ger viktiga bidrag till de lokala ekonomierna och till att bibehålla den sociala strukturen i kustsamhällena med tanke på att dessa bidrar med fler arbetstillfällen per fångad fiskmängd än andra fiskeflottsegment, särskilt i öområden och avlägsna kustområden.
3.
Europaparlamentet föreslår att sådan fiskeutrustning inte tillåts som hotar kustbeståndens hållbarhet och livskraften hos de delar av samhället som är beroende av fiskerisektorn.
a) Småskaligt kustfiske.
b) Fartygens längd.
c) Det avstånd från hemmahamnen inom vilket fartyget bedriver sin verksamhet, med hänsyn till medlemsstaternas olika geografiska och maritima förhållanden.
d) En maximitid under vilken fartygen är borta från hemmahamnen.
Europaparlamentet uppmanar kommissionen att skyndsamt föreslå sätt att harmonisera data om kustfisket i Europeiska unionen, så att särdragen i enskilda nationella och regionala fisken skyddas.
Europaparlamentet anser att det är viktigt att kustfiskare och samhällen som är beroende av kustfisket blir mer direkt delaktiga i förädling och handel för att stärka deras vinstunderlag och höja deras levnadsstandard.
Europaparlamentet uppmanar kommissionen att erkänna kustfiskets och det traditionella fiskets särskilda karaktär inom den gemensamma fiskeripolitiken, och att avgöra i hur hög grad de befintliga instrumenten är lämpade för att reagera på sektorns behov, samt anpassa dem på lämpligt sätt.
19.
I det här sammanhanget kräver Europaparlamentet vidare att åtgärderna ges erforderlig publicitet för att se till att alla berörda parter med lätthet har tillgång till heltäckande information om utbildningsmöjligheter.
37.
MOTIVERING
1.
INLEDNING
Kustfisket har en avgörande betydelse för hela kustekonomiers socioekonomiska överlevnad.
De har en viktig potentiell roll inom gemenskapens fiskeripolitik – men så är inte fallet i dag.
De har inte minst en mycket betydelsefull funktion för ett hållbart utnyttjande av fiskeresurserna i gemenskapens kustvatten.
Det saknas en särskild rättslig ram för kustfiskesektorn.
Därför står denna viktiga sektor helt utanför dagens gemenskapslagstiftning om fiske.
Denna situation gör att förutsättningarna för kustfiskeindustrin blir ogynnsamma och måste åtgärdas omgående.
På begäran av föredraganden och fiskeriutskottet har Europaparlamentet beställt en studie om sektorn i fråga.
Denna studie, med titeln ”Kustfiske och problem för fiskare som idkar kustfiske” , sammanställdes av Centro Tecnológico del Mar – Fundación Cetmar.
Den lades fram för utskottet vid en offentlig utfrågning i Bryssel den 24 november 2005.
Vid denna medverkade också framstående specialister från ett antal medlemsstater med presentationer.
På grundval av slutsatserna i den ovannämnda studien, experternas presentationer, ovärderliga bidrag från ledamöterna och slutsatserna från diskussionerna skall föredraganden inrikta sig på den aktuella situationen för kustfisket i EU.
Jag skall försöka identifiera de inbyggda svagheterna i sektorn och föreslå några möjliga lösningar som skulle kunna stärka sektorn betydligt, och inte bara bidra till att lokala ekonomier utvecklas utan också till att bibehålla kustsamhällenas sociala struktur.
2.
DEFINITION AV KUSTFISKE
I Europeiska gemenskapens lagstiftning definieras småskaligt kustfiske som fiskeriverksamhet som bedrivs av fartyg som är högst 12 meter långa och inte använder trålar.
”I denna förordning skall med ’småskaligt kustfiske’ avses fiske som bedrivs av fartyg med en total längd på under tolv meter” som inte använder den trålutrustning som omtalas i Tabell 2 i Bilaga 1 till kommissionens förordning (EG) nr 2090/98 av den 30 september 1998 om gemenskapens register över fiskefartyg
Artikel 11 i rådets förordning (EG) nr 2792/1999 av den 17 december 1999 om föreskrifter och villkor för gemenskapens strukturstöd inom fiskerisektorn. .
I praktiken använder emellertid varje medlemsstat sin egen definition.
Ett stort antal termer används för närvarande för att definiera sektorn, däribland hantverksmässigt fiske, småskaligt fiske och kustfiske .
Alla dessa termer tolkas olika i medlemsstaterna.
Tolkningarna varierar på grund av den nationella lagstiftningen, kulturella traditioner, typen av fiske och de nationella fiskeflottornas struktur.
Det är bara två medlemsstater som har rättsliga definitioner.
Olika typer av båtar kan användas för kustfiske – från mycket små fartyg som bara fiskar nära kusten till större fartyg som kan fiska mycket längre ut till havs.
Vilka värden som åsätts varje parameter varierar från land till land, och till och med från region till region.
Dessutom är parametrarna ofta inte klart definierade.
Gemenskapen behöver en koordinerad strategi för kustfisket.
Eftersom den här industrin uppfattas såsom verkande i ett klart heterogent sammanhang i varje medlemsstat anser föredraganden att en harmonisering av konceptet och en definition av småskaligt kustfiske bara kan uppnås genom EU‑lagstiftning.
Föredraganden anser emellertid också att EU måste ha en realistisk linje genom att tillåta avvikande definitioner i medlemsstaterna.
Framtida regelverk måste innehålla bestämmelser som gör sådana nationella anpassningar möjliga.
Några kriterier som kan användas i en gemensam definition är
a) hantverksmässigt fiske,
b) fartyg som återvänder till hamnen varje dag,
c) fartyg som bedriver fiske mindre än 20 km från sin hemmahamn.
3.
LAGSTIFTNING SOM PÅVERKAR KUSTFISKET
· Tillämpning av gemenskapsrätten
En av de grundläggande underliggande svårigheterna med att reglera kustfisket är att det helt saknas integration mellan EG:s bestämmelser och den nationella lagstiftningen.
Nästan alla EG‑bestämmelser avser högsjöfiske.
Ironiskt nog hänvisas det ofta i EG:s regelverk till den besvärliga ekonomiska situationen i fiskesektorn och till att olika kustbefolkningar är beroende av fisket.
Det är ju just dessa kustsamhällen som är mest beroende av kustfisket, men detta avspeglas inte i EG‑rätten.
· Kustfisket och den gemensamma fiskeripolitiken
Eftersom det inte finns någonting konkret i den befintliga gemenskapslagstiftningen som direkt kopplar kustfisket till en given geografisk eller maritim plats är fiske av det här slaget helt enkelt dömt att samexistera med andra större och mer kraftfulla kommersiella fartyg.
En av de få källor som tillsammans med kommissionens förordning (EG) nr 2090/98 av den 30 september 1998 om gemenskapens register över fiskefartyg ger en antydan om att små kustfartyg kan arbeta i kustvattnen under medlemsstaternas överinseende är artikel 9 i förordning (EG) nr 2371/2002 om bevarande och hållbart utnyttjande av fiskeresurserna inom ramen för den gemensamma fiskeripolitiken :
”Medlemsstaters åtgärder inom tolvmilsgränsen
1.
En medlemsstat får vidta icke ‑diskriminerande åtgärder för bevarande och förvaltning av fiskeriresurserna och för att minimera fiskets inverkan på bevarandet av de marina ekosystemen inom en gräns på 12 sjömil från dess baslinjer, förutsatt att gemenskapen inte har antagit åtgärder för bevarande och förvaltning särskilt för detta område.
Medlemsstatens åtgärder skall vara förenliga med de mål som fastställs i artikel 2 och får inte vara mindre stränga än gällande gemenskapslagstiftning.”
· Andra aspekter av förordning (EG) nr 2371/2002
Enligt förordningen undantas fartyg som är under 15 meter långa från kravet att installera system för fjärrövervakning och identifiering.
Detta är en karaktäristisk egenskap hos kustfisket som skiljer det från industriellt fiske och högsjöfiske.
Denna aspekt specificeras emellertid inte i förordningen.
I artikel 31 om regionala rådgivande nämnder nämns inte kustfiskets specifika natur alls.
Den handlar bara om ”havsområden” och ”fiskezoner” samt vattenbruk, men inte om olika slags fiskeverksamhet.
· Förordning (EG) nr 1421/2004
I förordning (EG) nr 1421/2004
Rådets förordning (EG) nr 1421/2004 av den 19 juli 2004 om ändring av förordning (EG) nr 2792/1999 om föreskrifter och villkor för gemenskapens strukturstöd inom fiskerisektorn. står det att ”skydd och utveckling av akvatiska resurser gäller inte enbart åtgärder till havs” , men skyddet för kustresurser genom kustfiske nämns långt ifrån och det görs inte någon specifik hänvisning till kustfisket i det här sammanhanget i förordningen.
4.
ATT ADMINISTRERA KUSTFISKET
Under utfrågningen beskrev några talare kustfiskesektorn som ”en smältdegel med många små företag”.
Andra talare sade att bristen på sammanslutningar och kooperativ för kustfiskare ”skapar en fragmentarisk undersektor till fiskeindustrin”.
I en del områden finns det en ökande fiskeansträngning av enskilda aktörer.
I andra områden, där antalet aktörer minskar, försöker man gå samman till större och mer effektiva enheter.
Det finns också en ökande specialisering på enskilda arter, det vill säga att sektorn är mindre generellt inriktad än tidigare.
Det finns inte så många organ som specifikt styr kustfisket.
Sektorn är också frånvarande eller helt underrepresenterad när det fattas beslut om fiskeripolitiken i gemenskapen, på nationell och regional nivå.
Med tanke på restriktionerna för tillträdet innanför tolvmilsgränsen är det kustmedlemsstaterna som har hela ansvaret för att administrera kustfisket inom ramen för den gemensamma fiskeripolitiken.
Därför har alla länder och regioner försökt utveckla sina egna administrativa strukturer.
Trots detta lider kustsektorn fortfarande av det allvarliga problemet med underrepresentation i de flesta instanser.
Utvecklingen av kooperativa styrelseformer i en del medlemsstater på den senaste tiden har haft positiva effekter på sektorn, något som också framhölls vid utfrågningen, vilka har skapat ett passande forum för diskussioner om de trender och de frågor som berör sektorn.
Som en av de inbjudna talarna vid utfrågningen sade: ”Nu är det avgörande att vi går från motsättningar till konsensus och från isolationism till gemenskap, så att kustfiskarna kan gå framåt tillsammans med samma vision.
Samarbetet bör så långt möjligt basera sig på ett frivilligt partnerskap.
Att koppla samman lokala fiskare och de organisationer som företräder dem är en av de högst prioriterade framtidsfrågorna.
En effektiv administration av fisket kan ge ett hållbart och bärkraftigt fiske och maximera de ekonomiska och sociala vinsterna.”
5.
SOCIOEKONOMISKA ASPEKTER
Den utpräglat traditionella kustfiskesektorn där sysselsättningsstrukturen brukade bygga på det lokala samhället och familjeband genomgår oroande förändringar.
En konsekvens av att fiskesamhällena åldras är att det blir allt svårare att modernisera fisket och införa nya, bättre metoder.
Följden är att kustfisket i dag ter sig allt mindre lockande för unga människor.
Tyvärr är utbildningsnivån i fiskesamhällena låg både vad gäller teoretisk och praktisk utbildning.
Yrkesutbildningen i sektorn är informell och traditionell utan några särskilda kurser eller utbildningsprogram.
Bristen på lämpliga utbildningsprogram är ett allvarligt hinder för sektorns utveckling.
Den begränsar flödet av relevant information till myndigheter och administrativa organ allvarligt.
I de flesta fall begränsar den sektorns deltagande i utformningen av de styråtgärder som berör den.
Den hindrar fiskarna att använda och dra nytta av den senaste och bästa tekniken.
Under utfrågningen var alla överens om att utbildning är avgörande för om denna viktiga sektor skall få den utveckling den behöver.
· Levnadsstandarder och sociala förhållanden
Beroendet av kustfisket är stort i de kustområden där fiskesamhällena finns.
Tyvärr kännetecknas dock sektorn generellt sett av låga inkomster för både kaptener och besättningar.
I flertalet fall betyder det osäkra anställningsförhållanden och hårda arbetsvillkor.
Det betyder också höga risker för arbetstagarna och låg social status.
Sektorn kännetecknas också av deltidsarbete.
För att kunna försörja sina familjer och hjälpa till att bevara och underhålla sin fiskeverksamhet tvingas fiskarna ofta komplettera sina inkomster med olika deltidsarbeten.
Det är oerhört svårt för fiskarna i kustfiskesektorn att få lån och ekonomiskt stöd.
Finansinstituten betraktar kustfisket som en högrisksektor.
Ovanstående punkter är några exempel på faktorer som gör det svårt för sektorn att få tillgång till finansiering.
· Kvinnorna och kustfisket
Det är uppenbart att kvinnornas roll i det europeiska fisket präglas av sektorns starkt traditionella natur, och mycket av det de gör sker på frivillig basis.
Parlamentet har tidigare, i och med sitt krav på en EU‑resolution om kvinnliga nätverk
Europaparlamentets resolution A6‑0341/2005 av den 30 november 2005 om kvinnliga nätverk: fiskeri, jordbruk och diversifiering. , tillstått att kvinnorna i fiskesektorn inte bara är aktiva inom förädling, upptagande och vattenbruk utan också inom marknadsföring, forskning, journalistik, administration, utbildning och representation i både fiske‑ och vattenbrukssektorerna.
Kvinnorna spelar en viktig roll i förädlingsindustrin, och i en del regioner är över 50 procent av de anställda kvinnor.
Kvinnorna kan i stor utsträckning bidra till fiskeberoende samhällens socioekonomiska utveckling, och dessa möjligheter måste nu skyndsamt tas tillvara.
Att inrikta sig på att integrera kvinnor i beslutsfattande organ och sammanslutningar kan vara ett första steg.
· Ekonomiska frågor
Några klara slutsatser från utfrågningen var att logistiken för marknadstillträde är besvärlig på grund av a) begränsad tillgång på lagringsutrymmen till lands, b) avståndet till marknaden, c) produkternas hållbarhet och d) de små aktörernas begränsade erfarenhet av marknadsföring och företagande.
Föredraganden instämmer i dessa slutsatser och anser att en omfattande fragmentering av avlastningspunkter för fångsterna allvarligt komplicerar kontroller, transporter och marknadsföring.
Fiskarna har ingen stark förhandlingsposition när det gäller produkternas försäljningspris och har svårt att göra sig gällande.
Avsaknaden av marknadsföringsstrukturer av kooperativt slag leder till betydande ekonomiska förluster för fiskarna.
I många fall är konsumentpriserna på kustfiskets produkter överdrivet höga, särskilt på grund av det stora antalet mellanhänder på vägen till marknaden.
De prisökningar som sker kommer aldrig producenterna/fiskarna till del.
· Konkurrens om resurser och arbetskraft
Man kan inte bortse ifrån att det finns olika slags fiskeverksamhet som konkurrerar om samma fisk och skaldjur i samma fysiska utrymme i samma kustområden.
Det finns konkurrens mellan fiskare som arbetar med samma slags fiskeutrustning.
Det finns konkurrens mellan fiskare som använder olika slags fiskeutrustning, till exempel mellan kusttrålare och mycket mindre fartyg.
En annan allvarlig aspekt som man måste ta hänsyn till är konkurrensen från verksamhet på uppgång som till exempel fritidsfisket.
Eftersom det inte finns någon formell ram ökar fritidsfisket spänningarna och skapar agg mot kommersiella användningar.
Om den här frågan inte hanteras på ett seriöst sätt och lösningar kommer fram är det mycket troligt att vi kommer att få se fler konflikter mellan fiskesektorn och andra som använder kusterna.
Föredraganden anser att användningen av områden till havs bör regleras genom att exploaterings‑ och åtkomsträttigheter tilldelas, till exempel genom att utvecklingen av viss verksamhet inskränks och licenser blir obligatoriska, för att motverka konkurrens om resurserna.
· Säkerhetsfrågor
Kustfisket bedrivs för närvarande med småskaliga fartyg som till största delen arbetar i närheten av kusten.
Ett antal åtgärder bör vidtas för att öka säkerheten ombord på dessa fartyg, med tanke på att många fartyg som är kortare än 12 meter är gamla eller omoderna.
Mot bakgrund av de betydande skillnaderna i säkerhet mellan högsjöfiske och småskaliga fiskeflottor är det fortfarande viktigt att reglera säkerheten på små fartyg.
Det koncept som beskrivs i detalj i Miguelezbetänkandet om Fiskeri: säkerhet och olycksorsaker
Europaparlamentets resolution A5‑0087/2001 av den 12 mars 2001 om Fiskeri: säkerhet och olycksorsaker. har antagits av fiskeriutskottet och parlamentet.
6.
SLUTSATSER
Det beror också på sociala förändringar och på ekonomiska aspekter som påverkar driftskostnaderna och skapar efterfrågan på produkterna.
Men det allra viktigaste är att det beror på om vi antar en lämplig EU‑lagstiftning som är utformad specifikt för sektorn i fråga.
Föredraganden vill understryka att vi måste
– erkänna vilken social och ekonomisk betydelse sektorn har,
– förbättra levnadsstandarden för de människor som är beroende av kustfisket,
– införa passande system för yrkesutbildning riktade till berörda grupper i kustfiskebefolkningen, inte minst för att ge bättre kunskaper i marknadsföring,
– locka unga människor till sektorn för att säkra kontinuiteten,
– uppmuntra integration av kvinnor i kustfiskesektorn,
– utveckla och modernisera kustfisket,
– ta fram nya sätt att saluföra produkterna och fullt ut integrera kustfiskarna i marknadsföringen,
– öka samarbetet och bygga ut kommunikationskanalerna mellan berörda organisationer och intressenter,
– integrera den nationella kustfiskeripolitiken med gemenskapspolitiken,
– ta fram åtgärder för att minimera effekterna av de ökade rörliga kostnader som följer av de mycket instabila bränslepriserna,
– införa regler för säkerheten ombord på små fartyg som bedriver kustfiske,
YTTRANDE från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
till fiskeriutskottet
över kustfiske och problem för fiskare som idkar kustfiske
( 2004/2264(INI) )
Föredragande:
Teresa Riera Madurell
FÖRSLAG
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män uppmanar fiskeriutskottet att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
EGT L 359, 19.12.1986, s.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att säkerställa kvinnornas fulla deltagande i kustfiskesamhällenas besluts-, representations- och rådgivningsorgan på europeisk, nationell och regional nivå.
ÄRENDETS GÅNG
Titel
Kustfiske och problem för fiskare som idkar kustfiske
Referensnummer
2004/2264(INI)
Ansvarigt utskott
PECH
Yttrande Tillkännagivande i kammaren
FEMM 13.1.2005
Förstärkt samarbete – tillkännagivande i kammaren
Föredragande av yttrande Utnämning
Teresa Riera Madurell 25.1.2005
Tidigare föredragande av yttrande
Behandling i utskott
5.10.2005
23.1.2006
0.0.0000
Antagande
24.1.2006
Slutomröstning: resultat
+:
–:
0:
22
Slutomröstning: närvarande ledamöter
Edit Bauer, Věra Flasarová, Claire Gibault, Lissy Gröner, Zita Gurmai, Piia-Noora Kauppi, Urszula Krupa, Pia Elda Locatelli, Marie Panayotopoulos-Cassiotou, Teresa Riera Madurell, Raül Romeva i Rueda, Amalia Sartori, Corien Wortmann-Kool, Anna Záborská
Slutomröstning: närvarande suppleanter
Anna Hedh, Mary Honeyball, Christa Klaß, Maria Martens, Zita Pleštinská, Zuzana Roithová, Heide Rühle, Bernadette Vergnaud
Slutomröstning: närvarande suppleanter (art.
178.2)
Anmärkningar (tillgängliga på ett enda språk)
ÄRENDETS GÅNG
Titel
Kustfiske och problem för fiskare som idkar kustfiske
Förfarandenummer
2004/2264(INI)
Ansvarigt utskott Tillstånd: tillkännagivande i kammaren
PECH 13.1.2005
Rådgivande utskott Tillkännagivande i kammaren
FEMM 13.1.2005
Inget yttrande avges Beslut
Förstärkt samarbete Tillkännagivande i kammaren
Föredragande Utnämning
Seán Ó Neachtain 25.11.2004
Tidigare föredragande
Behandling i utskott
23.11.2005
29.11.2005
20.3.2006
Antagande
19.4.2006
Slutomröstning: resultat
+:
–:
24
5
Slutomröstning: närvarande ledamöter
James Hugh Allister, Stavros Arnaoutakis, Elspeth Attwooll, Marie-Hélène Aubert, Iles Braghetto, Luis Manuel Capoulas Santos, David Casa, Paulo Casaca, Zdzisław Kazimierz Chmielewski, Carmen Fraga Estévez, Ioannis Gklavakis, Alfred Gomolka, Pedro Guerreiro, Ian Hudghton, Heinz Kindermann, Henrik Dam Kristensen, Albert Jan Maat, Willy Meyer Pleite, Rosa Miguélez Ramos, Philippe Morillon, Seán Ó Neachtain, Bernard Poignant, Struan Stevenson, Margie Sudre
Slutomröstning: närvarande suppleant(er)
Simon Coveney, Chris Davies
Slutomröstning: närvarande suppleant(er) (art.
178.2)
Carlos Carnero González, Salvador Garriga Polledo, Eugenijus Gentvilas, Antonio Masip Hidalgo
Ingivande
26.4.2006
Anmärkningar (tillgängliga på ett enda språk)
SLUTLIG VERSION
A6-0187/2006
*
BETÄNKANDE
om Republiken Österrikes, Republiken Finlands och Konungariket Sveriges initiativ inför antagandet av rådets rambeslut om ett europeiskt verkställighetsbeslut och överförande av dömda personer mellan Europeiska unionens medlemsstater
(7307/2005 – C6‑0139/2005 – 2005/0805(CNS))
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Föredragande:
Ioannis Varvitsiotis
PE 371.769v03-00
Teckenförklaring
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................34
ÄRENDETS GÅNG..................................................................................................................37
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om Republiken Österrikes, Republiken Finlands och Konungariket Sveriges initiativ inför antagandet av rådets rambeslut om ett europeiskt verkställighetsbeslut och överförande av dömda personer mellan Europeiska unionens medlemsstater
(7307/2005 – C6‑0139/2005 – 2005/0805(CNS) )
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
– med beaktande av Republiken Österrikes, Republiken Finlands och Konungariket Sveriges initiativ (7307/2005)
EUT C 150, 21.6.2005, s.
1. ,
– med beaktande av artiklarna 93 och 51 i arbetsordningen,
– med beaktande av betänkandet från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor ( A6‑0187/2006 ).
2.
Rådet uppmanas att på nytt höra Europaparlamentet om rådet har för avsikt att väsentligt ändra Republiken Österrikes, Republiken Finlands och Konungariket Sveriges initiativ.
Republiken Österrikes, Republiken Finlands och Konungariket Sveriges initiativ
Parlamentets ändringar
Ändringsförslag
1
Titeln
Rådets rambeslut om ett europeiskt verkställighetsbeslut och överförande av dömda personer mellan Europeiska unionens medlemsstater
Rådets rambeslut om tillämpning av principen om ömsesidigt erkännande på brottmålsdomar avseende frihetsstraff eller frihetsberövande åtgärder i syfte att verkställa dessa domar i Europeiska unionen
Motivering
Titeln på rambeslutet ändras på grund av de ändringar som gjorts i rådets arbetsgrupp och för att lägga tonvikten på dokumentets båda grundläggande aspekter, nämligen ömsesidigt erkännande och verkställande av frihetsstraff.
Erkännandet och verkställigheten bör inte ske på grundval av ett ”europeiskt verkställighetsbeslut” utan på grundval av domen och ett intyg.
Ändringsförslag
2
Skäl 5
(5) I förbindelserna mellan medlemsstaterna, som präglas av ett särskilt ömsesidigt förtroende för de övriga medlemsstaternas rättssystem, bör man gå längre än enligt befintliga instrument från Europarådet som rör överförande av verkställighet av straff.
Ett grundläggande åtagande bör fastställas för den verkställande staten att ta emot de av sina medborgare och de personer som är varaktigt lagligt bosatta på dess territorium, vilka i en annan medlemsstat slutligt dömts till frihetsstraff eller omfattas av beslut om frihetsberövande, oberoende av deras samtycke, såvida inte särskilda skäl för vägran föreligger .
(5) I förbindelserna mellan medlemsstaterna, som präglas av ett särskilt ömsesidigt förtroende för de övriga medlemsstaternas rättssystem, bör man gå längre än enligt befintliga instrument från Europarådet som rör överförande av verkställighet av straff och göra det möjligt för den verkställande staten att erkänna domar som avkunnats av myndigheterna i den utfärdande staten .
Trots att den dömda personen måste ges tillfredsställande skydd bör det inte längre vara nödvändigt att han eller hon medverkar i förfarandet genom att hans eller hennes samtycke krävs för att en dom skall översändas till en annan medlemsstat för erkännande och verkställighet av den ådömda påföljden .
Motivering
Syftet är att främja samarbetet när det gäller verkställandet av domar i brottmål.
Ändringsförslaget är i enlighet med 1997 års tilläggsprotokoll till Europarådets konvention från 1983, i vilken tillämpningsområdet för den dömda personens samtycke begränsas.
Ändringsförslag
3
Skäl 5a (nytt)
(5a) Det ömsesidiga förtroendet för det europeiska området för frihet, säkerhet och rättvisa i brottmål måste stärkas genom åtgärder på europeisk nivå som syftar till bättre harmonisering och ömsesidigt erkännande av domar i brottmål och genom införande av viss europeisk straffrättslig lagstiftning och praxis.
Motivering
Ändringsförslaget grundar sig på tanken om att främja en europeisk strafflagstiftning.
Ändringsförslag
4
Skäl 6
(6) Överförande av dömda personer till den stat där personen är medborgare , den stat där de är lagligen bosatta eller den stat till vilken personerna har nära anknytning för avtjänande av straffet främjar deras sociala återanpassning.
(6) Överförande av dömda personer till den stat där dessa är medborgare eller den stat där de är stadigvarande lagligt bosatta för avtjänande av straffet kommer att underlätta deras sociala återanpassning.
Motivering
Begreppet ”nära anknytning” är oklart och skulle behöva en omfattande definition.
Ändringsförslag
5
Skäl 7
(7) Detta rambeslut avser att stå i överensstämmelse med de grundläggande rättigheter och de principer som erkänns i artikel 6 i fördraget och återspeglas i Europeiska unionens stadga om de grundläggande rättigheterna, särskilt i kapitel VI i denna.
Inget i detta rambeslut bör tolkas som ett förbud att vägra verkställa ett beslut om det finns objektiva skäl att tro att påföljden syftar till att straffa en person på grundval av dennes kön, ras, religion, etniska ursprung, nationalitet, språk, politiska uppfattning eller sexuella läggning, eller att denna persons ställning kan skadas av något av dessa skäl.
(7) Detta rambeslut avser att stå i överensstämmelse med de grundläggande rättigheter och de principer som erkänns i artikel 6 i fördraget och återspeglas i Europeiska unionens stadga om de grundläggande rättigheterna, särskilt i kapitel VI i denna.
Inget i detta rambeslut bör tolkas som ett förbud att vägra verkställa ett beslut om det finns objektiva skäl att tro att påföljden syftar till att straffa en person på grundval av dennes kön, ras, religion, etniska ursprung, nationalitet, språk, politiska uppfattning eller sexuella läggning, eller att denna persons ställning kan skadas av något av dessa skäl.
Under förfarandet bör även bestämmelserna om processuella rättigheter i brottmål respekteras, såsom dessa anges i rådets rambeslut.
Motivering
På det här sättet garanteras ett mer fullödigt skydd av rättigheterna inom förfarandets ramar.
Ändringsförslag
6
a) europeiskt verkställighetsbeslut: ett beslut fattat av en behörig myndighet i en utfärdande stat som avser verkställighet av en slutlig påföljd som ådömts en fysisk person av en domstol i den staten ,
a) dom: ett beslut eller avgörande av en domstol i den utfärdande staten vilket vunnit laga kraft och innebär att en fysisk person ådöms en påföljd ,
(Om ändringen antas skall hela texten anpassas i överensstämmelse härmed.)
Motivering
Ändringsförslaget återspeglar de ändringar som gjorts under diskussionerna i rådets arbetsgrupp.
Ändringsförslag
7
b) påföljd: varje frihetsstraff eller frihetsberövande åtgärd som utdöms av en domstol efter straffrättsligt förfarande för en straffbar gärning för en angiven tid eller på obestämd tid ,
b) påföljd: varje frihetsstraff eller annan frihetsberövande åtgärd som utdöms under en begränsad eller obegränsad tid på grund av en straffbar gärning efter ett straffrättsligt förfarande ,
Motivering
Ändringsförslaget återspeglar de ändringar som gjorts under diskussionerna i rådets arbetsgrupp.
Ändringsförslag
8
c) utfärdande stat: den medlemsstat där ett europeiskt verkställighetsbeslut har utfärdats ,
c) utfärdande stat: den medlemsstat där en dom i den mening som avses i detta rambeslut har avkunnats ,
Motivering
Ändringsförslaget återspeglar de ändringar som gjorts under diskussionerna i rådets arbetsgrupp.
Ändringsförslag
9
d) verkställande stat: den medlemsstat till vilken ett europeiskt verkställighetsbeslut har översänts för verkställighet.
d) verkställande stat: den medlemsstat till vilken en dom har översänts för erkännande och verkställighet av den ådömda påföljden .
Motivering
Ändringsförslaget återspeglar de ändringar som gjorts under diskussionerna i rådets arbetsgrupp.
Ändringsförslag
10
2.
Utan att det påverkar tillämpningen av artikel 4 får varje medlemsstat, om organisationen av dess interna system gör det nödvändigt, utse en eller flera centrala myndigheter till att ansvara för det administrativa översändandet och mottagandet av ett europeiskt verkställighetsbeslut och att bistå de behöriga myndigheterna.
utgår
Motivering
Genom ändringsförslaget blir åtgärden mer effektiv och mindre byråkratisk.
Ändringsförslag
11
3.
3.
Rådets generalsekretariat skall hålla den erhållna informationen tillgänglig för alla berörda medlemsstater.
Motivering
Genom ändringsförslaget blir åtgärden mer effektiv och mindre byråkratisk.
Ändringsförslag
12
1.
1.
Syftet med detta rambeslut är att fastställa regler för medlemsstaternas erkännande av en dom och verkställande av den ådömda påföljden , oberoende av om verkställigheten redan inletts.
Motivering
Ändringsförslaget är en följd av de ändringar som gjorts i rådets arbetsgrupp och är avsett att lägga tonvikten på dokumentets båda grundläggande aspekter, nämligen ömsesidigt erkännande och verkställande av frihetsstraff.
Erkännandet och verkställigheten bör inte ske på grundval av ett ”europeiskt verkställighetsbeslut” utan på grundval av domen och ett intyg.
Ändringsförslag
13
Om utöver påföljden böter och/eller förverkande har utdömts, men ännu inte betalats, indrivits eller verkställts, skall detta inte hindra översändandet av en dom.
Motivering
Bestämmelsen ingick ursprungligen i artikel 4 i förslaget.
Ändringsförslag
14
Motivering
Ändringsförslag
15
Ändringsförslag
16
– Artikel 8: Erkännande och verkställighet av ett europeiskt verkställighetsbeslut
– Artikel 8: Erkännande och verkställighet av en dom
Motivering
Ändringsförslaget är en följd av de ändringar som gjorts i rådets arbetsgrupp.
Ändringsförslag
17
– Artikel 8: Erkännande och verkställighet av ett europeiskt verkställighetsbeslut
– Artikel 8: Erkännande och verkställighet av en dom
Motivering
Ändringsförslaget är en följd av de ändringar som gjorts i rådets arbetsgrupp.
Ändringsförslag
18
Den stat som utfärdat den europeiska arresteringsordern skall förse den verkställande staten med den information som ett europeiskt verkställighetsbeslut innehåller .
De behöriga myndigheterna skall kommunicera direkt med varandra i frågor som rör denna punkt.
Den stat som utfärdat den europeiska arresteringsordern skall förse den verkställande staten med domen tillsammans med ett intyg i enlighet med artikel 4 .
De behöriga myndigheterna skall kommunicera direkt med varandra i frågor som rör denna punkt.
Motivering
Ändringsförslaget är en följd av de ändringar som gjorts i rådets arbetsgrupp.
Ändringsförslag
19
Översändande av ett europeiskt verkställighetsbeslut
Översändande av en dom och ett intyg
Motivering
Ändringsförslaget är en följd av de ändringar som gjorts i rådets arbetsgrupp.
Ändringsförslag
20
-1. a) En dom tillsammans med ett intyg enligt denna artikel får översändas till en av följande medlemsstater:
i) Den stat där den dömda personen är medborgare eller stadigvarande lagligt bosatt.
ii) Den stat där den dömda personen är medborgare och till vilken han eller hon kommer att utvisas när han eller hon avtjänat sitt fängelsestraff på grund av domen eller ett administrativt beslut som fattas till följd av domen.
iii) Den stat där den dömda personen är medborgare eller stadigvarande lagligt bosatt och som har överlämnat honom eller henne till den utfärdande staten på grundval av en europeisk arresteringsorder med förbehåll att personen, efter att ha hörts, skall återsändas till den verkställande staten för vidare verkställighet av den påföljd som utdömts mot honom eller henne i den utfärdande staten.
iv) Den stat där den dömda personen befinner sig eller är medborgare i eller är stadigvarande lagligt bosatt och som samtycker till erkännande och verkställighet av påföljden.
v) Den stat där personen är stadigvarande lagligt bosatt, om inte han eller hon har förlorat eller kommer att förlora uppehållstillståndet på grund av domen eller ett administrativt beslut som fattas till följd av domen.
vi) Den stat som samtycker till översändandet av domen tillsammans med intyget för erkännande och verkställighet av den ådömda påföljden.
b) Innan domen översänds skall den behöriga myndigheten i den utfärdande staten särskilt överväga att på lämpligt sätt samråda med den behöriga myndigheten i den verkställande staten.
Samråd är obligatoriskt när domen, i enlighet med de kriterier som fastställs i punkt 1, kan översändas till två eller flera medlemsstater.
c) Den verkställande staten får på eget initiativ begära att den utfärdande staten översänder domen tillsammans med intyget.
Motivering
Detta är en mer objektiv definition av kriterierna för att sända över en dom till en annan medlemsstat.
Ändringsförslag
21
1.
I det sistnämnda fallet får översändandet av ett europeiskt verkställighetsbeslut övervägas endast med den dömda personens samtycke.
Den verkställande staten får även självmant uppmana den utfärdande staten att översända ett europeiskt verkställighetsbeslut.
Den dömda personen får även begära att den utfärdande eller verkställande statens behöriga myndigheter inleder ett förfarande enligt detta rambeslut .
1.
För att den påföljd som utdömts skall kunna erkännas och verkställas, skall den behöriga myndigheten i den utfärdande staten i enlighet med artikel 3a översända domen eller en bestyrkt kopia av den, tillsammans med intyget, direkt till den behöriga myndigheten i den verkställande staten, i form av en skriftlig uppteckning som skall möjliggöra för den verkställande staten att fastställa äktheten.
Originalet av domen, eller en bestyrkt kopia av den, och originalet av intyget skall på begäran översändas till den verkställande staten.
All officiell kommunikation skall också ske direkt mellan de nämnda behöriga myndigheterna .
Motivering
Samma sak gäller för andra liknande rättsliga åtgärder.
Ändringsförslag
22
2.
Ett europeiskt verkställighetsbeslut får inte översändas om personen mot vilken påföljden har utdömts är varaktigt lagligt bosatt i den utfärdande staten, såvida inte den dömda personen lämnar sitt samtycke till överföringen eller beslutet, eller ett administrativt beslut, som fattas till följd av detta innehåller ett avvisnings- eller utvisningsbeslut eller någon annan åtgärd, som innebär att personen inte tillåts stanna på den utfärdande statens territorium efter det att påföljden har avtjänats.
utgår
Motivering
Det bakomliggande syftet med den här punkten omfattas av artikel 3a.
Ändringsförslag
23
3.
Verkställandet av böterna i en annan medlemsstat skall grundas på relevanta bestämmelser på detta område med tillämpning mellan medlemsstaterna.
utgår
Motivering
Ändringsförslaget är en följd av de ändringar som gjorts i rådets arbetsgrupp.
Ändringsförslag
24
3a.
Intyget, för vilket ett standardformulär återges i bilaga A, skall vara undertecknat av den behöriga myndigheten i den utfärdande staten, vilken också skall intyga att dess innehåll är korrekt.
Motivering
Ändringsförslaget är en följd av de ändringar som gjorts i rådets arbetsgrupp.
Ändringsförslag
25
4.
Det europeiska verkställighetsbeslutet skall översändas av den behöriga myndigheten i den utfärdande staten direkt till den behöriga myndigheten i den verkställande staten, i form av en skriftlig uppteckning som skall möjliggöra för den verkställande staten att fastställa äktheten.
Allt officiellt informationsutbyte skall också ske direkt mellan de nämnda behöriga myndigheterna.
4.
Domen skall översändas av den behöriga myndigheten i den utfärdande staten direkt till den behöriga myndigheten i den verkställande staten, i form av en skriftlig uppteckning som skall möjliggöra för den verkställande staten att fastställa äktheten och som kan inbegripa uppgifter i någon form om den dömda personens tid i fängelset .
Allt officiellt informationsutbyte skall också ske direkt mellan de nämnda behöriga myndigheterna.
Motivering
Om två fångar avtjänar samma påföljd och överförs till sina ursprungsländer vid samma tidpunkt – och den ena fången har visat förbättring och uppträtt exemplariskt under denna tid medan den andra har uppfört sig illa och inte alls visat någon bättring och är i behov av ytterligare omsorg och rehabilitering – så är det enligt nuvarande lagstiftning förbjudet enligt lagen om skydd av personuppgifter att överföra rapporter om deras tid i fängelset från den utfärdande staten till den stat som tar emot dem.
Av det här följer att den mottagande staten inte kan veta vilken av fångarna som tryggt kan friges och vilken av dem som fortsättningsvis utgör en fara för samhället.
Ändringsförslag
26
5.
5.
Den utfärdande staten skall översända domen tillsammans med intyget till endast en verkställande stat åt gången.
Motivering
Ändringsförslaget är en följd av de ändringar som gjorts i rådets arbetsgrupp.
Ändringsförslag
27
6.
6.
Om den behöriga myndigheten i den verkställande staten inte är känd av den behöriga myndigheten i den utfärdande staten, skall den sistnämnda vidta alla nödvändiga efterforskningar via kontaktpunkterna i det europeiska rättsliga nätverk som inrättades genom rådets gemensamma åtgärd 98/428/RIF, för att erhålla information från den verkställande staten.
Motivering
Ändringsförslaget är en följd av de ändringar som gjorts i rådets arbetsgrupp.
Ändringsförslag
28
7.
utgår
Motivering
Kontakterna måste ske via de behöriga myndigheterna.
Ändringsförslag
29
Underrättelse till den dömda personen och dennes uppfattning
Underrättelse till den dömda personen och brottsoffren
Motivering
”Uppfattning” stryks eftersom det inte anger den praktiska konsekvensen av att ta hänsyn till den dömdes uppfattning när det gäller överföring och val av stat.
Ändringsförslaget är i enlighet med 1997 års tilläggsprotokoll till Europarådets konvention från 1983, i vilken tillämpningsområdet för den dömda personens samtycke begränsas.
Ändringsförslag
30
1.
En dömd person som befinner sig i den utfärdande staten skall om möjligt ges tillfälle till att muntligt eller skriftligt ange sin uppfattning innan ett europeiskt verkställighetsbeslut utfärdas.
Dennes uppfattning skall dock även i dessa fall beaktas när beslut fattas om huruvida ett europeiskt verkställighetsbeslut skall utfärdas och, i förekommande fall, till vilken verkställande stat det skall översändas.
1.
En dömd person som befinner sig i den utfärdande staten skall ges tillfälle till att muntligt eller skriftligt ange sin uppfattning innan ett europeiskt verkställighetsbeslut utfärdas.
Dennes uppfattning skall dock även i dessa fall beaktas när beslut fattas om huruvida ett europeiskt verkställighetsbeslut skall utfärdas och, i förekommande fall, till vilken verkställande stat det skall översändas.
Motivering
Den dömda personen skall alltid ges tillfälle att yttra sig, detta i enlighet med artikel 39 i Europarådets konvention från 1970 enligt vilken domaren innan ett utfärdandebeslut utfärdas skall ge den dömda personen möjlighet att ge uttryck för sin uppfattning.
Ändringsförslag
31
1a.
Brottsoffren skall också underrättas både om att det finns en ansökan om erkännande och verkställighet av en dom och om resultatet av förfarandet, inbegripet beslutet att överföra den dömda personen från den utfärdande staten till den verkställande staten.
Motivering
Den dömda personens brottsoffer skall också få möjlighet att underrättas om alla förfaranden som avser erkännande och verkställighet av den dömda personens dom i en annan medlemsstat.
Ändringsförslag
32
2.
En dömd person som befinner sig i den utfärdande staten skall underrättas av den behöriga myndigheten i denna stat om följderna av en överföring till den verkställande staten.
Om den dömda personen befinner sig i den verkställande staten skall underrättelsen lämnas av den behöriga myndigheten i den staten , om detta är motiverat i rättvisans intresse .
2.
En dömd person som befinner sig i den utfärdande staten skall underrättas av den behöriga myndigheten i denna stat om följderna av en överföring till den verkställande staten.
Om den dömda personen befinner sig i den verkställande staten skall underrättelsen lämnas av den behöriga myndigheten i den staten.
Motivering
Formuleringen ”om detta är motiverat i rättvisans intresse” är juridiskt vag.
Ändringsförslag
33
Artikel 6
1.
Det europeiska verkställighetsbeslutet skall innehålla den information som anges i formuläret i bilagan.
Den behöriga myndigheten i den utfärdande staten skall underteckna verkställighetsbeslutet och intyga att innehållet är korrekt.
2.
Det europeiska verkställighetsbeslutet skall översättas till det officiella språket eller ett av de officiella språken i den verkställande staten.
Motivering
Ändringsförslaget är en följd av de ändringar som gjorts i rådets arbetsgrupp och är avsett att lägga tonvikten på dokumentets båda grundläggande aspekter, nämligen ömsesidigt erkännande och verkställande av frihetsstraff.
Erkännandet och verkställigheten bör inte ske på grundval av ett ”europeiskt verkställighetsbeslut” utan på grundval av domen och ett intyg.
Ändringsförslag
34
Erkännande och verkställighet av ett europeiskt verkställighetsbeslut
Erkännande av domen och verkställighet av påföljden
Motivering
Ändringen föreslås för att texten skall överensstämma med den ändrade titeln på rambeslutet.
Ändringsförslag
35
1.
1.
Motivering
Ändringen föreslås för att texten skall överensstämma med den ändrade titeln på rambeslutet.
Ändringsförslag
36
2.
Om påföljdens längd är oförenlig med grundläggande principer i den verkställande statens lagstiftning, får den behöriga myndigheten i den verkställande staten besluta att anpassa påföljden till strängaste föreskrivna nivå för ett brott enligt den nationella lagstiftningen i denna stat.
2.
Om påföljdens längd är oförenlig med den verkställande statens lagstiftning, får den behöriga myndigheten i den verkställande staten, efter att ha hört den utfärdande staten, besluta att verkställa påföljden upp till den strängaste föreskrivna nivån för brottet enligt den nationella lagstiftningen i denna stat.
Motivering
Den verkställande staten kommer att sänka påföljden till den högsta påföljdsnivån för motsvarande brottskategori i enlighet med den verkställande statens lagstiftning.
Ändringsförslag
37
3.
Om påföljdens art är oförenlig med den verkställande statens lagstiftning, får den behöriga myndigheten i denna stat genom ett rättsligt eller administrativt beslut anpassa påföljden till ett straff eller en åtgärd som i dess egen lagstiftning föreskrivs för brott av samma typ.
Ett sådant straff eller en sådan åtgärd skall så nära som möjligt motsvara den påföljd som utdömts i den utfärdande staten, vilket innebär att påföljden inte kan omvandlas till bötesstraff.
Påföljden får inte innebära en skärpning av den påföljd som utdömts i den utfärdande staten.
3.
Om påföljdens art är oförenlig med den verkställande statens lagstiftning skall straffet eller åtgärden så nära som möjligt motsvara den påföljd som utdömts i den utfärdande staten, vilket innebär att påföljden inte kan omvandlas till bötesstraff.
Påföljden får inte innebära en skärpning eller sänkning av den påföljd som utdömts i den utfärdande staten.
Motivering
Påföljden enligt den verkställande statens lagstiftning bör hanteras särskilt försiktigt eftersom de påföljder som föreskrivs skiljer sig mellan medlemsstaterna.
Ändringsförslag
38
4.
Efter att ha informerats får den verkställande staten minska påföljden i den utsträckning som den utfärdande staten angett.
4.
Efter att ha informerats får den verkställande staten minska påföljden i den utsträckning som den utfärdande staten angett.
Motivering
I enlighet med de föreslagna ändringarna av artikel 7.
Ändringsförslag
39
1.
De behöriga myndigheterna i den verkställande staten får vägra att erkänna och verkställa ett europeiskt verkställighetsbeslut , om
1.
De behöriga myndigheterna i den verkställande staten får vägra att erkänna domen och verkställa påföljden , om
Ändringsförslag
40
a) den berörda personen har dömts för samma gärning i den verkställande staten eller i en annan stat än den utfärdande eller den verkställande staten, under förutsättning att beslutet i det senare fallet har verkställts, håller på att verkställas eller inte längre kan verkställas enligt den utfärdande statens lagstiftning ,
a) det intyg som avses i artikel 4 är ofullständigt eller uppenbarligen inte överensstämmer med domen ,
Motivering
Ändringsförslag
41
Motivering
-a) (nytt) För att säkerställa överensstämmelsen med artikel 3a.
Ändringsförslag
42
ab) verkställandet av påföljden skulle strida mot principen ne bis in idem,
Motivering
Detta är ett skäl för att vägra att erkänna eller verkställa ett beslut vid brott mot principen ne bis in idem.
Ändringsförslag
43
Motivering
Ändringen föreslås för att texten skall överensstämma med den ändrade titeln på rambeslutet.
Ändringsförslag
44
c) verkställigheten av beslutet har preskriberats enligt den verkställande statens lagstiftning såvida det europeiska verkställighetsbeslutet avser gärningar som omfattas av denna verkställande stats behörighet enligt dess egen lagstiftning,
c) verkställigheten av påföljden har preskriberats enligt den verkställande statens lagstiftning och om denna avser gärningar som omfattas av denna verkställande stats behörighet enligt dess egen lagstiftning,
Ändringsförslag
45
ca) det enligt lagen i den verkställande staten föreligger immunitet som gör det omöjligt att verkställa beslutet,
Ändringsförslag
46
d) det europeiska verkställighetsbeslutet har utfärdats för en fysisk person som enligt lagen i den verkställande staten på grund av sin ålder inte kan göras straffrättsligt ansvarig för de gärningar som det europeiska verkställighetsbeslutet avser,
d) påföljden har ådömts en person som enligt lagen i den verkställande staten på grund av sin ålder inte kan göras straffrättsligt ansvarig för de gärningar som domen avser,
Ändringsförslag
47
e) mindre än sex månader av strafftiden återstår att verkställa vid den tidpunkt då domen tas emot av den behöriga myndigheten i den verkställande staten ,
Motivering
Ändringsförslaget är i enlighet med artikel 7.
Minst sex månader i den verkställande staten stöder tanken om återanpassning.
Ändringsförslag
48
f) den berörda personen inte samtycker till översändandet av det europeiska verkställighetsbeslutet och beslutet avser verkställighet av en påföljd som ådömts i ett beslut som fattats i personens frånvaro, såvida den berörda personen inte personligen kallats eller på annat sätt underrättats om de rättsliga åtgärder som ledde till beslutet som fattades i personens frånvaro, eller om personen inte till en behörig myndighet har meddelat att han eller hon inte bestrider saken ,
f) domen meddelades i personens frånvaro, såvida det inte i intyget anges att personen kallats personligen eller via en behörig företrädare enligt nationell lagstiftning underrättats om tid och plats för de rättsliga förfaranden som ledde till att domen meddelades i personens frånvaro ,
Ändringsförslag
49
g) den fysiska person för vilken det europeiska verkställighetsbeslutet har utfärdats varken är medborgare i den verkställande staten eller är varaktigt lagligt bosatt där eller har nära anknytning till denna stat.
utgår
Ändringsförslag
50
2.
2.
Ändringsförslag
51
2a.
Erkännandet av domen får uppskjutas i den verkställande staten om det intyg som avses i artikel 4 är ofullständigt eller uppenbarligen inte överensstämmer med domen.
Motivering
Ändringsförslaget grundar sig på artikel 18 i rambeslutet om ett europeiskt verkställighetsbeslut.
Ändringsförslag
52
Beslut om ett europeiskt verkställighetsbeslut och tidsfrister
Motivering
Eftersom uttrycket ”europeiskt verkställighetsbeslut” ändrats i hela texten.
Ändringsförslag
53
1.
Den behöriga myndigheten i den verkställande staten skall snarast möjligt , dock senast tre veckor efter att ha tagit emot det europeiska verkställighetsbeslutet, besluta om dess verkställighet .
1.
Motivering
Tidsfristerna måste vara korta men realistiska.
Ändringsförslag
54
1a.
Ändringsförslag
55
1b.
Ändringsförslag
56
2a.
Om det i specifika fall inte går att fatta beslut om erkännande av domen och verkställighet av påföljden inom de tidsfrister som fastställs i punkterna 1a och 1b, skall den behöriga myndigheten i den verkställande staten utan dröjsmål underrätta den behöriga myndigheten i den utfärdande staten om detta samt om skälen till detta.
I ett sådant fall får tidsfristerna förlängas med ytterligare 30 dagar.
Motivering
Tidsfristerna måste vara korta men realistiska.
Ändringsförslag
57
1.
En person för vilken ett europeiskt verkställighetsbeslutet utfärdats och som befinner sig i den utfärdande staten skall överföras till den verkställande staten så snart som möjligt vid en tidpunkt som de berörda myndigheterna i den utfärdande och den verkställande staten skall komma överens om .
1.
En dömd person som befinner sig i den utfärdande staten skall överföras till den verkställande staten senast 30 dagar efter det att den verkställande staten har fattat det slutgiltiga beslutet om att erkänna domen och verkställa påföljden .
Motivering
Tidsfristerna måste vara korta men realistiska.
Ändringsförslag
58
2.
utgår
Ändringsförslag
59
3.
3.
Om oförutsedda omständigheter hindrar att personen överförs inom den tidsfrist som anges i punkt 1 , skall de behöriga myndigheterna i den verkställande och den utfärdande staten omedelbart kontakta varandra.
Överförandet skall äga rum så snart dessa omständigheter inte längre föreligger.
Den behöriga myndigheten i den utfärdande staten skall omedelbart informera den behöriga myndigheten i den verkställande staten och de skall komma överens om en ny tidpunkt för överförandet.
I så fall skall överförandet äga rum inom tio dagar från och med den nya tidpunkt som överenskommits.
Motivering
Ändringsförslag
60
1.
Varje medlemsstat skall tillåta transitering genom sitt territorium av en dömd person som överförs till den verkställande staten, förutsatt att medlemsstaten har fått uppgifter om
1.
Varje medlemsstat skall underrättas om transitering genom sitt territorium av en dömd person som överförs till den verkställande staten och erhålla en kopia av intyget från den utfärdande staten .
a) identitet och nationalitet på den person som är föremål för ett europeiskt verkställighetsbeslut ,
b) att det finns ett europeiskt verkställighetsbeslut ,
c) brottets art och brottsrubricering för det brott som ligger till grund för det europeiska verkställighetsbeslutet ,
d) beskrivning av brottets omständigheter, inklusive tidpunkt och plats .
Motivering
Information om, i stället för tillåtelse till transitering skulle göra det hela mindre byråkratiskt.
Ändringsförslag
61
2.
Transiteringsmedlemsstaten skall meddela sitt beslut, som skall fattas med prioritet senast en vecka efter mottagandet av framställningen enligt samma förfarande.
2.
Framställningen om transitering samt det intyg som avses i punkt 1 får översändas på varje sätt som gör det möjligt att få en skriftlig uppteckning.
Transiteringsmedlemsstaten skall meddela sitt beslut, som skall fattas med prioritet senast en vecka efter mottagandet av framställningen enligt samma förfarande.
Ändringsförslag
62
2a.
Transiteringsmedlemsstaten får hålla den dömda personen i fängsligt förvar endast under den tid som krävs för transitering genom dess territorium.
Ändringsförslag
63
3.
Om en icke planerad landning görs skall emellertid den utfärdande medlemsstaten lämna de uppgifter som avses i punkt 1.
3.
Vid transport med flyg utan planerad mellanlandning skall inte någon underrättelse om transitering krävas.
Om en icke planerad landning görs skall emellertid den utfärdande medlemsstaten lämna de uppgifter som avses i punkt 1 inom 48 timmar .
Ändringsförslag
64
1.
Det europeiska verkställighetsbeslutets verkställighet regleras av lagen i den verkställande staten på samma sätt som för påföljder utfärdade av den verkställande staten .
Myndigheterna i den verkställande staten skall med förbehåll för punkterna 2 och 3 ha behörighet att besluta om verkställighetsförfarandena och att fastställa alla åtgärder i samband därmed, inklusive grunderna för villkorlig frigivning.
1.
Verkställigheten av en påföljd regleras av lagen i den verkställande staten.
Myndigheterna i den verkställande staten skall med förbehåll för punkterna 2 och 3 ha behörighet att besluta om verkställighetsförfarandena och att fastställa alla åtgärder i samband därmed, inklusive grunderna för villkorlig frigivning.
Ändringsförslag
65
2.
2.
Från det frihetsstraff som totalt skall avtjänas i den verkställande staten skall den behöriga myndigheten i den verkställande staten göra avdrag motsvarande hela den period av frihetsstraffet som redan avtjänats av den dömda personen i samband med den påföljd som ligger till grund för domen .
Ändringsförslag
66
3.
3.
Såvida inte annat avtalats mellan den utfärdande och den verkställande staten får villkorlig frigivning beviljas endast om den dömda personen har avtjänat totalt minst hälften av påföljden i den utfärdande och den verkställande staten eller har avtjänat en påföljd under en viss tid i enlighet med bestämmelserna i den utfärdande och den verkställande statens lagstiftning .
Motivering
Europarådets expertgrupp för de europeiska konventionerna om brottmål påpekade i sitt yttrande av den 22 januari att fastställandet av ett minimitak för påföljden skulle skada flexibiliteten och hindra beslutsfattande i enlighet med de enskilda fallen.
Gruppen uttalade sig följaktligen för en lösning baserad på idén om en viss tidsperiod som är förenlig med rättvisans syften.
Ändringsförslag
67
1a.
Punkt 1 skall tillämpas på personer som överförs när de passerar genom tranisteringsmedlemsstater.
Motivering
Specialitetsbestämmelsen måste införas för att de dömda personernas rättigheter skall skyddas när kravet på deras samtycke tas bort.
Ändringsförslag
68
1.
Amnesti eller nåd får beviljas av den utfärdande staten och även av den verkställande staten.
1.
Amnesti eller nåd får beviljas av den utfärdande staten i samråd med den verkställande staten eller av den verkställande staten.
Motivering
Det är inte acceptabelt att den utfärdande staten har rätt att bevilja amnesti eller nåd om den dömda personen har överförts till den verkställande staten och den verkställande statens lagstiftning gäller.
Ändringsförslag
69
b) om ett beslut att inte erkänna och verkställa det europeiska verkställighetsbeslutet enligt artikel 9 och om skälen till beslutet,
b) om ett beslut att i enlighet med artikel 9 helt eller delvis inte erkänna domen och verkställa påföljden samt om skälen till beslutet,
Ändringsförslag
70
Motivering
Man måste vara särskilt försiktig när det gäller skillnaderna mellan medlemsstaterna i fråga om påföljder.
Ändringsförslag
71
Ändringsförslag
72
e) om att den berörda personen utan skäl underlåtit att börja avtjäna påföljden,
utgår
Ändringsförslag
73
ga) när domen väl har erkänts och godkänts.
Ändringsförslag
74
Artikel 17a
Språk
Intyget, för vilket ett standardformulär återges i bilagan, skall översättas till det officiella språket eller ett av de officiella språken i den verkställande staten.
Varje medlemsstat kan i samband med rambeslutets antagande eller vid en senare tidpunkt, i en förklaring som skall deponeras hos rådets generalsekretariat, förklara att den kommer att godta en översättning till ett eller flera andra av de officiella språken i unionen.
MOTIVERING
1.
Inledning
Detta är ett initiativ från Österrike, Finland och Sverige som syftar till att påskynda överföringen av dömda personer till en viss stat som dessa på något sätt har anknytning till och där det anses vara troligt att en optimal social återanpassning kan ske.
Rambeslutet ger en smidig mekanism för att en medlemsstat som personen i fråga är medborgare i, är bosatt i eller har nära band till skall kunna erkänna och verkställa domar som innebär frihetsberövande eller säkerhetsåtgärder (vid sinnesjukdom eller nedsatt tillräknelighet) och som en domstol i en annan medlemsstat har avkunnat.
Initiativet tar hänsyn till slutsatserna från Tammerfors och särskilt till det utökade ömsesidiga erkännandet av beslut i brottmål, uppmuntrandet av ömsesidig tillit mellan de nationella rättsliga myndigheterna och unionens utarbetande av en konsekvent straffrättslig politik för att på ett effektivt sätt bekämpa allvarliga brott i alla former, särskilt genom att fastställa minimipåföljder.
Enligt Europarådets konvention om överförande av dömda personer av den 21 mars 1983, som alla medlemsstater har ratificerat, kan dömda personer endast överföras till den stat där de är medborgare för att avtjäna återstoden av sina påföljder där, och endast om de själva och de berörda staterna samtycker till detta.
I tilläggsprotokollet till konventionen av den 18 december 1997, som man bör notera att inte alla medlemsstater har undertecknat, begränsas de dömda personernas utrymme för samtycke.
En första diskussion ägde rum i utskottet för medborgerliga fri‑ och rättigheter samt rättsliga och inrikes frågor den … och ett arbetsdokument delades ut.
2.
Syftet med förslaget
Den ursprungliga texten (7307/05 COPEN 54) har redan ändrats av den ansvariga arbetsgruppen i rådet, så att följande centrala punkter i dokumentet framkom:
· Kriterierna för att överföra en dömd person från en medlemsstat till en annan för att denne skall avtjäna återstoden av sin påföljd där är: a) medborgarskap tillsammans med laglig bosättning, b) stadigvarande laglig bosättning, och c) den stat som den dömde samtycker till att bli överförd till och till vilken han eller hon har nära anknytning.
När beslutet översänds till den verkställande staten tillåts den dömda personen att muntligt eller skriftligt framföra sin uppfattning om han eller hon inte har rätt att överklaga.
· En förteckning över 32 brott, identisk med den som återfinns i rambeslut 2002/584/RIF om en europeisk arresteringsorder, som skall medföra erkännande och verkställighet av beslut som innebär frihetsberövande utan kontroll av dubbel straffbarhet för gärningen.
Påföljden kan inte under några omständigheter omvandlas till ett bötesstraff och den får heller inte vara strängare än den påföljd som den utfärdande staten har utdömt.
· Skäl för att inte erkänna och inte verkställa ett beslut: a) intyget är inte ifyllt, b) kriterierna för överföring av den dömda personen är inte uppfyllda, c) brott mot principen om förbud mot dubbel lagföring, d) domen avser ett brott som inte finns med i förteckningen i artikel 7, e) preskription, f) asyl eller privilegier, g) personen har inget brottsansvar, samt h) det återstår mindre än fyra månader att avtjäna av påföljden.
3.
Föredragandens uppfattning
1.
Begreppet ”till vilken personerna har nära anknytning” måste klargöras, för de fall då beslutet bara översänds med den dömdes samtycke.
Det bör också göras en klar åtskillnad mellan kriterierna ”medborgarskap” och ”stadigvarande bosättning”.
2.
Begreppet ”uppfattning” (den dömda personens uppfattning, muntlig eller skriftlig) kan ses över eftersom det inte specificerar de praktiska konsekvenserna av att ta hänsyn till denna uppfattning i fråga om överföringen och valet av stat.
3.
Den dömda personens offer bör också kunna få information om beslutet att överföra personen i fråga till en annan medlemsstat, i enlighet med bestämmelserna i rådets rambeslut 2001/220/RIF av den 15 mars 2001 om brottsoffrets ställning i straffrättsliga förfaranden.
Särskild hänsyn bör tas till offrens utsatta position, eventuella skadeståndsprocesser och deras rätt att få information om utgången av processerna och delta personligen, en rätt som upphävs om den dömda personen överförs till ett annat land.
Brottsoffren bör således garanteras likabehandling och respekt för sin värdighet, och deras rättigheter och rättsliga intressen i processen bör tryggas.
4.
Det finns många invändningar mot att inkludera förteckningen över specifika brott.
Minimipåföljden bör fastställas till högst tre år, och man bör också se till att det återstår minst sex månader att avtjäna av påföljden i den verkställande staten.
Genom kontroll av dubbel straffbarhet undviker man överföringar i syfte att avtjäna påföljder för gärningar som inte definieras som brott i den stat personen överförs till.
5.
Man bör vara särskilt försiktig med att anpassa de utdömda påföljderna till lagen i den verkställande staten, med tanke på skillnaderna i preskribering av påföljder mellan medlemsstaterna.
6.
Det krävs för många uppgifter under överföringsförfarandet, t.ex. ”brottets art och brottsrubricering” och ”beskrivning av brottets omständigheter”.
Hela förfarandet är för byråkratiskt och formellt.
Dessutom har föredraganden invändningar mot att man talar om att en av EU:s medlemsstater ”tillåter” transitering genom sitt territorium av en dömd person, eftersom det handlar om ett enda stort område där det råder fri rörlighet för personer och där gränserna har avskaffats.
(Specialitetsprincipen bör eventuellt utvidgas till att omfatta de medlemsstater som den dömda personen passerar vid överföringen.)
7.
Specialitetsprincipen bör tryggas för att se till att den dömda personen inte ställs inför rätta för andra gärningar än dem som han avtjänar sin påföljd för, eftersom man strävar efter att minska de dömda personernas utrymme för samtycke.
8.
Det är inte acceptabelt att den utfärdande staten har rätt till amnesti, benådning eller förnyad prövning om den dömda personen har överförts till den verkställande staten och denna stats lagstiftning därför är tillämplig.
Möjligen efter samråd med den utfärdande staten.
9.
Diskussionsämne: tanken att främja europeisk straffrätt.
ÄRENDETS GÅNG
Titel
Republiken Österrikes, Republiken Finlands och Konungariket Sveriges initiativ inför antagandet av rådets rambeslut om ett europeiskt verkställighetsbeslut och överförande av dömda personer mellan Europeiska unionens medlemsstater
Referensnummer
7307/2005 – C6-0139/2005 – 2005/0805(CNS)
Begäran om samråd med parlamentet
18.5.2005
LIBE 26.5.2005
Inget yttrande avges Beslut
Ioannis Varvitsiotis 4.7.2005
Tidigare föredragande
Behandling i utskott
24.1.2006
20.3.2006
18.4.2006
Antagande
15.5.2006
Slutomröstning: resultat
+:
–:
0:
38
Slutomröstning: närvarande ledamöter
Alexander Alvaro, Roberta Angelilli, Edit Bauer, Johannes Blokland, Mihael Brejc, Kathalijne Maria Buitenweg, Maria Carlshamre, Giusto Catania, Carlos Coelho, Fausto Correia, Kinga Gál, Patrick Gaubert, Elly de Groen-Kouwenhoven, Ewa Klamt, Magda Kósáné Kovács, Barbara Kudrycka, Stavros Lambrinidis, Romano Maria La Russa, Sarah Ludford, Antonio Masip Hidalgo, Claude Moraes, Lapo Pistelli, Martine Roure, Inger Segelström, Antonio Tajani, Ioannis Varvitsiotis, Manfred Weber, Stefano Zappalà, Tatjana Ždanoka
Slutomröstning: närvarande suppleanter
Camiel Eurlings, Giovanni Claudio Fava, Sophia in 't Veld, Sylvia-Yvonne Kaufmann, Bill Newton Dunn, Marie-Line Reynaud
Slutomröstning: närvarande suppleanter (art.
178.2)
Panagiotis Beglitis, Emine Bozkurt, Pasqualina Napoletano
Ingivande
17.5.2006
Anmärkningar (tillgängliga på ett enda språk)
...
SLUTLIG VERSION
A6-0251/2006
***I
BETÄNKANDE
om förslaget till Europaparlamentets och rådets direktiv om begränsning av utsläppande på marknaden och användning av perfluoroktansulfonat (ändring av rådets direktiv 76/769/EEG)
(KOM(2005)0618 – C6‑0418/2005 – 2005/0244(COD))
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Föredragande:
Carl Schlyter
PE 372.192v02-00
Teckenförklaring
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................17
ÄRENDETS GÅNG..................................................................................................................21
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till Europaparlamentets och rådets direktiv om begränsning av utsläppande på marknaden och användning av perfluoroktansulfonat (ändring av rådets direktiv 76/769/EEG)
( KOM(2005)0618 – C6‑0418/2005 – 2005/0244(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2005)0618 )
Ännu ej offentliggjort i EUT. ,
– med beaktande av artikel 51 i arbetsordningen,
– med beaktande av betänkandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A6‑0251/2006 ).
Kommissionens förslag
Parlamentets ändringar
Ändringsförslag
1
TITELN
Förslag till Europaparlamentets och rådets direktiv om begränsning av utsläppande på marknaden och användning av perfluoroktansulfonat (ändring av rådets direktiv 76/769/EEG)
Förslag till Europaparlamentets och rådets direktiv om begränsning av utsläppande på marknaden och användning av perfluoroktansulfonat och perfluoroktansyra (ändring av rådets direktiv 76/769/EEG)
Motivering
Förenta staternas miljöskyddsbyrå EPA har funnit att perfluoroktansyra (PFOA) och dess salter ger upphov till liknande problem eftersom strukturen påminner om PFOS.
I en bedömning från 2002 fanns indikationer på systemisk toxicitet och carcinogenicitet, och bloddata visade att allmänheten i hög grad var utsatt.
Flera studier har visat att PFOA och dess salter dessutom är mycket persistenta i miljön samt att de inte är biologiskt nedbrytbara under normala miljöförhållanden.
PFOA är dessutom mycket persistent i människor, den metaboliseras inte och halveras först efter många år.
I detta direktiv bör det därför även införas begränsningar för PFOA och dess salter.
Ändringsförslag
2
SKÄL 1
(1) OECD har gjort en farobedömning mot bakgrund av den information som fanns tillgänglig i juli 2002.
Enligt bedömningen ger de potentiella riskerna med perfluoroktansulfonat (PFOS) skäl till oro.
(1) OECD har gjort en farobedömning mot bakgrund av den information som fanns tillgänglig i juli 2002.
Enligt bedömningen är perfluoroktansulfonat (PFOS) persistent, bioackumulerande och toxiskt för däggdjur och ger därför skäl till oro.
Motivering
PFOS viktigaste riskegenskaper enligt OECD:s farobedömning bör specificeras.
Ändringsförslag
3
SKÄL 1A (nytt)
(1a) Perfluoroktansyra (PFOA) och dess salter ger upphov till liknande problem eftersom strukturen påminner om PFOS.
Studier har visat att PFOA och dess salter har en potentiellt systemisk toxicitet och carcinogenicitet, och bloddata har visat att allmänheten i hög grad är utsatt för exponering.
PFOA och dess salter är mycket persistenta i miljön och är inte biologiskt nedbrytbara under normala miljöförhållanden.
PFOA är dessutom mycket persistent i människor, metaboliseras inte och halveras först efter flera år.
Den vetenskapliga rådgivande panelen vid Förenta staternas miljöskyddsbyrå har därför föreslagit att PFOA skall klassificeras som ett ämne som troligen är cancerogent för människor.
Motivering
Eftersom PFOS och PFOA är så lika bör även PFOA omfattas av detta direktiv.
Förenta staternas miljöskyddsbyrå EPA har bevisat att PFOA är mycket persistent och bioackumulerande.
I ett förslag till översyn av EPA:s utkast till riskbedömning föreslår den vetenskapliga rådgivande panelen att PFOA skall klassificeras som ett ämne som troligen är cancerogent för människor.
I februari 2006 röstade panelen för inbördes utvärdering för att godta rekommendationen att PFOA skall betraktas som ett ämne som troligen är cancerogent, i enlighet med panelens förslag till rapport från januari 2006.
Ändringsförslag
4
SKÄL 3
(3) Vetenskapliga kommittén för hälso- och miljörisker (SCHER) har rådfrågats.
Enligt SCHER behövs det fler vetenskapliga riskbedömningar av PFOS, men kommittén anser också att det kan bli nödvändigt med riskbegränsningsåtgärder för att undvika att tidigare användningar återupptas.
Enligt SCHER förefaller den nuvarande kritiska användningen inom flygindustrin, halvledarindustrin och den fotografiska industrin inte utgöra en relevant risk för miljön eller folkhälsan, om utsläppen i miljön och exponeringen på arbetsplatserna minskas.
När det gäller brandsläckningsskum anser SCHEER att hälso- och miljöriskerna med alternativ måste bedömas innan ett slutligt beslut fattas.
Beträffande förkromning bör det göras en bedömning av åtgärderna för att minska utsläppen .
(3) Vetenskapliga kommittén för hälso- och miljörisker (SCHER) har rådfrågats.
Den har funnit att PFOS är mycket persistent, mycket bioackumalerande och toxiskt och kan spridas i miljön över stora avstånd samt ha skadliga effekter.
PFOS uppfyller därför kriterierna för att betraktas som en långlivad organisk förorening enligt Stockholmskonventionen.
Enligt SCHER behövs det fler vetenskapliga riskbedömningar av PFOS, men kommittén anser också att det kan bli nödvändigt med riskbegränsningsåtgärder för att undvika att tidigare användningar återupptas.
Enligt SCHER förefaller den nuvarande kritiska användningen inom flygindustrin, halvledarindustrin och den fotografiska industrin inte utgöra en relevant risk för miljön eller folkhälsan, om utsläppen i miljön och exponeringen på arbetsplatserna minskas.
När det gäller brandsläckningsskum menar SCHER att hälso- och miljöriskerna med alternativ måste bedömas innan ett slutligt beslut fattas.
SCHER föreslår en villkorlig undantagsperiod på fem år för den fotografiska industrin och halvledarindustrin samt för brandsläckningsskum.
Beträffande förkromning föreslår SCHER omedelbara begränsningar .
Motivering
Enligt Vetenskapliga kommittén för hälso- och miljörisker (SCHER) uppfyller PFOS kriterierna för att betraktas som en långlivad organisk förorening.
SCHER föreslår en undantagsperiod på fem år för vissa användningar och undantagslösa begränsningar för förkromning.
Ändringsförslag
5
SKÄL 3A (nytt)
(3a) Både PFOS och PFOA uppfyller kriterierna för att klassificeras som farliga ämnen i enlighet med Europaparlamentets och rådets direktiv 2000/60/EG om upprättande av en ram för gemenskapens åtgärder på vattenpolitikens område 1 .
Enligt det direktivet är Europaparlamentet och rådet skyldiga att anta särskilda åtgärder mot vattenföroreningar.
För prioriterade farliga ämnen skall målet med sådana åtgärder vara att utsläpp och spill upphör eller successivt minskar.
Det är lämpligt att vidta sådana åtgärder för PFOS och PFOA.
_______________________
1 EGT L 327, 22.12.2000, s.
1.
1).
Motivering
PFOS och PFOA uppfyller helt klart kriterierna för att klassificeras som farliga ämnen enligt ramdirektivet om vatten.
Även om de ännu inte har förts upp i förteckningen över prioriterade farliga ämnen bör gemenskapen ändå behandla dem på samma sätt som prioriterade farliga ämnen.
Ändringsförslag
6
SKÄL 4
(4) För att skydda folkhälsan och miljön förefaller det därför nödvändigt att begränsa utsläppandet på marknaden och användningen av PFOS.
Det föreslagna direktivet omfattar största delen av exponeringsriskerna.
Andra smärre användningar av PFOS förefaller inte utgöra någon risk och är därför undantagna.
De kommer att undersökas ytterligare och bli föremål för en särskild konsekvensanalys .
(4) För att skydda folkhälsan och miljön är det därför nödvändigt att begränsa utsläppandet på marknaden och användningen av PFOS och PFOA s å att utsläpp och spill successivt kan minskas .
Undantag för nödvändig användning under ett övergångsstadium bör endast beviljas för användning i kontrollerade slutna system .
Motivering
Ändringsförslag
7
SKÄL 5
(5) Produkter innehållande PFOS bör också begränsas för att skydda miljön.
I detta direktiv bör endast nya produkter begränsas, och det bör därför inte gälla produkter som redan används eller produkter på andrahandsmarknaden.
(5) Varor innehållande PFOS och PFOA bör också begränsas för att skydda miljön.
I detta direktiv bör endast nya produkter begränsas , förutom när det gäller brandsläckningsskum , och det bör därför inte gälla produkter som redan används eller produkter på andrahandsmarknaden.
Medlemsstaterna bör emellertid vidta åtgärder för att förhindra ytterligare utsläpp från sådana produkter.
Motivering
Termen ”produkt” är för allmän och kan utgöra en hänvisning till ett ämne, en beredning eller en vara.
I denna bestämmelse åsyftas emellertid varor, vilka definieras i gemenskapens kemikalielagstiftning, och därför bör termen ”produkt” ersättas av den korrekta termen ”vara”.
Direktivets räckvidd bör utökas så att det även omfattar PFOA.
PFOS har använts i mycket större utsträckning under tidigare år, varför medlemsstaterna måste vidta åtgärder för att skydda människors hälsa mot varor som innehåller PFOS.
Ändringsförslag
8
SKÄL 5A (nytt)
(5a) Med tanke på de särskilda riskerna med PFOS och PFOA bör medlemsstaterna göra en inventering av användningen av PFOS och PFOA som sådana eller ingående i beredningar eller varor och vidta de åtgärder som krävs för att utsläpp och spill av PFOS och PFOA i miljön från de inventerade produkterna skall upphöra.
Motivering
PFOS infördes på marknaden på 1970‑talet.
År 2000 användes ca 500 ton PFOS i EU.
Den nuvarande användningen har sjunkit markant och utgör nu ca 12 ton per år.
Därför kan den s.k. tidigare användningen – som i praktiken fortfarande pågår – mycket väl utgöra den största utsläppskällan.
För att undvika att PFOS från dessa produkter släpps ut i miljön måste medlemsstaterna inventera samtliga produkter som innehåller PFOS och vidta de åtgärder som krävs för att undvika att dessa produkter släpper ut ännu mera PFOS i miljön.
I en sådan inventering bör även PFOA‑baserade produkter ingå.
Ändringsförslag
9
BILAGA, TABELLEN
Bilaga I, punkt XX, högerspalten, led 1 (direktiv 76/769/EEG)
1) Får inte släppas ut på marknaden eller användas som ämne eller beståndsdel i beredningar i en koncentration som är lika med eller högre än 0,1 viktprocent.
1) Får inte släppas ut på marknaden eller användas som ämne eller beståndsdel i beredningar i en koncentration som är lika med eller högre än 0,005 viktprocent.
Motivering
PFOS används på grund av sina särskilda resistenta egenskaper ofta som beläggning eller ytaktivt ämne och används då, i det stora flertalet av användningarna, i små koncentrationer som ligger långt under det normala tröskelvärdet på 0,1 viktprocent.
Det är allmänt känt att 0,1 viktprocent är ett olämpligt tröskelvärde.
Studier som svenska naturvårdsverket genomfört visar att man för att åstadkomma några märkbara begränsningar av dagens användningar av PFOS måste fastställa koncentrationsnivåerna till 0,005 viktprocent i syfte att täcka alla användningar av PFOS‑derivat.
Ändringsförslag
10
BILAGA, TABELLEN
Bilaga I, punkt XX, högerspalten, led 2 (direktiv 76/769/EEG)
2) Får inte släppas ut på marknaden i produkter eller delar av dem i en koncentration som är lika med eller högre än 0,1 viktprocent.
2) Får inte släppas ut på marknaden i varor eller delar av dem i en koncentration som är lika med eller högre än 0,005 viktprocent i ett homogent material som inte mekaniskt kan sönderdelas i olika material .
Motivering
PFOS används på grund av sina särskilda resistenta egenskaper ofta som beläggning eller ytaktivt ämne och används då, i det stora flertalet av användningarna, i små koncentrationer som ligger långt under det normala tröskelvärdet på 0,1 viktprocent.
Det är allmänt känt att 0,1 viktprocent är ett olämpligt tröskelvärde.
Studier som svenska naturvårdsverket genomfört visar att man för att åstadkomma några märkbara begränsningar av dagens användningar av PFOS måste fastställa koncentrationsnivåerna till 0,005 viktprocent i syfte att täcka alla användningar av PFOS‑derivat.
Ändringsförslag
11
BILAGA, TABELLEN
Bilaga I, punkt XX, högerspalten, led 3, strecksats 1 (direktiv 76/769/EEG)
– fotoresister eller antireflexbeläggning för fotolitografiska processer,
* Åtta år efter detta direktivs ikraftträdande.
1 Kommissionens direktiv 2001/59/EG av den 6 augusti 2001 om anpassning till tekniska framsteg för tjugoåttonde gången av rådets direktiv 67/548/EEG om tillnärmning av lagar och andra författningar om klassificering, förpackning och märkning av farliga ämnen (EGT L 225, 21.8.2001, s.
1).
Motivering
Bruket av PFOS i dessa kritiska användningar sker i noga övervakade slutna system och utgör en minimal risk för människors hälsa och miljön.
Ändringsförslag
12
BILAGA, TABELLEN
Bilaga I, punkt XX, högerspalten, led 3, strecksats 2 (direktiv 76/769/EEG)
– industriell ytbehandling av film, filmpapper eller fotoplåtar,
* Sex år efter det att detta direktiv har trätt i kraft.
Motivering
Det finns för närvarande ett litet antal användningar av PFOS-ämnen i bruk i samband med fotoframställning.
Dessa kemikalier har unika egenskaper under framställningen, användningen och hanteringen av vissa fotografiska produkter och i dagsläget finns det inte något alternativ till dem.
Ändringsförslag
13
BILAGA, TABELLEN
Bilaga I, punkt XX, högerspalten, led 3, strecksats 3 (direktiv 76/769/EEG)
– medel för att förhindra dimbildning vid förkromning,
utgår
Motivering
Ytbehandlingsindustrins användning av PFOS står för den överlägset största delen av utsläppen i miljön.
SCHER stöder en begränsning.
Användningen av PFOS i dekorativ förkromning kan ersättas genom att man byter ut Cr (VI) mot Cr (III) med betydande driftskostnadsbesparingar efter den inledande engångskostnaden.
Användningen av PFOS som medel för att förhindra dimbildning vid hård förkromning och plätering av plast kan ersättas av mekaniska alternativ för att förhindra dimbildning samt förbättrad ventilation.
Det finns därför inget skäl att undanta förkromning.
Ändringsförslag
14
BILAGA, TABELLEN
Bilaga I, punkt XX, högerspalten, led 3, strecksats 4 (direktiv 76/769/EEG)
– hydrauloljor inom flygindustrin,
(c) hydrauloljor inom flygindustrin fram till … * ,
* Tio år efter det att detta direktiv har trätt i kraft.
Motivering
För närvarande finns det inga alternativ till PFOS i hydrauloljor.
Det har påpekats att processen för att godkänna en ny olja för användning i kommersiell luftfart historiskt sett har tagit ungefär tio år från koncept till kommersiell tillverkning.
Det är därför rimligt att tillåta ett tioårigt undantag från utfasningen, så att det finns tillräckligt med tid för att ta fram alternativ.
Om inga säkrare alternativ har blivit tillgängliga kan det tidsbegränsade undantaget förlängas (se ändringsförslag 18).
Ändringsförslag
15
BILAGA, TABELLEN
Bilaga I, punkt XX, högerspalten, led 3, strecksats 5 (direktiv 76/769/EEG)
– brandsläckningsskum,
utgår
Motivering
Brandsläckningsskum som innehåller PFOS står för den överlägset största andelen produkter som innehåller PFOS.
PFOS används inte längre för att tillverka brandsläckningsskum.
Säkrare alternativ fria från organiska halogenföreningar finns redan att tillgå.
I det samråd med berörda parter som hölls i Förenade kungariket om ett nationellt förbud 2005 begärde alla brandkårsorganisationer ett omedelbart användningsstopp och säker avfallshantering.
Med tanke på hur farligt PFOS är kan det inte accepteras att det är tillåtet att använda det kvarvarande lagret (som skadar miljön och hälsan) trots att det finns säkrare alternativ.
Ändringsförslag
16
BILAGA, TABELLEN
Bilaga I, punkt XX, högerspalten, led 3, strecksats 6 (direktiv 76/769/EEG)
– kontrollerade slutna system där koncentrationen av PFOS som går ut i miljön är lägre än 1µg/kg och där utsläppet är lägre än 0,1 viktprocent av det PFOS som används i systemet.
* Sex år efter detta direktivs ikraftträdande.
Motivering
Det behövs en snävare definition av kontrollerade slutna system och en tidsfrist.
Ändringsförslag
17
BILAGA, TABELLEN
Bilaga I, punkt XX, högerspalten, led 3a (nytt) (direktiv 76/769/EEG)
* Datum för detta direktivs ikraftträdande.
** Arton månader efter detta direktivs ikraftträdande.
Motivering
Med tanke på hur farligt PFOS är kan det inte accepteras att det är tillåtet att använda det kvarvarande lagret (som skadar miljön och hälsan) trots att det finns säkrare alternativ.
Ändringsförslag
18
BILAGA, TABELLEN
Bilaga I, punkt XX, högerspalten, led 3b (nytt) (direktiv 76/769/EEG)
Motivering
Det bör gå att förlänga undantaget om tillverkarna kan visa att de trots att de har gjort allt vad de har kunnat inte har lyckats ta fram säkrare alternativ eller alternativa processer.
Ändringsförslag
19
BILAGA, TABELLEN
Bilaga I, punkt XX, högerspalten, led 3c (nytt) (direktiv 76/769/EEG)
(3c) Medlemsstaterna skall göra en inventering av användningen av PFOS som sådant eller ingående i beredningar eller varor.
Medlemsstaterna skall vidta de åtgärder som krävs för att utsläpp och spill av PFOS i miljön från de inventerade produkterna skall upphöra.
Motivering
Eftersom det endast är bilagan i direktiv 76/769/EEG som kommer att föras över till REACH måste alla tilläggsbestämmelser om utfasningen anges i bilagan.
PFOS infördes på marknaden på 1970‑talet.
År 2000 användes ca 500 ton PFOS i EU.
Den nuvarande användningen har sjunkit markant och utgör nu ca 12 ton per år.
Därför kan den s.k. tidigare användningen – som i praktiken fortfarande pågår – mycket väl utgöra den största utsläppskällan.
För att undvika att PFOS från dessa produkter släpps ut i miljön måste medlemsstaterna inventera samtliga produkter som innehåller PFOS och vidta de åtgärder som krävs för att undvika att dessa produkter släpper ut ännu mer PFOS i miljön.
BILAGA, TABELLEN
Bilaga I, punkt XXa (ny) (direktiv 76/769/EEG)
Vänsterspalten:
Högerspalten:
1) Får inte släppas ut på marknaden eller användas som ämne eller beståndsdel i beredningar i en koncentration som är lika med eller högre än 0,005 viktprocent efter … (*) .
2) Får inte släppas ut på marknaden i varor eller delar av varor i en koncentration som är lika med eller högre än 0,005 viktprocent i ett homogent material som inte mekaniskt kan sönderdelas i olika material efter … * .
3) Tillverkarna kan begära undantag från punkterna 1 och 2 före … ** .
Undantag skall beviljas för nödvändiga användningar för en begränsad tid och skall avgöras från fall till fall, om tillverkarna kan visa att de har gjort allt vad de har kunnat för att ta fram säkrare alternativ eller alternativa processer och att säkrare alternativ eller alternativa processer fortfarande saknas.
4) Medlemsstaterna skall upprätta en förteckning över användningar av PFOA som sådan eller ingående i beredningar eller varor.
* Tre år efter det att detta direktiv har trätt i kraft.
** Arton månader efter det att detta direktiv har trätt i kraft. ”
Motivering
På grund av de strukturella likheterna mellan PFOS och PFOA (perfluoroktansyra) bör även PFOA omfattas av detta direktiv.
MOTIVERING
”Allt vetenskapligt arbete är ofullbordat – oavsett om det bygger på observationer eller experiment.
Allt vetenskapligt arbete riskerar att omkullkastas eller förändras av nya vetenskapliga rön.
Detta ger oss emellertid inte frihet att bortse från den kunskap vi redan har, eller att skjuta upp de åtgärder som verkar krävas vid en viss tidpunkt.”
Sir Austin Bradford Hill, skrifter från Royal Society of Medicine, 1965
Inledning
De flesta av oss känner till de stora problemen inom klorindustrin.
Klorkemi står för en grupp ämnen som DDT, PCB:er och CFC:er som förstörde miljön.
Trots att problemen med dessa ämnen blev kända redan på 1960‑talet genom Rachel Carsons bok ”Tyst vår” [”Silent Spring”] tog det flera decennier att fasa ut dem på 1980‑ och 1990‑talen.
Men de finns fortfarande kvar: de förorenar vår miljö, näringskedjan och våra kroppar, skadar ozonlagret och bidrar till klimatförändringar – eftersom de är persistenta.
Många människor önskar att denna typ av industriell kemi kunde förpassas till historien.
Perfluoroktansulfonat (PFOS) – som kommissionens förslag handlar om – står för en relativt ny kategori av perfluorföreningar .
De är ett exempel på hur ett okontrollerat experimenterande med persistenta kemikalier har fortsatt trots ”klorerfarenheterna”.
PFOS står för ett dubbelt misslyckande: den gällande kemikalielagstiftningens oförmåga att skydda människors hälsa och miljön samt oförmågan att lära sig av historien.
Perfluorföreningar – och kemikalielagstiftningens misslyckande
Perfluorföreningar har fått en mängd tillämpningar i konsumentprodukter samt industriella tillämpningar tack vare sin stabilitet och sina avstötande egenskaper.
PFOS var en av huvudkomponenterna i en produkt som tillverkades för att skydda tyg från att få fläckar.
Enligt Vetenskapliga kommittén för hälso‑ och miljörisker (SCHER) är PFOS mycket persistent, mycket bioackumulerande och toxiskt.
PFOS – vars produktion startade på 1970‑talet – har nu blivit en allmänt förekommande förorening.
PFOS har hittats i en rad olika arter världen över – från isbjörn till albatross, från Arktis till mitt i Stilla havet.
I en blodprovsundersökning som WWF genomförde 2004 – i vilken 47 människor från 17 länder, däribland 39 ledamöter av Europaparlamentet, undersöktes – hittades PFOS och sex andra perfluorföreningar i var och en av de 47 försökspersonerna.
Det var kombinationen av PFOS‑föroreningar i en mängd olika arter, inklusive människan, plus oroande toxikologiska data som fick den ledande marknadsaktören att år 2000 självmant upphöra med sin tillverkning av PFOS.
I flera decennier var således användningen av PFOS helt oreglerad, ända till dess att irreversibel skada hade åsamkats: global förorening av ett ämne som är mycket persistent, mycket bioackumulerande och toxiskt.
Perfluorföreningar – och oförmågan att lära av historien
Fluor är en av fem halogener i det periodiska systemet.
Ytterligare två välkända halogener som används mycket i den kemiska industrin är brom och klor.
De delar mycket specifika egenskaper.
De är alla mycket reaktiva – men när de kombineras med en kolatom gör de molekylen mer persistent, och i många fall även mer bioackumulerande och toxisk.
Man hade en naiv förhoppning om att den kemiska industrin hade lärt sig sin läxa från de massiva och pågående miljöskador som orsakas av organiska klorföreningar och att den skulle undvika organisk kemi i samband med brom och fluor.
Tyvärr är det tvärtom.
Tillverkningen av perfluorföreningar startade på 1970‑talet och har ökat markant sedan dess – medan de viktigaste klorföreningarna fasades ut.
Lagstiftaren på efterkälken
Även om det är vanligt att lagstiftaren är sen och ofta begränsar ämnen först när de är på väg ut är PFOS ett extremt exempel på detta.
I detta fall var det den ledande marknadsaktören som insåg att PFOS höll på att bli en för stor risk och därför beslutade att upphöra med sin produktion 2000 – efter mer än 20 års tillverkning.
De behöriga myndigheterna i Förenade kungariket följde upp detta i EU och konstaterade en nationell utfasning för de flesta kvarvarande användningsområden 2004.
Fastän den ledande marknadsaktören även fasade ut sin tillverkning av perfluoroktansyra (PFOA), ett ämne som ger upphov till mycket likartade problem eftersom dess struktur påminner om PFOS, och fastän de största tillverkarna i Förenta staterna har åtagit sig att drastiskt minska utsläppen av PFOA och halterna av PFOA i slutprodukten tar kommissionen inte upp åtgärder angående PFOA i sitt förslag.
Föredraganden föreslår följande ändringar för att stärka kommissionen förslag:
1) Lägre utfasningströskel: Enligt SCHER finns PFOS‑kemikalier i produkter i en koncentration på mellan 0,001 procent och 50 procent.
Det administrativa standardtröskelvärde på 0,1 procent som kommissionen föreslår passar därför inte PFOS.
För att garantera att begränsningen blir effektiv måste tröskeln sänkas till 0,001 procent.
En bred majoritet i utskottet stödde en sänkning av tröskeln till 0,005 procent.
2) Strykning av tre undantag:
Vid vissa kromtillämpningar kan PFOS ersättas genom att Cr (VI) byts ut mot Cr (III), vilket leder till stora besparingar.
I samband med andra tillämpningar kan användningen av PFOS ersättas av mekaniska alternativ för att hindra dimbildning samt förbättrad ventilation.
Det finns därför inget skäl att undanta förkromning.
En bred majoritet i utskottet stödde detta tillvägagångssätt.
PFOS används inte längre vid tillverkningen av brandsläckningsskum.
Det finns stor tillgång på säkrare alternativ fria från organiska halogenföreningar.
Med tanke på hur farligt PFOS är kan det inte accepteras att kvarvarande lager används trots att det finns säkrare alternativ.
En överväldigande majoritet i utskottet stödde detta tillvägagångssätt och förordade en övergångsperiod för att ersätta befintliga lager.
Det är oacceptabelt med ett sådant undantag, särskilt i ospecifika allmänna ordalag.
En överväldigande majoritet i utskottet förordade en snävare definition och en tidsfrist.
3) Tidsbegränsning för de tre återstående undantagen, med möjlighet att förlänga undantaget för två av tillämpningarna: Undantag från utfasningen bör endast beviljas för en begränsad tid, så att alternativ uppmuntras.
Tidsfristerna bör fastställas från fall till fall.
För två av tillämpningarna kan det vara motiverat att tillåta att tidsfristen förlängs om tillverkarna kan visa att de har gjort allt vad de har kunnat för att ta fram säkrare alternativ eller alternativa processer, och att säkrare alternativ eller alternativa processer fortfarande saknas.
En överväldigande majoritet i utskottet stödde en förlängning av tidsfristen för alla undantag.
a.
Fotolitografi : Studier visar att processen för att ersätta PFOS i fotolitografi kommer att ta minst 3–4 år.
Det är därför rimligt att fastställa en tidsplan på fyra år för att fasa ut denna användning, med möjlighet att förlänga detta undantag i enlighet med beskrivningen ovan.
Detta undantag bör endast beviljas när användningen sker i kontrollerade slutna system i den mening som avses i EU:s kemikalielagstiftning.
En överväldigande majoritet i utskottet förordade en förlängd tidsram (8 år).
b.
Industriell ytbehandling av film : Mer än 80 procent av denna användning av PFOS har redan framgångsrikt ersatts av säkrare ämnen under de senaste tio åren.
Med tanke på ytterligare tekniska förändringar på grund av skiftet till digital fotografering är det rimligt att anta att de återstående användningsområdena kan ersättas inom fyra år.
En överväldigande majoritet i utskottet förordade en förlängd tidsram (6 år).
c.
Hydrauloljor inom flygindustrin : Det finns för närvarande inga alternativ till PFOS i hydrauloljor.
Processen för att godkänna en ny olja för användning i kommersiell luftfart har historiskt sett tagit ungefär tio år.
Det är därför rimligt att bevilja ett undantag på tio år från utfasningen – med möjlighet till förlängning (se ovan) – för att få mer tid att utveckla alternativ.
En överväldigande majoritet i utskottet stödde detta tillvägagångssätt.
4) Inventering av de PFOS ‑produkter som används: Med tanke på att PFOS‑tillverkningen sjönk kraftigt efter 2000 kan tidigare användningsområden – som i praktiken fortfarande existerar – mycket väl utgöra den största utsläppskällan.
För att undvika att PFOS från dessa produkter släpps ut i miljön bör medlemsstaterna göra en inventering av samtliga produkter som innehåller PFOS och vidta de åtgärder som krävs för att undvika att dessa släpper ut ännu mer PFOS i miljön.
En bred majoritet i utskottet instämde i detta tillvägagångssätt.
5) Tillägg av PFOA till utfasningens räckvidd: Perfluoroktansyra (PFOA) och dess salter ger upphov till liknande problem eftersom strukturen påminner om PFOS.
I en undersökning av Förenta staternas miljöskyddsbyrå (EPA) från 2002 gjordes bedömningen att det fanns tecken på systemisk toxicitet och carcinogenicitet, och bloddata visar att allmänheten i hög grad är utsatt för exponering.
Många studier har visat att PFOA och dess salter även är mycket persistenta i miljön och i människokroppen.
I detta direktiv bör man därför även föreskriva en utfasning av användningen av PFOA och dess salter senast tre år efter det att direktivet har trätt i kraft.
Med förbehåll för en begäran inom 18 månader kan tillverkarna beviljas undantag för nödvändig användning, om de kan visa att de har gjort allt vad de har kunnat för att utveckla säkrare alternativ eller alternativa processer, och att säkrare alternativ och alternativa processer fortfarande saknas.
I analogi med bestämmelserna för PFOS bör medlemsstaterna även göra en inventering av samtliga produkter som innehåller PFOA och vidta de åtgärder som krävs för att undvika att dessa produkter släpper ut ännu mer PFOS i miljön.
Detta tillvägagångssätt stöddes av en bred majoritet i utskottet.
Slutord
Eftersom de flesta perfluorföreningarna förekommer i små volymer, och på grund av den politiska kompromissen om REACH, tror föredraganden tyvärr att det kan ta lång tid innan REACH kan skydda människors hälsa och miljön mot andra perfluorföreningar, såvida inte specifika åtgärder vidtas mot dessa.
ÄRENDETS GÅNG
Titel
Förslag till Europaparlamentets och rådets direktiv om begränsning av utsläppande på marknaden och användning av perfluoroktansulfonat (ändring av rådets direktiv 76/769/EEG)
Referensnummer
KOM(2005)0618 – C6-0418/2005 – 2005/0244(COD)
Framläggande för parlamentet
5.12.2005
Ansvarigt utskott Tillkännagivande i kammaren
ENVI 13.12.2005
ITRE 13.12.2005
ITRE 21.2.2006
Carl Schlyter 21.2.2006
Tidigare föredragande
Förenklat förfarande – beslut
Behandling i utskott
30.5.2006
13.7.2006
Antagande
13.7.2006
Slutomröstning: resultat
+:
–:
54
1
Slutomröstning: närvarande ledamöter
Adamos Adamou, Georgs Andrejevs, Johannes Blokland, John Bowis, Frieda Brepoels, Dorette Corbey, Avril Doyle, Mojca Drčar Murko, Edite Estrela, Anne Ferreira, Karl-Heinz Florenz, Alessandro Foglietta, Matthias Groote, Françoise Grossetête, Cristina Gutiérrez-Cortines, Satu Hassi, Marie Anne Isler Béguin, Caroline Jackson, Dan Jørgensen, Christa Klaß, Eija-Riitta Korhola, Holger Krahmer, Urszula Krupa, Peter Liese, Linda McAvan, Marios Matsakis, Roberto Musacchio, Péter Olajos, Adriana Poli Bortone, Vittorio Prodi, Frédérique Ries, Guido Sacconi, Karin Scheele, Carl Schlyter, Horst Schnellhardt, Richard Seeber, Kathy Sinnott, Jonas Sjöstedt, Bogusław Sonik, María Sornosa Martínez, Antonios Trakatellis, Thomas Ulmer, Anja Weisgerber, Åsa Westlund, Anders Wijkman
Slutomröstning: närvarande suppleant(er)
Slutomröstning: närvarande suppleant(er) (art.
178.2)
Ingivande
19.7.2006
Anmärkningar (tillgängliga på ett enda språk)
SLUTLIG
A6-0326/2006
*
BETÄNKANDE
om förslaget till rådets beslut om ingående av ett avtal mellan Europeiska gemenskapen och Rumäniens regering om Rumäniens medverkan i den verksamhet som bedrivs av Europeiska centrumet för kontroll av narkotika och narkotikamissbruk
(KOM(2006)0256 – C6‑0321/2006 – 2006/0087(CNS))
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Föredragande:
Jean-Marie Cavada
PE 378.527v02-00
Teckenförklaring
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING............................................................................................................................6
ÄRENDETS GÅNG....................................................................................................................7
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till rådets beslut om ingående av ett avtal mellan Europeiska gemenskapen och Rumäniens regering om Rumäniens medverkan i den verksamhet som bedrivs av Europeiska centrumet för kontroll av narkotika och narkotikamissbruk
( KOM(2006)0256 – C6‑0321/2006 – 2006/0087CNS))
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
– med beaktande av förslaget till rådets beslut ( KOM(2006)0256 )
Ännu ej offentliggjort i EUT. ,
– med beaktande av förslaget till avtal mellan Europeiska gemenskapen och Republiken Rumäniens regering om Rumäniens medverkan i den verksamhet som bedrivs av Europeiska centrumet för kontroll av narkotika och narkotikamissbruk,
1.
MOTIVERING
Som kommissionen påpekar i sitt meddelande gjorde Europeiska rådet vid sitt möte i Luxemburg i december 1997 kandidatländernas deltagande i program och gemenskapsorgan till ett instrument för en förbättrad strategi inför anslutningen och angav samtidigt att det bör avgöras från fall till fall om kandidatländerna skall få delta eller inte.
Kommissionen har följaktligen förhandlat fram bilaterala avtal med Bulgarien, Rumänien och Turkiet som innebär ett stort antal fördelar, i synnerhet den fördelen att dessa länder genom avtalen får en möjlighet att lära känna beslutsprocessen inom Europeiska centrumet för kontroll av narkotika och narkotikamissbruk och medverka när centrumets arbetsprogram fastställs.
Föredraganden godkänner de tekniska och ekonomiska arrangemang som gäller för Bulgariens, Rumäniens och Turkiets medverkan i den verksamhet som bedrivs av centrumet.
Han rekommenderar därför att ingåendet av bilaterala avtal med Bulgarien, Rumänien och Turkiet bör godkännas utan ändringar så att länderna i fråga kan medverka i den verksamhet som bedrivs av Europeiska centrumet för kontroll av narkotika och narkotikamissbruk.
ÄRENDETS GÅNG
Titel
Förslag till rådets beslut om ingående av ett avtal mellan Europeiska gemenskapen och Rumäniens regering om Rumäniens medverkan i den verksamhet som bedrivs av Europeiska centrumet för kontroll av narkotika och narkotikamissbruk
Referensnummer
KOM(2006)0256 – C6‑0321/2006 – 2006/0087(CNS)
Begäran om samråd med parlamentet
27.9.2006
LIBE
BUDG
Jean-Marie Cavada 20.6.2006
Behandling i utskott
12.7.2006
4.10.2006
Antagande
4.10.2006
Ingivande
10.10.2006
SLUTLIG VERSION
A6-0329/2006
10.10.2006
BETÄNKANDE
om begäran om fastställelse av Mario Borghezios immunitet och privilegier
(2006/2151(IMM))
Utskottet för rättsliga frågor
Föredragande:
Maria Berger
PE 378.650v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT...........................................................3
MOTIVERING............................................................................................................................4
ÄRENDETS GÅNG....................................................................................................................9
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
om begäran om fastställelse av Mario Borghezios immunitet och privilegier
( 2006/2151(IMM) )
Europaparlamentet fattar detta beslut
– med beaktande av Mario Borghezios begäran om fastställelse av hans immunitet, med anledning av en skrivelsen daterad den 23 maj 2006 och tillkännagiven i kammaren den 1 juni 2006,
– med beaktande av EG-domstolens domar av den 12 maj 1964 och 10 juli 1986
Mål 101/63, Wagner mot Fohrmann och Krier, svensk specialutgåva I, s.
203 och mål 149/85, Wybot mot Faure m.fl., svensk specialutgåva VIII, s.
703. ,
– med beaktande av betänkandet från utskottet för rättsliga frågor ( A6‑0329/2006 ).
MOTIVERING
I begäran om fastställelse av immunitet hänvisar parlamentsledamoten Borghezio till en skrivelse som han fått från åklagarmyndigheten vid domstolen i Milano angående inledande av straffrättsliga förfaranden (artikel 369 och 369a i den italienska brottmålslagen) och avslutande av förundersökning (artikel 415a brottmålslagen).
Denna artikel har följande ordalydelse:
635, deturpa o imbratta cose mobili o immobili altrui è punito, a querela della persona offesa, con la multa fino a L. 200.000.
Se il fatto è commesso su cose di interesse storico o artistico ovunque siano ubicate o su immobili compresi nel perimetro dei centri storici, si applica la pena della reclusione fino a un anno o della multa fino a lire due milioni e si procede d'ufficio.
13, comma 2, della L. 08.10.97, n.
352.
Art.
639-bis.
631, 632, 633 e 636 si procede d'ufficio se si tratta di acque, terreni, fondi o edifici pubblici o destinati ad uso pubblico.” .
Den 25 januari 2005 skall Borghezio nämligen med en sprejburk ha skrivit orden ”skam över Forleo” på en trottoar framför justitiepalatset i Milano.
Borghezio åberopade framför allt att han under en demonstration med anledning av en terroristdom gett uttryck för sin åsikt genom att på trottoaren skriva ordet ”skam” med en sprejburk som han fått låna av en annan deltagare i demonstrationen.
På detta vis hade han endast gett uttryck för sin åsikt men inte avsiktligt gjort sig skyldig till någon skadegörelse.
I den mån det överhuvudtaget blivit några skador på trottoaren var dessa försumbara.
Att en sådan bagatell tas upp som ett brottmål visar enligt Borghezio att det handlar om fumus persecutionis , dvs. att syftet är att skada honom politiskt.
II.
TEXTER OCH ÖVERVÄGANDEN OM EUROPAPARLAMENTSLEDAMÖTERNAS IMMUNITET
1.
Artiklarna 9 och 10 i protokollet om Europeiska gemenskapernas immunitet och privilegier av den 8 april 1965 lyder som följer:
”9.
Europaparlamentets ledamöter får inte förhöras, kvarhållas eller lagföras på grund av yttranden de gjort eller röster de avlagt under utövandet av sitt ämbete.
10.
Under Europaparlamentets sessioner skall dess ledamöter
a) vad avser deras egen stats territorium, åtnjuta den immunitet som beviljas parlamentsledamöter i deras stat,
b) vad avser alla andra medlemsstaters territorium, inte få kvarhållas eller lagföras.
Immuniteten skall även vara tillämplig på ledamöterna under resan till och från Europaparlamentets mötesplats.
Immuniteten kan inte åberopas av en ledamot som tas på bar gärning och kan inte hindra Europaparlamentet att utöva sin rätt att upphäva en av dess ledamöters immunitet.”
2.
Parlamentets ledamöter får inte ställas till svars för röster de avlagt eller yttranden de gjort under utövandet av sitt mandat.
Ingen parlamentsledamot får utan att dennes kammare gett sitt samtycke utsättas för kroppsvisitation eller husrannsakan och inte omhändertas eller på annat sätt begränsas i sin personliga frihet eller hållas i fängsligt förvar, förutom vid verkställande av en lagakraftvunnen dom eller om ledamoten tas på bar gärning och ett gripande i sådana fall är påbjudet.
Vidare krävs kammarens samtycke för att parlamentsledamöters samtal eller meddelanden skall få avlyssnas eller fångas upp och för att deras post skall få beslagtas.
3.
Förfarandet i Europaparlamentet omfattas av bestämmelserna i artiklarna 6 och 7 i arbetsordningen.
Dessa lyder som följer:
”Artikel 6: Upphävande av immunitet
1.
Parlamentet skall vid utövandet av sina befogenheter i frågor som rör immunitet och privilegier i första hand försöka upprätthålla parlamentets integritet som en demokratisk lagstiftande församling och befästa ledamöternas oberoende när dessa fullgör sina åligganden.
/…/
3.
Varje begäran om fastställelse av immunitet och privilegier som en ledamot eller före detta ledamot lämnar in till talmannen skall tillkännages i kammaren och hänvisas till behörigt utskott.
/…/”
”Artikel 7: Immunitetsförfaranden
1.
Behörigt utskott skall utan dröjsmål, och i den ordning de inkommit, pröva varje begäran om upphävande av immunitet och varje begäran om fastställelse av immunitet eller privilegier.
2.
Utskottet skall lägga fram ett förslag till beslut, i vilket utskottet endast skall rekommendera huruvida en begäran om upphävande av immuniteten eller en begäran om fastställelse av immunitet och privilegier skall bifallas eller avslås.
3.
Utskottet kan uppmana den berörda myndigheten att förse utskottet med alla upplysningar och preciseringar som det anser sig behöva för att kunna ta ställning till om immuniteten bör upphävas eller fastställas.
De har rätt att låta sig företrädas av en annan ledamot.
/…/
6.
7.
Utskottet får emellertid under inga omständigheter uttala sig i skuldfrågan, eller på annat sätt yttra sig över ledamoten eller om det riktiga i att väcka åtal för de uttalanden eller handlingar som tillskrivs ledamoten, inte ens vid tillfällen där utskottet genom prövning av en begäran erhåller detaljerad kunskap i fallet.
/…/”
4.
Sedan sin första femåriga valperiod har Europaparlamentet i sitt arbete utvecklat vissa allmänna principer, som slutgiltigt erkändes genom en resolution av den 10 mars 1987
EGT C 99, 13.4.1987. s.
Syftet med den parlamentariska immuniteten
Den parlamentariska immuniteten är inget privilegium för de enskilda parlamentsledamöterna utan en garanti för parlamentets och dess ledamöters oberoende gentemot andra myndigheter.
Av denna princip följer att det inte handlar om tidpunkten för det påtalade brottet, som kan vara både innan och efter det att ledamoten valts in, utan endast om att skyddet av parlamentet som institution går före skyddet av dess ledamöter.
Till följd av parlamentets olika beslut har det uppstått en enhetlig definition av begreppet europeisk parlamentarisk immunitet, som i princip är oberoende av de regler som tillämpas i de nationella parlamenten.
På så vis undviks att ledamöterna behandlas olika beroende på vilken nationalitet de har.
Detta innebär att immuniteten i medlemsstaternas nationella rätt visserligen beaktas, men vid beslut om huruvida en ledamots immunitet skall upphävas tillämpar Europaparlamentet sina egna fasta principer.
Den parlamentariska immuniteten syftar till att skydda ledamöternas yttrandefrihet och frihet att föra politiska debatter.
Därför har parlamentets behöriga utskott alltid företrätt principen att immuniteten aldrig kan upphävas när de handlingar som ledamoten anklagas för hör till dennes politiska verksamhet eller har direkt koppling till denna.
Till detta räknas bland annat meningsyttringar som kan antas tillhöra ledamotens politiska verksamhet, exempelvis i samband med demonstrationer och offentliga sammankomster, i politiska publikationer, i pressen, i en bok, i TV, genom undertecknande av en politisk avhandling eller inför en domstol.
Till denna princip kommer även andra överväganden som talar mot respektive för ett upphävande av immuniteten, i synnerhet överväganden avseende fumus persecutionis , dvs. förmodandet att den straffrättsliga åtgärden har till syfte att skada ledamotens politiska verksamhet.
Enligt definitionen i motiveringen till Donnezbetänkandet innebär begreppet fumus persecutionis i stora drag att immuniteten inte kan upphävas när det finns anledning att misstänka att den rättsliga åtgärden syftar till att skada ledamotens politiska verksamhet.
Om exempelvis talan väcks av en politisk motståndare kommer immuniteten, fram till dess att motsatsen är bevisad, inte att upphävas om det kan antas att anklagelsen är ämnad att skada ledamoten i fråga i stället för att ge den drabbade gottgörelse.
Immuniteten upphävs inte heller om talan väcks under omständigheter där det är uppenbart att det gjorts enbart för att skada ledamoten.
III.
MOTIVERING TILL FÖRSLAGET TILL BESLUT
Utskottet för rättsliga frågor har ingående dryftat artiklarna 9 och 10 i protokollet och den immunitet och de privilegier som kan komma i fråga.
Utskottet började med att pröva om artikel 9 i protokollet är tillämplig.
Enligt artikel 9 har en ledamot absolut immunitet vad gäller yttranden som han eller hon gjort under utövandet av sitt ämbete.
Mario Borghezio hävdar att han genom att spreja ordet ”skam” på trottoaren framför justitiepalatset gett uttryck för en åsikt som är kopplad till hans ämbete som ledamot i Europaparlamentet.
Att spreja en text med en sprejburk kan i och för sig även vara en meningsyttring, men i det här fallet handlar det inte om meningsyttringen som sådan utan om den skadegörelse som sprejen på trottoaren orsakat.
Vad gäller tillämpningen av artikel 10 första stycket a i protokollet om immunitet och privilegier synes det inte finnas några skäl att anta att det rör sig om fumus persecutionis .
Det finns inga faktorer som talar för att anklagelsen mot Mario Borghezio syftade till att skada hans verksamhet som ledamot i Europaparlamentet.
Man kan utgå ifrån att en sprejaktion som utförts av en annan italiensk medborgare under liknande omständigheter skulle ha beivrats på samma sätt.
IV.
SLUTSATSER
På grundval av ovanstående överväganden och efter att ha prövat argumenten för och emot fastställelse av immunitet rekommenderar utskottet för rättsliga frågor att Mario Borghezios begäran om fastställelse av immunitet avslås.
ÄRENDETS GÅNG
Titel
Begäran om fastställelse av Mario Borghezios immunitet och privilegier
Förfarandenummer
2006/2151(IMM)
Mario Borghezio 23.5.2006 1.6.2006
Ansvarigt utskott Tillkännagivande i kammaren
JURI 1.6.2006
Föredragande Utnämning
Maria Berger 12.6.2006
Tidigare föredragande
Behandling i utskott
12.9.2006
Antagande
3.10.2006
Slutomröstning: resultat
+:
–:
0:
17 1 0
Slutomröstning: närvarande ledamöter
Maria Berger, Carlo Casini, Rosa Díez González, Bert Doorn, Monica Frassoni, Giuseppe Gargani, Klaus-Heiner Lehne, Katalin Lévai, Antonio López-Istúriz White, Hans-Peter Mayer, Aloyzas Sakalas, Francesco Enrico Speroni, Diana Wallis, Rainer Wieland, Tadeusz Zwiefka
Slutomröstning: närvarande suppleant(er)
Jean-Paul Gauzès, Luis de Grandes Pascual, Kurt Lechner, Marie Panayotopoulos-Cassiotou
Slutomröstning: närvarande suppleant(er) (art.
178.2)
Ingivande
10.10.2006
Anmärkningar (tillgängliga på ett enda språk)
...
SLUTLIG VERSION
A6-0442/2006
om nomineringen av Nadezhda Sandolova till uppdraget som ledamot av revisionsrätten
(C6‑0411/2006 – 2006/0811(CNS))
Budgetkontrollutskottet
Föredragande:
José Javier Pomés Ruiz
PE 380.959v03-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
BILAGA 1 : CURRICULUM VITAE OF NADEZHDA SANDOLOVA
BILAGA 2: REPLIES OF NADEZHDA SANDOLOVA TO THE QUESTIONNAIRE
ÄRENDETS GÅNG
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
om nomineringen av Nadezhda Sandolova till uppdraget som ledamot av revisionsrätten
( C6‑0411/2006 – 2006/0811(CNS) )
– med beaktande av artikel 101 i arbetsordningen,
– med beaktande av betänkande från budgetkontrollutskottet ( A6‑0442/2006 ).
BILAGA 1 : CURRICULUM VITAE OF Nadezhda Sandolova
1.
Family name: Sandolova
2.
Forenames: Nadezhda
3.
Date of birth: 17 April, 1956
4.
Nationality: Bulgarian
5.
Education: Higher
Institution
Higher Economic University
Karl Marx, Sofia, Bulgaria
Date: from (month/year): to (month/year)
1976-1980
Degree(s) or Diploma(s) obtained:
M.Sc., Planning, Management and Balance
7.
Language skills: (increasing competence from 1 to 5)
Language
Reading
Speaking
Writing
Bulgarian
5
5
5
German
5
5
5
English
5
5
4
Russian
5
5
5
8.
Membership of professional bodies: N/A
9.
10.
Key qualifications: – audit of the National Central Bank
– audit of state debt
– other specific audits
11.
Experience in foreign postings:
1.Date
2.Date
From 16 April 2004 to the present
From May 2005
to the present
1.Country
2.Country
Paris , France
Norway , Oslo
1.Company
2.Company
Council of Europe Development Bank
INTOSAI Development
Institute
1.Position
2.Position
Member of the Auditing Board
Consultant ASOSAI Training program
12.
Professional Experience Record:
Date: from (month/year) to (month/year)
November 1995 to April 2005
Location
Sofia
Company
National Audit Office
Position
Member of the Board, Head of Specific Audits Department, Liaison Officer
Description
Audit of the National Central Bank, audit of state debt, audit of the Fund for Guaranteeing Bank Deposits, audit of the Bulgarian Agency for Export Insurance, audit of privatisation, audit of state guaranteed credits
Date: from (month/year) to (month/year)
May 1991-Nov 1995
Location
Sofia
Company
Ministry of Industry
Position
Head of Department
Description
Analysis of the debt of state enterprises, granting credits to state enterprises and relations with International Financial Institutions
Date: from (month/year) to (month/year)
1993-1995
Location
Sofia
Company
Sofia Bank Ltd.
Position
Member of the Board of Directors
Description
Management
Date: from (month/year) to (month/year)
1988-to the present
Location
Sofia
Company
St Kliment Ohridski Sofia University
Position
Chief Research Assistant and Lecturer , Faculty of Economics
Description
Teaching micro and macroeconomics ; Public control;
has more than 30 publications in the field of economic reforms
Date: from (month/year) to (month/year)
1980-1986
Location
Sofia
Company
Research Institute of Economics of Construction
Position
Research worker
Description
Financial and economic analysis of construction
BILAGA 2: REPLIES OF Nadezhda SANDOLOVA TO THE QUESTIONNAIRE
PROFESSIONAL EXPERIENCE
1.
Please highlight the main aspects of your professional experience in public finance, management, management auditing.
Most of all, I would like to highlight that my educational background, as well as my professional experience, were entirely orientated to the matters of management, public finance and control.
The main motive in my professional development in these strongly interwoven areas has always been the principle of constant self-improvement through becoming acquainted with the international experience and modern standards and practices.
Some of the main aspects of my experience in the area of management are:
- my activity as a head of division in the Ministry of Industry from 1991 to 1994, where I had the chance to practically take part in the reform of the Bulgarian economy and its setting to act in the conditions of the market.
My functions at that time were the negotiation of the first loans from the World Bank, the relations of our country with the International Monetary Fund, as well as the implementation of any possible measures on the part of the government for the effective use of the consigned credit resource;
- my activity as a member of the Managing Board of one of the largest state banks of that time, from 1993 to 1995.
This position not only gave me a good insight into the reforms at the bank and industrial sectors, but it also enriched my experience of management decisions and work in a collegiate management body.
As main aspects of my professional experience in the area of control and management control in particular, I would point out my activity as a member of National Audit Office (NAO) of the Republic of Bulgaria in the period 1995-2005.
In 1995 the Bulgarian Parliament adopted a decision to reestablish the NAO again on the basis of a new law, after its activity had been stopped for more than 45 years.
I would define these ten years not only as an accumulation of management and audit experience, but also as the biggest challenge in my professional experience.
The establishment of a supreme audit institution, the selection and training of auditors, the study and introduction of international experience in its work, is a process of simultaneous reformation of external audit and its implementation into practice.
From 1998 to 2005 I was Liaison Officer of the Bulgarian National Audit Office.
During these years I took part in the regular meetings of Liaison Officers and in the meetings of the Heads of SAI’s of the countries applying for EU membership and the ECA, as well as in the preparation of the documents for our mutual work with the European Court of Auditors.
In 2001 I was in charge of the self-assessment group of the Contact Committee.
Lastly, but also of great importance, I would like to mention that for all the years, from 1988 until the present moment, I taught at the Faculty of Economy of ‘St.
Kliment Ohridski ’ University of Sofia, in the area of macroeconomics and public finance, with the full awareness that education is the best investment for the future development of a country.
2.
What are the three most important decisions to which you have been party in your professional life?
I would express my opinion that in the management process all decisions are important because they give rise to definite responsibilities and consequences.
But I would mention some of the decisions that I have made during my activity which were a kind of a challenge for me and have brought to positive results in the practice of the institution that I have worked for.
1.
The decision to lead the first audit of the relations between the Central Bank and the state budget and the first audit of State Debt of the Republic of Bulgaria.
For the successful realisation of both audits I am extremely grateful to the European Court of Auditors and also to the Court of Auditors of the Federal Republic of Germany for the support and exchanged experience.
Within the Contact Committee of the Heads of the EU candidate country SAIs and the ECA , the Bulgarian NAO received extremely effective and crucial support in methodological and practical way for the development of audit practices and the introduction of internationally accepted auditing standards.
The joint audit which was carried out, between the Bulgarian National Audit Office and the German Court of Audit and the Court of Audit of Spain in the area of State Debt led to public recognition that the Bulgarian NAO has reached a European professional level in this particular area of auditing.
2.
My decision to develop a methodology and to carry out the first self-assessment of a supreme audit institution, the example being with the Bulgarian National Office in the year 2000.
This decision of mine was motivated and supported by the Contact Committee and SIGMA.
The results were reported at a meeting held in Sofia of the Heads of EU candidate country SAIs and some MS SAIs in 2001, and this practice was evaluated as a leading one in this area.
I have the copyrights for the methodology of self-assessment.
3.
Lastly, but of equal importance, I would like to point out my decision from last year to accept the invitation of IDI INTOSAI to participate as a leading consultant in the development and conduct of a course for state debt auditing, which is designed in Russian and is designed especially for practical use within the countries of the Commonwealth of Independent States (CIS) and Mongolia.
The course should reflect in an adequate way the auditing standards of INTOSAI.
On this year’s annual meeting of the INTOSAI’s Public Debt Committee, a very high grade was given to the content, conduction and contribution of the course for the improvement of audit practices in these countries.
INDEPENDENCE
3.
The Treaty stipulates that the Members of the Court of Auditors shall be “completely independent” in the performance of their duties.
How would you apply this obligation to your prospective duties?
“Completely independent” is stipulated in Article 247 of the Treaty and specified in the Staff Regulations.
More detailed explanation about the supreme audit institutions’ independence is explained in the Lima Declaration.
According to this and in compliance with the internationally accepted standards, the Court of Auditors and its Members should enjoy:
- Institutional independence
- Operational independence
- Financial independence and
- Political independence.
As a Member of the Court I would base my activities and audit opinions only on facts, dates, evidence, audit standards and my professional knowledge and experience.
I must not seek nor take instructions or advice from any government or from any other body.
I will do my best to avoid any incompatibility and I will apply the Court’s policies in respect of independence.
4.
Have you received a discharge for the management duties you carried out previously, if such a procedure applies?
Yes, I have.
I have not received an individual discharge but as a Member of collegiate management bodies which were discharged according to the Bulgarian legal procedures I have.
The procedures were applied as follows:
- From 1993 to 1995 being a Member of the Board of Directors of one of the biggest Bulgarian Trade Banks – Sofia Bank, I received a discharge at the end of every financial year by the Shareholders’ Meeting with the adoption of an Annual Report.
The discharging procedure was stipulated in the Bulgarian Trade Banks Law.
-From 1995 to 2005 being a Member of the National Audit Office of Bulgaria I received a discharge at the end of every budget year by the Parliament with the adoption of the Annual Activity Report of the NAO.
The discharging procedure was stipulated in the National Audit Office Law and Parliament Rules.
5.
Do you have any business or financial holdings or any other commitments, which might conflict, with your prospective duties?
Are you prepared to disclose all your financial interests and other commitments to the President of the Court and make them public?
In case you are involved in any current legal proceedings, would you please give details?
I do not have any business or any financial holdings or any other commitments, which might conflict with my prospective duties.
During my entire working period I have worked only in State Administration and State Bodies.
Since April 2003 I have been a Member of the Auditing Board of the Council of Europe Development Bank (CEB).
I was appointed to this position by the Bulgarian Government and by the CEB Authorities for a 3-year-mandate, which will end in March 2007.
All my prospective commitments consist of not more than one week work in Paris until the end of my mandate.
It is no problem for me to terminate my mandate immediately.
I am absolutely ready to disclose all my financial interests to the President of the Court and to make them public at any time.
I am not involved in any current legal proceedings.
6.
Are you prepared to step down from any elected office and to give up any active function with responsibilities in a political party after your appointment as Court Member?
Yes, I do.
I do not have any such appointments.
I have never been a member of any political party nor have I ever had any active functions with political responsibilities.
7.
How would you deal with a major irregularity or even fraud and/or corruption case involving actors in the Member State of your origin?
No matter what the origin of the actor is, I would always strictly follow the auditing standards with all my respect to the equal rights and obligations of each Member State, taking into account all existing Treaty regulations concerning dealing with protection of the financial interests of the Community against irregularities, fraud and corruption.
In cases of potential fraud, I will follow the procedures described in ECA’s decision 97/2004 and other rules of the Court, which relate to internal investigations.
I would adopt a neutral position irrespective of the country in which an audit or investigation is taking place.
I will do my best to deal with the cases without being influenced by my own origin.
PERFORMANCE OF DUTIES
8.
What should be the main features of a sound financial management culture in any public service?
Sound financial management culture in a public service, whether belonging to the Community or not, in my opinion should be a management culture plus high quality management systems, which can provide the necessary guarantees that resources are used in the best possible way.
Within such systems there must be an unambiguous allocation of responsibilities in relation to the implementation of policies and programs, as well as the achievement of clearly defined objectives.
The classical principles of good financial management are economy, effectiveness and efficiency.
As the most important main features of a sound financial management culture should be mentioned:
1.Those suitable for within the bodies – clearly defined objectives, accountability, high quality of information and internal communication systems, precise definition of the competences and responsibilities (based on written internal rules), improvement of the management capacity, active human resources management, good communication between different levels in the management structure, efficient internal control and internal audit systems, etc.
2.
Those suitable for between the bodies – effective information and communication system, preventing overlaps in function and responsibilities, clear legal framework, etc.
3.
Those suitable for guaranteeing the quality of the management systems – availability of effective external audit, well-defined interaction between internal control, internal audit and external audit, transparency, quality of reporting, etc.
The modern sound financial management culture should use the instruments of prevention and risk analysis and should be able to improve and to develop itself in accordance to the fast changing environment.
9.
In its last Monitoring Report on Romania and Bulgaria, the Commission indicates delays in these countries’ administrations in setting up proper systems of financial control, including ex-ante control, independent internal and external audit.
What measures should receive priority?
In the last Monitoring Report on Bulgaria it is said “In the area of financial control, progress has been made with regard to the extended Decentralised Implementation System (EDIS) accreditation process for some of the structures concerned although efforts at capacity building for implementing the Structural Funds in particular need to be reinforced.
However, no accreditation has taken place yet”.
In the last Monitoring Report (September 2006), the only finding related to Bulgaria is the delay in the implementation and harmonization of EDIS.
But Bulgaria currently faces the following challenges.
These are the challenges in the area which require proper measures in the near future:
- Implementation of the newly adopted laws on financial management and control and internal audit in the public sector.
Till this moment it has led to great structural changes in the public bodies which have to follow the new requirements and to improve the quality of the internal control.
In all ministries which will conduct operational programmes, special training and a preparation are going on.
There is a special support and advisory activities provided by SIGMA.
- Guaranteeing the independence of the NAO in the Constitution and the focus on performance audits as a key factor for public funds management.
In the existing Constitution the independence of the NAO is not formulated well enough.
The NAO has not the power to control the state-owned enterprises and this limits its capacity to audit the use of money till the end beneficiaries.
The NAO should initiate changes in its Act aiming to extend its audit field.
Concerning performance audit and the implementation of its results, the NAO can activate its relationships with the Budgetary Commission in Parliament.
- Developing the CHU as a driver of the changes in the PIFC system, further implementation of the concept of financial management and control,
better understanding of the principle of management accountability by the managers in the public sector.
- Increased support by managers to the newly established internal audit functions.
The managers should take measures to optimize the internal institutional conditions in order to ensure the functioning of the new internal control’s responsibilities.
They should apply strong criteria concerning the professional abilities of the internal control staff.
- Establishment of External Audit Committees in the public sector organizations in order to strengthen the independence of the internal audit function.
These Audit Committees can provide external assurance as to the quality and the independence of the internal control activities.
10.
According to the Treaty the Court shall assist Parliament in exercising its powers of control over the implementation of the budget.
How would you describe your duties with regard to reporting to the European Parliament and its Committee on Budgetary Control, in particular?
As a member of the European Court of Auditors I can only answer that I will strictly follow the Treaty and the rules by assisting Parliament in exercising its powers of control over the implementation of the budget.
But based on my professional experience related to the Reporting of the Bulgarian National Audit Office to the Parliament, I can underline some points in the relationships between both of them, as it follows:
- it is very important that the reports and the opinions of the Audit Office are materially accurate , based on adequate, relevant and reliable information and at the same time they are understandable;
- the rapporteur - the member of the Audit Office must be capable to explain and to discuss all findings and recommendations in the report with the Members of the Budgetary Commission and must be able to answer all their questions in an atmosphere of mutual respect.
- in my opinion it was a good practice in Bulgaria to have regular meetings with the Budget Commission.
These meetings gave us the opportunity to discuss some very important topics concerning the budgetary legislation and spending the budget money in some particular areas.
In general, my understanding is that the most efficient way to assist Parliament, no matter which it is, in exercising its powers of control over the implementation of the budget is to work in dialogue and cooperation developing a culture of mutual trust and respect.
11.
What do you think is the added value of performance audit and how should the findings be incorporated in the management?
According to the Financial Regulation, EU funds should be managed based on the principles of economy, efficiency and effectiveness.
The European Court of Auditors carries out performance audits on important and specific topics and based on their results presents special reports to the Commission on Budgetary Control.
Performance audit is a modern tool to assess whether public funds have been used with economy, efficiency and effectiveness.
We could say that this type of audit is a huge step forward in the development and contribution of control.
It is the first to go beyond the tradition and practice of merely reviewing the accounts and the quality of the financial records of the underlying transactions.
On the one hand, performance audit provides taxpayers with a clear assessment of how and on what their money has been spent.
On the other hand, as a new audit technique it can largely contribute to improving the management of public institutions and to reducing the risks of public resources being spent in an ineffective way.
The Bulgarian National Audit Office (BNAO) has been applying the techniques of performance auditing since the year 2000 and has in practice materialised its positive impact.
For this accomplishment, the BNAO is particularly grateful to the UK National Audit Office for providing training of audit staff for the applying of this new type of audit in Bulgaria through a 2-year Twinning project.
Carrying our performance audit is a challenging task.
The difficulties are rooted primarily in the fact that the results are dependent on the auditors’ professional judgment; it is not always possible to quantify the findings.
In contrast to financial audit, there are no standardised audit criteria set be legislation and regulation, suitable for all audits.
Instead, unique criteria need to be developed for each individual audit.
I would like to point out several very important principles that should be observed if auditors are to add value by this type of audit, and that the findings and recommendations serve as a basis for improving the management of public institutions.
These are:
· The auditors should be knowledgeable about the nature and the activity of the audited entity, i.e. this entails tolerance during the audit and full understanding of the subject matter;
· The criteria for risk assessment, evaluation of the internal controls and measuring the effectiveness should be developed jointly and in agreement with the auditee;
· The audit findings should be formulated in an atmosphere of understanding and tolerance together with the auditee’s management, and should be fully supported with evidence and not solely with analytical considerations;
· The recommendations should also be discussed in advance and correctly understood by the auditee in order to guarantee their positive impact.
If such a complex subject matter could be summed up, two major principles would be outlined: the better formulated the objectives are, the easier the auditor’s work would be.
And last but not least, if performance audit is to reach its objectives, it should be viewed as a dialogue, as a sign of sound financial management.
12.
How could the cooperation improve between the Court of Auditors, the National Audit Institutions and the European Parliament (Committee on Budgetary Control) concerning the audit of the EU budget?
I know that this question is high on the EU agenda.
I will try to answer it using my experience and my knowledge of the statutory requirements, the procedures and standards of audit of the EU budget.
1.
According to the Treaty, only the European Court of Auditors (ECA) has the power to give an independent opinion on the financial statements and to report on issues of sound financial management and to provide an annual statement of assurance (DAS) on the legality and regularity of the transactions underlying the accounts as well as on the reliability of the accounts.
The national Supreme Audit Institutions (SAIs) are the external audit bodies which fulfill their mandates by their respective constitutions and report to the National Parliaments.
There is no shared responsibility for the audit of the EU budget between the European Court of Auditors and the SAIs.
2.
I think that the question concerns the future development of the whole control system at the European level.
Undoubtedly the following principles should be achieved: “a number of conditions must be met to set up a model where one level of control feeds the next level”, clear legislation and definition of rules and responsibilities, and efficiency which balances between cost and benefit.
3.
The Treaty states that the European Court of Auditors and the Supreme Audit Institutions of the Member States are to co-operate in a spirit of trust while maintaining their respective independence.
In his speech at the ECOFIN Council, Brussels, 7 November, 2006, Mr.
Hubert Weber, President of the European Court of Auditors said that “the Court remains committed to continuing its close cooperation with the national audit bodies of the European Union.
In practice this entails operational support for the Court’s on-the-spot audits, the exchange of professional information and knowledge, the joint development of practical and technical support.”
Having in mind the existing statutory requirements and the fact the over 76% of the European money is being managed by the national administrations in the Member States, and that the Court’s 2005 Annual Report on the implementation of the EU budget contains yet again a substantially critical opinion on its implementation in the part of the legality and regularity of underlying transactions in majority of EU expenditure under shared management .
I consider the following appropriate.
1.
The national supreme audit institutions should contribute, in a most effective way, to the reforming and development of the financial management and internal control systems in their countries; acquire powers and sufficient experience to audit EU funds so as to act as a guarantor of their proper implementation.
For example, in 2003, an audit department specialised in audits of pre-accession funds was set up in the Bulgarian National Audit Office.
The results of these audits are reported to the Bulgarian Parliament, following which they are sent to the ECA for information.
2.
The ECA, within the Contact Committee of the Heads of SAIs of the EU Member States, to continue its support for the MS SAIs in several very important aspects:
· Methodological and technical support with a view to improving the quality of external audit in the EU field; ability of the MS SAIs to produce national SAI reports on the management of EU funds to be presented to the national parliaments;
· Systematic support so that the management systems in the Member States are able to provide adequate and reconciled data in respect of the spending of the European budgetary funds.
According to “Redesigning accountability structures and control activities in the EU”, a draft working document of 07.09.2006, Committee on Budgetary Control: “Qualified information can only be provided if audits are carried out according to standards jointly developed by the Commission and the national audit institutions.”
It would be beneficial if the ECA would support this process.
· Creation of legal and practical possibilities for carrying our joint audits in the critical areas.
I have experience in such an audit and am convinced that this form of co-operation is particularly effective.
It is likely that my thoughts on the subject do not cover all possible measures.
Practice will always be a richer and truer basis for taking the correct management decisions on the basis of a dialog between the relevant authorities.
OTHER QUESTIONS
13.
Would you withdraw your candidacy if Parliament’s opinion on your appointment as Member of the Court were unfavourable?
Taking into account that this hearing, as a part of the adoption procedure, has a very important role to guarantee my professional abilities and their compatibility with the criteria of holding a post, if the Parliament’s opinion is unfavourable I would immediately withdraw my candidacy.
ÄRENDETS GÅNG
Titel
Nominering av Nadezhda Sandolova till uppdraget som ledamot av revisionsrätten
Referensnummer
C6‑0411/2006 – 2006/0811(CNS)
Begäran om samråd med parlamentet
7.11.2006
CONT 29.11.2006
José Javier Pomés Ruiz 23.10.2006
Behandling i utskott
28.11.2006
Antagande
28.11.2006
Slutomröstning: närvarande ledamöter
Inés Ayala Sender, Herbert Bösch, Paul van Buitenen, Simon Busuttil, Mogens N.J. Camre, Paulo Casaca, Szabolcs Fazakas, Markus Ferber, Christofer Fjellner, Ingeborg Gräßle, Ona Juknevičienė, Rodi Kratsa-Tsagaropoulou, Dan Jørgensen, Nils Lundgren, Edith Mastenbroek, Jan Mulder, José Javier Pomés Ruiz, Brian Simpson, Bart Staes, Kyösti Virrankoski
Slutomröstning: närvarande suppleanter
Daniel Caspary, Bárbara Dührkop Dührkop, Salvador Garriga Polledo, Edit Herczog, Eija-Riitta Korhola, Albert Jan Maat, Ashley Mote
Slutomröstning: närvarande suppleanter (art.
178.2)
Toine Manders
Ingivande
30.11.2006
Anmärkningar (tillgängliga på ett enda språk)
SLUTLIG VERSION
A6-0067/2007
om Kosovos framtid och EU:s roll
(2006/2267(INI))
Utskottet för utrikesfrågor
Föredragande:
Joost Lagendijk
PE 384.211v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
YTTRANDE FRÅN UTSKOTTET FÖR INTERNATIONELL HANDEL...............................12
ÄRENDETS GÅNG..................................................................................................................15
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om Kosovos framtid och EU:s roll
( 2006/2267(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av resolution 1244 från Förenta nationernas säkerhetsråd av den 10 juni 1999,
– med beaktande av rapporten från den särskilda representanten för FN:s generalsekreterare om en omfattande översyn av hur standarderna genomförs, framlagd inför FN:s säkerhetsråd den 7 oktober 2005,
– med beaktande av FN:s säkerhetsråds beslut av den 24 oktober 2005 om att stöda generalsekreterarens förslag om att inleda samtal om Kosovos status,
– med beaktande av utnämningen den 14 november 2005 av Martti Ahtisaari till Förenta nationernas generalsekreterares särskilda sändebud för processen avseende Kosovos framtida status,
– med beaktande av kontaktgruppens slutsatser av den 31 januari 2006 där det understryks att problemet Kosovo är speciellt till sin karaktär – vilket enligt dessa slutsatser beror på Jugoslaviens upplösning och de därpå följande konflikterna, den etniska rensningen och händelserna 1999 samt den långa perioden av internationell förvaltning i enlighet med säkerhetsrådets resolution 1244 (1999) – och där en snabb förhandlingslösning på frågan efterlyses som bästa väg att följa,
– med beaktande av ordförandeskapets slutsatser från Europeiska rådets möte den 14‑15 december 2006 som fullt ut ställer sig bakom Ahtisaaris ansträngningar att finna en lösning på dödläget och som bekräftar unionens beredskap att spela en viktig roll när den framtida lösningen skall förverkligas,
– med beaktande av det särskilda sändebudets slutrapport/rekommendationer om ... av den....,
– med beaktande av artikel 45 i arbetsordningen,
– med beaktande av betänkandet från utskottet för utrikesfrågor och yttrandet från utskottet för internationell handel ( A6‑0067/2007 ), och av följande skäl:
C. Händelserna i mars 2004 måste fördömas men visar att spänningarna mellan de albanska och serbiska samfunden i Kosovo lever kvar och att det är nödvändigt att finna en lösning som garanterar dessa båda folkgruppers och andra etniska gruppers rättigheter, såsom framgår av publikationer från OSSE, Europarådet och andra organisationer som bedriver verksamhet för att skydda minoriteter.
D. Ett avgörande i frågan om Kosovos framtida status kommer att bidra till utvecklingen av dess ekonomi och framväxten av en mogen politisk kultur och ett tolerant samhälle utan segregering.
F. Den slutliga lösningen kan inte dikteras av hot om en radikalisering i Kosovo eller i Serbien utan måste vara resultatet av en lösning som beaktar alla berörda parters intressen.
G. Ytterligare dröjsmål med att fastställa Kosovos status kan få negativa konsekvenser för den känsliga och spända situation som redan råder.
H. Händelserna 1999, den långvariga internationella interimsförvaltningen samt utvecklingen och den gradvisa konsolideringen av Kosovos interimsinstitutioner för självstyre har skapat en mycket speciell situation som gör tanken på att Kosovo på nytt skulle införlivas med Serbien föga realistisk.
I. Förbindelserna mellan Kosovo och Serbien utmärks av att de kulturella, religiösa och ekonomiska banden mellan dem är intima och därför bör de vidareutvecklas i en anda av partnerskap och god grannsämja, vilket ligger i hela Kosovos och Serbiens befolknings intresse.
J. Bristen på förtroende mellan olika etniska grupper, den labila situation som fortsättningsvis råder och behovet av att vidareutveckla och befästa demokratiska multietniska institutioner i Kosovo kräver en fortsatt internationell närvaro under överskådlig framtid.
K. Det internationella samfundet bör fortsätta att investera i utbildningssystemet, särskilt i ljuset av de stora utmaningar som den yngre generationen i Kosovo står inför.
L. Med tanke på Kosovos strategiska läge måste Europeiska unionen spela en central roll när det gäller att övervaka, garantera och underlätta genomförandet av en lösning på frågan om Kosovos status samt bistå vid inrättandet och konsolideringen av demokratiska institutioner i Kosovo, varvid Europaparlamentet påtar sig ett övervakningsansvar.
M. EU:s bidrag måste emellertid göras beroende av att vissa minimikrav i överenskommelsen uppfylls.
N. Lösningen på frågan om den slutgiltiga statusen måste överensstämma med EU:s principer, det vill säga förutse en konstitutionell ram som är förenlig med Kosovos europeiska perspektiv och tillåta unionen att fullt ut utnyttja de instrument som står till förfogande.
– ger Kosovo tillgång till internationella finansorganisationer och således möjlighet till ekonomisk återhämtning och till att skapa förutsättningar för att inrätta arbetstillfällen,
– förutser en internationell närvaro för att upprätthålla Kosovos mångetniska karaktär och tillvarata den serbiska befolkningsgruppens och romerbefolkningens samt andra etniska gruppers intressen och säkerhet,
– tillhandahåller internationellt stöd för att utveckla effektiva och oberoende institutioner för hela Kosovos befolkning, vilka fungerar i överensstämmelse med rättsstatsprincipen och de demokratiska grundreglerna,
– förverkliga Kosovos önskan om att integreras i Europa, vilket med tiden kommer att göra det möjligt för landet att med sina grannländer ingå ett ömsesidigt beroende.
– en klar definition av rollen och uppdraget för den internationella civila och säkerhetsrelaterade närvaron,
– klara bestämmelser om decentralisering som garanterar väsentlig autonomi inom nyckelområden som utbildning, hälsa och lokal säkerhet och, när det gäller de serbiska kommunerna, tillåter direkta men transparenta förbindelser med Belgrad; dessa bestämmelser måste vara ekonomiskt hållbara och får inte underminera ett enhetligt Kosovos budgetära, verkställande och lagstiftningsmässiga privilegier,
– full respekt för de mänskliga rättigheterna, däribland en skyldighet att i författningen säkerställa minoriteters och flyktingars vitala intressen samt adekvata mekanismer för att tillvarata dessa intressen,
– skydd av alla kulturella och religiösa platser,
– bestämmelser om inrättandet av en lättutrustad, multietnisk intern säkerhetsstyrka för Kosovo, vars verksamhets räckvidd, möjligheter och funktioner är begränsade och som verkar under strikt övervakning av den Natoledda Kosovostyrkan Kfor,
– internationella garantier för att alla grannstaters territoriella integritet respekteras.
Europaparlamentet välkomnar därför det faktum att Ahtisaaris förslag innebär en omfattande autonomi för serbiska och andra samfund, inklusive en vittgående kommunal autonomi i linje med europeiska principer om subsidiaritet och självstyre.
– genomföra villkoren för lösningen,
– utveckla en autonom, etniskt balanserad, institutionell, administrativ, juridisk och politisk kapacitet,
– göra framsteg när det gäller att efterleva FN:s standarder och EU:s riktmärken för stabilisering och associering.
Europaparlamentet understryker att det internationella samfundet måste ha direkta befogenheter att vidta korrigerande och, i vissa fall, ställföreträdande åtgärder, bland annat på följande viktiga områden
– skydd av minoriteters livsviktiga intressen,
– beskydd av känsliga platser,
– säkerhet,
– rättsväsendet och rättsutövningen i vidare mening, särskilt i kampen mot organiserad brottslighet.
Europaparlamentet uppmärksammar behovet av ett rättvist utbildningssystem som är tillgängligt för alla och som ser till att romiska och ashkali elever undervisas delvis på sitt modersmål för att på detta sätt stärka dessa minoritetsgruppers identitet och kultur.
Europaparlamentet är berett att ställa de kompletterande resurser till förfogande som krävs för att finansiera EU:s framtida involvering i Kosovo i syfte att förverkliga lösningen om Kosovos status och stöda Kosovos EU-perspektiv, detta under förutsättning att
– den lösning av statusfrågan som stöds av FN:s säkerhetsråd vederbörligen tar hänsyn till unionens gemensamma ståndpunkt,
– tillräckligt samråd äger rum på förhand avseende räckvidden, målen, medlen och formaliteterna för ett sådant uppdrag, så att parlamentet tillförsäkras om att resurserna står i proportion till uppgifterna,
– de kompletterande finansiella resurserna beviljas i enlighet med villkoren i det interinstitutionella avtalet om budgetdisciplin och sund ekonomisk förvaltning av den 14 juni 2006
EUT C 139, 14.6.2006, s.
1. , och
– utveckling av ett kosovanskt medborgarskapsbegrepp som uttryckligen utgår från regionens flerspråkiga och multietniska karaktär och som samtidigt ger fullt erkännande åt de olika folkgrupper som tillsammans utgör Kosovos befolkning,
– allvarligt och konstruktivt arbete för att skapa ett multietniskt, mångkulturellt, mångreligiöst och tolerant land och samhälle där samtliga etniska gruppers rättigheter respekteras.
27.
Europaparlamentet upprepar att stabiliserings- och associeringsprocessen bland annat kommer att stärka Kosovos ekonomiska förbindelser med medlemsstaterna och med landets grannar på västra Balkan och underlätta stabiliseringsprocessen i regionen.
37.
39.
YTTRANDE FRÅN UTSKOTTET FÖR INTERNATIONELL HANDEL
till utskottet för utrikesfrågor
över Kosovos framtid och EU:s roll
( 2006/2267(INI) )
Föredragande:
Erika Mann
FÖRSLAG
Utskottet för internationell handel uppmanar utskottet för utrikesfrågor att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet påminner om att en lyckosam utgång av den reformprocess som nu pågår kommer att få marknaden att fungera väl igen, stimulera ekonomisk tillväxt och bidra till att vidmakthålla den politiska stabiliteten i regionen.
ÄRENDETS GÅNG
Titel
Kosovos framtid och EU:s roll
Referensnummer
2006/2267(INI)
Ansvarigt utskott
AFET
Behandling i utskott
Antagande
26
Francisco Assis, Jean-Pierre Audy, Enrique Barón Crespo, Daniel Caspary, Christofer Fjellner, Béla Glattfelder, Jacky Henin, Syed Kamall, Sajjad Karim, Erika Mann, David Martin, Javier Moreno Sánchez, Caroline Lucas, Georgios Papastamkos, Peter Šťastný, Robert Sturdy, Gianluca Susta, Johan Van Hecke, Zbigniew Zaleski
Slutomröstning: närvarande suppleanter
Panagiotis Beglitis, Małgorzata Handzlik, Jens Holm, Jörg Leichtfried, Eugenijus Maldeikis
Slutomröstning: närvarande suppleanter (art.
178.2)
Ignasi Guardans Cambó, Pia Elda Locatelli
Anmärkningar (tillgängliga på ett enda språk)
ÄRENDETS GÅNG
Titel
Kosovos framtid och EU:s roll
Förfarandenummer
2006/2267(INI)
Ansvarigt utskott Tillstånd: tillkännagivande i kammaren
Föredragande Utnämning
Behandling i utskott
Antagande
+:
–:
56
7
3
Slutomröstning: närvarande ledamöter
Roberta Alma Anastase, Christopher Beazley, Angelika Beer, Panagiotis Beglitis, Bastiaan Belder, André Brie, Véronique De Keyser, Giorgos Dimitrakopoulos, Hélène Flautre, Hanna Foltyn-Kubicka, Michael Gahler, Jas Gawronski, Bronisław Geremek, Maciej Marian Giertych, Ana Maria Gomes, Klaus Hänsch, Jelko Kacin, Ioannis Kasoulides, Bogdan Klich, Joost Lagendijk, Vytautas Landsbergis, Emilio Menéndez del Valle, Willy Meyer Pleite, Francisco José Millán Mon, Pasqualina Napoletano, Annemie Neyts-Uyttebroeck, Raimon Obiols i Germà, Cem Özdemir, Janusz Onyszkiewicz, Justas Vincas Paleckis, Alojz Peterle, Tobias Pflüger, Bernd Posselt, Raül Romeva i Rueda, Libor Rouček, Katrin Saks, José Ignacio Salafranca Sánchez-Neyra, Jacek Saryusz-Wolski, György Schöpflin, István Szent-Iványi, Antonio Tajani, Charles Tannock, Josef Zieleniec
Slutomröstning: närvarande suppleant(er)
Laima Liucija Andrikienė, Maria Badia I Cutchet, Giulietto Chiesa, Ryszard Czarnecki, Alexandra Dobolyi, Árpád Duka-Zólyomi, Glyn Ford, Lilli Gruber, Tunne Kelam, Evgeni Kirilov, Jaromír Kohlíček, Antonio López-Istúriz White, Sarah Ludford, Erik Meijer, Doris Pack, Antonyia Parvanova, Lapo Pistelli, Frédérique Ries, Aloyzas Sakalas, Anders Samuelsen, Adrian Severin, Csaba Sándor Tabajdi
Slutomröstning: närvarande suppleant(er) (art.
178.2)
Miloš Koterec
Ingivande
SLUTLIG VERSION
A6-0078/2007
*
BETÄNKANDE
om förslaget till rådets beslut om ändring av beslut 2004/585/EG om inrättande av regionala rådgivande nämnder inom ramen för den gemensamma fiskeripolitiken
(KOM(2006)0732 – C6‑0051/2007 – 2006/0240(CNS))
Fiskeriutskottet
Föredragande:
Elspeth Attwooll
PE 384.344v03-00
Teckenförklaring
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING............................................................................................................................6
ÄRENDETS GÅNG....................................................................................................................7
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till rådets beslut om ändring av beslut 2004/585/EG om inrättande av regionala rådgivande nämnder inom ramen för den gemensamma fiskeripolitiken
( KOM(2006)0732 – C6‑0051/2007 – 2006/0240(CNS) )
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till rådet ( KOM(2006)0732 )
Ännu ej offentliggjort i EUT. ,
– med beaktande av artikel 37 i EG-fördraget, i enlighet med vilken rådet har hört parlamentet ( C6‑0051/2007 ),
– med beaktande av artikel 51 i arbetsordningen,
– med beaktande av betänkandet från fiskeriutskottet ( A6‑0078/2007 ).
MOTIVERING
Kommissionens förslag syftar till att ge arbetet inom de regionala rådgivande nämnderna en bättre grund genom att förbättra villkoren för finansieringen av dem.
Detta skall genomföras på så sätt att nämnderna integreras i budgeten, vilket innebär a) att gemenskapens bidrag inte längre behöver minskas successivt och b) att de omfattas av en enda redovisningsmetod i stället för av två separata metoder som för närvarande.
Förslaget är mycket välkommet.
Parlamentet har konsekvent stött ett ökat engagemang av parterna i utvecklingen av den gemensamma fiskeripolitiken.
Det tillstyrkte principen om regionaliserade insatser i beslutsprocessen i sin resolution från 2001 om kommissionens grönbok om den framtida gemensamma fiskeripolitiken
Betänkande av Ó Neachtain, 2003/0238(CNS) , ( KOM(2003)0607 ), EUT L 256, 3.8.2004, s.
17–22. .
I det senare dokumentet, liksom vid flera andra tillfällen därefter, efterlyste parlamentet emellertid en finansieringsnivå och en finansieringsmetod som är tillräckliga för att nämnderna skall kunna fungera effektivt och kontinuerligt.
För närvarande fungerar fyra av de sju planerade regionala rådgivande nämnderna fullt ut, medan de övriga sannolikt kommer att tas i bruk inom en nära framtid.
Dessutom har en gemensam kommitté inrättats för att samordna nämndernas verksamhet.
Kommissionen har mottagit rekommendationer och råd vid mer än 80 tillfällen, och de regionala rådgivande nämnderna har även gett ett värdefullt bidrag till diskussionerna inom parlamentets fiskeriutskott.
Åtgärder bör således vidtas för att säkra nämndernas finansiella bärkraft på lång sikt.
För att undvika osäkerhet bör man ange att förslaget inte inverkar på några andra aspekter av de regionala rådgivande nämndernas sammansättning och arbete.
Detta kommer att bli föremål för en översyn som offentliggörs senare i år, vilket fiskeriutskottet motser med intresse.
ÄRENDETS GÅNG
Titel
Ändring av beslut 2004/585/EG om inrättande av regionala rådgivande nämnder inom ramen för den gemensamma fiskeripolitiken
Referensnummer
KOM(2006)0732 – C6-0051/2007 – 2006/0240(CNS)
Begäran om samråd med parlamentet
19.1.2007
Ansvarigt utskott
Tillkännagivande i kammaren
PECH
1.2.2007
Rådgivande utskott
Tillkännagivande i kammaren
BUDG
1.2.2007
Inget yttrande avges
Beslut
BUDG
14.2.2007
Föredragande
Utnämning
Elspeth Attwooll
9.1.2007
Behandling i utskott
25.1.2007
27.2.2007
Antagande
22.3.2007
Slutomröstning: resultat
+:
–:
0:
26
1
Slutomröstning: närvarande ledamöter
Jim Allister, Alfonso Andria, Stavros Arnaoutakis, Elspeth Attwooll, Marie-Hélène Aubert, Iles Braghetto, Luis Manuel Capoulas Santos, Paulo Casaca, Zdzisław Kazimierz Chmielewski, Emanuel Jardim Fernandes, Carmen Fraga Estévez, Duarte Freitas, Ioannis Gklavakis, Pedro Guerreiro, Ian Hudghton, Heinz Kindermann, Rosa Miguélez Ramos, Marianne Mikko, Philippe Morillon, Seán Ó Neachtain, Willi Piecyk, Struan Stevenson, Catherine Stihler, Daniel Varela Suanzes-Carpegna
Slutomröstning: närvarande suppleanter
Vincenzo Aita, Ole Christensen, Jan Mulder, Thomas Wise
Ingivande
27.3.2007
SLUTLIG VERSION
A6-0082/2007
*
BETÄNKANDE
om förslaget till rådets beslut om anpassning av bestämmelserna om domstolen på de områden som omfattas av avdelning IV i tredje delen av fördraget om upprättandet av Europeiska gemenskapen
(KOM(2006)0346 – C6‑0304/2006 – 2006/0808(CNS))
Utskottet för rättsliga frågor
Föredragande:
József Szájer
PE 382.638v03-00
Teckenförklaring
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING............................................................................................................................6
ÄRENDETS GÅNG....................................................................................................................9
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till rådets beslut om anpassning av bestämmelserna om domstolen på de områden som omfattas av avdelning IV i tredje delen av fördraget om upprättandet av Europeiska gemenskapen
( KOM(2006)0346 – C6‑0304/2006 – 2006/0808(CNS) )
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
– med beaktande av förslaget till rådets beslut, som utgör en bilaga till kommissionens meddelande ( KOM(2006)0346 – C6-0304/2006 ),
– med beaktande av artikel 51 i arbetsordningen,
– med beaktande av betänkandet från utskottet för rättsliga frågor ( A6‑0082/2007 ).
1.
Europaparlamentet begär att medlingsförfarandet enligt den gemensamma förklaringen av den 4 mars 1975 inleds om rådet har för avsikt att avvika från den text som parlamentet har godkänt.
MOTIVERING
Utvärdering
Enligt EG-domstolen är förhandsavgöranden ”av avgörande betydelse för att den genom fördraget tillkomna rätten behåller sin karaktär av gemenskapsrätt” och ”har som ändamål att under alla omständigheter säkerställa att denna rätt har samma verkan i alla gemenskapens stater
Mål 166/73 Rheinmühlen mot.
Artikel 234 ger EG-domstolen behörighet att meddela förhandsavgöranden beträffande tolkningen eller giltigheten av rättsakter som beslutats av gemenskapens institutioner.
När det gäller rättligt samarbete i civilrättsliga frågor sett ur utskottet för rättsliga frågors behörighetsperspektiv och i synnerhet internationell privaträtt, kan man konstatera att införlivandet av konventionerna i gemenskapslagstiftningen samt erkännandet och verkställigheten av domar i civil- och handelsrättsliga mål samt i äktenskapsmål enligt förordningarna nr 44/2001 och nr 1347/2000 utgör ett steg tillbaka i utvecklingen jämfört med de tidigare protokollen till dessa konventioner, som tilldelar lagstiftningsansvar för förhandsavgöranden även till appellationsdomstolar och inte enbart till domstolar som utgör högsta instans
Se Lenaerts, Arts, Maselis, Bray (ed.), Procedural Law of the European Union , Sweet & Maxwell, London, 2006, at 22-001. .
Artikel 67:
1.
Rådet skall under en övergångsperiod av fem år efter Amsterdamfördragets ikraftträdande besluta enhälligt på förslag av kommissionen eller på initiativ av en medlemsstat och efter att ha hört Europaparlamentet.
2.
Efter denna femårsperiod skall rådet.
- besluta på förslag av kommissionen; kommissionen skall pröva varje begäran från en medlemsstat om att kommissionen skall lägga fram ett förslag för rådet,
- efter att ha hört Europaparlamentet enhälligt besluta i syfte att låta alla eller delar av de områden som omfattas av denna avdelning regleras av förfarandet i artikel 251 och att anpassa bestämmelserna om domstolens behörighet. skall tillämpas för att göra artikel 68 otillämplig.
Således kan domstolen tillämpa standardbestämmelserna i artikel 234 utan att rätten att begära förhandsavgöranden begränsas enbart till domstolar i högsta instans.
Förslaget innebär att
· enhetlig tillämpning och tolkning av gemenskapslagstiftningen garanteras
· det rättsliga skyddet, på områden som är särskilt känsliga när det gäller grundläggande rättigheter, stärks
· den försvagning av rättskyddet, som Amsterdamfördraget medfört på det civilrättsliga området, som omfattas av artikel 65, kan åtgärdas
· gemenskapens rättssystem kan fungera normalt på detta område.
Rent konkret bidrar förslaget till att främja enhetlig tolkning och tillämpning av gemenskapslagstiftningen och en enhetlig ordning för rättsligt skydd inom de områden som omfattas av avdelning IV i EG-fördraget.
Tillämpas förfarandet för förhandsavgöranden fullt ut på avdelning IV skulle detta stärka det rättsliga skyddet för de berörda personerna.
För närvarande kan en person som anser att hans grundläggande rättigheter kränkts genom en gemenskapsakt, som antagits i enlighet med avdelning IV, enbart förelägga EG-domstolen ett ärende för förhandsavgörande om alla överklagandemöjligheter på det nationella planet uttömts dvs. att ärendet tagits upp i högsta instans.
Kostnaderna för ett sådant förfarande kan avskräcka många parter och därigenom kan rättssäkerheten komma att bli lidande.
Det är tveksamt om de nuvarande förhållandena är förenliga med unionens åligganden enligt Europakonventionen om skydd för de mänskliga rättigheterna.
Om förslaget antas kommer även nationella domstolar att i första instans kunna begära förhandsavgörande.
Det bör betonas att kommissionen har poängterat att det ökade antalet ärenden avseende begäran om förhandsavgöranden inom detta område inte kommer att öka domstolens arbete i orimlig omfattning om man litar till att de medel som avsatts för det interna arbetet och de nya möjligheter som skapas genom Nicefördraget, som påskyndat förfarandet
Vid tillämpning av påskyndat förfarande för meddelande av förhandsavgöranden kan domstolens ordförande i undantagsfall besluta, på begäran av den nationella domstolen och på förslag från den föredragande domaren och efter att generaladvokaten hörts, att det påskyndade förfarandet skall tillämpas då det kan konstateras i enlighet med nämnda omständigheter att beslut om en begäran som ställts till domstolen är ytterst brådskande.
Ordföranden fastställer omedelbart datumet för överläggningarna som meddelas alla berörda parter, som kan inge redogörelser i ärendet eller skriftliga synpunkter inom en tidsfrist på minst 15 dagar. , tillämpas på ett effektivt sätt.
Vidare föreslår domstolen att det införs en ny form av förfarande – ett påskyndat förfarande för förhandsavgöranden – som skulle möjliggöra att ett ärende behandlas ännu snabbare än vad som är fallet vid det påskyndade förfarandet.
Enligt detta förfarande skulle ärenden som kräver en ytterst snabb behandling kunna hänförs till en särskild instans som skulle tillämpa ett förenklat förfarande men med eventuell möjlighet till att ärendet behandlas på nytt.
Sammanfattning
Med hänvisning till ovanstående bör kommissionens förslag förordas och parlamentets begäran till rådet om att upphäva de begränsningar av EG-domstolens befogenheter som hänför sig till avdelning IV i fördraget återupprepas.
Se P6_TA-PROV(2006)0525 , Cavada. ”.
Det är nödvändigt att aktivera den övergångsklausul som avses i artikel 67 för att komma till rätta med de demokratiska brister som fortfarande präglar området för frihet, säkerhet och rättvisa och utvidga omfattningen av det rättsliga skyddet inom de känsliga områden som omfattas av avdelning IV i EG-fördraget med hänvisning till gemenskapsinstitutionernas växande befogenheter.
ÄRENDETS GÅNG
Titel
Anpassning av bestämmelserna i avdelning IV i EG-fördraget om domstolens behörighet
Referensnummer
KOM(2006)0346 - C6-0304/2006 - 2006/0808(CNS)
Begäran om samråd med parlamentet
20.9.2006
Ansvarigt utskott
Tillkännagivande i kammaren
JURI
28.9.2006
Rådgivande utskott
Tillkännagivande i kammaren
LIBE
28.9.2006
Inget yttrande avges
Beslut
LIBE
19.12.2006
Föredragande
Utnämning
József Szájer
2.10.2006
Behandling i utskott
27.2.2007
Antagande
20.3.2007
Slutomröstning: resultat
+:
–:
0:
26
Slutomröstning: närvarande ledamöter
Marek Aleksander Czarnecki, Cristian Dumitrescu, Monica Frassoni, Giuseppe Gargani, Klaus-Heiner Lehne, Katalin Lévai, Antonio Masip Hidalgo, Hans-Peter Mayer, Manuel Medina Ortega, Aloyzas Sakalas, Francesco Enrico Speroni, Rainer Wieland, Jaroslav Zvěřina, Tadeusz Zwiefka
Slutomröstning: närvarande suppleanter
Mogens N.J. Camre, Nicole Fontaine, Janelly Fourtou, Jean-Paul Gauzès, Eva Lichtenberger, Arlene McCarthy, Marie Panayotopoulos-Cassiotou, Michel Rocard, Gabriele Stauner, József Szájer, Jacques Toubon
Slutomröstning: närvarande suppleanter (art.
178.2)
Toine Manders
SLUTLIG VERSION
A6-0084/2007
BETÄNKANDE
om avtal om ekonomiskt partnerskap
(2005/2246(INI))
Utskottet för internationell handel
Föredragande:
Robert Sturdy
PE 376.650v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING..........................................................................................................................13
ÄRENDETS GÅNG..................................................................................................................17
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om avtal om ekonomiskt partnerskap
( 2005/2246(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av sina resolutioner av den 13 december 2001 om Europaparlamentets resolution om WTO:s möte i Qatar
EGT C 177 E, 25.7.2002, s.
290. , av den 25 september 2003 om WTO:s femte ministerkonferens i Cancún
EUT C 77 E, 26.3.2004, s.
393. , av den 12 maj 2005 om utvärderingen av Doharundan efter beslutet av WTO:s allmänna råd av den 1 augusti 2004
EUT C 92 E, 20.4.2006, s.
397. , av den 6 juli 2005 om en allmän uppmaning till kamp mot fattigdom: Förpassa fattigdomen till historien
EUT C 157 E, 6.7.2006, s.
397. , av den 1 december 2005 om förberedelserna inför WTO:s sjätte ministerkonferens i Hongkong
EUT C 285 E, 22.11.2006, s.
32. , av den 23 mars 2006 om utvecklingspåverkan av avtalen om ekonomiskt partnerskap
EUT C 292 E, 1.12.2006, s.
121. , av den 4 april 2006 om bedömningen av Doharundan efter WTO:s ministerkonferens i Hongkong
EUT C 293 E, 2.12.2006, s.
155. , av den 1 juni 2006 om handel och fattigdom: Utformning av en handelspolitik som maximerar handelns bidrag till fattigdomslindringen
Antagna texter, P6_TA(2006)0242 . samt av den 7 september 2006 om beslutet att tills vidare skjuta upp förhandlingarna om utvecklingsagendan från Doha
Antagna texter, P6_TA(2006)0350 . ,
– med beaktande av den gemensamma parlamentariska AVS­‑EG-församlingens resolution av den 23 november 2006, som antogs i Barbados, om översynen av förhandlingarna om avtalen om ekonomiskt partnerskap,
– med beaktande av förklaringen från Kapstaden som enhälligt antogs av den gemensamma parlamentariska AVS‑EU-församlingen den 21 mars 2002, och i vilken det uppmanas till inrättandet av riktmärken för utvecklingen som kan användas för att utvärdera hur handelsöverläggningarna mellan AVS och EU framskrider och deras resultat,
– med beaktande av deklarationen från 2006 års årliga parlamentariska konferens om WTO, vilken antogs den 2 december 2006 i Genève,
– med beaktande av sin ståndpunkt av den 9 mars 2005 om förslaget till rådets förordning om tillämpning av Allmänna preferenssystemet
EUT C 320 E, 15.12.2005, s.
145. ,
– med beaktande av rådets förordning (EG) nr 980/2005 av den 27 juni 2005 om tillämpning av Allmänna preferenssystemet
EUT L 169, 30.6.2005, s.
1. ,
– med beaktande av partnerskapsavtalet mellan medlemmarna i gruppen av stater i Afrika, Västindien och Stillahavsområdet, å ena sidan, och Europeiska gemenskapen och dess medlemsstater, å andra sidan, undertecknat i Cotonou den 23 juni 2000 (Cotonouavtalet),
– med beaktande av rådets (allmänna frågor och yttre förbindelser) slutsatser av den 10 och 11 april 2006 och den 16 oktober 2006 samt Europeiska rådets slutsatser av den 15 och 16 juni 2006,
– med beaktande av meddelandet från kommissionen till rådet, Europaparlamentet, Europeiska ekonomiska och sociala kommittén och regionkommittén med förslag till gemensam förklaring från rådet, Europaparlamentet och kommissionen: Europeiska unionens utvecklingspolitik – Dokument om europeiskt samförstånd ( KOM(2005)0311 ),
– med beaktande av kommissionens arbetsdokument med titeln ”Handels‑ och utvecklingsaspekter av EPA‑förhandlingarna” ( SEK(2005)1459 ),
– med beaktande av allmänna tull‑ och handelsavtalet (GATT), särskilt dess artikel XXIV,
– med beaktande av förklaringen från WTO:s fjärde ministerkonferens, som antogs den 14 november 2001 i Doha,
– med beaktande av beslutet i WTO:s allmänna råd av den 1 augusti 2004,
– med beaktande av förklaringen från WTO:s sjätte ministerkonferens, som antogs den 18 december 2005 i Hongkong,
– med beaktande av rapporten och rekommendationerna från arbetsgruppen för handelsrelaterat bistånd, som antogs av WTO:s allmänna råd den 10 oktober 2006,
– med beaktande av Sutherlandrapporten om WTO:s framtid,
– med beaktande av FN:s millenniedeklaration av den 8 september 2000, i vilken millennieutvecklingsmålen formuleras som kriterier vilka kollektivt upprättats av det internationella samfundet för att utrota fattigdomen,
– med beaktande av resultaten från FN:s världstoppmöte 2005,
– med beaktande av rapporten ”Investing in Development: A Practical Plan to Achieve the Millennium Development Goals” från FN:s arbetsgrupp för millennieprojektet som letts av professor Jeffrey Sachs,
– med beaktande av kommunikén av den 8 juli 2005 från G8‑mötet i Gleneagles,
– med beaktande av rapporten från FN:s konferens för handel och utveckling (UNCTAD) – ”Least Developed Countries 2006: Developing Productive Capacities”,
– med beaktande av den ekonomiska rapporten om Afrika 2004 ”Unlocking Africa’s Trade Potential” från FN:s ekonomiska kommission för Afrika,
– med beaktande av AVS riktlinjer för förhandlingarna om avtalet om ekonomiskt partnerskap, vilka antogs av AVS ministerråd den 27 juni 2002 i Punta Cana (Dominikanska republiken), och beslutet om förhandlingarna om ekonomiska partnerskap och deltagande i det internationella handelssystemet, som antogs vid det tredje toppmötet med stats‑ och regeringscheferna i AVS den 19 juli 2002 i Nadi (Fiji),
– med beaktande av deklarationen från det fjärde toppmötet med stats‑ och regeringscheferna för AVS‑länderna den 23–24 juni 2004 i Maputo, Moçambique, med avseende på den ekonomiska utvecklingsdimensionen,
– med beaktande av deklarationen från det 81:a sammanträdet med AVS‑ministerråd i Bryssel den 21–22 juni 2005,
– med beaktande av beslut nr 2/LXXXIII/06 från det 83:e sammanträdet med AVS‑ministerråd i Port Moresby (Papua Nya Guinea) den 28–31 maj 2006,
– med beaktande av deklarationen från det femte toppmötet med stats‑ och regeringscheferna i AVS‑länderna i Khartoum (Sudan) den 8 december 2006,
– med beaktande av artikel 45 i arbetsordningen,
– med beaktande av betänkandet från utskottet för internationell handel ( A6‑0084/2007 ), och av följande skäl:
A. EU:s nuvarande handelsförbindelser med AVS‑länderna – som ger dem förmånstillträde till EU:s marknader på icke‑ömsesidig grund – uppfyller inte Världshandelsorganisationens (WTO) regler.
B. I Cotonouavtalet beskrivs parternas överenskommelse om att ingå nya WTO-kompatibla handelsarrangemang, successivt avlägsna handelshinder mellan sig och fördjupa samarbetet inom alla områden som är relevanta för handeln och utvecklingen.
C. Förhandlingarna går inte framåt i samma takt i de sex regionerna, vilket leder till oro för att de inte kommer att slutföras i alla regioner före 2007 års utgång.
D. Det finns en utbredd oro för att förhandlingarna inte har avancerat så långt som de borde ha gjort vid detta skede i förhandlingsprocessen.
E. En viktig orsak till dröjsmålet har varit att båda sidor har misslyckats med att lägga fram och svara på förslag i tid.
F. Ännu ett formellt WTO‑undantag skulle vara politiskt kostsamt och svårt att uppnå.
G. I många AVS‑länder har informationen om och involveringen i processen för avtal om ekonomiskt partnerskap på landsnivå varit oroväckande låg.
H. Bristen på framsteg i förhandlingarna om utvecklingsagendan från Doha i WTO försvårar förhandlingarna om avtal om ekonomiskt partnerskap.
I. Båda parterna är överens om att ”utvecklingsdimensionen” är central för avtal om ekonomiskt partnerskap, men förhandlarna har hittills inte lyckats komma överens om en gemensam definition av begreppet.
J. Det är mycket viktigt att avtalen om ekonomiskt partnerskap bidrar till en hållbar social och ekonomisk utveckling och lindring av fattigdomen i AVS‑länderna.
K. I en allt mer globaliserad värld är det oundvikligt att handelsförmånerna urholkas.
M. En ökad ömsesidighet mellan EU och AVS bör främja AVS‑ländernas konkurrenskraft, men det kommer sannolikt att skada konkurrenssvaga industrier och bräckliga ekonomier.
N. Avtal om ekonomiskt partnerskap utformas inte alltid så att de stämmer överens med befintliga regionala arrangemang för ekonomisk integration.
O. Jordbruket är utvecklingsmotorn för de flesta AVS‑länder, och för att avtalen om ekonomiskt partnerskap skall kunna bli ett utvecklingsredskap måste de behandla de utmaningar som jordbruket i AVS‑länderna står inför.
Q. En ökning av den inomregionala handeln, som avtalen om ekonomiskt partnerskap syftar till, hindras av svaga infrastrukturer inom regionerna och många andra handelshinder än tullar.
R. De regionala förberedande arbetsgruppernas misslyckande med att spela den roll som man avsåg har förhindrat förhandlingarna och gett upphov till frågor om den framtida effektiviteten hos de övervakningsmekanismer som är kopplade till avtalen om ekonomiskt partnerskap.
S. Bristen på information vid analysen av AVS‑ekonomierna har gjort det mycket svårt att genomföra fullständiga konsekvensanalyser av avtalen om ekonomiskt partnerskap.
T. Förbättrade handelsregler måste följas av ökat stöd för handelsrelaterat bistånd.
U. Det handelsrelaterade biståndet syftar till att stödja utvecklingsländernas förmåga att utnyttja nya handelsmöjligheter.
V. Man måste finna en lösning på problemet med anpassningskostnader i samband med förberedelserna inför och genomförandet av de avregleringar som krävs som en del av avtalen om ekonomiskt partnerskap.
W. Enligt artikel 37.4 i Cotonouavtalet krävs en formell och omfattande översyn av de arrangemang som planeras för alla länder för att se till att ingen ytterligare tid behövs för förberedelser eller förhandlingar.
2.
Europaparlamentet bekräftar på nytt sin inställning att om avtalen om ekonomiskt partnerskap utformas på rätt sätt kan de ge nytt liv åt handelsförbindelserna mellan AVS och EU, främja AVS‑ländernas ekonomiska diversifiering och regionala integration samt minska fattigdomen i AVS‑länderna.
Parlamentet betonar att ”Dokument om europeiskt samförstånd” (förklaringen om utvecklingspolitik), särskilt punkt 36, ger vägledning åt förhandlarna i samband med avtalen om ekonomiskt partnerskap.
Europaparlamentet uttrycker sin oro över den långsamma förhandlingstakten och den brist på påtagliga framsteg som följer av den, med många kritiska problem som fortfarande återstår att diskutera eller avtala om.
Europaparlamentet uppmanar kommissionen att göra sitt yttersta för att förhandlingarna om utvecklingsagendan från Doha skall kunna återupptas och för att se till att avregleringsavtalen främjar utvecklingen i fattiga länder.
Europaparlamentet inser att förmånstillträde till marknaderna inte har varit ett tillräckligt verktyg i sig självt för att utveckla AVS‑länderna och understryker att man, för att uppnå det målet, måste vidta kompletterande åtgärder som stärker AVS‑ländernas konkurrenskraft.
28.
Europaparlamentet påminner om att AVS‑länderna ofta är starkt beroende av råvaror och uppmanar EU att utveckla effektivare biståndsinstrument för anpassning och diversifiering av produktionen, samt för utveckling av bearbetningsindustri och små och medelstora företag i AVS‑länderna.
Europaparlamentet uppmanar kommissionen och AVS‑länderna att se översynen av avtalen om ekonomiskt partnerskap som en möjlighet att öppet diskutera hindren för att slutföra förhandlingarna och lägga fram detaljerade förslag för att komma förbi dem.
37.
Europaparlamentet påminner om AVS‑ländernas krav i ett antal olika forum om alternativ till avtal om ekonomiskt partnerskap, men noterar bristen på officiella krav från AVS‑länderna i enlighet med artikel 37.6 i Cotonouavtalet.
38.
Europaparlamentet uppmanar kommissionen att lägga fram förslag till de alternativ inriktade på utveckling som erbjuder mer än bara marknadstillträde, såsom fallet är med ”Allt utom vapen” och GSP+.
40.
Europaparlamentet kräver ett tvistlösningssystem för avtal om ekonomiskt partnerskap som är tillräckligt enkelt och kostnadseffektivt för att snabbt kunna tas i bruk om parterna inte uppfyller sina åtaganden.
Europaparlamentet uppmanar kommissionen att ta initiativ till och mobilisera internationellt bistånd för att revidera eller klargöra artikel XXIV i GATT‑avtalet i fråga om frihandelsavtal mellan parter med olika utvecklingsnivå.
Europaparlamentet kräver inrättandet av en parlamentarisk tillsynskommitté för avtal om ekonomiskt partnerskap – inom den gemensamma parlamentariska AVS‑EG församlingen och inte som ytterligare en institution – för att offentligt övervaka och se över hur genomförandet av avtalen om ekonomiskt partnerskap påverkar handel och utveckling, göra utvecklingspolitiken mer sammanhängande och utarbeta mekanismer som garanterar ansvarsskyldighet och regelbunden rapportering om hur avtalen om ekonomiskt partnerskap bidrar till en rättvis och hållbar utveckling.
MOTIVERING
Syftet med detta betänkande har varit att det skall vara konstruktivt, realistiskt och balanserat.
Föredraganden har försökt att fokusera på verkligheten att avtal om ekonomiskt partnerskap mellan EU och AVS‑länderna kommer att ingås, att WTO‑förenligheten är viktig och ”att åstadkomma en hållbar utveckling och att uppnå en gradvis integrering av AVS‑staterna i världsekonomin, minska och på sikt utrota fattigdomen”
En stor del av debatten om handel och utveckling är polariserad.
År av diskussioner om fördelarna med avregleringen och den fria handeln har inte bidragit till att föra förhandlingarna framåt.
Trots att dessa debatter är intressanta är det viktigt att rikta uppmärksamheten mot hur de vackra orden i Cotonouavtalet skall införas i avtalen om ekonomiskt partnerskap.
När det gäller handel och utveckling ligger problemet i detaljerna.
Förhandlingarna om avtal om ekonomiskt partnerskap har kännetecknats av misstro och meningsskiljaktigheter om hur handeln skall göras till ett ”utvecklingsverktyg”.
Misstag har begåtts i inställningen till och genomförandet av förhandlingar som är omfattande och ambitiösa.
Rösterna hos dem som kommer att påverkas av avtalen om ekonomiskt partnerskap har inte alltid blivit tillräckligt hörda, och effekterna av avtal om ekonomiskt partnerskap på AVS‑länderna har inte alltid kvantifierats helt.
Svårigheter
Svårigheterna med att förhandla fram ett ”partnerskapsavtal” mellan sådana ojämlika partner i kontroversiella och komplexa frågor är uppenbara.
Bristen på detaljerad ekonomisk information och begränsningar av kapaciteten i AVS‑länderna har, tillsammans med EU:s institutionella stelhet – där GD Bistånd inom Europeiska kommissionen är ansvarigt för medlen medan GD Handel är ansvarigt för förhandlingarna – bidragit till en förhandlingsmiljö som skiljer sig mycket från ett konventionellt frihandelsavtal.
Kommissionens oförmåga att göra ”utvecklingsdimensionen” tillräckligt central för förhandlingarna om avtal om ekonomiskt partnerskap har varit ett betydande hinder för framstegen i samtalen om avtal om ekonomiskt partnerskap.
AVS‑ländernas oförmåga att i detalj beskriva vad de vill ha i ”utvecklingsdimensionen” utöver begäran om ytterligare finansiering för vilken ingen kostnadsberäkning har gjorts har gjort det svårt för berörda parter att hålla kommissionen ansvarig i kravet på ”utvecklingsfrämjande avtal om ekonomiskt partnerskap”.
Det beror särskilt på att de instrument som inrättas för att se till att förhandlingarna om avtal om ekonomiskt partnerskap är ”utvecklingsfrämjande” antingen inte har fungerat eller har saknat trovärdighet.
Om den omständigheten att kommissionen protesterar över att AVS‑länderna alltid bara ber om mer finansiering, medan AVS‑länderna klagar över att kommissionen inte förstår deras behov, låter som ett dysfunktionellt äktenskap beror det troligen på att detta är ett partnerskap med kommunikationsproblem.
Intrycket kvarstår att EU tvingar igenom frihandelsavtal som kommer att skada AVS‑länderna genom att säga en sak officiellt och en annan privat.
Tidigare erfarenheter i många AVS‑länder har lett till en skeptisk inställning till huruvida att göra det som givarländerna vill kommer att minska fattigdomen.
Program för avreglering av handel under 1980‑ och 1990‑talen i många AVS‑länder uppfattades i dessa länder inte som den stora framgång som internationella organisationer och givarländernas regeringar hade fått dem att tro att de skulle bli.
Varje avtal om ekonomiskt partnerskap som undertecknas av en regional grupp måste vara politiskt önskvärt på både kort och lång sikt.
Löftet om ekonomiska fördelar i en avlägsen framtid kommer inte att räcka om intrycket kvarstår att avtal om ekonomiskt partnerskap kräver avreglering utan fördelar som inte redan är tillgängliga för de minst utvecklade länderna enligt avtal om ekonomiskt partnerskap.
Positiva förslag
Handelssamtalen går vanligen långsamt framåt fram till precis före den deadline då saker och ting plötsligt börjar hända.
I detta fall kommer denna taktik inte att vara användbar eftersom fördelarna måste vara tydliga innan avtal om ekonomiskt partnerskap ingås för att skingra oron för att AVS‑länderna manövreras ut i utbyte mot en stor check med återvunna pengar.
Det är rätt av AVS‑länderna att ifrågasätta huruvida kommissionens förslag kommer att bidra till deras utveckling på det sätt som de vill och huruvida löftena om ytterligare ekonomiskt bistånd verkligen är utöver detta.
Om avtal om ekonomiskt partnerskap skall kunna ingås med framgång måste det dock finnas ett större engagemang i och ansvarstagande för resultatet av förhandlingarna om avtal om ekonomiskt partnerskap än vad som har varit fallet med processen.
Föredraganden anser att en parlamentarisk tillsynskommitté för avtal om ekonomiskt partnerskap skulle bidra till detta mål, och den gemensamma parlamentariska AVS‑EG‑församlingen utgör den lämpliga miljön för denna tillsyn.
Den är ett forum som behöver ett syfte, medan avtalen om ekonomiskt partnerskap är ett partnerskap med demokratiska problem som rör ansvar och trovärdighet.
Den omständigheten att den gemensamma parlamentariska församlingen är knuten till Cotonouavtalet, som kommer att upphöra 2020 – men den parlamentariska tillsynen över avtalen om ekonomiskt partnerskap skulle inte göra det – kan tyda på att ytterligare en institution bör skapas.
Det skulle inte vara ett effektivt utnyttjande av resurser.
Ytterligare resurser
Det är tydligt att ytterligare resurser kommer att behövas för att hantera effekterna av förändringar som inleds i avtalen om ekonomiskt partnerskap.
Upptrappningen av underlättandet av handel, tekniskt bistånd och stöd till AVS‑producenterna för att uppfylla EU‑standarderna måste vara tillräckligt omfattande för att kvitta förlusterna från tullintäkter och hjälpa AVS‑länderna att utnyttja tillträdet till marknaden.
I första hand kräver detta ett större arbete för att se till att medel som redan har utlovats spenderas snabbt och effektivt.
Förbättringar av EUF‑förfarandena (Europeiska utvecklingsfonden) bör prioriteras tillsammans med begäran om mer pengar.
EU måste hållas ansvarigt för allt sitt utvecklingsbistånd och kan inte utlova ogrundade belopp över ospecificerade tidsperioder utan tydliga mål.
EU måste emellertid arbeta för att se till att mer bistånd ges till projekt som kommer att öka AVS‑ländernas konkurrenskraft och tillväxt utan att minska utgifterna för hälsa och utbildning.
Slutsatser
Detta betänkande ger en påminnelse i tid till kommissionen om att tidsfristen fram till den 1 januari 2008 närmar sig snabbt, och det återstår en oroväckande stor mängd arbete.
Allvarliga frågor om förmågan och viljan hos många AVS‑länder att genomföra de ambitiösa förslagen från kommissionen kommer sannolikt inte att besvaras före utgången av 2007.
Att granskningen inte var ”inkluderande och konsulterande med alla berörda parter inbegripet icke‑statliga aktörer och parlamentsledamöter”
Krav som framfördes av AVS‑rådet i Port Moresby. gör en andra Europaparlamentets resolution där oro uttrycks över de långsamma framstegen i samtalen ännu mer brådskande, särskilt med avseende på tidsfristen.
I alla regioner anses detta mål som bäst vara mycket ambitiöst.
Även om det inte ligger i någons intresse att tvinga fram ett avtal kommer fokuseringen på ännu ett WTO‑avstående inte att lösa de bakomliggande problem som har gjort framstegen i förhandlingarna om avtalen om ekonomiskt partnerskap så svåra redan från början.
När det gäller tidsfristen behövs en balans, precis som för utfasningen av avregleringen.
På WTO‑nivå vet ingen vad som kommer att hända om sex helt nya avtal om ekonomiskt partnerskap inte träder in i den internationella handelns värld den 1 januari 2008.
Om vissa regioner behöver mer tid anser föredraganden att AVS‑ländernas export till EU inte bör skadas i väntan på en slutgiltig lösning.
Förhandlarna måste fortsätta med förhandlingarna för att nå en ömsesidigt gynnsam lösning om avtalen om ekonomiskt partnerskap som kommer att bidra till AVS‑ländernas utveckling.
Avtalen om ekonomiskt partnerskap måste vara ett äkta partnerskap om de skall kunna fungera.
ÄRENDETS GÅNG
Titel
Avtal om ekonomiskt partnerskap
Förfarandenummer
2005/2246(INI)
INTA 15.12.2005
Rådgivande utskott Tillkännagivande i kammaren
Inget yttrande avges Beslut
Robert Sturdy 11.10.2005
Tidigare föredragande
Behandling i utskott
3.10.2006
23.1.2007
27.2.2007
Antagande
21.3.2007
Slutomröstning: resultat
+:
–:
21
6
Slutomröstning: närvarande ledamöter
Kader Arif, Graham Booth, Carlos Carnero González, Christofer Fjellner, Béla Glattfelder, Eduard Raul Hellvig, Jacky Henin, Syed Kamall, Ģirts Valdis Kristovskis, Caroline Lucas, Marusya Ivanova Lyubcheva, Erika Mann, David Martin, Georgios Papastamkos, Godelieve Quisthoudt-Rowohl, Tokia Saïfi, Peter Šťastný, Robert Sturdy, Daniel Varela Suanzes-Carpegna, Zbigniew Zaleski
Slutomröstning: närvarande suppleant(er)
Jean-Pierre Audy, Panagiotis Beglitis, Danutė Budreikaitė, Albert Deß, Elisa Ferreira, Małgorzata Handzlik, Jens Holm, Eugenijus Maldeikis, Zuzana Roithová
Slutomröstning: närvarande suppleant(er) (art.
178.2)
Sepp Kusstatscher, Corien Wortmann-Kool
Ingivande
27.3.2007
Anmärkningar (tillgängliga på ett enda språk)
SLUTLIG VERSION
A6-0096/2007
BETÄNKANDE
om den framtida regionalpolitikens bidrag till Europeiska unionens innovativa kapacitet
(2006/2104(INI))
Utskottet för regional utveckling
Föredragande:
Mieczysław Edmund Janowski
PE 382.399v04-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING..........................................................................................................................15
YTTRANDE från budgetutskottet ............................................................................18
ÄRENDETS GÅNG..................................................................................................................21
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om den framtida regionalpolitikens bidrag till Europeiska unionens innovativa kapacitet
( 2006/2104(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av artiklarna 2, 3, 158, 159 och 160 i EG-fördraget,
– med beaktande av rådets förordning (EG) nr 1083/2006 av den 11 juli 2006 om allmänna bestämmelser för Europeiska regionala utvecklingsfonden, Europeiska socialfonden och Sammanhållningsfonden
EUT L 210, 31.7.2006, s.
25. samt rättelsen till denna
EUT L 239, 1.9.2006, s.
248. ,
– med beaktande av rådets förordning (EG) nr 1084/2006 av den 11 juli 2006 om inrättande av Sammanhållningsfonden
EUT L 210, 31.7.2006, s.
79. ,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1080/2006 av den 5 juli 2006 om Europeiska regionala utvecklingsfonden
EUT L 210, 31.7.2006, s.
1. ,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1081/2006 av den 5 juli 2006 om Europeiska socialfonden
EUT L 210, 31.7.2006, s.
12. ,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1082/2006 av den 5 juli 2006 om en europeisk gruppering för territoriellt samarbete (EGTS)
EUT L 210, 31.7.2006, s.
19. ,
– med beaktande av rådets beslut av den 6 oktober 2006 om gemenskapens strategiska riktlinjer för sammanhållningen (2006/702/EG)
EUT L 291, 21.10.2006, s.
11. ,
– med beaktande Europaparlamentets och rådets beslut nr 1982/2006/EG av den 18 december 2006 om Europeiska gemenskapens sjunde ramprogram för verksamhet inom området forskning, teknisk utveckling och demonstration (2007–2013)
EUT L 412, 30.12.2006, s.
1. ,
– med beaktande Europaparlamentets och rådets beslut (EG) nr 1639/2006 av den 24 oktober 2006 om att upprätta ett ramprogram för konkurrenskraft och innovation (2007–2013)
EUT L 310, 9.11.2006, s.
15.
– med beaktande av sin resolution av den 10 mars 2005 om Europaparlamentets resolution om vetenskap och teknik – politiska riktlinjer för forskningsstöd i Europeiska unionen
EUT C 320, 15.12.2005, s.
259. ,
– med beaktande av kommissionens meddelande ”En sammanhållningspolitik för att stödja tillväxt och sysselsättning: Gemenskapens strategiska riktlinjer för perioden 2007–2013” ( KOM(2005)0299 ),
– med beaktande av kommissionens meddelande till rådet, Europaparlamentet, Europeiska ekonomiska och sociala kommittén samt Regionkommittén ”Kunskap i praktiken: en brett upplagd innovationsstrategi för EU” ( KOM(2006)0502 ),
– med beaktande av kommissionens meddelande till rådet, Europaparlamentet, Europeiska ekonomiska och sociala kommittén samt Regionkommittén ”Mer forskning och innovation – Att investera i tillväxt och sysselsättning: En gemensam strategi” ( KOM(2005)0488 ),
– med beaktande av kommissionens meddelande till rådet och Europaparlamentet ”Sammanhållningspolitiken och städerna: städernas och tätorternas bidrag till tillväxt och sysselsättning i regionerna” ( KOM(2006)0385 ),
– med beaktande av kommissionens meddelande ”Tredje framstegsrapporten om sammanhållningen: Mot nytt partnerskap för tillväxt, sysselsättning och sammanhållning” ( KOM(2005)0192 ),
– med beaktande av slutsatserna från Europeiska rådets möte i Lissabon den 23‑24 mars 2000,
- med beaktande av den europeiska stadgan för småföretag som antogs vid Europeiska rådets möte i Feira den 19-20 juni 2000,
– med beaktande av kommissionens meddelande inför europeiska rådets vårmöte 2006 ”Dags att lägga in en högre växel.
Ett nytt partnerskap för tillväxt och sysselsättning” ( KOM(2006)0030 ),
– med beaktande av kommissionens meddelande till Europeiska rådet (det informella mötet den 20 oktober 2006 i Lahtis, Finland) ”Ett innovationsvänligt, modernt Europa” ( KOM(2006)0589 ),
– med beaktande av kommissionens meddelande till europeiska rådet ”Europeiska tekniska institutet: nästa steg mot inrättandet” ( KOM(2006)0276 ),
– med beaktande av kommissionens meddelande ”Regioner för ekonomisk förändring” ( KOM(2006)0675 ),
- med beaktande av rapporten från den oberoende expertgruppen för forskning och utveckling under ledning av Esko Aho med titeln ”Creating an Innovative Europe” (januari 2006), slutrapporten om främjandet av den regionala potentialen för forskning från Europeiska rådgivande forskningskommittén (ERAB) med titeln ”Stimulating regional potential for research and innovation” (november 2005) och kommissionens rapport om innovativa strategier och åtgärder med titeln ”Innovative strategies and actions: results of 15 years of regional experimentation” (oktober 2005),
– med beaktande av European Innovation Progress Report 2006 (TrendChart),
– med beaktande av Regionkommitténs ståndpunkter och yttranden,
– med beaktande av artikel 45 i arbetsordningen,
– med beaktande av betänkandet från utskottet för regional utveckling ( A6‑0096/2007 ), och av följande skäl:
B. Investeringar i sig är inte någon garanti för utveckling men blir, om lämplig politik förs och tillväxtinriktade åtgärder stöds, oumbärliga medel för att utveckling verkligen skall komma till stånd.
C. En ökad innovativ kapacitet bör kunna minska skillnaderna mellan enskilda regioner och därmed till att förverkliga principerna om social solidaritet och harmonisk utveckling.
F. Innovation inom Europeiska unionen bör ses som en dynamisk och interaktiv process där olika aktörer deltar, bland annat regionala och lokala aktörer, i enlighet med subsidiaritetsprincipen.
H. Vissa åtgärder kräver stora finansiella investeringar, medan andra bara behöver nyskapande idéer och/eller att det skapas goda och begripliga lagar som också respekteras.
J. Ungefär 60–70 procent av gemenskapens direktiv genomförs på regional och lokal nivå.
K. Strukturfonderna måste utnyttjas på ett flexibelt sätt så att enskilda regioners specifika kvaliteter kan utnyttjas.
M. Små och medelstora företag spelar en viktig roll för att bygga upp EU:s innovativa kapacitet, bland annat genom det flexibla och snabba sätt på vilket de anammar ny teknik och nya styrformer.
O. Utvecklingen av sektorn för hållbar energi är en av de största utmaningarna för EU.
P. Jordbruket är också en del av ekonomin i vid bemärkelse.
Q. En betydande del, nämligen närmare 70 procent, av medlemsstaternas inkomster kommer från tjänster.
R. De demografiska prognoserna för EU (låga födelsetal och en åldrande befolkning) är en social utmaning för EU och skapar stora möjligheter för innovativa åtgärder i medlemsstaterna, inbegripet tjänstesektorn.
S. Det är viktigt att skapa lämpliga infrastrukturvillkor för transporter, telekommunikationer och informationsnätverk.
V. Innovation är en av Europeiska unionens tre prioriteringar som ingår i de strategiska riktlinjerna (2007-2013).
Politik för humankapital, utbildning, vetenskap och forskning
Europaparlamentet uppmanar kommissionen, rådet och lokala myndigheter att främja forskningsprojekt där resultaten får praktiska tillämpningar och därmed bidrar till regional utveckling.
I syfte att stärka innovationsandan riktar Europaparlamentet en begäran till kommissionen, medlemsstaterna, Regionkommittén och regionala myndigheter att det regionala och lokala samhället skall involveras systematiskt genom en flerriktad stärkning av dialogen med samhället, och särskilt med näringslivskretsar, i enlighet med ”bottom-up”-principen.
8.
(a) administrativ information (på alla nivåer) så att man via Internet kan underlätta huvuddelen av alla myndighetsärenden, inklusive dem som gäller ekonomisk verksamhet.
(b) vetenskaplig, ekonomisk, rättslig och kulturell information, med respekt för upphovsrätten (mer tillgängliga e-bibliotek).
Europaparlamentet uppmanar kommissionen, medlemsstaterna och lokala och regionala myndigheter att se till att alla medborgare har tillgång till sådan information och att uppgifterna i så hög grad som möjligt utförs med hjälp av IKT, något som är särskilt viktigt för personer vars personliga eller yrkesmässiga situation kräver distansarbete eller distansstudier och för dem som själva väljer att arbeta hemma, särskilt de som tar hand om barn, personer med funktionshinder och anhörigvårdare.
Europaparlamentet erkänner nödvändigheten av att skapa innovationsgrupper och innovationsområden på regional nivå och att via nätverk knyta dem samman med motsvarande strukturer i andra regioner och medlemsstater eller tredjeländer.
Europaparlamentet uppmanar kommissionen att utarbeta en strategi för att skapa en öppen, gemensam och konkurrenskraftig europeisk arbetsmarknad för vetenskapsmän och medlemsstaterna och regionala myndigheter att införa denna strategi så att forskare får möjlighet att utvecklas yrkesmässigt genom lämpliga karriärutsikter och åtgärder för underlättad rörlighet.
Ekonomisk politik, energipolitik och finansiella och administrativa verktyg
Europaparlamentet rekommenderar att nationella, regionala och lokala myndigheter vidtar innovativa åtgärder inom tjänstesektorn i vid bemärkelse, inbegripet allmännyttiga tjänster.
Europaparlamentet uppmanar kommissionen, medlemsstaterna och regionala myndigheter att inte bara fokusera på stora projekt och spetsforskningsenheter utan också uppmärksamma mindre projekt i mindre gynnande regioner och skapa anpassade mikrokreditmekanismer.
Europaparlamentet uppmanar medlemsstaterna och kommissionen, i syfte att stoppa den avfolkning av vissa regioner som beror på strukturella nackdelar (såsom fattigdom och arbetslöshet) att på ett effektivare sätt genomföra politiken för utjämning mellan regionerna med beaktande av utvecklingen av innovationer i de regionala ekonomierna, något som skulle stärka gemenskapens innovativa kapacitet och bidra till att uppnå verklig territoriell sammanhållning.
Europaparlamentet uppmanar medlemsstaterna och regionala myndigheter, med tanke på att huvuddelen av EU:s medborgare bor i städer och tätorter och samtidigt den roll dessa spelar som lokala och regionala innovationscentra, att stödja en långsiktig fysisk planering, att skapa lämpliga villkor för ett rationellt och harmoniskt utnyttjande av städernas yta och en hållbar utveckling av dessa, med beaktande av behov såsom ekonomisk utkomst, bostäder och rekreationsmöjligheter, samtidigt som miljön skyddas.
Med tanke på att landbygden, där ungefär 20 procent av gemenskapens befolkning bor, är av strategisk betydelse för EU:s livsmedelsförsörjning, uppmanar Europaparlamentet kommissionen, medlemsstaterna och regionala myndigheter att knyta frågan om produktion och bearbetning av livsmedelsprodukter till innovationspolitiken, liksom landsbygdsbefolkningens levnadsvillkor.
God praxis och konsolidering av innovationspolitiken
Europaparlamentet hoppas att denna resolution kommer att visa på det intresse som städer och regioner har för regional utveckling och tillväxt och att den kommer att bidra till debatten om den årliga rapporteringen av medlemsstaternas krav inom ramen för Lissabonstrategin.
MOTIVERING
Europeiska unionens regionalpolitik bör koppla samman två grundläggande frågor, gemenskapens sammanhållning och behovet av innovationsfrämjande verksamhet.
Under perioden för budgetramen 2007–2013 skall medel från Europeiska regionala utvecklingsfonden, Sammanhållningsfonden och Europeiska socialfonden bidra till att tre grundläggande mål uppnås: konvergens, konkurrenskraft och europeiskt territoriellt samarbete.
Tack vare dessa medel bör gemenskapens regionalpolitik inriktas inte bara på att utjämna skillnaderna i utveckling mellan olika områden inom EU utan också på att öka hela gemenskapens kapacitet för innovativa åtgärder på alla områden.
Vi bör således inte förspilla våra medborgares tid, pengar eller kreativa möjligheter.
Vad som behövs är en lämplig anda och en förståelse så att innovationer inte blir någon exklusiv domän för vetenskapsmän, forskare, uppfinnare, industrimän, affärsmän och politiker.
Framför allt i lokala och regionala sammanhang måste folk känna att innovationer är något för alla, att de kan förbättra deras livsvillkor och livskvalitet.
Därför måste man klart och tydligt understryka att innovationsfrämjande verksamhet är ett måste för EU som helhet, enskilda medlemsstater och samtliga regioner.
Man bör vara medveten om att de medel som EU sammantaget disponerar för närvarande utgör endast cirka 1 procent av gemenskapens BNP.
Utan motsvarande engagemang från medlemsstaterna (och naturligtvis också pengar) kommer innovation endast att bli ett tjusigt slagord, ett ord som låter lika i våra språk då det härstammar från det latinska innovatio .
Det är således hög tid att gå från deklarationer och åtaganden till konkret handling, för innovation är inte ett självändamål.
Innovation bör omfatta den praktiska helhetsutformningen av verksamhet som syftar till en verklig sammanhållning inom gemenskapen när det gäller vetenskap, utbildning och forskning, konstruktion och teknik, juridik och organisation, förvaltning och administration, ekonomi och handel, energi och miljö.
Innovativa lösningar behövs också för sociala problem, hälsovårdsproblem, och frågan om tillgång till kultur.
Var och en av dessa aspekter har sin regionala dimension.
Grunden för all verksamhet som gemenskapen liksom medlemsstaterna och regionerna bedriver bör vara människans välfärd i vid bemärkelse.
Investeringar i människor bör därför ligga i centrum för gemenskapens verksamhet, dvs. skapandet av lämpliga villkor för deras utveckling, bland annat tillgång till utbildning, så att man kan dra nytta av deras intellektuella potential och kreativa förmåga.
Vi måste dessutom utnyttja de positiva erfarenheter som Europas folk samlat under många generationer.
Detta är den grundläggande källan till vår europeiska framgång i den internationella konkurrensen.
Således behövs såväl långtgående, innovativa tankar från många européer som konkreta, innovativa åtgärder.
Det är så mycket nödvändigare som Europas demografiska situation är på väg bli dramatisk.
Inför de nuvarande utmaningarna satte EU genom Lissabonstrategin upp målet att bli världens mest konkurrenskraftiga ekonomi.
Detta skall uppnås bland annat genom att öka utgifterna för forskning och utveckling (FoU) till 3 procent av BNP.
För närvarande är det bara två EU‑länder som uppnår denna nivå - Sverige och Finland.
Lika stora skillnader när det gäller FoU‑investeringar kan ses på regional nivå.
Enligt tillgänglig statistik uppnår 21 av 254 regioner (EU-25) denna nivå.
För att de nya målen i sammanhållningspolitiken skall uppnås är det nödvändigt med aktivare insatser på regional och lokal nivå för att uppnå målen i Lissabonstrategin.
Den innovationsfrämjande politiken, oavsett om det är på EU-, medlemsstats- eller regionnivå, måste vi se i en dynamisk kontext, dvs. ta i beaktande att även andra utvecklas.
Europeiska unionen är en av de två ledande ekonomierna i världen.
BNP i hela EU ligger mycket nära USA:s BNP (12,5 biljoner USD, enligt uppgift från Världsbanken).
EU har dock hittills hamnat efter sina största rivaler när det gäller investeringar i kunskapsekonomin.
Vi bör studera hur Kina och Indien förhåller sig till detta problem.
Enligt tillgängliga uppgifter är EU:s investeringar i forskning 1,96 procent av BNP (2,59 procent av BNP i USA, 12,0 procent av BNP i Japan).
För att Lissabonstrategins mål (även efter dess uppdatering från juli 2005) verkligen skall uppnås är det nödvändigt med ett heltäckande tillvägagångssätt för detta problem, även inom den nya regionalpolitiken.
Denna ståndpunkt återspeglas i kommissionens meddelande av den 13 september 2006 ”Kunskap i praktiken: en brett upplagd innovationsstrategi för EU”.
Där specificeras 10 punkter som har särskild betydelse för den förnyade Lissabonstrategin när det gäller tillväxt och sysselsättning.
Det kan vara värt att påminna om detta citat från meddelandet: ”Det viktigaste ansvaret för att främja innovation vilar ofta på den regionala nivån.
Regionerna bör därför vara delaktiga i utarbetandet och genomförandet av de nationella reformprogrammen, bl.a. genom att de utformar sina egna regionala innovationsstrategier.
Ytterligare satsningar bör göras för att underlätta politiskt lärande och utbyte av bra lösningar mellan medlemsstaterna.
Färdplanen för ett mer innovativt Europa måste således också ha en regional dimension.
Och var det än är möjligt bör affärsänglars verksamhet bidra till större innovationsfrämjande effekter av den politik som förs på lokal och regional nivå.
I detta betänkande har ansträngningar gjorts för att ta hänsyn till ett så vitt spektrum som möjligt av ömsesidiga kopplingar mellan gemenskapens regionalpolitik och dess innovativa potential.
Många källor och synpunkter från företrädare från kommissionen och Regionkommittén har beaktats.
Det kan vara värt att notera att ganska olika åsikter kommer till uttryck i denna fråga.
Ett exempel är det manifest i nio punkter om innovation som den oberoende informationstjänsten Science Business publicerade i november 2006 och som berör relationerna mellan näringslivet och universitetsvärlden.
YTTRANDE från budgetutskottet
till utskottet för regional utveckling
över den framtida regionalpolitikens bidrag till EU:s innovativa kapacitet
( 2006/2104(INI) )
Föredragande:
Nathalie Griesbeck
FÖRSLAG
Budgetutskottet uppmanar utskottet för regional utveckling att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet uttrycker oro över att anslagen till forskning och utveckling inte är tillräckliga för att tillfredsställa unionens verkliga behov så att dess konkurrenskraft kan säkras, även om Europeiska unionens organ erkänner att främjandet av innovationer är av väsentlig betydelse.
Europaparlamentet erkänner nödvändigheten av att skapa innovationsgrupper och innovationsområden på regional nivå och att via nätverk knyta dem samman med motsvarande strukturer i andra regioner och medlemsstater eller tredjeländer.
ÄRENDETS GÅNG
Titel
Den framtida regionalpolitikens bidrag till EU:s innovativa kapacitet
Referensnummer
2006/2104(INI)
Ansvarigt utskott
REGI
BUDG 18.5.2006
Förstärkt samarbete – tillkännagivande i kammaren
Föredragande av yttrande Utnämning
Nathalie Griesbeck 20.9.2004
Tidigare föredragande av yttrande
Behandling i utskott
25.1.2007
Antagande
25.1.2007
Slutomröstning: resultat
+:
–:
0:
29
Slutomröstning: närvarande ledamöter
Slutomröstning: närvarande suppleanter
Paul Rübig, Hans-Peter Martin
Slutomröstning: närvarande suppleanter (art.
178.2)
Anmärkningar (tillgängliga på ett enda språk)
...
ÄRENDETS GÅNG
Titel
Den framtida regionalpolitikens bidrag till Europeiska unionens innovativa kapacitet
Förfarandenummer
2006/2104(INI)
REGI 18.5.2006
BUDG 18.5.2006
Inget yttrande avges Beslut
Mieczysław Edmund Janowski 2.5.2006
Tidigare föredragande
Behandling i utskott
21.6.2006
4.10.2006
23.1.2007
Antagande
20.3.2007
Slutomröstning: resultat
+:
–:
43
4
Slutomröstning: närvarande ledamöter
Alfonso Andria, Stavros Arnaoutakis, Elspeth Attwooll, Tiberiu Bărbuleţiu, Jean Marie Beaupuy, Rolf Berend, Jana Bobošíková, Vasile Dîncu, Gerardo Galeote, Iratxe García Pérez, Eugenijus Gentvilas, Pedro Guerreiro, Gábor Harangozó, Marian Harkin, Mieczysław Edmund Janowski, Gisela Kallenbach, Tunne Kelam, Evgeni Kirilov, Sérgio Marques, Miguel Angel Martínez Martínez, Yiannakis Matsis, Miroslav Mikolášik, Jan Olbrycht, Maria Petre, Markus Pieper, Wojciech Roszkowski, Elisabeth Schroedter, Stefan Sofianski, Grażyna Staniszewska, Catherine Stihler, Kyriacos Triantaphyllides, Oldřich Vlasák, Vladimír Železný
Slutomröstning: närvarande suppleant(er)
Jan Březina, Brigitte Douay, Den Dover, Emanuel Jardim Fernandes, Dariusz Maciej Grabowski, Ljudmila Novak, Mirosław Mariusz Piotrowski, Zita Pleštinská, Christa Prets, Toomas Savi, László Surján, Károly Ferenc Szabó, Nikolaos Vakalis
Slutomröstning: närvarande suppleant(er) (art.
178.2)
Věra Flasarová
Ingivande
30.3.2007
Anmärkningar (tillgängliga på ett enda språk)
SLUTLIG VERSION
A6-0184/2007
***II
ANDRABEHANDLINGS-REKOMMENDATION
om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets beslut om inrättande av ett andra gemenskapsprogram för åtgärder på hälsoområdet (2007–2013)
(16369/2/2006 – C6‑0100/2007 – 2005/0042A(COD))
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Föredragande:
Antonios Trakatellis
PE 386.560v02-00
Teckenförklaring
* Samrådsförfarandet
majoritet av de avgivna rösterna
**I Samarbetsförfarandet (första behandlingen)
majoritet av de avgivna rösterna
**II Samarbetsförfarandet (andra behandlingen)
*** Samtyckesförfarandet
majoritet av parlamentets samtliga ledamöter utom i de fall som avses i artiklarna 105, 107, 161 och 300 i EG-fördraget och artikel 7 i EU-fördraget
***I Medbeslutandeförfarandet (första behandlingen)
majoritet av de avgivna rösterna
***II Medbeslutandeförfarandet (andra behandlingen)
***III Medbeslutandeförfarandet (tredje behandlingen)
majoritet av de avgivna rösterna för att godkänna det gemensamma utkastet
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................15
ÄRENDETS GÅNG..................................................................................................................17
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets beslut om inrättande av ett andra gemenskapsprogram för åtgärder på hälsoområdet (2007–2013)
(16369/2/2006 – C6‑0100/2007 – 2005/0042A(COD) )
(Medbeslutandeförfarandet: andra behandlingen)
Europaparlamentet utfärdar denna resolution
– med beaktande av rådets gemensamma ståndpunkt (16369/2/2006 – C6‑0100/2007 ),
– med beaktande av parlamentets ståndpunkt vid första behandlingen av ärendet
EUT C 291 E, 30.11.2006, s.
372. , en behandling som avsåg kommissionens förslag till Europaparlamentet och rådet ( KOM(2005)0015 )
Ännu ej offentliggjort i EUT. ,
– med beaktande av kommissionens ändrade förslag ( KOM(2006)0234 )
Ännu ej offentliggjort i EUT. ,
– med beaktande av artikel 62 i arbetsordningen,
– med beaktande av andrabehandlingsrekommendationen från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A6‑0184/2007 ).
1.
Rådets gemensamma ståndpunkt
Parlamentets ändringar
Ändringsförslag
1
Skäl 7
(7) Åtta vanliga orsaker till dödlighet och sjuklighet relaterade till icke smittsamma sjukdomar i WHO:s europeiska region är hjärt och kärlsjukdomar, neurologiska och psykiatriska störningar, cancer, sjukdomar i matsmältningsorganen, sjukdomar i andningsorganen, sjukdomar i sinnesorganen, muskuloskelettala sjukdomar och diabetes mellitus.
(7) Åtta vanliga orsaker till dödlighet och sjuklighet relaterade till icke smittsamma sjukdomar i WHO:s europeiska region är hjärt‑ och kärlsjukdomar, neurologiska och psykiatriska störningar, cancer, sjukdomar i matsmältningsorganen, sjukdomar i andningsorganen, sjukdomar i sinnesorganen, muskuloskelettala sjukdomar och diabetes mellitus.
I enlighet med detta bör kommissionen under detta programs löptid lägga fram förslag till rekommendationer från rådet om prevention, diagnos och kontroll av stora sjukdomar.
Motivering
Här återinförs ändringsförslag 105 från första behandlingen.
Om man utbyter bästa praxis i fråga om större sjukdomar i hela Europa kommer detta otvivelaktigt att ge ett mervärde till de nationella hälsostrategierna.
Det är också motiverat med insatser från EU:s sida av effektivitetsskäl och på grund av att man kan minska skillnaderna mellan medlemsstaterna genom att göra de nationella strategierna mer enhetliga.
Till de stora sjukdomarna i Europa hör bland annat hjärt- och kärlsjukdomar, cancer, diabetes och sinnessjukdom.
Ändringsförslag
2
Skäl 10
(10) Programmet bör bygga på resultaten från det tidigare programmet för gemenskapsåtgärder på folkhälsoområdet (2003–2008).
Det bör bidra till en hög fysisk och psykisk hälsonivå och ökad jämlikhet i hälsofrågor i hela gemenskapen genom att insatserna inriktas på att förbättra folkhälsan, förebygga ohälsa och sjukdomar samt undanröja faror för människors hälsa i syfte att bekämpa sjuklighet och förtida dödlighet.
(10) Programmet bör bygga på resultaten från det tidigare programmet för gemenskapsåtgärder på folkhälsoområdet (2003–2008).
Motivering
Programmet bör stärka kapaciteten att ge medborgarna information om hälsofrågor och på så sätt bredda deras kunskaper och valmöjligheter.
Ändringsförslag
3
Skäl 18
(18) Bästa praxis är viktigt eftersom hälsofrämjande och förebyggande åtgärder bör mätas i ändamålsenlighet och effektivitet och inte enbart utifrån ekonomiska hänsyn.
Bästa praxis och de senaste metoderna för att behandla sjukdomar och skador bör främjas så att ytterligare hälsoförluster förhindras och europeiska nätverk av referenscentrum för specifika sjukdomar bör utvecklas.
(18) Bästa praxis är viktigt eftersom hälsofrämjande och förebyggande åtgärder bör mätas i ändamålsenlighet och effektivitet och inte enbart utifrån ekonomiska hänsyn.
Bästa praxis och de senaste metoderna för att behandla sjukdomar och skador bör främjas så att ytterligare hälsoförluster förhindras och europeiska nätverk av referenscentrum för specifika sjukdomar bör utvecklas.
Det är även viktigt att främja goda alternativ som kan vara att föredra av sociala, religiösa eller andra individuella skäl.
Motivering
Det är viktigt att beakta att sjukvården i dag är så bra att man på grund av sociala, religiösa eller andra individuella preferenser kanske väljer en behandlingsmetod som objektivt inte är exakt lika bra som en annan.
Det kan handla om att en som är döende i cancer hellre vill vara nära sina anhöriga än förlänga livslängden eller om att personer av religiösa skäl väljer att inte acceptera bloddonation.
Ändringsförslag
4
(23a) Det behövs en helhetsbetonad och mångsidig syn på folkhälsa, varför även kompletterande och alternativ medicin bör omfattas av de insatser som stöds av programmet.
Motivering
Ändringsförslag 145 från första behandlingen.
Miljontals EU-medborgare utnyttjar kompletterande och alternativ medicin.
Det är viktigt med en helhetsbetonad och mångsidig syn i programmet och att kompletterande och alternativ medicin tas med i dess verksamheter.
Ändringsförslag
5
Skäl 25
(25) I detta beslut fastställs, för hela den tid programmet pågår, en finansieringsram som under det årliga budgetförfarandet utgör den särskilda referensen för budgetmyndigheten enligt punkt 37 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning.
(25) I detta beslut fastställs, för hela den tid programmet pågår, en finansieringsram som under det årliga budgetförfarandet utgör den särskilda referensen för budgetmyndigheten enligt punkt 37 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning.
Vid utarbetandet av det preliminära budgetförslaget förbinder sig den budgetansvariga myndigheten och kommissionen att inte avvika från detta med mer än fem procent under hela den tid programmet gäller, om inte nya objektiva långsiktiga omständigheter uppstår, vilka uttryckligen och exakt skall anges, varvid det bör tas hänsyn till de resultat som uppnåtts vid genomförandet av programmet, framför allt utgående från utvärderingarna.
Alla ökningar till följd av sådana variationer bör förbli inom det tak som finns för den ifrågavarande budgetrubriken.
Motivering
Eftersom budgeten bantats ner måste alla möjligheter som det interinstitutionella avtalet erbjuder undersökas och utnyttjas för att programmet skall få ökade anslag vid det årliga budgetförfarandet.
Ändringsförslag
6
Skäl 25a (nytt)
(25a) Den budgetansvariga myndigheten kan besluta om ändringar i kommissionens årliga programplanering, som tjänar endast som vägledning, och öka åtagande- och betalningsbemyndigandena under de första två eller tre åren av perioden, eventuellt tillsammans med en övervakningsklausul av det slag det stadgas om i det interinstitutionella avtalet.
Motivering
Eftersom budgeten bantats ner måste alla möjligheter som det interinstitutionella avtalet erbjuder undersökas och utnyttjas för att programmet skall få ökade anslag vid det årliga budgetförfarandet.
Ändringsförslag
7
Skäl 25b (nytt)
Motivering
Eftersom budgeten för programmet bantats ner måste alla möjligheter som det interinstitutionella avtalet erbjuder undersökas.
Ändringsförslag
8
Skäl 27
(27) EU:s investeringar i folkhälsa och hälsorelaterade projekt måste öka.
I detta hänseende bör medlemsstaterna uppmuntras att prioritera bättre folkhälsa i sina nationella program.
Det behövs en större medvetenhet om möjligheterna till EU‑finansiering på hälsoområdet.
Medlemsstaterna bör uppmuntras att utbyta erfarenheter av finansiering på hälsoområdet genom strukturfonderna.
(27) EU:s investeringar i folkhälsa och hälsorelaterade projekt måste öka.
I detta hänseende uppmuntras medlemsstaterna att prioritera bättre folkhälsa i sina nationella program.
Det behövs en större medvetenhet om möjligheterna till EU‑finansiering på hälsoområdet.
Medlemsstaterna bör uppmuntras att utbyta erfarenheter av finansiering på hälsoområdet genom strukturfonderna.
Motivering
Eftersom allt stöd från gemenskapen bygger på medfinansiering har medlemsstaterna ansvaret för att delta i finansieringen av hälsofrämjandet.
Ändringsförslag
9
– Främja hälsa.
– Främja åtgärder som leder till hälsosammare levnadsvanor och bidra till minskad ojämlikhet i fråga om hälsa.
Motivering
Här återinsätts kommissionens ursprungliga förslag och dessutom en del av ändringsförslag 50 vid första behandlingen.
Ändringsförslag
10
1.
Finansieringsramen för genomförande av programmet för den tidsperiod som anges i artikel 1 skall vara 365 600 000 EUR .
1.
Finansieringsramen för genomförande av programmet för den tidsperiod som anges i artikel 1 skall vara 402 160 000 EUR .
Motivering
Meningen med den föreslagna tioprocentiga ökningen är att i viss mån korrigera den drastiska budgetnedskärningen.
Vid första behandlingen föreslog parlamentet en budget på 1 500 miljoner EUR.
Nu bör man ta modell av exemplet med LIFE+, där parlamentet också antog en ökning av budgeten vid andra behandlingen, och ställa nödvändiga anslag till förfogande genom att använda den marginal som finns i rubriken 3b.
Ändringsförslag
11
2.
De årliga anslagen skall godkännas av budgetmyndigheten inom ramen för budgetramen.
2.
De årliga anslagen skall godkännas av budgetmyndigheten inom ramen för budgetramen och stå i överensstämmelse med den flexibilitet i lagstiftningen som erbjuds av punkt 37 i det interinstitutionella avtalet, samt flexibilitetsinstrumentet enligt punkt 27 i detta avtal och den halvtidsöversyn som föreskrivs i förklaring 3 till detta avtal .
Motivering
Gemenskapens anslag till hälsoprogrammet är ojämnt fördelade jämfört med anslagen till de övriga fleråriga programmen och därför måste anslagen till hälsoprogrammet utökas i enlighet med flexibiliteten i lagstiftningen, flexibilitetsinstrumentet och halvtidsöversynen av finansieringsramen.
Ändringsförslag
12
3.
Det ekonomiska stödet kan utges av gemenskapen tillsammans med en eller flera medlemsstater eller av gemenskapen tillsammans med de behöriga myndigheterna i andra deltagande länder, om detta är lämpligt med tanke på det mål som skall uppnås.
I detta fall skall gemenskapens stöd vara högst 50 %, utom för åtgärder med exceptionellt stort nyttovärde, varvid gemenskapens stöd skall uppgå till högst 70 %.
Gemenskapens stöd kan tilldelas ett offentligt eller icke vinstdrivande organ som den berörda medlemsstaten eller behöriga myndigheten har utsett genom ett öppet förfarande och som kommissionen har godkänt.
3.
Det ekonomiska stödet kan utges av gemenskapen tillsammans med en eller flera medlemsstater eller av gemenskapen tillsammans med de behöriga myndigheterna i andra deltagande länder, om detta är lämpligt med tanke på det mål som skall uppnås.
I detta fall skall gemenskapens stöd vara högst 50 %, utom för åtgärder med exceptionellt stort nyttovärde, varvid gemenskapens stöd skall uppgå till högst 70 %.
Gemenskapens stöd kan tilldelas ett offentligt eller icke vinstdrivande organ som den berörda medlemsstaten eller behöriga myndigheten har utsett genom ett öppet förfarande och som kommissionen har godkänt.
Detta gemenskapsstöd skall utgå på grundval av de kriterier för patient- och konsumentorganisationer som Europeiska läkemedelsmyndigheten har fastställt.
Motivering
Här återinsätts ändringsförslag 54 från första behandlingen.
Ändringsförslag
13
Bilaga, punkt 2.1.2.
2.1.2.
Stödja initiativ för att fastställa orsakerna till, hantera och minska ojämlikheter i hälsa inom och mellan medlemsstaterna, bland annat sådana ojämlikheter som har samband med könsskillnader, för att bidra till välstånd och sammanhållning; främja investeringar i hälsa i samarbete med annan gemenskapspolitik och andra gemenskapsfonder; öka solidariteten mellan nationella hälso‑ och sjukvårdssystem genom att stödja samarbete i frågor som gäller gränsöverskridande vård.
2.1.2.
Stödja initiativ för att fastställa orsakerna till, hantera och minska ojämlikheter i hälsa inom och mellan medlemsstaterna, bland annat sådana ojämlikheter som har samband med könsskillnader, för att bidra till välstånd och sammanhållning; främja investeringar i hälsa i samarbete med annan gemenskapspolitik och andra gemenskapsfonder; öka solidariteten mellan nationella hälso‑ och sjukvårdssystem genom att stödja samarbete i frågor som gäller gränsöverskridande vård och patienternas rörlighet .
Motivering
I bilagan bör patienternas rörlighet uttryckligen nämnas.
Här återinsätts delar av ändringsförslag 114 från första behandlingen.
Ändringsförslag
14
Bilaga, punkt 2.1.2a. (ny)
2.1.2a.
Bekräfta att patienterna har rättigheter även i egenskap av sjukvårdskonsumenter.
Motivering
Patienter i EU är i dag friskare och mer välinformerade än någonsin.
Sjukvården har förändrats, så den blivit mer professionell och innefattar ett bredare spektrum av aktörer.
Patienten har i dag inte enbart ett behov av skydd utan även ett behov av att kunna utnyttja de medicinska landvinningarna och mångfalden inom vårdsektorn, vilket bör återspeglas i lagstiftningen när det gäller framför allt information och rätt till valfrihet i vården.
Ändringsförslag
15
Bilaga, punkt 2.2.1.
2.2.1.
Påverka hälsans bestämningsfaktorer för att främja och förbättra fysisk och psykisk hälsa, genom att skapa förutsättningar för en hälsosam livsstil och förebygga sjukdomar; vidta åtgärder i fråga om nyckelfaktorer som kost, fysisk aktivitet och sexuell hälsa och i fråga om missbruksrelaterade bestämningsfaktorer, till exempel tobak, alkohol och droger, med tonvikten på nyckelmiljöer som skolor och arbetsplatser, och under hela livscykeln.
2.2.3.
Motivering
Ändringsförslag 87 från första behandlingen.
Detta klargörande syftar till att säkra att åtgärder för att påverka hälsans bestämningsfaktorer inbegriper insatser för att bekämpa beroende av receptbelagda läkemedel, som är en viktig bestämningsfaktor för hälsan.
Ändringsförslag
16
Bilaga, punkt 2.2.3.
2.2.3.
Stödja åtgärder som avser hälsoeffekterna av mer allmänna miljörelaterade och socioekonomiska bestämningsfaktorer.
2.2.3.
Åtgärda hälsoeffekterna av mer allmänna miljörelaterade och socioekonomiska bestämningsfaktorer , framför allt kvaliteten på inomhusluft och exponering för toxiska kemikalier .
Motivering
Det behövs en mer kraftfull formulering i fråga om miljö och hälsa, i stil med ändringsförslag 93 från första behandlingen.
Ändringsförslag
17
Bilaga, punkt 3.1.1a. (ny)
3.1.1a.
Upprätta ett system inom gemenskapen för samarbete kring referenscentrum till förmån för utökad tillämpning av god praxis i medlemsstaterna.
Motivering
Även om målet med hälsovårdssystem inte längre finns med bör stöd till samarbete mellan befintliga referenscentrum tas med i bilagan.
Här återinsätts kommissionens ursprungliga förslag och delar av ändringsförslag 116 från första behandlingen.
Ändringsförslag
18
Bilaga, punkt 3.2.1.
3.2.1.
Fortsätta utvecklingen av ett hållbart system för hälsoövervakning med mekanismer för att samla in uppgifter och information, med lämpliga indikatorer; samla in uppgifter om hälsotillstånd och hälsostrategier; utveckla, som en del av gemenskapens statistikprogram, den statistiska delen av detta system.
3.2.1.
Fortsätta utvecklingen av ett hållbart system för hälsoövervakning med mekanismer för att samla in uppgifter och information, med lämpliga indikatorer; samla in uppgifter om hälsotillstånd och hälsostrategier; inrätta ett europatäckande register över större sjukdomar (t.ex. cancer) åtminstone över livmoderhalscancer, bröstcancer och tjocktarms- och ändtarmscancer, utgående från uppgifter som samlats in vid genomförandet av rådets förordning om cancerscreening; samt utveckla metoder och upprätthålla databaser; utveckla, tillsammans med gemenskapens statistikprogram, den statistiska delen av detta system.
Motivering
Här återinsätts delar av ändringsförslag 126 från första behandlingen i ändrad form.
MOTIVERING
Bakgrund
Våren 2005 lade kommissionen fram ett förslag till ett gemensamt hälso- och konsumentskyddsprogram för perioden 2007–2013 och framhöll då, att det skulle medföra synergivinster både inom förvaltningen och politiken om man slog samman två rätt små program till ett enda stort program.
Det borde även anslås tillräckliga medel för programmet, nämligen 1 203 miljoner EUR, för att det skulle gå att genomföra åtgärderna på folkhälsans och konsumentskyddets område.
Europaparlamentet ställde inte upp bakom tanken på ett gemensamt program för två helt annorlunda sektorer inom politiken, utan beslutade att spjälka upp programmet i två delar, nämligen hälsoprogrammet och konsumentskyddsprogrammet.
Budgeten spjälkades också upp, utgående från den traditionella fördelningen mellan områdena hälsa och konsumentskydd.
När parlamentet antog programmen vid första behandlingen lät parlamentet den ursprungliga budgeten för konsumentskyddsprogrammet kvarstå och ökade avsevärt budgeten för hälsoprogrammet (från 969 miljoner EUR till 1 500 miljoner EUR).
Avsikten var att ge rådet och kommissionen en klar fingervisning om vad parlamentet prioriterade.
Budgetarna för de nya fleråriga programmen inom alla politikområden ingick i förhandlingarna om den nya finansieringsramen för 2007–2013.
Kompromissen mellan medlemsstaterna i december 2005 ledde till att flera politikområden fick avsevärt lägre anslag än vad kommissionen ursprungligen föreslagit.
Det här kunde Europaparlamentet delvis rätta till vid förhandlingarna med rådet våren 2006, men somliga politikområden drabbades värre av uppgörelsen än andra.
Ett av de politikområden som drabbades hårdast var folkhälsan och hälsoprogrammet blev det största offret.
Den ursprungliga budgeten på 969 miljoner EUR som föreslagits av kommissionen och som parlamentet plussat på till 1 500 miljoner EUR bantades ner till bara 365,6 miljoner EUR.
Alltså fick kommissionen lov att slimma ner programmet när den framlade sitt reviderade förslag efter parlamentets första behandling och uppgörelsen om finansieringsramen.
Föredraganden tog med stöd av skuggföredragandena vara på alla möjligheter att rätta till situationen.
Alla försök stupade dock på rådets motstånd, fastän det finländska ordförandeskapet nog visade prov på viss god vilja vid förhandlingarna med parlamentet.
Mot slutet av november 2006 nådde rådet fram till en politisk överenskommelse om hälsoprogrammet för 2007–2013 och antog då i mångt och mycket texten i kommissionens reviderade förslag, också budgeten.
Frågor inför andra behandlingen
Föredraganden håller med om att vi inte precis har särskilt mycket svängrum i budgethänseende.
Han påpekar dock att finansieringsramen låter oss flexa litet grann med marginalerna för varje rubrik och det gör också det årliga budgetförfarandet.
Då man tänker på hur viktigt hälsoprogrammet är har man all orsak att aktivt undersöka och utnyttja de möjligheter som står till buds.
Själva texten behöver också ses över.
I dagens läge, när budgeten bantats ner, är det uppenbarligen inte längre vettigt att anta en väldigt detaljerad förteckning över åtgärder i samband med programmet.
Men ändå måste man få ordning på några av de punkter som parlamentet tog upp vid första behandlingen.
Till exempel syftet med programmet.
Vid första behandlingen tyckte parlamentet det var väldigt viktigt att programmet uttryckligen skulle ta itu med ojämlikheter i fråga om hälsa.
Alltså bör det här också finnas med i programmets syften och mål.
Parlamentet ville också ha kriterier för vilka icke-statliga organisationer som kunde få direkt stöd enligt programmet, exaktare beskrivningar av åtgärderna inom områdena miljö och hälsa, ett system inom gemenskapen för samarbete kring referenscentrum samt ett europatäckande register över sådana cancerformer som omfattas av rådets rekommendation om screening för cancer.
Föredraganden har tagit med motsvarande ändringsförslag i sitt förslag till rekommendation.
Med tanke på hur bred samsyn det råder om dessa ändringar i parlamentet borde rådet visa prov på flexibilitet ifall rådet inte vill att frågan skall gå till förlikning.
ÄRENDETS GÅNG
Titel
Gemenskapens handlingsprogram inom hälsoområdet (2007-2013)
Referensnummer
16369/2/2006 – C6-0100/2007 – 2005/0042A(COD)
Parlamentets första behandling – P ‑nummer
16.3.2006 T6-0093/2006
Kommissionens förslag
KOM(2005)0115 - C6-0097/2005
Kommissionens ändrade förslag
KOM(2006)0234
Mottagande av den gemensamma ståndpunkten: tillkännagivande i kammaren
29.3.2007
Ansvarigt utskott
Tillkännagivande i kammaren
ENVI
29.3.2007
Föredragande
Utnämning
Antonios Trakatellis
24.5.2005
Behandling i utskott
11.4.2007
Antagande
8.5.2007
Slutomröstning: resultat
+:
–:
0:
42
1
Slutomröstning: närvarande ledamöter
Adamos Adamou, Georgs Andrejevs, Margrete Auken, Irena Belohorská, Johannes Blokland, John Bowis, Frieda Brepoels, Martin Callanan, Dorette Corbey, Chris Davies, Avril Doyle, Mojca Drčar Murko, Jill Evans, Satu Hassi, Gyula Hegyi, Jens Holm, Marie Anne Isler Béguin, Dan Jørgensen, Christa Klaß, Urszula Krupa, Marie-Noëlle Lienemann, Peter Liese, Linda McAvan, Alexandru-Ioan Morţun, Roberto Musacchio, Riitta Myller, Péter Olajos, Miroslav Ouzký, Daciana Octavia Sârbu, Karin Scheele, Carl Schlyter, Horst Schnellhardt, Kathy Sinnott, Antonios Trakatellis, Thomas Ulmer, Anja Weisgerber, Åsa Westlund, Anders Wijkman, Glenis Willmott
Slutomröstning: närvarande suppleanter
SLUTLIG VERSION
A6-0287/2007
20.7.2007
BETÄNKANDE
Föredragande:
Britta Thomsen
PE 388.641v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING..........................................................................................................................15
YTTRANDE från utskottet för miljö, folkhälsa och livsmedelssäkerhet 19
YTTRANDE från utskottet för regional utveckling ...................................26
YTTRANDE från utskottet för internationell handel ...............................31
YTTRANDE från utskottet för jordbruk och landsbygdens utveckling 35
ÄRENDETS GÅNG..................................................................................................................39
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om en färdplan för förnybar energi i Europa
( 2007/2090(INI) )
Europaparlamentet utfärdar denna resolution,
– med beaktande av kommissionens meddelande – En energipolitik för Europa ( KOM(2007)0001 ),
– med beaktande av kommissionens meddelande – Färdplan för förnybar energi ( KOM(2006)0848 ),
– med beaktande av kommissionens meddelande – Rapport om framsteg för förnybar energi ( KOM(2006)0849 ),
– med beaktande av kommissionens meddelande – Lägesrapport om biodrivmedel ( KOM(2006)0845 ),
– med beaktande av ordförandeskapets slutsatser från Europeiska rådets möte den 8–9 mars 2007 om Europeiska rådets stöd till ”Europeiska rådets handlingsplan (2007–2009) – En energipolitik för Europa” (7224/07),
– med beaktande av kommissionens arbetsdokument – Färdplan för förnybar energi – ( SEK(2006)1720 /2), som åtföljer färdplanen för förnybar energi,
– med beaktande av konsekvensanalysen ( SEK(2006)1719 /2), som åtföljer färdplanen för förnybar energi,
– med beaktande av kommissionens arbetsdokument – Lägesrapport om biodrivmedel – ( SEK(2006)1721 /2), som åtföljer kommissionens meddelande ( KOM(2006)0845 ),
– med beaktande av sin resolution av den 14 december 2006 om en europeisk strategi för en hållbar, konkurrenskraftig och trygg energiförsörjning – Grönbok
Antagna texter, P6_TA(2006)0603 . ,
– med beaktande av sin resolution av den 14 december 2006 om en strategi för biomassa och biobränsle
Antagna texter, P6_TA(2006)0604 . ,
– med beaktande av sin resolution av den 1 juni 2006 om effektivare energiutnyttjande eller hur man kan göra mer med mindre – Grönbok
Antagna texter, P6_TA(2006)0243 . ,
– med beaktande av sin resolution av den 23 mars 2006 om tryggad energiförsörjning i Europeiska unionen
Antagna texter, P6_TA(2006)0110 . ,
– med beaktande av sin resolution av den 14 februari 2006 om användning av förnybara energikällor för uppvärmning och nedkylning
Antagna texter , P6_TA(2006)0058 . ,
– med beaktande av sin resolution av den 29 september 2005 om andelen förnybar energi i EU och förslag på konkreta åtgärder
EUT C 227 E, 21.9.2006, s.
599. ,
– med beaktande av sin ståndpunkt fastställd vid andra behandlingen den 13 april 2005 inför antagandet av Europaparlamentets och rådets direktiv om upprättande av en ram för att fastställa krav på ekodesign för energianvändande produkter,
– med beaktande av sin ståndpunkt fastställd vid andra behandlingen den 18 december 2003 inför antagandet av Europaparlamentets och rådets direktiv om främjande av kraftvärme på grundval av efterfrågan på nyttiggjord värme på den inre marknaden för energi,
– med beaktande av sin ståndpunkt fastställd vid andra behandlingen den 12 mars 2003 inför antagandet av Europaparlamentets och rådets direktiv om främjande av användningen av biodrivmedel eller andra förnybara drivmedel
EUT C 61 E, 10.3.2004, s.
260. ,
– med beaktande av sin ståndpunkt fastställd vid andra behandlingen den 4 juli 2001 inför antagandet av Europaparlamentets och rådets direktiv om främjande av el producerad från förnybara energikällor på den inre marknaden för el
EGT C 65 E, 14.3.2002, s.
113. ,
– med beaktande av artikel 45 i arbetsordningen,
– med beaktande av betänkandet från utskottet för industrifrågor, forskning och energi och yttrandena från utskottet för internationell handel, utskottet för miljö, folkhälsa och livsmedelssäkerhet, utskottet för regional utveckling och utskottet för jordbruk och landsbygdens utveckling ( A6‑0287/2007 ), och av följande skäl:
A. Vid Europeiska rådets vårmöte i mars 2007 antogs ett bindande mål på 20 procent för andelen förnybar energi av all energikonsumtion i EU senast 2020.
B. Detta mål utgör ett stort steg framåt mot en hållbar europeisk energipolitik som tryggar energiförsörjningen och säkrar konkurrenskraftig energi från förnybara energikällor till ett rimligt pris.
C. I sin resolution av den 14 december 2006 efterlyste Europaparlamentet ambitiösa bindande sektorsmål om att andelen förnybar energi 2020 skall uppgå till 25 procent av primärenergin, och föreslog en färdplan för hur andelen förnybar energi 2040 skall uppgå till 50 procent.
D. Förnybara energikällor, inklusive vattenkraft, har historiskt sett spelat en viktig roll för EU:s elförsörjning.
F. Direktiven för att främja förnybara energikällor på elområdet har lett till eller stärkt hållbar utveckling på detta område i alla medlemsstater.
I. Det finns inga rättsliga bestämmelser om förnybara energikällor för uppvärmning och nedkylning.
J. Förnybara energikällor är ett viktigt inslag i en hållbar energimix och bidrar till
a) minskat importberoende och större variation i bränslemixen,
b) lägre utsläpp av koldioxid och andra ämnen,
c) utveckling av ny och innovativ teknik,
d) sysselsättning och regional utveckling.
K. Marknadsutvecklingen för förnybara energikällor varierar mycket mellan medlemsstaterna, vilket i första hand inte beror på skillnader i potential, utan snarare på olika, och i några fall olämpliga, politiska och rättsliga villkor samt i många fall orimliga administrativa hinder för projektgenomförande.
M. Att uppnå målet att förbättra energieffektiviteten med 20 procent till 2020 är en förutsättning för att kunna nå målet om 20 procent förnybar energi.
N. Främjandet av en marknad för förnybara energikällor kommer att bidra till att nå de reviderade Lissabonmålen genom att öka sysselsättningen och medlemsstaternas och EU:s forsknings‑ och innovationsinsatser.
P. Transportbränslen utgör en betydande och ökande källa till koldioxidutsläpp samtidigt som de även är den huvudsakliga orsaken till luftföroreningar i stadsområden.
Q. Hållbara lösningar på utmaningarna på energiområdet kan nås genom ökad användning av förnybar energi , större förbättringar av energieffektivitet, energibesparingar och teknisk innovation när det gäller klimatvänlig användning av lokala energikällor.
R. Inom uppvärmning och kylning finns en unik möjlighet att använda inte bara förnybar energi utan även överskottsvärme från elproduktion, industri och avfallsförbränning för att på så sätt minska användningen av fossila bränslen och begränsa koldioxidutsläppen.
S. Det är nödvändigt både att garantera att unionens medborgare har en trygg, högkvalitativ energiförsörjning och att skydda miljön, i enlighet med skyldigheten att tillhandahålla allmänna och samhällsomfattande tjänster.
T. Genomförandet av gemenskapens befintliga regelverk för energisektorn är bristfälligt, särskilt när det gäller förnybara energikällor något som på lång sikt undergräver investerarnas förtroende.
U. Utdragna tillståndsförfaranden för projekt för förnybar energi, kraftledningar och distributionsnät står i vägen för en snabb utveckling av förnybara energikällor.
V. Särskilt i fråga om biodrivmedel kan bristen på tydliga miljömässiga och sociala skyddsmekanismer få betydande negativa konsekvenser, såsom en ökad regnskogsskövling utan någon märkbar minskning av växthusgasutsläppen.
Europaparlamentet uppmanar kommissionen att senast 2007 lägga fram ett förslag om en rättslig ram för förnybar energi som skall antas genom medbeslutandeförfarandet med artikel 175.1 i EG-fördraget som rättslig grund.
2.
Europaparlamentet uppmanar kommissionen att i sitt kommande förslag till översyn av systemet för handel med utsläppsrätter säkra en bättre fungerande internalisering av externa kostnader för energiproduktion genom att utsläppsrätterna auktioneras ut för att skapa lika villkor för förnybar energi och garantera att priset blir korrekt.
Europaparlamentet betonar vikten av att utarbeta och genomföra handlingsplaner för förnybar energi på gemenskapsnivå och nationell nivå, och understryker att dessa planer bör bidra till att skapa en verklig gemensam energipolitik för EU.
Europaparlamentet beklagar att man fortfarande inom EU kan notera ett alltför ringa intresse hos de regionala och lokala myndigheterna för utbyggnad och användning av förnybar energi.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att bidra till att skapa ett marknadsklimat som gynnar förnybara energikällor genom att det aktivt främjar decentraliserad produktion och användning av förnybar energi.
Europaparlamentet uppmanar kommissionen att se till att gemenskapslagstiftningen om förnybar energi och de nationella handlingsplanerna innehåller kriterier och bestämmelser som gör det möjligt att undvika konflikter mellan olika användare av biomassa.
Den inre marknaden och nätinfrastrukturen
Europaparlamentet anser att öppet, rättvist och prioriterat tillträde till näten är en nödvändig förutsättning för en framgångsrik integration och expansion av elproduktionen från förnybara energikällor, och att rutinerna för nättillträde och planering bör förenklas och harmoniseras ytterligare, med beaktande av utvecklingen av tekniken för förnybar energi och dess oregelbundna flöde för att undvika att de nationella näten destabiliseras.
Europaparlamentet uppmanar till ökade insatser för att samordna EU‑omfattande planeringsförfaranden och webbplatser om förnybar energi och ordentliga sammanlänkningar av näten.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att bidra till att det skapas en gynnsam marknadsmiljö för förnybar energi, där det också bör ingå att man avskaffar snedvridande subventioner och proaktivt använder den offentliga upphandlingen inom EU, så att man på det sättet kan bidra till att få ned kostnaderna för både energieffektiv teknik och teknik som bygger på förnybar energi.
Europaparlamentet begär att man skall se över eventuell befintlig gemenskapslagstiftning som hindrar utvecklingen av EU:s energipolitiska prioriteringar, inbegripet den framtida utvecklingen av storskaliga tidvattenprojekt.
Europaparlamentet välkomnar Europeiska investeringsbankens stöd till förnybar energi i form av förmånliga krediter och uppmanar kommissionen att stödja den typen av finansiering och uppmuntra den i den offentliga och privata sektorn där det finns ett intresse av satsningar på att utveckla förnybar energi.
Europaparlamentet uppmanar kommissionen att påskynda det omfattande antagandet i alla medlemsstater av bestämmelser om bästa praxis som gör det obligatoriskt, åtminstone i befintliga och avsevärt renoverade eller nya byggnader, att en minimiandel av värmebehovet tillgodoses genom värme från förnybara energikällor, vilket redan är fallet i allt fler regioner och kommuner.
Transport och biodrivmedel
Europaparlamentet uppmanar kommissionen att sträva efter ett samarbete med WTO och liknande internationella organisationer för att garantera internationell acceptans för specifika hållbarhetskriterier och certifieringssystemet, och på så sätt öka den hållbara produktionen av biobränsle runtom i världen och skapa lika villkor för alla.
Europaparlamentet uppmanar medlemsstaterna att undersöka möjligheterna till förnybara energikällor i sina olika regioner för att varje land skall kunna utnyttja de möjligheter som finns så väl som möjligt och på sätt uppmuntra regionerna att använda förnybara energikällor.
Europaparlamentet uppmanar medlemsstaterna att med hjälp av den öppna samordningsmetoden söka efter och jämföra exempel på bästa metoder för att främja produktion och användning av biomassa och biobränslen.
MOTIVERING
En färdplan för förnybar energi
EU står vid en vändpunkt.
Det budskap som föredraganden främst vill lyfta fram i detta betänkande är vikten av att skapa en lämplig ram för denna europeiska satsning.
Målet för förnybar energi kan därför inte betraktas som skilt från de andra målen för genomförandet av en inre marknad för el, målet att nå en energieffektivitetspotential på 20 procent och översynen av handeln med utsläppsrätter för koldioxid.
Alla dessa mål är förbundna med varandra och EU:s främsta prioritering är därför att skapa en lämplig rättslig ram och förmå medlemsstaterna att genomföra den lagstiftning och de beslut som redan har antagits.
EU måste garantera ett långsiktigt perspektiv som uppmuntrar investerarna att engagera sig i denna omfattande satsning.
Dessa nödvändiga förutsättningar måste uppfyllas för att EU skall kunna nå de politiska målen för ökad försörjningstrygghet, minskning av koldioxidutsläppen och skapande av nya arbetstillfällen.
Samtidigt är det viktigt att utforma en energipolitik som bygger på solidaritet med utvecklingsländerna, där 1,6 miljarder personer inte har tillgång till energi.
Energisektorn kan inte längre bara betraktas som en energileverantör, utan måste även vara en aktör och samarbetspartner för att lösa problemen med miljön, klimatet och trygg energiförsörjning.
Nationella handlingsplaner
Föredraganden stöder kommissionens förslag om att de enskilda medlemsstaternas andel av förnybar energi skall fastställas i de nationella handlingsplanerna.
Det finns emellertid fallgropar med denna strategi som man måste vara medveten om vid utformandet och genomförandet av de individuella planerna:
1) En gemensam europeisk energipolitik
För det första är det viktigt att betona att de nationella målen inte får överskugga den dominerande ambitionen att utforma en gemensam energipolitik för EU.
Det är först och främst viktigt att utvidga den gemensamma europeiska rättsliga ramen för förnybar energi och för uppfyllandet av EU:s klimat‑ och energimål.
Detta innebär att kommissionens förslag om en rättslig ram för förnybar energi måste omfatta översyner av direktivet om el från förnybara energikällor, biodrivmedelsdirektivet och ett förslag om en rättslig ram för förnybar energi inom kylnings‑ och uppvärmningssektorn.
Samtidigt måste de befintliga direktiven för det faktiska genomförandet av den inre marknaden för el genomföras (se även nedan).
2) Rättvis fördelning av bördan
För det andra är den största utmaningen att se till att alla medlemsstater bidrar till att nå det ambitiösa målet på 20 procent förnybar energi och 20 procents energieffektivitet till 2020.
Hittills har endast ett fåtal mycket aktiva medlemsstater bidragit till utvecklingen av förnybar energi i EU.
Föredraganden anser därför att kommissionen måste ges en central roll i arbetet med samordning, kvalitetssäkring och övervakning av de olika ländernas insatser.
Dessutom skall medlemsstaterna vara skyldiga att lämna regelbundna rapporter så att kommissionen fortlöpande kan ingripa om de enskilda medlemsstaterna inte uppfyller sina skyldigheter.
Kommissionen måste kunna kontrollera att de nationella handlingsplanerna uppfyller kraven och ha rätt att avslå dem om det inte finns tillräcklig dokumentation om utvecklingen av förnybar energi i förhållande till de nationella målen och där det inte är klart dokumenterat hur systemoperatörerna förväntas genomföra sådan utveckling och hur de nödvändiga investeringarna skall finansieras.
Föredraganden föreslår att bördan skall delas på grundval av en objektiv beräkning av de olika ländernas potential för förnybar energi.
Därför är det fel att hävda att ett land skall klara sig billigare undan bara för att det har stora resurser av förnybar energi om potentialen för förnybar energi fortfarande är stor.
Det är följaktligen viktigt att se till att tekniken anpassas till de lokala förhållandena.
Föredraganden är oroad över vissa medlemsstaters inställning att särskild hänsyn skall tas till länder med en låg kolenergimix.
Syftet med att anta mål för förnybar energi måste vara att främja förnybara energikällor och inte bara energikällor med lågt kolinnehåll i allmän bemärkelse.
Fördelarna med förnybar energi för EU handlar inte bara om att minska koldioxidutsläppen utan handlar minst lika mycket om den energi som EU kan producera, och därigenom både minska beroendet av energiimport och bidra till att skapa arbetstillfällen och tillväxt i EU.
Det finns särskild anledning att vara uppmärksam på följderna av en eventuell minskning av de relevanta målen till under 20 procent för de största medlemsstaterna.
Om detta till exempel skulle beslutas för de fem största medlemsstaterna kommer det att innebära – eftersom de svarar för så mycket som 60 procent av energikonsumtionen – att en oproportionerligt stor andel av förnybar energi kommer att krävas av de övriga länderna för att nå EU:s övergripande mål på 20 procent.
3) Metoden för att beräkna bidraget från teknik för förnybar energi
Det finns ett särskilt problem med den statistiska metoden för att beräkna bidraget från de olika teknikerna för förnybar energi.
Den metod som används av Eurostat för att beräkna bidraget från de olika teknikerna för förnybar energi innebär, som kommissionen påpekar i ”Färdplan för förnybar energi”, att den el som kommer från vindkraft och solenergi straffas i förhållande till elen från biomassa.
Detta beror på att bidraget från biomassa beräknas på grundval av biomassans energiinnehåll innan den omvandlas till el genom förbränning i en kraftstation.
Omvandlingsprocessen medför en betydande förlust på cirka 60 procent som inte dras av i beräkningen av biomassans bidrag.
Vindkraft och solenergi beräknas på grundval av energiinnehållet i den el som genereras.
Det faktum att förlusten under omvandlingsprocessen inte räknas med ger biomassa en orättvis fördel framför vind‑ och solenergi.
Denna ofördelaktiga situation orsakar i synnerhet problem för de länder där andelen vindkraft eller solenergi av elproduktionen är särskilt hög.
Kommissionen bör överväga denna problematiska fråga i samband med att den lägger fram sitt förslag till direktiv om förnybar energi.
När det gäller de nationella handlingsplanerna är föredraganden slutligen oroad för huruvida kommissionen, och i synnerhet generaldirektoratet för energi och transport, har tillräckligt med personal för att klara av det mycket omfattande genomförande‑ och övervakningsarbetet.
Parlamentet måste i starkast möjliga ordalag vädja om att nödvändig personal rekryteras för att garantera att de högt ställda målen och planerna inte läggs på hyllan och glöms bort.
Den inre marknaden
För att målet på 20 procent förnybar energi skall kunna nås måste villkoren för tillträde till elöverföringsnäten för förnybara energikällor förbättras.
Detta kräver att den inre marknaden för energi fungerar bra, med ett öppet, icke‑diskriminerande och effektivt nättillträde för förnybar energi, och nätet måste samtidigt vara tillräckligt utvecklat för att kunna klara stora kvantiteter el från förnybara energikällor.
Föredraganden anser att en uppdelning av ägarskapet för de systemansvariga för överföringssystemen från de kommersiella verksamheterna är den bästa garantin för att producenter av förnybar energi inte kommer att diskrimineras när det gäller nättillträde.
Stödordningar
Föredraganden anser att samordnade stödsystem på EU‑nivå är det slutliga målet, men marknaden är inte redo för detta i nuläget.
Å ena sidan är det viktigt att först kunna garantera fullt genomförande av den inre marknaden för el och att det råder rättvisa och lika villkor för el från alla energikällor, och å andra sidan måste ett system som garanterar teknisk mångfald utformas, så att de tekniker som fortfarande bara befinner sig på experimentstadiet men som har potential på lång sikt inte trängs ut från marknaden i förtid.
För att en inre marknad för förnybar energi skall kunna inrättas är det även viktigt att ta hänsyn till de skilda egenskaperna hos förnybar energi, särskilt skillnaderna mellan bränsleenergi och producerad energi, se avsnittet om metoder ovan.
Annars kommer marknadsfördelarna för länder som t.ex. har stor potential för biomassa eller för sol- eller vindenergi skilja sig stort sinsemellan.
Transportsektorn och förnybar energi
Föredraganden instämmer i kommissionens bedömning om att biodrivmedel för närvarande utgör en stor möjlighet för att öka andelen förnybar energi inom transportsektorn.
Samtidigt anser föredraganden emellertid att det är viktigt att betona behovet av att tillämpa en allsidig strategi för transportsektorn, så att den ökade inriktningen på biodrivmedel inte minskar pressen på sektorn för att utveckla effektivare bilar och på de politiska målen för att bygga ut kollektivtrafiken, samt övergången från vägtransporter till tåg- och sjötransporter.
Ett system som främjar de mest genomförbara biodrivmedelsteknikerna, t.ex. genom certifiering, måste införas.
Systemet bör omfatta både koldioxid‑ och energiöversyner, samt andra miljöeffekter, t.ex. minskad biologisk mångfald.
Systemet måste garantera att det finns effektiva incitament för att främja de tekniker som ger de bästa resultaten enligt dessa översyner.
Samtidigt är det viktigt att se till att certifieringssystemet inte blir ett tekniskt hinder för handeln med tredjeländer.
Främjandet av biodrivmedel får inte leda till att ett nytt system för jordbruksstöd i EU införs, genom att till exempel utestänga konkurrenter från tredjeländer från EU:s marknader.
EU får inte återgå till en protektionistisk politik till försvar för trångsynta sektoriella intressen.
Tendenserna i livsmedelspriserna måste följas noggrant och det är viktigt att se till att det finns lämpliga incitament för att garantera att produktionen av biodrivmedel inte leder till höjningar av livsmedelspriserna och har negativa effekter för befolkningarna i utvecklingsländer.
Den sociala dimensionen
Föredraganden anser att det är viktigt att energipolitikens sociala dimension alltid inbegrips tillsammans med miljödimensionen, säkerhetspolitiska överväganden och ekonomiska perspektiv.
Alla måste ha tillgång till energi, och införandet av förnybar energi får inte orsaka prisökningar som gör att konsumenterna inte har råd att köpa energi för uppvärmning eller el.
Man kan inte förutsätta att marknaden skall lösa detta problem, så EU måste vara redo att stödja de särskilt sårbara grupperna i samhället, som påverkas särskilt starkt av ökande energipriser.
Samtidigt vill föredraganden dock framhålla att betoningen på förnybar energi kommer att skapa möjligheter till arbetstillfällen och tillväxt även i avlägset belägna och mindre bemedlade regioner inom EU.
YTTRANDE från utskottet för miljö, folkhälsa och livsmedelssäkerhet
till utskottet för industrifrågor, forskning och energi
över en färdplan för förnybar energi i Europa
( 2007/2090(INI) )
Föredragande:
Vittorio Prodi
FÖRSLAG
Utskottet för miljö, folkhälsa och livsmedelssäkerhet uppmanar utskottet för industrifrågor, forskning och energi att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
6.
Vidare vidhåller parlamentet att det bör läggas fram ett lagstiftningsförslag för EU-målet på grundval av artikel 175.1 i EG-fördraget, så att både rådet och Europaparlamentet odelat skall kunna medverka.
Europaparlamentet upprepar sitt krav på ett direktiv om främjande av förnybara energikällor inom uppvärmnings- och kylningssektorn, eftersom detta är ett område med avsevärda möjligheter som skulle kunna förverkligas på kort tid och till relativt låga kostnader.
Europaparlamentet betonar framför allt att det måste anläggas mindre och decentraliserade försörjningsstrukturer för att man skall kunna nå målet med en drastisk ökning av andelen lokalproducerad ren energi och påpekar vilka möjligheter kraftvärme och jordvärme erbjuder i detta hänseende.
Europaparlamentet pekar även på behovet av avsevärda investeringar i forskning och utveckling för att främja EU:s innovationskapacitet på området förnybar energi, med beaktande av redan befintliga teknikplattformar.
a) Bidra till att nuvarande mål och framtida, mer ambitiösa mål, kan nås.
b) Stämma överens med principerna för den inre marknaden för el.
c) Ingå som ett led i ett systematiskt arbete för utbyggnad av förnybara energikällor, där det tas hänsyn till särdragen hos de enskilda formerna av förnybar energi, liksom också till geografiska särdrag och olika former av teknik.
d) Effektivt främja användningen av förnybara energikällor och samtidigt vara enkelt och så effektivt som möjligt, framför allt ur kostnadssynvinkel.
e) Internalisera de externa kostnaderna för samtliga energikällor.
f) Tillhandahålla tillräckligt långa övergångstider för de nationella stimulanssystemen, så att inte investerarnas förtroende tar skada.
Parlamentet anser att det i samband med dessa kriterier kunde vara på sin plats med enhetliga gemenskapsrättsliga bestämmelser om inmatningssystem, men att man också kunde tänka sig en modell med kvoter eller anbudsförfaranden, under förutsättning att de svagheter som framkommit hos sådana modeller i somliga medlemsstater går att avhjälpa.
Europaparlamentet påpekar att det brännbara avfallet till 60 procent brukar bestå av förnybart material och efterlyser därför att sådant avfall skall omvandlas till gas och att den energi som alstras vid förbränningen av gasen skall tas till vara på ett miljöriktigt hållbart sätt.
Europaparlamentet uppmanar även kommissionen och medlemsstaterna att öka insatserna till förmån för omvandlingen av biomassa till gas, eftersom biomassa skulle kunna utnyttjas som källmaterial för att framställa syntetiskt flytande fordonsbränsle.
34.
ÄRENDETS GÅNG
Titel
En färdplan för förnybar energi i Europa
Förfarandenummer
2007/2090(INI)
Ansvarigt utskott
ITRE
ENVI 26.4.2007
Förstärkt samarbete – tillkännagivande i kammaren
Föredragande av yttrande Utnämning
Vittorio Prodi 27.3.2007
Tidigare föredragande av yttrande
Behandling i utskott
7.5.2007
Antagande
5.6.2007
Slutomröstning: resultat
+:
–:
0:
56
Slutomröstning: närvarande ledamöter
Adamos Adamou, Georgs Andrejevs, Margrete Auken, Liam Aylward, Irena Belohorská, Johannes Blokland, John Bowis, Hiltrud Breyer, Martin Callanan, Dorette Corbey, Chris Davies, Avril Doyle, Mojca Drčar Murko, Edite Estrela, Jill Evans, Anne Ferreira, Karl-Heinz Florenz, Matthias Groote, Caroline Jackson, Dan Jørgensen, Christa Klaß, Eija-Riitta Korhola, Holger Krahmer, Urszula Krupa, Peter Liese, Jules Maaten, Linda McAvan, Alexandru-Ioan Morţun, Riitta Myller, Péter Olajos, Miroslav Ouzký, Antonyia Parvanova, Vittorio Prodi, Frédérique Ries, Guido Sacconi, Daciana Octavia Sârbu, Karin Scheele, Carl Schlyter, Richard Seeber, María Sornosa Martínez, Antonios Trakatellis, Evangelia Tzampazi, Thomas Ulmer, Anja Weisgerber, Glenis Willmott
Slutomröstning: närvarande suppleanter
Iles Braghetto, Kathalijne Maria Buitenweg, Milan Gaľa, Genowefa Grabowska, Erna Hennicot-Schoepges, Karsten Friedrich Hoppenstedt, Miroslav Mikolášik, Claude Turmes
Slutomröstning: närvarande suppleanter (art.
178.2)
Agustín Díaz de Mera García Consuegra, Christopher Heaton-Harris, Syed Kamall
Anmärkningar (tillgängliga på ett enda språk)
...
14.6.2007
över en färdplan för förnybar energi i Europa
Föredragande:
Marian Harkin
FÖRSLAG
Utskottet för regional utveckling uppmanar utskottet för industrifrågor, forskning och energi att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet uttrycker sin besvikelse över att kommissionen inte bättre kopplar samman utvecklingen av förnybara energikällor med dess inverkan på arbetsmarknadsstrukturen, på utbudet av utbildning och yrkesutbildning liksom på utvecklingen av industriförbindelserna.
Europaparlamentet uppmanar kommissionen att göra det obligatoriskt att när detta är tekniskt möjligt använda sig av samproduktion när förnybar energi produceras från biomassa och att undersöka vilken påverkan projekt med vedpannor har på den lokala och hållbara utvecklingen på området för virke, med tanke på att denna sektor spelar en särskilt stor roll för värderingen av olika regioner och för ekonomins livskraft på landsbygden.
Europaparlamentet uppmanar rådet och Europeiska kommissionen att förutom att utveckla lagstiftningen och förbättra tekniken ägna särskild uppmärksamhet åt vad som krävs för att lyckas, dvs. ett starkt engagemang från de lokala och regionala myndigheterna och från samtliga samhällsaktörer.
Europaparlamentet kräver att subsidiaritetsprincipen skall beaktas till fullo och att lokala och regionala myndigheter skall utarbeta lokala energiplaner som omfattar energibesparing, energieffektivitet och en ökad användning av förnybar energi.
Europaparlamentet uppmanar medlemsstaterna att uppmuntra myndigheterna att tillhandahålla ekonomiska incitament, uppmuntra utbildning, innovation och forskning och utveckling inom området för förnybara energikällor och att utöka innovationsmöjligheterna för företagen.
Europaparlamentet uppmanar medlemsstaterna och kommissionen att genom territoriellt samarbete främja utvecklingen av regionala nätverk för alternativa och förnybara energikällor för konsumenter och slutanvändare.
Europaparlamentet uppmanar medlemsstaterna, vilka hittills har gjort stora investeringar i gamla energiformer, att se till att det investeras tillräckligt, både privat och offentligt, i förnybara energikällor när det gäller forskning och utrustning.
ÄRENDETS GÅNG
Titel
En färdplan för förnybar energi i Europa
Förfarandenummer
2007/2090(INI)
Ansvarigt utskott
ITRE
Yttrande Tillkännagivande i kammaren
REGI 26.4.2007
Förstärkt samarbete – tillkännagivande i kammaren
Föredragande av yttrande Utnämning
Marian Harkin 12.4.2007
Tidigare föredragande av yttrande
Behandling i utskott
2.5.2007
Antagande
7.6.2007
Slutomröstning: resultat
+:
–:
0:
45
Slutomröstning: närvarande ledamöter
Stavros Arnaoutakis, Elspeth Attwooll, Jean Marie Beaupuy, Bernadette Bourzai, Wolfgang Bulfon, Antonio De Blasio, Vasile Dîncu, Gerardo Galeote, Iratxe García Pérez, Eugenijus Gentvilas, Ambroise Guellec, Zita Gurmai, Gábor Harangozó, Filiz Husmenova, Mieczysław Edmund Janowski, Gisela Kallenbach, Tunne Kelam, Evgeni Kirilov, Miloš Koterec, Constanze Angela Krehl, Jamila Madeira, Sérgio Marques, Yiannakis Matsis, Miroslav Mikolášik, James Nicholson, Lambert van Nistelrooij, Jan Olbrycht, Maria Petre, Wojciech Roszkowski, Elisabeth Schroedter, Dimitar Stoyanov, Kyriacos Triantaphyllides, Vladimír Železný
Slutomröstning: närvarande suppleanter
Jan Březina, Den Dover, Mojca Drčar Murko, Lidia Joanna Geringer de Oedenberg, Ljudmila Novak, Francisca Pleguezuelos Aguilar, Zita Pleštinská, Samuli Pohjamo, Christa Prets, Toomas Savi, Gheorghe Vergil Şerbu, László Surján
Slutomröstning: närvarande suppleanter (art.
178.2)
YTTRANDE från utskottet för internationell handel
till utskottet för industrifrågor, forskning och energi
över en färdplan för förnybar energi i Europa
( 2007/2090(INI) )
Föredragande:
Sajjad Karim
FÖRSLAG
Utskottet för internationell handel uppmanar utskottet för industrifrågor, forskning och energi att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet uppmanar kommissionen att säkra en rättvis internationell handel med biodiesel inom ramen för WTO, och att vidta åtgärder mot en snedvridning av den europeiska marknaden som beror på högsubventionerad export av biodiesel från tredjeländer.
ÄRENDETS GÅNG
Titel
En färdplan för förnybar energi i Europa
Förfarandenummer
2007/2090(INI)
Ansvarigt utskott
ITRE
Förstärkt samarbete – tillkännagivande i kammaren
Föredragande av yttrande Utnämning
Behandling i utskott
Antagande
Slutomröstning: resultat
+:
–:
0:
12
1
Slutomröstning: närvarande ledamöter
Carlos Carnero González, Daniel Caspary, Françoise Castex, Christofer Fjellner, Béla Glattfelder, Eduard Raul Hellvig, Jacky Henin, Sajjad Karim, Erika Mann, Vural Öger, Georgios Papastamkos, Tokia Saïfi, Corien Wortmann-Kool
Slutomröstning: närvarande suppleanter
Slutomröstning: närvarande suppleanter (art.
178.2)
YTTRANDE från utskottet för jordbruk och landsbygdens utveckling
till utskottet för industrifrågor, forskning och energi
över ”En färdplan för förnybar energi i Europa”
( 2007/2090(INI) )
Föredragande:
Willem Schuth
FÖRSLAG
Europaparlamentet betonar att framställning och import av biobränslen endast får ske på två villkor, nämligen att EU:s energiberoende inte ökar och att det hela sker långsiktigt.
Europaparlamentet uppmanar med eftertryck kommissionen och medlemsstaterna att snabbt omvandla det bindande, övergripande målet på 20 procent till konkreta, bindande nationella mål.
ÄRENDETS GÅNG
Titel
”En färdplan för förnybar energi i Europa”
Förfarandenummer
2007/2090(INI)
Ansvarigt utskott
ITRE
AGRI 26.4.2007
Förstärkt samarbete – tillkännagivande i kammaren
Föredragande av yttrande Utnämning
Willem Schuth 27.2.2007
Tidigare föredragande av yttrande
Behandling i utskott
7.5.2007
5.6.2007
Antagande
5.6.2007
Slutomröstning: resultat
+:
–:
0:
29
1
Slutomröstning: närvarande ledamöter
Vincenzo Aita, Peter Baco, Niels Busk, Luis Manuel Capoulas Santos, Giuseppe Castiglione, Albert Deß, Ioannis Gklavakis, Lutz Goepel, Bogdan Golik, Friedrich-Wilhelm Graefe zu Baringdorf, Esther Herranz García, Atilla Béla Ladislau Kelemen, Heinz Kindermann, Véronique Mathieu, Mairead McGuinness, Rosa Miguélez Ramos, Neil Parish, Radu Podgorean, Agnes Schierhuber, Willem Schuth, Czesław Adam Siekierski, Csaba Sándor Tabajdi, Marc Tarabella, Donato Tommaso Veraldi, Andrzej Tomasz Zapałowski
Slutomröstning: närvarande suppleanter
Béla Glattfelder, Milan Horáček, Jan Mulder, Markus Pieper, Zdzisław Zbigniew Podkański
Slutomröstning: närvarande suppleanter (art.
178.2)
Anmärkningar (tillgängliga på ett enda språk)
ÄRENDETS GÅNG
Titel
En färdplan för förnybar energi i Europa
Förfarandenummer
2007/2090(INI)
26.4.2007
26.4.2007
8.5.2007
DEVE
Förstärkt samarbete Tillkännagivande i kammaren
Föredragande Utnämning
Britta Thomsen
Tidigare föredragande
Behandling i utskott
11.4.2007
5.6.2007
25.6.2007
Antagande
9.7.2007
Slutomröstning: resultat
+:
–:
36
1
Slutomröstning: närvarande ledamöter
John Attard-Montalto, Pilar del Castillo Vera, Jorgo Chatzimarkakis, Giles Chichester, David Hammerstein, Den Dover, Nicole Fontaine, Norbert Glante, Umberto Guidoni, Fiona Hall, Rebecca Harms, Erna Hennicot-Schoepges, Mary Honeyball, Ján Hudacký, Romano Maria La Russa, Anne Laperrouze, Angelika Niebler, Reino Paasilinna, Atanas Paparizov, Aldo Patriciello, Herbert Reul, Miloslav Ransdorf, Vladimír Remek, Mechtild Rothe, Paul Rübig, Andres Tarand, Britta Thomsen, Catherine Trautmann, Claude Turmes.
Slutomröstning: närvarande suppleant(er)
Pilar Ayuso, Avril Doyle, Göran Färm, Neena Gill, Edit Herczog, Lambert van Nistelrooij, Hannes Swoboda
Slutomröstning: närvarande suppleant(er) (art.
178.2)
Maria Badia i Cutchet
Ingivande
20.7.2007
Anmärkningar (tillgängliga på ett enda språk)
A6-0347/2007
***I
BETÄNKANDE
om förslaget till Europaparlamentets och rådets direktiv om upprättande av en ram för gemenskapens åtgärder för att uppnå en hållbar användning av bekämpningsmedel
(KOM(2006)0373 – C6‑0246/2006 – 2006/0132(COD))
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
Föredragande:
Christa Klaß
Rådgivande utskotts föredragande (*):
Michl Ebner , utskottet för jordbruk och landsbygdens utveckling
(*) Förfarande med associerade utskott – artikel 47 i arbetsordningen
PE 386.502v04-00
Teckenförklaring
* Samrådsförfarandet
majoritet av de avgivna rösterna
**I Samarbetsförfarandet (första behandlingen)
majoritet av de avgivna rösterna
**II Samarbetsförfarandet (andra behandlingen)
*** Samtyckesförfarandet
majoritet av parlamentets samtliga ledamöter utom i de fall som avses i artiklarna 105, 107, 161 och 300 i EG-fördraget och artikel 7 i EU-fördraget
***I Medbeslutandeförfarandet (första behandlingen)
majoritet av de avgivna rösterna
***II Medbeslutandeförfarandet (andra behandlingen)
***III Medbeslutandeförfarandet (tredje behandlingen)
majoritet av de avgivna rösterna för att godkänna det gemensamma utkastet
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................69
Yttrande från utskottet för rättsliga frågor om den föreslagna rättsliga grunden 71
YTTRANDE från utskottet för industrifrågor, forskning och energi 76
YTTRANDE från utskottet för jordbruk och landsbygdens utveckling (*) 85
ÄRENDETS GÅNG................................................................................................................118
(*) Förfarande med associerade utskott – artikel 47 i arbetsordningen
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till Europaparlamentets och rådets direktiv om upprättande av en ram för gemenskapens åtgärder för att uppnå en hållbar användning av bekämpningsmedel
( KOM(2006)0373 – C6‑0246/2006 – 2006/0132(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2006)0373 )
Ännu ej offentliggjort i EUT. ,
– med beaktande av yttrandet från utskottet för rättsliga frågor om den föreslagna rättsliga grunden,
– med beaktande av artiklarna 51 och 35 i arbetsordningen,
– med beaktande av betänkandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet och yttrandena från utskottet för industrifrågor, forskning och energi och utskottet för jordbruk och landsbygdens utveckling ( A6‑0347/2007 ).
Kommissionens förslag
Parlamentets ändringar
Ändringsförslag
1
Beaktandeled 1
Motivering
Syftet med direktivet är att minska bekämpningsmedlens effekt på människors hälsa och miljön.
Både människors hälsa och miljön bör nämnas som rättslig grund för direktivet.
Ändringsförslag
2
Skäl 1
(1) I överensstämmelse med artiklarna 2 och 7 i Europaparlamentets och rådets beslut nr 1600/2002/EG av den 22 juli 2002 om fastställande av gemenskapens sjätte miljöhandlingsprogram bör det upprättas en gemensam rättslig ram för att få till stånd en hållbar användning av bekämpningsmedel.
(1) I överensstämmelse med artiklarna 2 och 7 i Europaparlamentets och rådets beslut nr 1600/2002/EG av den 22 juli 2002 om fastställande av gemenskapens sjätte miljöhandlingsprogram bör det , med hänsyn tagen till försiktighetsprincipen, upprättas en gemensam rättslig ram för att få till stånd en hållbar användning av bekämpningsmedel.
Ändringsförslag
3
Skäl 2
(2) De åtgärder som föreskrivs i detta direktiv bör komplettera och inte påverka åtgärder enligt annan närliggande gemenskapslagstiftning, särskilt förordning (EG) nr […] om växtskyddsmedel, Europaparlamentets och rådets direktiv 2000/60/EG av den 23 oktober 2000 om upprättande av en ram för gemenskapens åtgärder på vattenpolitikens område och Europaparlamentets och rådets förordning (EG) nr 396/2005 av den 23 februari 2005 om gränsvärden för bekämpningsmedelsrester i eller på livsmedel och foder av vegetabiliskt och animaliskt ursprung och om ändring av rådets direktiv 91/414/EEG.
(2) De åtgärder som föreskrivs i detta direktiv bör komplettera och inte påverka åtgärder enligt annan närliggande gemenskapslagstiftning, särskilt förordning (EG) nr […] om växtskyddsmedel, Europaparlamentets och rådets direktiv 2000/60/EG av den 23 oktober 2000 om upprättande av en ram för gemenskapens åtgärder på vattenpolitikens område , Europaparlamentets och rådets förordning (EG) nr 396/2005 av den 23 februari 2005 om gränsvärden för bekämpningsmedelsrester i eller på livsmedel och foder av vegetabiliskt och animaliskt ursprung och om ändring av rådets direktiv 91/414/EEG samt livsmedelslagstiftningens bestämmelser som grundar sig på Europaparlamentets och rådets förordning (EG) nr 178/2002 av den 28 januari 2002 om allmänna principer och krav för livsmedelslagstiftning, om inrättande av Europeiska myndigheten för livsmedelssäkerhet och om förfaranden i frågor som gäller livsmedelssäkerhet 1 .
_______
1 E G T L 31, 1.2.2002, s.
1.
Förordningen senast ändrad genom kommissionens förordning (EG) nr 575/2006 (EUT L 100, 8.4.2006, s.
3).
Motivering
Genom tillägget införs en hänvisning till relevant livsmedelslagstiftning.
Ändringsförslag
4
Skäl 3
(3) För att underlätta genomförandet av detta direktiv bör medlemsstaterna använda nationella handlingsplaner i syfte att fastställa mål för minskning av risker, inbegripet faror, och beroendet av bekämpningsmedelsanvändning och främja icke-kemiska växtskyddsalternativ .
De nationella handlingsplanerna kan samordnas med genomförandeplaner enligt annan närliggande gemenskapslagstiftning och användas för att gruppera samman mål som skall nås enligt annan gemenskapslagstiftning om bekämpningsmedel.
(3) För att underlätta genomförandet av detta direktiv bör medlemsstaterna använda nationella handlingsplaner i syfte att fastställa kvantitativa mål , riktmärken, tidsplaner och indikatorer för förebyggande av både hälso- och miljörisker , utarbeta tidsplaner och indikatorer för bekämpningsmedelsanvändningens risker och intensitet, ange de ekonomiska resurserna och budgetposterna för genomförande av detta inom utsatt tid och främja och uppmuntra ibruktagandet av icke-kemiska växtskyddsmetoder .
De nationella handlingsplanerna bör samordnas med genomförandeplaner enligt annan närliggande gemenskapslagstiftning och användas för att gruppera samman mål som skall nås enligt annan gemenskapslagstiftning om bekämpningsmedel.
Motivering
När det gäller människors hälsa bör riskerna förebyggas helt och inte bara minskas.
Det måste vara klart för medlemsstaterna att syftet med målen i de nationella handlingsplanerna är att ta itu med både hälso- och miljörisker förknippade med användningen av bekämpningsmedel.
Om kravet på att främja icke-kemiska växtskyddsmetoder inte åtföljs av en genuin önskan i medlemsstaterna att uppmuntra ibruktagandet uppnås eventuellt inte detta mål.
Ändringsförslag
5
Skäl 4
(4) Informationsutbytet om de mål och åtgärder som medlemsstaterna fastställer i sina nationella handlingsplaner är en mycket viktig faktor för att nå målen för detta direktiv.
Därför bör medlemsstaterna uppmanas att regelbundet lämna rapporter till kommissionen och övriga medlemsstater, särskilt om genomförandet och resultatet av nationella handlingsplaner och gjorda erfarenheter.
(4) Informationsutbytet om de mål som uppnåtts och de åtgärdsområden som medlemsstaterna fastställer i sina nationella handlingsplaner är en mycket viktig faktor för att nå målen för detta direktiv.
Därför bör medlemsstaterna uppmanas att regelbundet lämna rapporter till kommissionen och övriga medlemsstater, särskilt om genomförandet och resultatet av nationella handlingsplaner och gjorda erfarenheter.
Motivering
I samband med informationsutbyte mellan medlemsstaterna är det inte de mål som fastställts utan i stället de mål som uppnåtts som är viktiga vad avser de åtgärder som vidtagits av medlemsstaterna.
Ändringsförslag
6
Skäl 6
(6) Det är önskvärt att medlemsstaterna inrättar system för utbildning av distributörer, rådgivare och yrkesmässiga användare av bekämpningsmedel så att de som använder eller kommer att använda bekämpningsmedel är fullt medvetna om möjliga hälso- och miljörisker och om lämpliga åtgärder för att minska riskerna så mycket som möjligt.
Utbildningar för yrkesmässiga användare kan samordnas med utbildningar som anordnas inom ramen för rådets förordning (EG) nr 1698/2005 av den 20 september 2005 om stöd för landsbygdsutveckling från Europeiska jordbruksfonden för landsbygdsutveckling (EJFLU).
(6) Det är önskvärt att medlemsstaterna inrättar system för utbildning och fortbildning av distributörer, rådgivare och yrkesmässiga användare av bekämpningsmedel så att de som använder eller kommer att använda bekämpningsmedel är fullt medvetna om möjliga hälso- och miljörisker och om lämpliga åtgärder för att minska riskerna så mycket som möjligt.
Utbildningar för yrkesmässiga användare bör samordnas med utbildningar som anordnas inom ramen för rådets förordning (EG) nr 1698/2005 av den 20 september 2005 om stöd för landsbygdsutveckling från Europeiska jordbruksfonden för landsbygdsutveckling (EJFLU).
Motivering
Man bör föreskriva utbildnings- och fortbildningsåtgärder för distributörer, rådgivare och yrkesmässiga användare av växtskyddsmedel.
Användarnas och säljarnas sakkunskap är nödvändig för att produkterna ska kunna användas korrekt och fylla avsedd funktion.
Ändringsförslag
7
Skäl 6a (nytt)
(6a) Användningen av olagliga växtskyddsmedel äventyrar den hållbara användningen av bekämpningsmedel och utgör en avsevärd risk för miljön och för människors och djurs hälsa.
Detta problem bör åtgärdas omedelbart.
Motivering
Förfalskningar och olaglig handel med växtskyddsmedel i Europa är ett stort och snabbt växande problem.
Detta problem undergräver alla eventuella strategier för hållbarhet genom att det äventyrar konsumenternas och jordbrukarnas hälsa, skadar miljön och förorsakar avsevärda ekonomiska och anseendemässiga skador för jordbrukarna, livsmedelskedjan, regeringar och växtskyddsindustrin.
Ändringsförslag
8
Skäl 7
(7) Konsumenterna och allmänheten bör , särskilt genom medierna, men även genom informationskampanjer, information som lämnas via detaljhandlare och andra lämpliga åtgärder, få kunskaper om de risker som är förknippade med användning av bekämpningsmedel , särskilt deras akuta och kroniska hälsoeffekter samt deras miljöeffekter på kort och lång sikt, och förses med information om icke-kemiska alternativ .
Medlemsstaterna bör övervaka och samla in uppgifter om effekterna av bekämpningsmedelsanvändning, inbegripet förgiftningsfall, samt främja långsiktiga forskningsprogram om effekterna av bekämpningsmedelsanvändning .
Motivering
Detta ändringsförslag tydliggör att konsumenterna och allmänheten bör informeras om bekämpningsmedlens akuta och kroniska effekter på människors hälsa och miljörisker och negativa effekter förknippade med användningen av bekämpningsmedel.
Det effektivaste sättet att informera allmänheten är genom medierna.
Detta skulle möjliggöra för människor att få den kunskap som behövs för att fatta välgrundade beslut och handla kunnigt när det gäller att skydda hälsan och den omgivande miljön.
Ändringsförslag
9
Skäl 9
Motivering
Nödvändigt förtydligande.
Ändringsförslag
10
Skäl 10
(10) Flygbesprutning av bekämpningsmedel kan ge betydande negativ påverkan på människors hälsa och på miljön, särskilt genom vindavdrift.
Det bör därför införas ett generellt förbud mot flygbesprutning, med möjlighet att medge undantag om det innebär klara fördelar och ger miljövinster jämfört med andra spridningsmetoder eller om lämpliga alternativ saknas.
(10) Flygbesprutning av bekämpningsmedel kan ge betydande negativ påverkan på människors hälsa och på miljön, särskilt genom vindavdrift.
Det bör därför införas ett generellt förbud mot flygbesprutning, med möjlighet att medge undantag om lämpliga alternativ saknas , om den bästa tillgängliga tekniken används för att minska avdrift (t.ex. avdriftsreducerande munstycken) och om boendes eller andra närvarande personers hälsa inte påverkas .
Motivering
Flygbesprutning ger inga miljövinster jämfört med andra spridningsmetoder.
Det bör inte vara möjligt att medge undantag i områden där boende och andra närvarande personer kan påverkas, exempelvis tättbefolkade landsbygdsområden, eller nära områden som används av allmänheten och av känsliga grupper, såsom skolor.
Ändringsförslag
11
Skäl 11
(11) Vattenmiljön är särskilt känslig för bekämpningsmedel.
Det är därför nödvändigt att ägna särskild uppmärksamhet åt att undvika förorening av ytvatten och grundvatten genom lämpliga åtgärder, exempelvis att skapa buffertzoner eller plantera häckar längs ytvatten för att minska vattnets exponering för vindavdrift.
Buffertzonernas omfattning bör bland annat avgöras av markförhållanden, klimat, vattendragets storlek och det aktuella områdets jordbruksförhållanden.
Användning av bekämpningsmedel i områden som används som dricksvattentäkt, på eller längs transportleder, t.ex. järnvägslinjer, på hårdgjorda eller mycket genomsläppliga ytor kan leda till högre risker för förorening av vattenmiljön.
I sådana områden bör därför användning av bekämpningsmedel begränsas så långt som möjligt, eller eventuellt undvikas helt.
(11) Vattenmiljön är särskilt känslig för bekämpningsmedel.
Det är därför nödvändigt att ägna särskild uppmärksamhet åt att undvika förorening av ytvatten och grundvatten genom lämpliga åtgärder, exempelvis att skapa buffertzoner eller plantera häckar längs ytvatten för att minska vattnets exponering för vindavdrift.
Buffertzonernas omfattning bör bland annat avgöras av markförhållanden, geologiska och topografiska förhållanden, klimat, vattendragets storlek och det aktuella områdets jordbruksförhållanden.
Användning av bekämpningsmedel i områden som används som dricksvattentäkt, på eller längs transportleder, t.ex. järnvägslinjer, på hårdgjorda eller mycket genomsläppliga ytor kan leda till högre risker för förorening av vattenmiljön.
I sådana områden bör därför användning av bekämpningsmedel begränsas så långt som möjligt, eller eventuellt undvikas helt.
Motivering
Wmywanie pestycydów sięga czasem głębiej niż występujący profil glebowy, dlatego nie tylko sama gleba warunkuje wymiary stref buforowych, ale podłoże skalne (tzw. skała macierzysta).
Gleby w Europie wykształcone są na różnych skałach macierzystych (np:. na wapieniach, piaskach, glinach, lessach, torfach), które różnią się zdolnościami absorpcyjnym.
Dlatego podłoże skalne będzie decydowało o wielkości stref buforowych.
Rzeźba terenu, w tym ekspozycja, nachylenie stoku warunkuje procesy wymywania i spłukiwania, zwłaszcza po ulewach ekstremalnych – przemieszczania cząstek gleby wraz ze stosowanym nawozami, środkami ochrony roślin, w tym pestycydami do niższych części stoku wykorzystywanego rolniczo lub do zbiorników wód powierzchniowych.
Ändringsförslag
12
Skäl 12
(12) Användning av bekämpningsmedel kan vara särskilt farlig i mycket känsliga områden, exempelvis Natura 2000‑områden som är skyddade enligt rådets direktiv 79/409/EEG av den 2 april 1979 om bevarande av vilda fåglar och rådets direktiv 92/43/EEG av den 21 maj 1992 om bevarande av livsmiljöer samt vilda djur och växter.
På andra platser, exempelvis allmänna parker, sportanläggningar och lekplatser för barn, innebär det stora risker om allmänheten exponeras för bekämpningsmedel.
Användning av bekämpningsmedel i dessa områden bör därför begränsas så långt som möjligt, eller eventuellt undvikas helt .
(12) Användning av bekämpningsmedel kan vara särskilt farlig i mycket känsliga områden, exempelvis Natura 2000‑områden som är skyddade enligt rådets direktiv 79/409/EEG av den 2 april 1979 om bevarande av vilda fåglar och rådets direktiv 92/43/EEG av den 21 maj 1992 om bevarande av livsmiljöer samt vilda djur och växter.
De bevarandeåtgärder som är nödvändiga för att uppnå naturskyddsmålen bör vidtas i enlighet med dessa direktiv.
På andra platser, exempelvis bostadsområden, allmänna parker, idrotts- och fritidsområden, skolgårdar och lekplatser för barn samt i närheten av anläggningar för allmän sjukvård (kliniker, sjukhus, rehabiliteringscenter, hälsohem, vårdhem) , innebär det stora risker om allmänheten exponeras för bekämpningsmedel.
I och omkring dessa områden måste därför användning av bekämpningsmedel förbjudas och icke ‑kemiska alternativ användas .
Motivering
Natura 2000-områdena, som för tillfället omfattar över 15 procent av gemenskapens landområden, inbegriper ett stort antal jordbruks- eller skogsbruksområden, i vilka användning av växtskyddsmedel inte strider mot bevarandemålen.
Trots detta är det lämpligt att genom en motsvarande hänvisning påminna om rättsakterna inom naturskyddslagstiftningen.
Kommissionen har erkänt att exponering för bekämpningsmedel i områden som används av allmänheten innebär stora risker.
Med tanke på de akuta och kroniska negativa effekter på hälsan som exponering för bekämpningsmedel kan förorsaka bör därför användningen av bekämpningsmedel förbjudas i och omkring alla områden där allmänheten kan utsättas för exponering (särskilt om de berörda personerna riskerar att utsättas för exponering under en lång tid, såsom personer som bor nära de behandlade områdena), särskilt, men inte uteslutande, för att skydda känsliga befolkningsgrupper.
Ändringsförslag
13
Skäl 14
(14) Om alla lantbrukare tillämpar allmänna standarder för integrerat växtskydd skulle det leda till en mer riktad användning av alla tillgängliga bekämpningsmetoder, däribland bekämpningsmedel.
Detta skulle därför bidra till att ytterligare minska riskerna för människors hälsa och för miljön.
Medlemsstaterna bör främja jordbruk med liten användning av bekämpningsmedel, särskilt integrerat växtskydd, och skapa nödvändiga förutsättningar för tillämpning av integrerat växtskydd.
Medlemsstaterna bör också uppmuntra användning av grödspecifika standarder för integrerat växtskydd.
(14) Om alla lantbrukare tillämpar allmänna och grödspecifika standarder för integrerat växtskydd skulle det leda till en mer riktad användning av alla tillgängliga bekämpningsmetoder, däribland bekämpningsmedel.
Detta skulle därför bidra till att ytterligare minska riskerna för människors hälsa och för miljön och till att minska användningen av bekämpningsmedel .
Medlemsstaterna bör främja jordbruk med liten användning av bekämpningsmedel, särskilt allmänna och grödspecifika standarder för integrerat växtskydd och en ökning av den andel mark som används för ekologiskt jordbruk , och skapa nödvändiga förutsättningar för tillämpning av integrerat växtskydd.
Medlemsstaterna bör också tillämpa bindande grödspecifika standarder för integrerat växtskydd.
Medlemsstaterna bör använda ekonomiska styrmedel för att främja integrerat växtskydd, för att tillhandahålla lantbrukarna rådgivning och utbildning och för att minska riskerna med bekämpningsmedelsanvändning.
En avgift på bekämpningsmedel bör vara en av åtgärderna för att finansiera tillämpningen av allmänna och grödspecifika metoder för integrerat växtskydd samt ökningen av den andel mark som används för ekologiskt jordbruk.
Motivering
Främjandet av icke-kemiska metoder bör inte begränsas till allmänna standarder för integrerat växtskydd utan det bör också omfatta ekologiskt jordbruk och grödspecifika standarder för integrerat växtskydd.
En skatt eller avgift på bekämpningsmedel har visat sig vara ett framgångsrikt sätt att finansiera åtgärder för minskning av bekämpningsmedel i många europeiska länder.
Medlemsstaterna bör kunna välja mellan olika skatte- eller avgiftssystem så att de kan välja ett system som bäst motsvarar deras behov.
Ekonomiska styrmedel brukar vara det effektivaste sättet att minska riskerna för miljön.
Ändringsförslag
14
Skäl 14a (nytt)
(14a) Principen om att förorenaren betalar bör tillämpas med avseende på kostnaderna i samband med genomförandet av detta direktiv.
Medlemsstaterna bör därför överväga att införa en avgift på bekämpningsmedel i syfte att finansiera genomförandet av sina nationella handlingsplaner.
Motivering
Producenternas ansvar för bekämpningsmedelsanvändningens externa kostnader bör ökas.
En avgift eller skatt på bekämpningsmedel bör vara en möjlighet för medlemsstaterna att uppnå en minskad användning och skapa specifika inkomster i syfte att täcka kostnaderna i samband med de nationella handlingsplanerna.
Ändringsförslag
15
Skäl 15
(15) Det är nödvändigt att mäta de framsteg som görs när det gäller att minska de risker och negativa effekter som bekämpningsmedelsanvändningen innebär för människors hälsa och för miljön.
De harmoniserade riskindikatorer som behövs för detta kommer att fastställas på gemenskapsnivå.
Medlemsstaterna bör använda dessa indikatorer för riskhantering på nationell nivå och för rapportering, och kommissionen bör beräkna indikatorer för att utvärdera framsteg på gemenskapsnivå.
Fram till dess att gemensamma indikatorer blir tillgängliga bör medlemsstaterna ha rätt att använda nationella indikatorer.
(15) Det är nödvändigt att mäta de framsteg som görs när det gäller att förebygga användningen av bekämpningsmedel och de risker och negativa effekter som bekämpningsmedelsanvändningen innebär för människors hälsa och för miljön.
De harmoniserade användnings- och riskindikatorer som behövs för detta kommer att fastställas på gemenskapsnivå.
Medlemsstaterna bör använda dessa indikatorer för att minska användningen av bekämpningsmedel och minska riskerna på nationell nivå och för rapportering, och kommissionen bör beräkna indikatorer för att utvärdera framsteg på gemenskapsnivå.
Fram till dess att gemensamma indikatorer blir tillgängliga bör medlemsstaterna ha rätt att använda nationella indikatorer , som bör överensstämma med kraven i detta direktiv och avse både hälso- och miljörisker förknippade med användningen av bekämpningsmedel .
Allmänheten, liksom alla andra berörda parter, bör delta i utvecklingen och fastställandet av nationella indikatorer.
Detta inbegriper ett krav på allmänhetens fulla tillgång till information som stöd för allmänhetens deltagande .
Bestämmelser om allmänhetens rätt att delta fullt ut och ha tillgång till information bör införas .
Motivering
Verktyg för att mäta vilka framsteg som gjorts när det gäller att minska användningen av och riskerna med bekämpningsmedel kommer att hjälpa medlemsstaterna att uppnå de mål som ställts upp inom ramen för gemenskapens sjätte miljöhandlingsprogram, nämligen att ”minska påverkan av bekämpningsmedel för människors hälsa och miljön och, mer allmänt, åstadkomma en mer hållbar användning av bekämpningsmedel samt en betydande total minskning av riskerna och av användningen av bekämpningsmedel”.
När det gäller människors hälsa bör riskerna och de negativa effekterna förebyggas helt och inte endast minskas.
Det bör göras klart för medlemsstaterna att de nationella indikatorerna avser både hälso- och miljörisker förknippade med användningen av bekämpningsmedel.
Det bör också vara klart för medlemsstaterna vilka kraven är för allmänhetens deltagande i utvecklingen och ändringen av nationella indikatorer och i deras mekanismer, i syfte att följa andan i direktiv 2003/35/EG, där allmänhetens deltagande fastställs.
Ändringsförslag
16
Skäl 15a (nytt)
(15a) Som ett led i tillämpningen av principen om att förorenaren betalar bör kommissionen pröva i vad mån tillverkarna av växtskyddsmedel och/eller de verksamma ämnen som ingår i dem bör medverka vid behandling och avhjälpande av skador på människors hälsa och miljön vilka kan uppkomma till följd av att växtskyddsmedel används.
Motivering
Såsom fallet också är inom andra områden av gemenskapens hälso- och miljöpolitik bör tillverkarens ansvar gälla även för växtskyddsmedel och de verksamma ämnena i dem.
Ändringsförslag
17
Skäl 19
(19) De åtgärder som krävs för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter 1 .
__________
1 EGT L 184, 17.7.1999, s.
23.
__________
1 EGT L 184, 17.7.1999, s.
23 .
Beslutet ändrat genom beslut 2006/512/EG (EUT L 200, 22.7.2006, s.
11) .
Motivering
Detta ändringsförslag är nödvändigt för att anpassa texten till bestämmelserna i det nya beslutet om kommittéförfarandet.
Ändringsförslag
18
Artikel 1
Genom detta direktiv upprättas en ram för att uppnå en mer hållbar användning av bekämpningsmedel genom att de risker och effekter som användningen av bekämpningsmedel innebär för människors hälsa och på miljön minskas på ett sätt som är förenligt med ett tillräckligt växtskydd .
Genom detta direktiv upprättas en ram för att uppnå en mer hållbar användning av bekämpningsmedel genom att användningen av bekämpningsmedel och de risker och effekter som användningen av bekämpningsmedel innebär för människors hälsa och på miljön minskas i enlighet med försiktighetsprincipen och genom att främjandet och användningen av icke-kemiska växtskyddsmetoder uppmuntras .
Motivering
Ändringsförslaget syftar till att säkerställa förenlighet med den temainriktade strategin för hållbar användning av bekämpningsmedel och förslaget till förordning om utsläppande av växtskyddsmedel på marknaden.
I den mån icke-kemiska alternativ är tillgängliga på marknaden till ett fördelaktigt pris bör de användas i stället för bekämpningsmedel.
Ändringsförslag
19
1.
Detta direktiv skall tillämpas på bekämpningsmedel i form av växtskyddsmedel enligt definitionen i förordning (EG) nr […] om utsläppande av växtskyddsmedel på marknaden.
1.
Detta direktiv skall tillämpas på bekämpningsmedel i form av
a) växtskyddsmedel enligt definitionen i förordning (EG) nr […] om utsläppande av växtskyddsmedel på marknaden , vilka används i jordbruket och i annan verksamhet,
__________
1 EGT L 123, 24.4.1998, s.
1.
Direktivet senast ändrat genom kommissionens direktiv 2006/140/EG (EUT L 414, 30.12.2006, s.
78).
Motivering
Produkter som används för bekämpning av skadedjur är väldigt lika växtskyddsmedel.
De kan innehålla samma verksamma ämnen som växtskyddsmedel och ibland förekomma i identiska beredningar (t.ex. kan rodenticider omfattas av de båda rättsakterna beroende på om de används som växtskyddsmedel eller för att skydda hygienen eller folkhälsan).
Även spridningsmetoderna kan vara mycket lika, t.ex. sprids vissa insekticider för folkhälsoändamål enligt biociddirektivet genom flygbesprutning, precis som vissa växtskyddsmedel.
Vissa produkter för bekämpning av skadedjur används inomhus (t.ex. insektsmedel) och kan därför leda till att människor utsätts för direkt exponering.
Åtgärderna måste omfatta användning både i jordbruket och i annan verksamhet.
Ändringsförslag
20
2.
Detta direktiv skall tillämpas utan att det påverkar tillämpningen av annan närliggande gemenskapslagstiftning.
2.
Detta direktiv skall tillämpas utan att det påverkar tillämpningen av annan närliggande gemenskapslagstiftning eller eventuella nationella skatteåtgärder som främjar användningen av mindre skadliga bekämpningsmedel .
Motivering
Det måste vara upp till medlemsstaterna att främja en mer hållbar användning av bekämpningsmedel genom skatteåtgärder om de så önskar.
Ändringsförslag
21
2a.
Medlemsstaterna får bevilja bidrag eller vidta skatteåtgärder för att främja användningen av mindre skadliga växtskyddsmedel.
Motivering
Det måste vara upp till medlemsstaterna att främja en mer hållbar användning av bekämpningsmedel genom skatteåtgärder om de så önskar.
Ändringsförslag
22
2b.
Åtgärderna i detta direktiv får inte hindra medlemsstaterna från att tillämpa försiktighetsprincipen vid begränsning av eller förbud mot användningen av bekämpningsmedel.
Ändringsförslag
23
b) yrkesmässig användare: en fysisk eller juridisk person som använder bekämpningsmedel i sin yrkesmässiga verksamhet , inbegripet operatörer, tekniker, arbetsgivare, egenföretagare både inom och utanför jordbrukssektorn .
Till användarna hör även golfbanor, tennisbanor och andra fritidsanläggningar, allmänna parker och infrastrukturområden såsom parkeringsplatser, vägar, järnvägar och liknande.
Motivering
I den engelska texten används uttrycket ”professional user”.
Den tyska översättningen ”gewerblicher Anwender” är felaktig.
Direktivet bör inte rikta sig enbart till lant brukare utan också till alla andra som använder växtskyddsmedel.
Ändringsförslag
24
(d) rådgivare: en fysisk eller juridisk person som ger råd om användningen av bekämpningsmedel , inbegripet privata rådgivningsföretag, handelsagenter, livsmedelsproducenter och detaljhandlare om tillämpligt .
d) rådgivare: en fysisk eller juridisk person som besitter en av medlemsstaterna fastställd utbildningsnivå och som därigenom är behörig att ge råd om användningen av bekämpningsmedel och i det sammanhanget följer de metoder som är godkända i det land där bekämpningsmedlet tillverkas samt gemenskapens gränsvärden för bekämpningsmedelsrester .
Ändringsförslag
25
e) utrustning för spridning av bekämpningsmedel: en apparat som är särskilt utformad för spridning av bekämpningsmedel eller produkter som innehåller bekämpningsmedel.
e) utrustning för spridning av bekämpningsmedel: en apparat som används för spridning av bekämpningsmedel eller produkter som innehåller bekämpningsmedel.
Motivering
Apparaterna måste inte vara utformade enkom för att användas vid växtskyddet för att de ska kunna användas för sådana ändamål.
Därför behövs det en annan lydelse.
Ändringsförslag
26
g) flygbesprutning: all spridning av bekämpningsmedel med flygplan eller helikopter .
g) flygbesprutning: all spridning av bekämpningsmedel med luftfartyg .
Motivering
Den nuvarande definitionen av flygbesprutning omfattar inte alla möjligheter till spridning av bekämpningsmedel från luften.
Bekämpningsmedel kan spridas med andra luftfartyg än flygplan och helikoptrar.
Ändringsförslag
27
ia) icke-kemiska växtskydds- och odlingsmetoder: användning av bekämpnings- och växtskyddstekniker som inte baserar sig på kemiska egenskaper.
Icke-kemiska växtskydds- och odlingsmetoder inbegriper växelbruk, fysisk och mekanisk bekämpning och naturlig rovdjursbekämpning.
Motivering
Det enda fungerande sättet att undanröja bekämpningsmedlens negativa effekter för folkhälsan, djur, vilda djur och växter och miljön i allmänhet är att anta ett förebyggande och verkligen hållbart tillvägagångssätt genom att prioritera icke-kemiska växtskydds- och odlingsmetoder.
Detta skulle vara mer i linje med målen för hållbart växtskydd, eftersom beroendet av komplexa kemikalier avsedda att döda växter, insekter eller andra former av liv inte kan klassificeras som hållbart.
Ändringsförslag
28
ib) användningsfrekvens: indikator som visar hur många gånger jordbruksmark i genomsnitt får behandlas med den föreskrivna dosen och som beräknas baserat på sammanlagda försäljningsmängder av varje bekämpningsmedel.
Motivering
La fréquence de traitement ou la fréquence de l'application (FA) est calculée en divisant le volume vendu pour chaque produit particulier ou substance active par le dosage recommandé par hectare pour un usage particulier.
Les résultats de ces calculs pour chaque pesticide et récolte sont divisés par le nombre total d’hectares en culture.
,
SA est la quantité vendue de produit formulé individuel ou de substances actives par an.
SD est la dose standard définie pour chaque produit formulé individuel ou les substances actives pour chaque récolte/type de récolte (dose recommandée par l’Etat Membre ou si absent, dose recommandée par le fabricant).
AGRA est la surface totale des terres arables.
Ändringsförslag
29
(ic) bekämpningsmedel: växtskyddsmedel enligt förordning (EG) nr […] om utsläppande av växtskyddsmedel på marknaden.
Motivering
I texten refererar man ömsom till ”bekämpningsmedel”, ömsom till ”växtskyddsmedel”.
För att undvika oklarheter och garantera rättslig visshet är det viktigt att definiera termen ”bekämpningsmedel”.
Ändringsförslag
30
id) minskning av användningen: en minskning av spridningen av bekämpningsmedel som inte nödvändigtvis är beroende av volymen.
Motivering
This amendment brings the Directive in line with the objective of use reduction and clarifies that use reduction is not linked to a decrease in the volume of pesticides but rather to the decrease in the number or rate of applications to the levels necessary to crop protection.
Treatment frequency index is a reliable use indicator already in use in some Member States, including Denmark.
Ändringsförslag
31
ie) index för behandlingsfrekvens: indexet baserar sig på den fastställda standarddos av det verksamma ämnet per hektar som behövs för en behandling mot skadegöraren i fråga.
Därför är det inte nödvändigtvis beroende av volymen, och det kan användas för att utvärdera minskningen av användningen.
Motivering
This amendment brings the Directive in line with the objective of use reduction and clarifies that use reduction is not linked to a decrease in the volume of pesticides but rather to the decrease in the number or rate of applications to the levels necessary to crop protection.
Treatment frequency index is a reliable use indicator already in use in some Member States, including Denmark.
Ändringsförslag
32
Nationella handlingsplaner för att minska risker och beroendet av bekämpningsmedel
Nationella handlingsplaner för att minska risker och användningen av bekämpningsmedel
Ändringsförslag
33
-1.
Inom ett år efter detta direktivs ikraftträdande ska medlemsstaterna i enlighet med bilaga IIa anta en bakgrundsrapport i syfte att fastställa nationella trender när det gäller användning av bekämpningsmedel och risker samt de prioriterade områden och grödor som ska tas upp i den nationella handlingsplanen.
Ändringsförslag
34
1.
Medlemsstaterna skall anta nationella handlingsplaner för att fastställa mål , åtgärder och tidtabeller för minskning av risker , inbegripet faror, och beroendet av bekämpningsmedel.
1.
Medlemsstaterna skall senast ett år efter detta direktivs ikraftträdande och efter samråd med lantbruks-, vinodlar- och miljöorganisationer samt näringslivet och andra berörda sektorer anta nationella handlingsplaner för att fastställa mål och indikatorer för minskning av risker och användningen av bekämpningsmedel inom 5 år och 10 år från basåret.
EU:s mål ska vara att minska behandlingsfrekvensen med 25 procent inom 5 år från basåret och med 50 procent inom 10 år.
Medlemsstaterna ska fastställa sina nationella mål med beaktande av EU:s mål och befintliga nationella minskningsmål.
De nationella handlingsplanerna kan också omfatta regionala planer, i syfte att beakta särskilda lokala förhållanden .
Vid sidan om ett allmänt mål för minskad användning som anges i form av ett index för behandlingsfrekvens ska de nationella handlingsplanerna åtminstone omfatta specifika mål för minskad användning för följande ämnen:
a) För verksamma ämnen som inger mycket stora betänkligheter (enligt definitionen i artikel 57 i Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 om registrering, utvärdering, godkännande och begränsning av kemikalier (Reach) 1 ) ska minskningsmålet vara en minskning på minst 50 procent i förhållande till indexet för behandlingsfrekvens , beräknat för år 2005 , före utgången av 2013, om inte medlemsstaten kan bevisa att den redan har uppnått ett jämförbart eller högre mål baserat på ett annat referensår från perioden 1995–2004.
______
1 EUT L 396, 30.12.2006, s.
1.
Motivering
Genom detta ändringsförslag införs tydliga tidtabeller för utarbetandet av nationella handlingsplaner.
Dessutom är kvantitativa minskningsmål en viktig del av varje program för minskning av risker och användning.
Detta ändringsförslag klargör att det behövs tydliga indikatorer och mål i de nationella handlingsplanerna.
För att de nationella handlingsplanerna ska bli effektiva och realistiska måste de utarbetas i samarbete med berörda parter.
Det är viktigt att de negativa aspekterna i samband med användningen av bekämpningsmedel minimeras.
Dessutom är det viktigt att de nationella handlingsplanerna också får bygga på de mål som tagits med i ramdirektivet om vatten.
Ändringsförslag
35
De nationella handlingsplanerna ska omfatta integrerat växtskydd i den mening som avses i artikel 13 och ska ge företräde åt icke-kemiska växtskyddsåtgärder.
Motivering
Integrerat växtskydd bör stimuleras.
Ändringsförslag
36
När medlemsstaterna upprättar och ändrar sina nationella handlingsplaner skall de ta hänsyn till de planerade åtgärdernas sociala, ekonomiska och miljömässiga effekter.
Minimikrav för de nationella handlingsplanerna anges i det vägledande dokumentet i bilaga IIb.
Motivering
Genom ändringsförslaget kopplas de nationella handlingsplanerna till ramdirektivets bestämmelser.
Även konsekvenserna för folkhälsan kan studeras.
Det enda fungerande sättet att undanröja bekämpningsmedlens negativa effekter för människors och djurs hälsa och miljön är att anta ett förebyggande tillvägagångssätt tillsammans med en brett upplagd övergång till faktiskt hållbara icke-kemiska växtskydds- och odlingsmetoder.
Detta skulle vara mer i linje med målen för hållbart växtskydd.
Ändringsförslag
37
1a.
Basåret ska vara den genomsnittliga användningen och de genomsnittliga riskerna under de tre sista kalenderåren före detta direktivs ikraftträdande.
Motivering
Detta ändringsförslag klargör att det behövs tydliga indikatorer och mål i de nationella handlingsplanerna.
Ändringsförslag
38
1b.
De nationella handlingsplanerna ska i nödvändig utsträckning innehålla information om de aspekter som anges i artiklarna 5–13.
I dessa planer ska hänsyn tas till planer som upprättats enligt andra gemenskapsbestämmelser om användning av växtskyddsmedel, t.ex. åtgärdsplaner enligt direktiv 2000/60/EG.
Åtgärderna i de nationella handlingsplanerna får i synnerhet vara lagstiftningsåtgärder, skatteåtgärder eller frivilliga åtgärder som ska grundas på resultaten av relevanta riskbedömningar.
Motivering
I direktivet bör åtminstone minimikrav på innehållet anges, eller vilka aspekter som ska kontrolleras då planerna upprättas.
Frågan om när det krävs ytterligare lagstiftning, stödåtgärder, skatteåtgärder eller andra åtgärder bör avgöras av medlemsstaterna.
Ändringsförslag
39
1c.
De nationella handlingsplanerna ska omfatta integrerat växtskydd i den mening som avses i artikel 13 och ge företräde åt icke-kemiska växtskyddsåtgärder samt uppmuntra lant brukare som väljer att använda icke ‑kemiska växtskyddsmedel.
Ändringsförslag
40
1d.
Kommissionen ska vartannat år sammanställa en rapport med resultaten från genomförandet av de nationella handlingsplanerna.
Ändringsförslag
41
Motivering
En regelbunden översyn av de nationella handlingsplanerna och regler för ett integrerat växtskydd är avgörande för att användningen av bekämpningsmedel och dess risker verkligen ska kunna minskas.
Ändringsförslag
42
De nationella handlingsplanerna skall ses över minst vart femte år och alla ändringar av de nationella handlingsplanerna skall utan onödigt dröjsmål rapporteras till kommissionen.
De nationella handlingsplanerna skall ses över minst vart tredje år och uppdateras beroende på om målen uppnåtts.
Översynen ska även omfatta en analys av om riskerna i handlingsplanen har beaktats på lämpligt sätt eller om de måste omprövas.
Alla ändringar av de nationella handlingsplanerna och de viktigaste resultaten av översynen skall utan onödigt dröjsmål rapporteras till kommissionen.
Kommissionen ska upprätta en Internetportal genom vilken allmänheten informeras om de nationella handlingsplanerna, eventuella ändringar och väsentliga resultat av genomförandet.
Motivering
En regelbunden översyn av de nationella handlingsplanerna och genomförandet av grödspecifikt integrerat växtskydd är grundläggande för att man ska kunna minska användningen och riskerna.
Bestämmelserna om översynen måste preciseras.
På grund av de olika lokala förhållanden som gäller för användningen av växtskyddsmedel bör också regionala planer beaktas.
Allmänhetens medverkan är en väsentlig del av de nationella handlingsplanerna.
Därför är det lämpligt att göra planer, ändringar och resultat av genomförandet tillgängliga genom en Internetportal.
Ändringsförslag
43
3.
Kommissionen skall göra all relevant information som meddelas i enlighet med punkt 2 tillgänglig för tredjeländer.
3.
Kommissionen skall göra all information som meddelas i enlighet med punkt 2 tillgänglig för tredjeländer och för allmänheten .
Motivering
Allmänheten har rätt att vara informerad i frågor som rör dess hälsa och miljön och bör vara fullt involverad i utarbetandet, utvecklingen, genomförandet, övervakningen och ändringen av de nationella handlingsplanerna och deras mekanismer i linje med andan i direktiv 2003/35/EG, där det föreskrivs om allmänhetens deltagande.
Informationen om de nationella handlingsplanerna bör göras tillgänglig via Internet på Europeiska kommissionens webbplats.
Ändringsförslag
44
3a.
Medlemsstaterna ska på en webbplats offentliggöra den information som meddelas enligt punkt 2.
Motivering
Av tydlighets- och insynsskäl bör allmänheten ha tillgång till denna typ av information, vilket även gör det möjligt för allmänheten att delta vid utarbetandet samt omprövning och övervakning av de nationella handlingsplanerna.
Ändringsförslag
45
4.
De bestämmelser om allmänhetens deltagande som anges i artikel 2 i direktiv 2003/35/EG skall tillämpas vid utarbetande och ändring av de nationella handlingsplanerna.
4.
De bestämmelser om allmänhetens deltagande som anges i artikel 2 i direktiv 2003/35/EG skall tillämpas vid utarbetande av den nationella bakgrundsrapporten, samt vid utarbetande och ändring av de nationella handlingsplanerna.
Alla berörda parter och den bredare allmänheten ska rådfrågas om alla aspekter av den nationella bakgrundsrapporten och de nationella handlingsplanerna, inbegripet utarbetande, utveckling, genomförande, mekanismer, övervakning och ändringar.
En balanserad representation av berörda parter, inbegripet dem som utsätts för negativa effekter till följd av användningen, ska säkerställas.
Motivering
Ändringsförslaget syftar till att säkerställa allmänhetens deltagande i utarbetandet av de nationella bakgrundsrapporterna och de nationella handlingsplanerna i enlighet med direktiv 2003/35/EG, där det föreskrivs om allmänhetens deltagande.
Ändringsförslag
46
4a.
Medlemsstaterna ska införa en finansieringsmekanism för genomförandet av de nationella handlingsplanerna , vilken bekostas via system med skatt eller avgifter på bekämpningsmedel.
Motivering
Skatte- och avgiftssystem har visat sig vara ett bra sätt att minska bekämpningsmedlen i vissa europeiska länder.
Sådana system bör införas i hela EU och bör kunna finansiera åtgärderna för att minska riskerna och användningen av bekämpningsmedel inom ramen för de nationella handlingsplanerna samt ett effektivt system för övervakning och information om planernas resultat.
Medlemsstaterna bör kunna välja det finansieringssystem som passar landets behov bäst.
Ändringsförslag
47
4b.
Medlemsstaterna ska öka sina ansträngningar att begränsa och förebygga olaglig användning av växtskyddsmedel, i samarbete med berörda parter.
Medlemsstaterna ska regelbundet rapportera om befintliga kontroller avseende olaglig användning.
Motivering
En grundläggande förutsättning för hållbar användning av växtskyddsmedel är att befintliga rättsliga krav tillämpas och efterlevs till fullo.
Nationella myndigheter bör därför noggrannare kontrollera att befintlig lagstiftning efterlevs och effektivare tillämpa befintliga krav på övervakning och efterlevnad.
Ändringsförslag
48
1.
Medlemsstaterna skall se till att alla yrkesmässiga användare, distributörer och rådgivare har tillgång till lämplig utbildning.
1.
Medlemsstaterna skall se till att alla yrkesmässiga användare, distributörer och rådgivare har tillgång till lämplig fristående utbildning eller fortbildning som inbegriper regelbunden uppdatering när det gäller ny tillgänglig information om hållbar och korrekt användning av växtskyddsmedel och som motsvarar de berördas ansvarsnivå och deras specifika roll inom integrerat växtskydd .
Därför ska minimikrav för denna utbildning och fortbildning införas på gemenskapsnivå.
Motivering
I många fall beror förorening av miljön och jordbruksprodukter med bekämpningsmedel på bristande sakkunskap.
Yrkesmässiga användare, distributörer och rådgivare bör uppdateras med den relevanta information som finns att tillgå.
Det är mycket viktigt att utbildning anordnas oberoende av vissa aktörers ekonomiska intressen.
Detta utesluter dock inte möjligheten att anlita sakkunniga från industrin eller icke-statliga organisationer.
Medlemsstaterna kan även uppfylla grundkraven enligt detta direktiv genom att erbjuda relevant utbildning.
När det gäller personer som redan har motsvarande utbildning kan det räcka med fördjupade studier av enskilda aspekter.
Minimikrav ger ökad kvalitet på utbildningen och underlättar informationsutbytet mellan olika användare i medlemsstaterna.
Ändringsförslag
49
Utbildningen skall vara utformad på ett sådant sätt att den ger tillräcklig kunskap om de ämnen som anges i bilaga I.
Utbildningen eller fortbildningen skall vara utformad på ett sådant sätt att den ger tillräcklig kunskap om de ämnen som anges i bilaga I.
Motivering
Medlemsstaterna bör även bidra till att de grundläggande kraven i detta direktiv uppfylls genom tillhandahållande av motsvarande utbildning och fortbildning.
När det gäller personer som redan har motsvarande utbildning kan det räcka med fördjupade studier av enskilda aspekter.
Ändringsförslag
50
1a.
Medlemsstaterna ska se till att yrkesmässiga användare, distributörer och rådgivare är medvetna om förekomsten av och riskerna med olagliga (förfalskade) växtskyddsmedel, och att de får lämplig utbildning för att kunna identifiera sådana produkter.
Motivering
Förfalskningar och olaglig handel med växtskyddsmedel inom EU är ett stort problem.
Det är viktigt att göra yrkesmässiga användare och distributörer medvetna om detta när det gäller att hantera problemet med olaglig handel med växtskyddsmedel.
Ändringsförslag
51
2.
2.
Motivering
Ändringsförslaget läggs fram eftersom tidsfristen måste vara förenlig med den tidsfrist som gäller vid upprättandet av de nationella handlingsplanerna.
Ändringsförslaget gör det möjligt att fastställa villkoren för utfärdande och tillbakadragande av intygen.
Ändringsförslag
52
3.
3.
Motivering
Medlemsstaterna bör även bidra till att de grundläggande kraven i detta direktiv uppfylls genom tillhandahållande av motsvarande utbildning och fortbildning.
När det gäller personer som redan har motsvarande utbildning kan det räcka med fördjupade studier av enskilda aspekter.
Ändringsförslag
53
Innehavarna av de intyg som avses i bilaga 1 ska delta i fortbildningsåtgärder när ansvariga nationella myndigheter anser detta vara nödvändigt.
Ändringsförslag
54
1.
1.
Intyget får vara högst 7 år gammalt.
Motivering
(661 tecken) Distributörer som säljer växtskyddsmedel måste vidta tillräckliga åtgärder för att se till att kunderna vid försäljning får tillräcklig information om korrekt användning, eventuella risker, korrekt lagring, hantering, spridning samt bortskaffande av växtskyddsmedel.
Pesticides users should be aware of the health risks of their use.
Therefore information must be provided at the point of sale, and not only in relation to those pesticides classified as toxic or very toxic, as all pesticides are deliberately designed to be toxic and so can pose hazards for human health.
Therefore, anyone who purchases pesticides, as well as those who use them, whether professional or non-professional, must be made aware of the risks and potential adverse health impacts of pesticide use.
Ändringsförslag
55
2.
2.
Ändringsförslag
56
3.
Medlemsstaterna skall ålägga distributörer som släpper ut bekämpningsmedel för icke yrkesmässig användning på marknaden att lämna allmän information om riskerna med bekämpningsmedelsanvändning, särskilt om faror, exponering, korrekt lagring, hantering och spridning samt bortskaffande.
3.
Medlemsstaterna skall ålägga distributörer som släpper ut bekämpningsmedel för icke yrkesmässig användning på marknaden att lämna allmän information om riskerna med och de möjliga negativa hälso- och miljöeffekterna av bekämpningsmedelsanvändning, särskilt om faror, exponering, korrekt lagring, hantering och spridning samt bortskaffande.
Detta gäller också för försäljning via Internet.
Motivering
Distributörer som säljer bekämpningsmedel måste vidta tillräckliga åtgärder för att se till att kunderna vid försäljning får tillräcklig information om korrekt användning, eventuella risker, korrekt lagring, hantering, spridning samt bortskaffande av bekämpningsmedel.
Både yrkesmässiga och icke yrkesmässiga användare av bekämpningsmedel måste vara fullt informerade om riskerna med och de möjliga negativa hälso- och miljöeffekterna av bekämpningsmedelsanvändning.
Ändringsförslag
57
Motivering
Åtgärderna bör i stället fastställas inom två år.
Ändringsförslag
58
3a.
Medlemsstaterna ska se till att befintliga åtgärder för inspektion och efterlevnadskontroll genomförs fullt ut för att säkerställa att olagliga (förfalskade) bekämpningsmedel inte saluförs.
Motivering
Bättre efterlevnadskontroll beträffande befintlig lagstiftning är grundläggande när det gäller att ta itu med problemet med förfalskning av och olaglig handel med bekämpningsmedel.
Ändringsförslag
59
Artikel 7
Informationsprogram
Informationsprogram , övervakning och forskning
Medlemsstaterna skall stödja informationsprogram riktade till allmänheten och underlätta allmänhetens tillgång till information om bekämpningsmedel, särskilt när det gäller hälso- och miljöeffekter och icke-kemiska alternativ.
1.
Medlemsstaterna skall stödja informationsprogram riktade till allmänheten och underlätta allmänhetens tillgång till information om riskerna med bekämpningsmedelsanvändning och möjliga akuta och kroniska hälso- och miljöeffekter till följd av bekämpningsmedelsanvändning.
Allmänheten ska även förses med information om den roll som bekämpningsmedel spelar i jordbruk och livsmedelsproduktion , om ansvarsfull användning av bekämpningsmedel, om faror och om icke-kemiska alternativ.
1a.
Medlemsstaterna ska upprätta bindande system för insamling av information om akuta och kroniska fall av bekämpningsmedelsförgiftning, särskilt bland bekämpningsmedelsoperatörer, arbetare, boende och alla andra befolkningsgrupper som riskerar att regelbundet exponeras för bekämpningsmedel.
1b.
Medlemsstaterna ska regelbundet övervaka och samla in information om indikatorarter som exponerats för bekämpningsmedel och om bekämpningsmedel i miljön, såsom i söt - och havsvatten, mark och luft, och regelbundet rapportera om denna information till kommissionen.
1c.
Medlemsstaterna ska genomföra långsiktiga forskningsprogram rörande specifika situationer där bekämpningsmedel har förknippats med effekter på människors hälsa och miljön, inbegripet studier om högriskgrupper, biologisk mångfald och kombinerade effekter.
1d.
I syfte att öka informationens jämförbarhet ska kommissionen i samarbete med medlemsstaterna inom tre år efter det att detta direktiv har trätt i kraft utveckla ett strategiskt vägledande dokument om övervakning och kartläggning av bekämpningsmedelsanvändningens effekter på människors hälsa och miljön.
Motivering
Genom ändringsförslaget ser man till att de planerade informationsprogrammen riktade till allmänheten inte bara tar upp riskerna med användning av bekämpningsmedel.
För närvarande är det i första hand riskerna med bekämpningsmedel som tas upp offentligt.
Man borde även sträva efter att objektivt redogöra för bekämpningsmedelsanvändningens nödvändighet och hållbarhet samt för dess betydelse inom dagens livsmedelsproduktion, såsom det anges i ändringsförslaget.
Informationsprogrammen bör också omfatta bekämpningsmedlens kroniska hälsoeffekter.
I medlemsstaterna måste det bedrivas övervakning och forskning för att man ska kunna samla in information och beräkna bekämpningsmedlens hälso- och miljöeffekter.
Ett rapporteringssystem finns redan i EU när det gäller bekämpningsmedelsrester i livsmedel, men det finns inget system för att övervaka förgiftningsfall och miljöeffekter som förorsakats av bekämpningsmedel.
Ändringsförslag
60
1.
Medlemsstaterna skall se till att utrustning och tillbehör för spridning av bekämpningsmedel i yrkesmässig användning inspekteras med jämna mellanrum.
1.
Medlemsstaterna skall se till att utrustning och tillbehör för spridning av bekämpningsmedel i yrkesmässig användning blir föremål för obligatoriska inspektioner med jämna mellanrum , minst vart femte år .
Motivering
Ett maximalt tidsintervall för kontroll av besprutningsutrustning måste fastställas.
Det är oerhört viktigt att bekämpningsmedel hanteras under betryggande former.
Kravet på obligatoriska inspektioner gör det möjligt att övervaka genomförandet av direktivet, framför allt inom området säkerhet.
Ändringsförslag
61
3.
3.
Obligatoriska inspektioner ska därefter äga rum minst vart femte år .
Motivering
I kommissionens förslag behandlas denna fråga inte alls.
Ändringsförslag
62
5.
5.
Motivering
Detta ändringsförslag är nödvändigt i syfte att anpassa texten till bestämmelserna i det nya beslutet om kommittéförfarandet.
Ändringsförslag
63
3.
Medlemsstaterna skall utse de myndigheter som är behöriga att medge undantag och skall informera kommissionen om detta.
3.
Medlemsstaterna skall utse de myndigheter som är behöriga att övervaka flygbesprutningar och skall informera kommissionen om detta.
Ändringsförslag
64
4.
Undantag får medges endast om följande villkor är uppfyllda:
4.
Undantag får medges endast om följande villkor är uppfyllda:
(a) Det får inte finnas några lämpliga alternativ, eller också skall det innebära klara fördelar i form av minskad påverkan på hälsa och miljö jämfört med markbaserad spridning av bekämpningsmedel.
(a) Det får inte finnas några lämpliga alternativ, eller också skall det innebära klara fördelar i form av minskad påverkan på människors hälsa och på miljön jämfört med markbaserad spridning av bekämpningsmedel.
(b) De bekämpningsmedel som används skall vara uttryckligen tillåtna för flygbesprutning.
(b) De bekämpningsmedel som används skall vara uttryckligen tillåtna för flygbesprutning ; ämnen som klassificeras som mycket giftiga (R50) för vattenorganismer ska inte tillåtas för flygbesprutning .
(ca) Flygbesprutning ska meddelas i förväg till behörig myndighet och godkännas av denna.
I tillståndet skall anges vilka åtgärder som är nödvändiga för att varna boende och andra närvarande personer och för att skydda miljön i närheten av det besprutade området.
(cb) Alla nödvändiga åtgärder ska vidtas för att i god tid varna boende och andra närvarande personer och för att skydda miljön i närheten av det besprutade området.
(cc) Det område som ska besprutas får inte ligga i närheten av allmänna områden eller bostadsområden, och boendes eller andra närvarande personers hälsa får inte påverkas.
(cd) Luftfartyget ska vara utrustat med bästa tillgängliga teknik för att minska vindavdrift (t.ex. avdriftsreducerande munstycken); vid användning av helikoptrar ska helikopterns sprutbommar vara försedda med injektionsmunstycken för att minska vindavdriften.
(ce) De sociala, ekonomiska och miljömässiga fördelarna ska uppväga de möjliga effekterna på boendes och andra närvarande personers hälsa.
Motivering
Flygbesprutning är i vissa situationer och områden och i fråga om vissa grödor (växternas höjd, angripna områden, epidemier) nödvändig som spridningsteknik.
Målet bör vara att införa obyråkratiska och hanterliga bestämmelser för flygbesprutning.
Särskilt i krissituationer måste man reagera snabbt på akuta skadegörarangrepp.
Man bör iaktta särskild varsamhet när ämnen tillåts för flygbesprutning.
Ändringsförslag
65
5.
En yrkesmässig användare som vill sprida bekämpningsmedel genom flygbesprutning skall lämna in en begäran till den behöriga myndigheten tillsammans med uppgifter som styrker att de villkor som anges i punkt 4 är uppfyllda.
5.
En yrkesmässig användare som vill sprida bekämpningsmedel genom flygbesprutning skall lämna in en begäran till den behöriga myndigheten tillsammans med uppgifter som styrker att de villkor som anges i punkt 4 är uppfyllda.
Anmälan ska innehålla information om besprutningstiden och om de mängder och typer av bekämpningsmedel som sprids.
Motivering
Allmänheten bör vara fullt informerad om besprutningstiden och om de mängder och typer av bekämpningsmedel som sprids för att kunna skydda sig mot exponeringsrisken.
Ändringsförslag
66
6.
De behöriga myndigheterna skall föra register över de undantag som medges.
6.
De behöriga myndigheterna skall föra register över de undantag som medges och göra dem tillgängliga för allmänheten .
Motivering
Allmänheten bör ha tillgång till information, och de behöriga myndigheterna bör göra informationen tillgänglig.
(Frédérique Ries)
Ändringsförslag
67
Artikel 9a (ny)
Artikel 9a
Markspridning
Lantbrukarna ska före användning av produkten informera eventuella grannar som kan exponeras för vindavdriften och som har begärt att bli informerade genom ett centraliserat informations- eller signalsystem.
Motivering
I den föregående artikeln om flygbesprutning anges bestämmelser med syfte att varna boende och andra närvarande personer.
Liknande bestämmelser bör fastställas för markspridning för att de boende ska varnas.
Numreringen ändras framöver.
Ändringsförslag
68
1.
Medlemsstaterna skall, om bekämpningsmedel används i närheten av vatten, se till att företräde ges åt
1.
Medlemsstaterna skall, om bekämpningsmedel används i närheten av vatten , särskilt förekomster av dricksvatten , se till att företräde ges åt
Motivering
Vattendrag som används som dricksvattentäkter är av grundläggande betydelse för samhället, och därför bör dessa vattendrag särskilt skyddas.
Ändringsförslag
69
(a) produkter som inte är farliga för vattenmiljön,
(a) produkter för vilka risken att hamna i vattenmiljön inte är stor ,
Motivering
Särskilt bör vattenförekomster som används som dricksvattentäkter skyddas för att man ska kunna uppnå målen i artikel 7 i ramdirektivet för vatten, som berör skyddet av vattenförekomster som används som dricksvattentäkter, samt värdet 0,1 mikrogram/liter, som fastställts i direktivet om dricksvatten.
Ändringsförslag
70
2.
2.
Motivering
Buffertzonerna bör vara minst 10 meter breda för att garantera ett allmänt minimiskydd för vattendrag och vattenförekomster.
Även om buffertzoner är nödvändiga räcker de ändå inte till för att lösa problemet med de olika vägar genom vilka bekämpningsmedlen hamnar i vatten.
De kommer inte nödvändigtvis att förebygga läckage genom dräneringsdiken eller ytavrinning, som är en av de främsta vägarna.
Ändringsförslag
71
Buffertzonernas omfattning skall fastställas på grundval av riskerna för förorening och det aktuella områdets jordbruksförhållanden .
Buffertzonernas omfattning skall fastställas på grundval av riskerna för förorening och det aktuella områdets jordbruks- och klimatförhållanden .
Motivering
Inte endast jordbruksförhållandena utan även klimatförhållandena bör tas i betraktande.
Ändringsförslag
72
Motivering
Buffertzonerna bör vara minst 10 meter breda för att garantera ett allmänt minimiskydd för vattendrag och vattenförekomster.
Även om buffertzoner är nödvändiga räcker de ändå inte till för att lösa problemet med de olika vägar genom vilka bekämpningsmedlen hamnar i vatten.
De kommer inte nödvändigtvis att förebygga läckage genom dräneringsdiken eller ytavrinning, som är en av de främsta vägarna.
Ändringsförslag
73
3.
3.
Medlemsstaterna skall se till att lämpliga åtgärder vidtas för att begränsa vindavdrift och långväga transport av bekämpningsmedel, åtminstone i högväxande grödor, inbegripet odlingar av frukt, vin och humle, i direkt anslutning till eller i närheten av ett vattendrag , genom att se till att användning av bekämpningsmedel i sådana områden förbjuds och icke-kemiska alternativ används .
Motivering
Bekämpningsmedel har visat sig spridas över avsevärda avstånd vilket kan resultera i att vattendrag riskerar att förorenas genom ett antal olika källor.
I syfte att undvika förorening av vattenmiljön bör man därför införa kraftfulla åtgärder.
Ändringsförslag
74
4.
4.
Medlemsstaterna skall se till att spridning av bekämpningsmedel begränsas så långt som möjligt eller undviks helt på och längs vägar, järnvägslinjer, genomsläpplig mark, sluttningar och annan infrastruktur nära ytvatten eller grundvatten, och på hårdgjorda ytor med hög risk för avrinning till ytvatten eller avloppssystem.
I alla dessa områden ska användning av icke-kemiska alternativ främjas .
Motivering
I porösa jordarter tränger olika ämnen och avloppsvatten lätt ned i djupare liggande jordlager.
Exempelvis på sandjordar tränger ämnen som är lösta i vatten lättare ned i djupare liggande jordlager, till skillnad från hur det förhåller sig på lerjordar, som är föga genomsläppliga.
Branta sluttningar underlättar utsköljning och avrinning framför allt efter häftiga regn, så att markpartiklar tillsammans med de gödnings- och växtskyddsmedel inklusive bekämpningsmedel som använts sprids till jordbruksmarker längre ned på sluttningarna eller till ytvatten.
I syfte att helt undvika förorening av dessa områden bör icke-kemiska alternativ användas.
Ändringsförslag
75
(a) Användning av bekämpningsmedel skall förbjudas eller begränsas till det absolut nödvändiga i områden som används av allmänheten eller av känsliga befolkningsgrupper, åtminstone parker, offentliga trädgårdar, sportanläggningar och lekplatser.
(a) Användning av bekämpningsmedel skall förbjudas i alla områden som används av allmänheten eller av känsliga befolkningsgrupper, åtminstone i bostadsområden, parker, offentliga trädgårdar, idrotts- och fritidsområden, skolgårdar och lekplatser samt i närheten av anläggningar för allmän sjukvård (kliniker, sjukhus, rehabiliteringscenter, hälsohem, vårdhem), och även i omfattande zoner – också kring ovannämnda områden – där besprutning ska vara förbjuden, framför allt, men inte enbart, för att skydda känsliga befolkningsgrupper, såsom spädbarn, barn, gravida kvinnor, äldre personer och personer som sedan tidigare har problem med hälsan och eventuellt går på medicin .
Motivering
Besprutning bör vara förbjuden i sådana områden som används av allmänheten, framför allt av känsliga befolkningsgrupper, såsom barn, i likhet med de regler som antagits exempelvis för gräsmattor i Kanada.
I andra känsliga områden bör besprutning vara förbjuden eller strikt begränsad.
Kring områden som används av allmänheten och framför allt av känsliga befolkningsgrupper bör det inrättas omfattande zoner där besprutning är förbjuden.
Kring skolor kan dessa zoner vara upp till fyra kilometer breda, såsom fallet är på vissa håll i Förenta staterna.
Idrottsområden fungerar ofta också som fritidsområden.
Semester- och fritidsanläggningar tjänar också idrottens behov.
Sådana platser bör vara fria från föroreningar, och de människor som vistas där bör inte exponeras för bekämpningsmedel.
Platser med anläggningar för allmän sjukvård (kliniker, sjukhus, sanatorier, rehabiliteringscenter, vårdhem etc.) bör skyddas från bekämpningsmedels skadliga inverkan.
Alla till buds stående medel bör användas för att inte allmänheten i onödan ska exponeras för bekämpningsmedel.
Ändringsförslag
76
(b) Användning av bekämpningsmedel skall förbjudas eller begränsas i särskilda bevarandeområden och andra områden som utsetts i syfte att fastställa nödvändiga bevarandeåtgärder enligt artiklarna 3 och 4 i direktiv 79/409/EEG och artiklarna 6, 10 och 12 i direktiv 92/43/EEG.
(b) Användning av bekämpningsmedel skall förbjudas eller strikt begränsas i bevarandeområden och andra områden som utsetts i syfte att fastställa nödvändiga bevarandeåtgärder enligt artiklarna 3 och 4 i direktiv 79/409/EEG och artiklarna 6, 10 och 12 i direktiv 92/43/EEG.
Motivering
Ändringsförslag
77
b) Användning av bekämpningsmedel skall förbjudas eller begränsas i särskilda bevarandeområden och andra områden som utsetts i syfte att fastställa nödvändiga bevarandeåtgärder enligt artiklarna 3 och 4 i direktiv 79/409/EEG och artiklarna 6, 10 och 12 i direktiv 92/43/EEG.
Ett förbud eller en begränsning enligt b får grundas på resultaten av relevanta riskbedömningar.
Ett förbud eller en begränsning ska grundas på resultaten av relevanta riskbedömningar.
Motivering
Det är viktigt att man verkligen kontrollerar känsliga områden (med tanke på vilda växter och djur eller känsliga grupper, såsom barn) för att se om användningen av bekämpningsmedel bör minskas eller till och med förbjudas.
Man måste bestämma detta från fall till fall och utifrån en riskbedömning.
Ändringsförslag
78
1.
Medlemsstaterna skall vidta de åtgärder som behövs för att säkerställa att följande arbetsmoment inte medför risk för människors hälsa eller säkerhet eller för miljön:
1.
Medlemsstaterna skall inom ramen för de nationella handlingsplanerna vidta de åtgärder som enligt relevanta riskbedömningar behövs för att säkerställa att följande arbetsmoment utförda av användare inte medför risk för människors hälsa eller säkerhet eller för miljön:
(a) Lagring, hantering, utspädning och blandning av bekämpningsmedel före spridning.
(a) Säker lagring, hantering, utspädning och blandning av bekämpningsmedel före spridning.
(b) Hantering av förpackningar för och rester av bekämpningsmedel.
(b) Säker hantering av förpackningar för och rester av bekämpningsmedel.
(c) Behandling av kvarvarande vätskor efter spridning.
(c) Behandling av kvarvarande vätskor efter spridning.
(d) Rengöring av utrustning som använts för spridning.
(d) Iordningställande, hantering, rengöring och lagring av utrustning som använts för spridning samt tillbehör, bland annat kemikalier och utrustning för besprutning .
Motivering
Det är nödvändigt med korrekt hantering och säker lagring av avfall från bekämpningsmedel för att man ska kunna minimera riskerna för förorening med bekämpningsmedel.
De föreslagna åtgärderna bör integreras i de nationella handlingsplanerna.
Det är främst fråga om att de befintliga bestämmelserna genom ändamålsenliga insatser ska genomföras i praktiken.
Det finns gott om föreskrifter i medlemsstaterna.
Det bör klargöras att kommissionens föreslagna åtgärd är utan betydelse för privat användning.
Ändringsförslag
79
3.
3.
Medlemsstaterna skall inom ramen för de nationella handlingsplanerna vidta de åtgärder som enligt relevanta riskbedömningar behövs för att man ska kunna se till att lagringsplatser för bekämpningsmedel utformas på ett sådant sätt att oönskade utsläpp undviks.
Motivering
Se motiveringen till ändringsförslag 46.
Ändringsförslag
80
1.
Medlemsstaterna skall vidta alla åtgärder som behövs för att främja jordbruk med små insatser av bekämpningsmedel, däribland integrerat växtskydd, och för att säkerställa att yrkesmässiga användare av bekämpningsmedel går över till en mer miljövänlig användning av alla tillgängliga växtskyddsåtgärder, företrädesvis lågriskalternativ om sådana kan användas och i annat fall produkter som, av de produkter som är tillgängliga för samma skadegörarproblem, ger minst påverkan på människors hälsa och på miljön.
1.
Medlemsstaterna skall vidta alla åtgärder , bland dem också ekonomiska styrmedel, som behövs för att främja jordbruk med små insatser av bekämpningsmedel, däribland integrerat växtskydd, och för att säkerställa att yrkesmässiga användare av bekämpningsmedel så snart som möjligt går över till en mer miljövänlig användning av alla tillgängliga växtskyddsåtgärder, företrädesvis lågriskalternativ om sådana kan användas och i annat fall produkter som, av de produkter som är tillgängliga för samma skadegörarproblem, ger minst påverkan på människors hälsa och på miljön.
Kommissionen ska lägga fram ett förslag om ett gemenskapsomfattande system för bekämpningsmedelsskatt.
Motivering
Ekonomiska styrmedel brukar vara det effektivaste sättet att minska riskerna för miljön.
Med hjälp av ett gemenskapsomfattande system för bekämpningsmedelsskatt går det att åstadkomma balans på marknaden för bekämpningsmedel inom EU och förebygga olaglig handel.
Det är viktigt att yrkesmässiga användare av bekämpningsmedel så snart som möjligt går över till en mer miljöriktig användning av de olika växtskyddsåtgärder som finns att tillgå.
Ändringsförslag
81
1a.
Motivering
Medlemsstaterna ska främja en mer hållbar och miljövänlig användning av bekämpningsmedel.
Det är dessutom viktigt att det finns en tydligare koppling mellan detta direktiv och förslaget till förordning om utsläppande av växtskyddsmedel på marknaden.
Ändringsförslag
82
2.
2.
Medlemsstaterna skall skapa eller stödja skapandet av alla nödvändiga förutsättningar för tillämpning av integrerat växtskydd och icke-kemiska växtskydds- och odlingsmetoder, och för varje enskild gröda beskriva bästa praxis för integrerat växtskydd , varvid icke-kemiska växtskyddsåtgärder ska ges företräde .
Motivering
EU Directive 91/414/EEC requires that a pesticide shall not be approved unless it has been established that there will be “no harmful effect” on humans or animals.
Priority should be given to non-chemical and natural methods of pest management as the only truly preventative and sustainable solution which is obviously more in line with the objectives for sustainable crop protection, than the reliance on complex chemicals designed to kill plants, insects or other forms of life, which cannot be classified as sustainable.
Member States need to promote and encourage the widespread adoption of non-chemical alternatives to plant protection.
Bästa praxis för icke-kemiska växtskyddsåtgärder hjälper yrkesmässiga användare att välja miljöriktigt i fråga om växtskydd och växtskyddsmedel.
Ändringsförslag
83
3.
3.
Medlemsstaterna skall särskilt se till att lantbrukare har tillgång till system, inbegripet utbildning enligt artikel 5, och verktyg för övervakning av skadegörare och för beslutsfattande samt till rådgivningstjänster om icke-kemiska växtskydds- och odlingsmetoder .
Motivering
Se motiveringen till artikel 13.1 och 13.2.
Ändringsförslag
84
4.
4.
Medlemsstaterna skall, senast den 30 juni 2011 , rapportera till kommissionen om genomförandet av punkterna 2 och 3 och särskilt om huruvida de nödvändiga förutsättningarna för tillämpning av integrerat växtskydd finns.
Motivering
Standarderna för integrerat växtskydd bör tillämpas snabbare än vad kommissionen föreskrivit.
Ändringsförslag
85
4a.
Minimikraven för utveckling av allmänna och grödspecifika standarder för integrerat växtskydd fastställs i bilaga IIc.
Ändringsförslag
86
5.
5.
Motivering
Det ska skapas enhetliga kriterier i EU för god yrkespraxis inom växtskydd och för ett integrerat växtskydd.
Kriterierna i fråga anges närmare i bilaga IIc, i syfte att underlätta genomförandet i medlemsstaterna.
Anpassningar till den vetenskapliga och tekniska utvecklingen bör göras i enlighet med bestämmelserna i det nya beslutet om kommittéförfarandet.
Ändringsförslag
87
6.
6.
Medlemsstaterna skall införa lämpliga incitament , också åtgärder för utbildning och finansiering, för att stödja användare när det gäller att tillämpa gröd- eller sektorspecifika riktlinjer för integrerat växtskydd vilka tar hänsyn till de allmänna kriterier som anges i bilaga IIc.
Sådana riktlinjer får också utarbetas av organisationer för yrkesmässiga användare.
Medlemsstaterna ska i sina nationella handlingsplaner enligt artikel 4 hänvisa till lämpliga riktlinjer .
Motivering
Det ska skapas enhetliga kriterier i EU för god yrkespraxis inom växtskydd och för ett integrerat växtskydd.
Kriterierna i fråga anges närmare i bilaga IIc, i syfte att underlätta genomförandet i medlemsstaterna.
Anpassningar till den vetenskapliga och tekniska utvecklingen bör göras i enlighet med bestämmelserna i det nya beslutet om kommittéförfarandet.
Utbildningsprogram och tillräckligt ekonomiskt stöd är en förutsättning för integrerat växtskydd och ekologiskt jordbruk.
Ändringsförslag
88
7.
7.
De allmänna standarderna för integrerat växtskydd skall utarbetas i enlighet med det förfarande som anges i artikel 52 i förordning (EG) nr […] , under offentligt deltagande från berörda parters sida .
Motivering
Deltagandet är av vikt med tanke på att standarderna för integrerat växtskydd allmänt ska accepteras.
Ändringsförslag
89
8a.
I syfte att införa grödspecifika metoder inom ramen för integrerat växtskydd och bidra till utvecklingen av ekologiskt jordbruk ska medlemsstaterna inrätta ett lämpligt finansieringssystem som bygger på beskattning av bekämpningsmedel.
Motivering
Skatter har visat sig vara ett bra sätt att minska användningen av bekämpningsmedel i ett antal av EU:s medlemsstater.
Medlemsstaterna måste kunna välja det lämpligaste skattesystemet efter behov.
Ändringsförslag
90
1.
Medlemsstaterna får, fram till dess att indikatorerna har fastställts, fortsätta att använda befintliga nationella indikatorer eller fastställa andra lämpliga indikatorer.
1.
Det ska råda krav på att allmänheten, vid sidan om alla andra berörda parter, deltar i utarbetandet och fastställandet av nationella indikatorer.
Detta förutsätter också att allmänheten får obegränsad tillgång till information för att kunna delta .
Motivering
Detta ändringsförslag är nödvändigt i syfte att anpassa texten till bestämmelserna i det nya beslutet om kommittéförfarandet.
Användningsindikatorer och mål i fråga om användningen bör fastställas vid sidan om riskindikatorer och mål i fråga om riskerna.
Det måste göras klart för medlemsstaterna att de nationella indikatorerna ska stå i förhållande till de risker för både hälsa och miljö som användningen av bekämpningsmedel innebär.
Det måste också göras klart för medlemsstaterna vilka krav som gäller i fråga om allmänhetens deltagande då de nationella indikatorerna utarbetas och fastställs samt då de tillämpas och ändras, för att man i detta sammanhang ska följa andan i direktiv 2003/35/EG om allmänhetens deltagande.
Ändringsförslag
91
a) Beräkning av gemensamma och harmoniserade riskindikatorer på nationell nivå.
a) Beräkning av gemensamma och harmoniserade risk- och användningsindikatorer på nationell nivå.
Ändringsförslag
92
Motivering
Man bör även fokusera på ovannämnda frågor eftersom också dessa frågor påverkar riskindikatorerna för användningen av växtskyddsmedel.
Ändringsförslag
93
c) Fastställande av prioriterade verksamma ämnen, prioriterade grödor, ohållbara metoder som kräver särskild uppmärksamhet eller goda metoder som kan användas som förebilder för att uppnå målen för detta direktiv när det gäller att minska risker och beroendet av växtskyddsmedel .
c) Fastställande av prioriterade verksamma ämnen, prioriterade grödor, ohållbara metoder som kräver särskild uppmärksamhet eller goda metoder som kan användas som förebilder för att uppnå målen för detta direktiv när det gäller att förebygga risker och faror både för hälsan och för miljön och beroendet av bekämpningsmedel; arbete för att främja och uppmuntra ibruktagandet av icke-kemiska växtskyddsmetoder .
Motivering
Risker för människors hälsa måste förebyggas helt och hållet och inte bara minskas.
Det här står i överensstämmelse med tidigare ändringsförslag.
Ändringsförslag
94
ca) Utvärdering och anpassning av de nationella handlingsplanerna.
Ändringsförslag
95
3.
3.
Medlemsstaterna skall meddela kommissionen och övriga medlemsstater resultaten av de utvärderingar som gjorts enligt punkt 2 och göra dem tillgängliga för allmänheten .
Motivering
Ändringsförslag
96
4.
4.
Motivering
Användningsindikatorer och mål i fråga om användningen bör fastställas vid sidan om riskindikatorer och mål i fråga om riskerna.
Ändringsförslag
97
Motivering
Ändringsförslag
98
5.
5.
Motivering
Ändringsförslag
99
5a.
När uppgifter samlas in ska man se till att gemenskapens lant brukare och vinodlare inte belastas med ytterligare dokumentationsskyldigheter eller orimliga anmälnings- eller rapporteringsskyldigheter.
Motivering
Lantbrukarna och vinodlarna omfattas redan av en bred dokumentations- och rapporteringsskyldighet.
Om det i framtiden utarbetas en förordning med statistik för växtskyddsmedel bör man se till att det inte uppstår ytterligare, orimliga anmälnings-, rapporterings- eller dokumentationsskyldigheter för lantbrukarna och vinodlarna.
Ändringsförslag
100
Rapportering
Bokföring och rapportering
-1.
De som bedriver handel med bekämpningsmedel ska bok föra alla bekämpningsmedel och all utrustning för spridning av bekämpningsmedel som de mottagit, sålt, levererat eller på annat sätt avhänt sig under en tid av två år.
Motivering
Dessa krav på bokföring gäller redan för personer som bedriver verksamhet med bekämpningsmedel och följer EUREPGAP-standarden eller de standarder för integrerat växtskydd som lantbrukarföreningar och lantbruksandelslag runtom i Europa ställer sig bakom.
Ändringsförslag
101
Artikel 15
Kommissionen skall regelbundet lämna en rapport till Europaparlamentet och rådet om framstegen i genomförandet av detta direktiv, vid behov tillsammans med förslag till ändringar.
Kommissionen skall vart tredje år lämna en rapport till Europaparlamentet och rådet om framstegen i genomförandet av detta direktiv och en utvärdering av de nationella handlingsplanerna , vid behov tillsammans med förslag till ändringar.
Medlemsstaterna ska årligen rapportera till kommissionen om sina nationella handlingsplaner .
Motivering
Regelbundna rapporter om hur genomförandet fortskridit är en förutsättning för ett framgångsrikt arbete.
På det här sättet kommer medlemsstaterna att kunna utbyta information sinsemellan, och kommissionen kommer att kunna utvärdera de nationella handlingsplanerna och, vid behov, tillämpningen av ändringarna.
Ändringsförslag
102
Artikel 15a (ny)
Artikel 15a
Utbyte av information och bästa praxis
Kommissionen ska inrätta en plattform för utbyte av information och bästa praxis om hållbar användning av bekämpningsmedel och om integrerat växtskydd.
Motivering
Utbyte av information och bästa praxis mellan medlemsstaterna och andra berörda parter ingår som ett viktigt led i främjandet av hållbar användning av bekämpningsmedel och integrerat växtskydd.
Detta innebär att upptäckter och iakttagelser som redan gjorts inte måste göras på nytt.
Befintliga initiativ (såsom European Initiative for Sustainable Development in Agriculture) skulle kunna inkluderas.
Ändringsförslag
103
2.
När det hänvisas till denna punkt skall artiklarna 3 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
2.
3.
Motivering
Detta ändringsförslag är nödvändigt för att anpassa texten till bestämmelserna i det nya beslutet om kommittéförfarandet.
Ändringsförslag
104
a) utarbetande av ett harmoniserat system inbegripet en lämplig databas för att samla in och lagra all information om riskindikatorer för bekämpningsmedel och för att göra denna information tillgänglig för behöriga myndigheter, andra berörda parter och allmänheten,
a) utarbetande av ett harmoniserat system inbegripet en lämplig databas för att samla in och lagra all information om risk- och användningsindikatorer för bekämpningsmedel och för att göra denna information tillgänglig för behöriga myndigheter, andra berörda parter och allmänheten,
Ändringsförslag
105
Motivering
Ändringsförslag
106
Bilaga I, rubriken och inledningen
Utbildningsprogram
Utbildningsprogram skall utformas på ett sådant sätt att de ger tillräcklig kunskap om följande:
Utbildnings- och fortbildningsprogram skall utformas på ett sådant sätt att de ger tillräcklig kunskap om följande:
Motivering
Genom detta ändringsförslag anpassas bilaga I till bestämmelserna i artikel 5 (jfr ändringsförslaget till artikel 5).
Ändringsförslag
107
All tillämplig lagstiftning om bekämpningsmedel och deras användning , märkning av bekämpningsmedel och märkningssystem, bekämpningsmedelsterminologi, samt säkerhet, toxicitet och ekotoxicitet i samband med bekämpningsmedel .
Motivering
Förbättringar i utbildningsprogrammen.
Ändringsförslag
108
Bilaga I, led 2, led a
a) risker för människor (operatörer, boende, andra närvarande personer, personer som ger sig in i behandlade områden och personer som hanterar eller äter behandlade produkter) och hur dessa förvärras av faktorer som rökning,
a) risker för människor (operatörer, boende, andra närvarande personer, personer som ger sig in i behandlade områden och personer som hanterar eller äter behandlade produkter) och alla potentiella akuta och kroniska skadeverkningar på hälsan till följd av långvarig exponering och hur dessa förvärras av faktorer som rökning , födointag eller underlåtenhet att använda lämplig skyddsutrustning ,
Motivering
De som använder bekämpningsmedel måste vara fullt medvetna om de risker och de potentiella akuta och kroniska skadeverkningar på hälsan till följd av långvarig exponering som användningen är förenad med.
Ändringsförslag
109
Bilaga I, led 2, led b
b) symptom på bekämpningsmedelsförgiftning och första hjälpen-åtgärder,
b) symptom på bekämpningsmedelsförgiftning och första hjälpen-åtgärder samt symptom på kronisk påverkan av hälsan ,
Motivering
Ändringsförslag
110
Bilaga I, led 2, led c
c) risker för icke-målväxter, nyttiga insekter, vilda djur och växter, biologisk mångfald och miljön i stort.
c) risker för icke-målväxter, nyttiga insekter, vilda djur och växter, biologisk mångfald och miljön i stort , med särskild hänsyn tagen till skadeverkningarna vid användning av bekämpningsmedel inom jordbruket, såsom förlust av naturliga fiender och minskad insektspollination .
Motivering
Användningen av bekämpningsmedel medför ett flertal externa kostnader för jordbruket, och därför bör de kunskaper man på senare tid fått om dessa skadeverkningar tas med i utbildningsprogrammen.
Ändringsförslag
111
Motivering
Ibland används bekämpningsmedel rent ”kosmetiskt”, det vill säga utan anknytning till någon bestämd skadegörare eller några bestämda sjukdomar, och då handlar det inte längre om växtskydd.
Med hänsyn tagen till de erkända riskerna och de akuta och kroniska skadeverkningarna på människors hälsa, vilka mera ingående beskrivits i konsekvensanalysen av den temainriktade strategin, bör medlemsstaterna vinnlägga sig om att främja och uppmuntra en brett upplagd övergång till icke-kemiska växtskydds- och odlingsmetoder.
Ändringsförslag
112
Introduktion till jämförande bedömning på användarnivå för att hjälpa yrkesmässiga användare att göra de lämpligaste valen mellan alla godkända medel för ett visst skadegörarproblem i en given situation.
Motivering
Ändringsförslag
113
Åtgärder för att minimera riskerna för människor, icke-målarter och miljön: säkra arbetsmetoder för lagring, hantering och blandning av bekämpningsmedel samt för bortskaffande av tomma förpackningar, annat förorenat material och bekämpningsmedelsrester (även bulkblandningar) i koncentrerad eller utspädd form; rekommenderat sätt att begränsa operatörens exponering (personlig skyddsutrustning).
Motivering
Var och en som använder bekämpningsmedel måste vara fullt medveten om alla potentiella exponeringsfaktorer med därtill hörande risker, detta med tanke på både sin egen hälsa och hälsan hos andra personer som kan komma att exponeras, framför allt personer som bor i närheten av besprutade fält.
Ändringsförslag
114
Metoder för att förbereda spridningsutrustning för arbete, inbegripet kalibrering, och för handhavande med minsta möjliga risker för användaren, andra personer, icke-målarter bland djur och växter, den biologiska mångfalden och miljön.
Motivering
Det måste tydligare framhållas att också vattentillgångarna behöver skydd.
Man måste också se till att det vidtas åtgärder i händelse av extrema väderleksförhållanden och om bekämpningsmedel kan läcka ut i vattenförekomster.
Vädret har en mycket kraftig inverkan på föroreningsnivån.
Om marken är våt är risken mycket större för att bekämpningsmedel kommer att rinna av med vattnet.
Häftigt regn kan kännbart öka risken för avrinning både från gårdstunen och från åkrarna.
Ändringsförslag
115
Användning och underhåll av spridningsutrustning och särskilda spruttekniker (t.ex. lågvolymssprutning, avdriftsreducerande munstycken) mål för den tekniska kontrollen av sprutor i bruk och metoder för att förbättra duschkvaliteten.
Ändringsförslag
116
Nödåtgärder för att skydda människors hälsa , miljön och vattentillgångarna vid oavsiktligt spill , förorening och extrema väderleksförhållanden med åtföljande risk för att bekämpningsmedel läcker ut .
Motivering
Det måste tydligare framhållas att också vattentillgångarna behöver skydd.
Man måste också se till att det vidtas åtgärder i händelse av extrema väderleksförhållanden och om bekämpningsmedel kan läcka ut i vattnet.
Vädret har en mycket kraftig inverkan på föroreningsnivån.
Om marken är våt är risken mycket större för att bekämpningsmedel kommer att rinna av med vattnet.
Häftigt regn kan kännbart öka risken för avrinning både från gårdstunen och från åkrarna.
Ändringsförslag
117
Bilaga I, led 10a (nytt)
Motivering
I ramdirektivet om vatten ingår krav på att ytvattnet, grundvattnet och bevarandet av livsmiljöer och arter som är direkt beroende av vatten samt förekomster av dricksvatten ska ägnas särskild omsorg.
Detta måste fastställas för utbildningsprogrammen så att de som yrkesmässigt använder bekämpningsmedel liksom också distributörer och rådgivare blir medvetna om dessa behov.
Ändringsförslag
118
Bilaga I, led 10b (nytt)
a) Bekämpning av skadegörare inom jordbruket.
b) Bekämpning av skadegörare inom skogsbruket.
c) Utsädesbehandling.
d) Bekämpning av skadegörare i vattenmiljö.
e) Bekämpning av skadegörare i anslutning till allmän väg .
f) Bekämpning av skadegörare av folkhälsoskäl.
g) Bekämpning av gnagare.
Ändringsförslag
119
Bilaga I, led 10c (nytt)
Motivering
I programmen bör det som ett led i bästa praxis även ingå en utveckling av kunskapen om riskbedömning, under hänsynstagande till de lokala förhållandena.
Ändringsförslag
120
Bilaga IIa (ny)
Bilaga IIa
Minimiinslag i nationella bakgrundsrapporter
Del A: Föreskrivna inslag i inledande nationella utredningar av minskad användning av bekämpningsmedel.
Beskrivning av aktuella förhållanden:
• Uppgifter om produktion, import, export, försäljning och distribution av bekämpningsmedel.
• Aktuella trender inom förbrukningen av bekämpningsmedel (totala mängden ingredienser som använts, respektive mängder bekämpningsmedel som använts vid olika tillämpningar på alla större grödor och utanför jordbruket, framför allt på allmänna platser, beräkning av index över behandlingsfrekvens).
• Beskrivning av hur de aktuella trenderna inom användningen av bekämpningsmedel påverkar miljön, livsmedelskedjan och människors hälsa, utgående från data som insamlats via befintliga program för övervakning.
• Översikt av aktuell lagstiftning och politiska styrmedel samt deras effektivitet.
• Utvärdering av behovet av bekämpningsmedel.
• Luckor som konstaterats i ovannämnda uppgifter.
Scenarier för minskad användning av bekämpningsmedel:
• En minskning av användningen på 30 procent och 50 procent, mätt enligt index över behandlingsfrekvens.
Konsekvensbedömning av de olika scenarierna:
• Konsekvenser för miljön (också i fråga om energi förbrukning och växthusgaser).
• Konsekvenser för folkhälsan (arbetare, boende, närvarande personer, resthalter i livsmedel).
• Konsekvenser för jordbruksproduktionen.
• Kostnader och nytta i ekonomiskt hänseende (också i fråga om minskade dolda kostnader) för de olika scenarierna.
Identifiering och bedömning av vad som behövs för att genomföra scenarierna :
• Konsekvenserna av de inslag som angivits i direktivet när det gäller att uppnå minskad användning av bekämpningsmedel.
• Vilka ytterligare vetenskapliga data som behövs och hur de ska samlas in, till exempel genom ytterligare övervakningskapacitet och forskningsanläggningar.
• Vilken ytterligare kapacitet som behövs för att minska användningen av bekämpningsmedel, till exempel arbete till förmån för ett mera extensivt jordbruk och inspektörer som har till uppgift att övervaka användningen.
• Möjliga sätt att finansiera genomförandet av de olika scenarierna, bland annat avgifter.
Slutsatser:
• Uppnåbara mål för minskad användning av bekämpningsmedel, både för enskilda grödor och för ändamål utanför jordbruket samt på landsomfattande nivå, varvid målen ska motsvara åtminstone de obligatoriska mål för minskning som fastställts i artikel 6 och syfta till att användningen ska minska ytterligare med tiden.
Del B: Föreskrivna inslag i kommande nationella utredningar gällande minskad användning av bekämpningsmedel.
• Utvärdering av erfarenheterna från de första tre åren gällande genomförandet av programmet för minskad användning av bekämpningsmedel.
• I övrigt: som ovan.
Fastställande av nya mål för nästa period.
Motivering
Denna nya bilaga behövs som ett vägledande dokument för medlemsstaterna när de ska utarbeta de nationella bakgrundsrapporterna, och för att medlemsstaternas rapporter och kommissionens utvärdering av situationen inom EU ska kunna göras enhetliga.
Ändringsförslag
121
Bilaga IIb (ny)
Bilaga IIb
Minimiinslag i de nationella handlingsplanerna för minskning av riskerna med och användningen av bekämpningsmedel
Kvalitativa och kvantitativa mål:
• Interi ms mål för minskning av riskerna och användningen, mätt med index över behandlingsfrekvensen.
• Mål för särskilda målgrupper , såsom offentliga myndigheter och lantbrukare, eller särskilda användningar, exempelvis i anslutning till allmän väg .
• Mål för minskad användning i områden som är känsliga för bekämpningsmedel.
• Mål för gradvis bortskaffande av bekämpningsmedel och resthalter av dem ur grundvatten och andra miljömedier.
• Mål för problemgrödor och/eller problemregioner.
Övervakning av användningen:
• Åtgärder för ett garanterat genomförande av praxis för integrerat växtskydd.
• Förbud mot spridning av bekämpningsmedel nära dricksvattentäkter eller i områden som är känsliga för bekämpningsmedel, såsom naturområden och buffertzoner.
• Förbud mot spridning av bekämpningsmedel i områden med stora exponeringsrisker, såsom skolor, parker och andra allmänna platser, vägkanter etc.
Forskning och informationsspridning:
• Forskning kring icke-kemiska alternativ till bekämpningsmedel.
• Demonstrationsprogram om hur användningen av bekämpningsmedel kan minskas med hjälp av icke-kemiska växtskyddsmetoder och växtskyddssystem.
• Utbildning av jordbrukskonsulenter i frågor som rör icke-kemiska växtskyddsmetoder och växtskyddssystem.
• Forskning kring frågan hur användningen av bekämpningsmedel kan minskas med hjälp av bättre utrustning, metoder och system för besprutning.
Information, utbildning och yrkesutbildning:
• Utbildning för alla som hanterar bekämpningsmedel om vilka risker dessa medför för hälsan samt om icke-kemiska växtskyddsmetoder och växtskyddssystem.
• Vägledning för dem som hanterar bekämpningsmedel, exempelvis om lagringen och hanteringen av dessa medel.
Utrustning för spridning av bekämpningsmedel:
• Inspektioner av utrustning som används.
Ekonomiska styrmedel:
• Ekonomiskt stöd till genomförandet av standarder och praxis i samband med integrerat växtskydd.
• Ekonomiskt stöd till andra sätt att minska användningen av bekämpningsmedel.
• Ökad användning av mekanismer för tvärvillkor.
Motivering
Denna nya bilaga behövs för att medlemsstaterna ska få vägledning vid genomförandet av sina nationella handlingsplaner och när det gäller att uppnå enhetlighet bland medlemsstaterna.
Ändringsförslag
122
Bilaga IIc (ny)
Bilaga IIc
Inslag i allmänna och grödspecifika kriterier för integrerat växtskydd
I det integrerade växtskyddet ska åtminstone följande allmänna kriterier ingå:
(a) Bland de olika till buds stående alternativen för att hindra och/eller utrota skadegörare ska framför allt följande användas eller stödjas:
• Optimalt växelbruk så att balans mellan markorganismerna uppnås och jorden bevaras i sunt skick, så att skadegörare i marken inte kommer åt att sprida sig och rökbehandling eller annan kemikaliebehandling av marken inte behövs.
• Åstadkommande av hälsosam jordmån för grödorna, exempelvis genom att öka den procentuella halten organiskt material i jorden, begränsa plöjningsdjupet, förebygga erosion och ha bästa möjliga växtföljd.
• Lämplig odlingsteknik, såsom falsk såbädd, tidpunkter för sådden, såddtäthet, undersådd, sådd i förband med optimalt avstånd, plöjning med reducerad bearbetning, hygienåtgärder, gallring.
• Odlingsväxter som är så resistenta och tåliga som möjligt samt godkänt/certifierat utsäde och plantmaterial.
• Väl avvägda gödselgivor utgående från uppgifter om vilka näringsämnen som redan finns i marken samt om jordarterna; kalkning och bevattning/dränering för att minska mottagligheten för skadegörare och sjukdomar.
Användning av grundvatten för bevattningsändamål ska undvikas.
• Åtgärder för att inte skadliga organismer ska spridas via maskiner och utrustning.
• Åtgärder för att skydda viktiga nyttoorganismer och öka deras antal, såsom användning av ekologiska infrastrukturer på och utanför produktionsställena, samt minimikrav på arealuttag och plantering av sådana växter som drar till sig naturliga fiender till skadegörare.
(b) Skadliga organismer ska övervakas med hjälp av lämpliga metoder och verktyg.
Dessa ska omfatta vetenskapligt underbyggda system för varning, prognos och tidig diagnos, i de fall sådana finns att tillgå, samt rådgivare med fackmannainsikter, av det slag som tillhandahålls från statligt och privat håll.
(c) Yrkesmässiga användare ska utgående från resultaten av övervakningen fatta beslut om huruvida och i så fall när växtskyddsåtgärder ska vidtas.
Fasta och vetenskapligt välunderbyggda tröskelvärden är väsentliga med tanke på beslutsfattandet.
Innan någon behandling inleds ska hänsyn tas till vilka tröskelvärden för skadegörare som eventuellt definierats för regionen i fråga.
(d) Biologiska, fysiska, mekaniska och andra icke-kemiska metoder ska alltid när det är möjligt ges företräde framför kemiska metoder.
Ogräsbekämpning ska ske genom mekanisk rensning eller med hjälp av andra icke-kemiska metoder, såsom värmebehandling.
Undantag får tillåtas endast om ogynnsam väderlek under en längre tid förhindrat mekanisk rensning.
(e) Växtskyddsmedel som används ska vara så målspecifika som möjligt och ha minsta möjliga biverkningar för människors hälsa och miljön; bland växtskyddsmedel av detta slag märks extrakt från växter och träd samt mineralämnen för att motverka svamp.
(f) Yrkesmässiga användare ska begränsa användningen av växtskyddsmedel och andra ingrepp till vad som är nödvändigt, exempelvis genom minskade doser, minskad spridningsfrekvens eller partiell spridning och därvid ta hänsyn till att riskerna för växtligheten ska förbli acceptabla och att insatserna av växtskyddsmedel inte får öka risken för att populationerna av skadliga organismer ska utveckla resistens.
(g) I de fall då risken för resistens mot ett växtskyddsmedel är känd och när förekomsten av skadliga organismer kräver att växtskyddsmedel vid upprepade tillfällen används på någon gröda ska tillgängliga strategier mot resistens användas, så att växtskyddsmedlen inte förlorar sin verkan.
I detta sammanhang får flera olika växtskyddsmedel med olika verkningssätt användas parallellt.
(h) Yrkesmässiga användare ska, utgående från varje enskild åker, bok föra de växtskyddsmedel som använt s .
De ska, utgående från denna bokföring och från övervakningen av de skadliga organismerna, undersöka nyttan med de växtskyddsåtgärder som använts.
Motivering
Definition av integrerat växtskydd.
MOTIVERING
Bakgrund
Genom beslutet om antagandet av sjätte miljöhandlingsprogrammet bekräftade Europaparlamentet och rådet att hälso- och miljöeffekterna av växtskyddsmedel måste minskas ytterligare.
De framhöll vikten av att uppnå en mer hållbar användning av bekämpningsmedel och föreslog en tvådelad strategi:
- Fullständigt genomförande och lämplig översyn av gällande lagstiftning.
- Utarbetande av en temainriktad strategi för hållbar användning av bekämpningsmedel.
I meddelandet ”Temainriktad strategi för hållbar användning av bekämpningsmedel” ( KOM(2006)0372 ) redogör kommissionen för de olika åtgärder som skulle kunna ingå i strategin.
Föreliggande förslag till direktiv ska bidra till genomförandet av den temainriktade strategin och inrättandet av en ram för åtgärder för hållbar användning av växtskyddsmedel.
Tillämp ningsområde
Föredraganden anser att titeln på det förslag till direktiv som har lagts fram kan missförstås.
Som kommissionen själv medger gäller förslaget till direktiv bestämmelser om en särskild grupp bekämpningsmedel, nämligen växtskyddsmedel.
Av det skälet bör begreppet ”bekämpningsmedel” i hela texten till direktivet ersättas med ”växtskyddsmedel”.
Detta bör uttryckligen klargöras i hela texten till direktivet.
Det är inte uteslutet att tillämpningsområdet kan komma att utvidgas vid ett senare tillfälle, men detta bör i så fall ske i samråd med Europaparlamentet.
Målsättning
Föredraganden anser att direktivet i enlighet med föreskrifterna i det sjätte miljöhandlingsprogrammet och den temainriktade strategin för hållbar användning av bekämpningsmedel främst måste handla om att minska de risker för och effekter på miljön och människors hälsa som användning av växtskyddsmedel medför.
De åtgärder som vidtas måste dock vara rimliga.
Detta innebär att de fördelar som användningen av växtskyddsmedel ger emellertid också måste beaktas med hänsyn till produktionens kvalitet och vinstmaximering.
Nationella handlingsplaner
Föredraganden delar kommissionens uppfattning att det främst bör vara en fråga för medlemsstaterna att inom ramen för de nationella handlingsplanerna bidra till att minska riskerna med användning av växtskyddsmedel.
Endast på detta sätt kan lämplig hänsyn tas till olika lokala förhållanden och faktorer.
Expertis och information
Föredraganden anser att yrkesmässiga användare, distributörer och rådgivare genom utbildnings- och fortbildningsåtgärder bör förbättra sina kunskaper om hur växtskyddsmedel hanteras på rätt sätt.
Allmänheten bör genom motsvarande program på lämpligt sätt informeras om hur växtskyddsmedel hanteras korrekt.
Tekniska bestämmelser
Utrustning och tillbehör för spridning av bekämpningsmedel bör inspekteras med jämna mellanrum.
Föredraganden anser att medlemsstaterna på vissa, klart definierade villkor ska få fastställa bestämmelser för flygbesprutning.
Vattenmiljön
I ramdirektivet om vatten föreskrivs grundläggande bestämmelser och åtgärder för att skydda vattenmiljön.
Vid genomförandet av ramdirektivet om vatten krävs dock att användning av växtskyddsmedel uppmärksammas särskilt.
I de nationella handlingsplanerna måste därför klart och tydligt fastställas vad som ska beaktas vid användning av växtskyddsmedel, också när det gäller spridning, buffertzoner och lagring i vattendrag och vattenskyddsområden.
God yrkesmässig praxis för växtskydd och integrerat växtskydd
De kriterier som fastställs i bilagorna III och IV beskriver inom vilka ramar god yrkesmässig praxis för växtskydd och integrerat växtskydd kan röra sig i Europeiska unionen.
I god yrkesmässig praxis för växtskydd ska det fastställas vilka grundkrav som ska uppfyllas av den som genomför åtgärder för växtskydd.
Med beaktande av de regionala förhållandena (t.ex. jordbruk, väderförhållanden och ekologi) ska medlemsstaterna eller yrkesförbund formulera odlings- eller sektorspecifika riktlinjer för integrerat växtskydd på grundval av de allmänna kriterierna i bilaga IV för integrerat växtskydd.
Det integrerade växtskyddet är förebilden för växtskyddet i Europeiska unionen och därmed även innovationsmotorn för växtskyddet.
Det integrerade växtskyddet kan också omfatta åtgärder med större ekonomiska risker för att minska användning av växtskyddsmedel och minska de risker som användningen medför.
Tillämpningen av dessa riktlinjer är frivillig och kan främjas genom särskilda stimulansåtgärder.
Inom vissa tidsintervall ska man kontrollera huruvida de allmänna kriterierna för god yrkesmässig praxis för växtskydd och de allmänna kriterierna för integrerat växtskydd ska anpassas i förhållande till läget inom vetenskapen och tekniken samt de allmänna framstegen.
Motsvarande anpassningar ska göras inom ramen för kommittéförfarandet.
Medlemsstaternas rapporter kommer att vara viktiga utgångspunkter för en diskussion om bilagorna.
Genom den tvådelade strategin säkerställs att det alltid går att göra mer för miljön och i förekommande fall få kompensation för sådana insatser.
Å andra sidan kommer god yrkesmässig praxis att främja arbete som sker i enlighet med principerna för integrerat växtskydd.
Yttrande från utskottet för rättsliga frågor om den föreslagna rättsliga grunden
Miroslav Ouzký
Ordförande
Utskottet för miljö, folkhälsa och livsmedelssäkerhet
BRYSSEL
Ärende: Yttrande över den rättsliga grunden för Europaparlamentets och rådets direktiv om upprättande av en ram för gemenskapens åtgärder för att uppnå en hållbar användning av bekämpningsmedel ( KOM(2006)0373 – C6‑0246/2006 – 2006/0132(COD) )
Vid utskottssammanträdet den 12 september 2007 behandlade utskottet detta ärende.
Bakgrund
Artikel 152
1.
En hög hälsoskyddsnivå för människor skall säkerställas vid utformning och genomförande av all gemenskapspolitik och alla gemenskapsåtgärder.
Gemenskapens insatser, som skall komplettera den nationella politiken, skall inriktas på att förbättra folkhälsan, förebygga ohälsa och sjukdomar hos människor och undanröja faror för människors hälsa.
Sådana insatser skall innefatta kamp mot de stora folksjukdomarna genom att främja forskning om deras orsaker, hur de överförs och hur de kan förebyggas samt hälsoupplysning och hälsoundervisning.
Gemenskapen skall komplettera medlemsstaternas insatser för att minska narkotikarelaterade hälsoskador, inklusive upplysning och förebyggande verksamhet.
2.
Gemenskapen skall främja samarbete mellan medlemsstaterna på de områden som avses i denna artikel och vid behov stödja deras insatser.
Medlemsstaterna skall i samverkan med kommissionen inbördes samordna sin politik och sina program på de områden som avses i punkt 1.
Kommissionen kan i nära kontakt med medlemsstaterna ta lämpliga initiativ för att främja en sådan samordning.
3.
Gemenskapen och medlemsstaterna skall främja samarbetet med tredje land och behöriga internationella organisationer på folkhälsans område.
4.
Rådet skall, enligt förfarandet i artikel 251 och efter att ha hört Ekonomiska och sociala kommittén samt Regionkommittén, bidra till att de mål som anges i denna artikel uppnås genom att
a) besluta om åtgärder för att fastställa höga kvalitets- och säkerhetsstandarder i fråga om organ och ämnen av mänskligt ursprung, blod och blodderivat; dessa åtgärder skall inte hindra någon medlemsstat från att upprätthålla eller införa strängare skyddsåtgärder,
b) med undantag från artikel 37 besluta om sådana åtgärder på veterinär- och växtskyddsområdet som direkt syftar till att skydda folkhälsan,
c) besluta om stimulansåtgärder som är utformade för att skydda och förbättra människors hälsa, dock utan att dessa åtgärder får omfatta någon harmonisering av medlemsstaternas lagar eller andra författningar.
Rådet kan också med kvalificerad majoritet på förslag av kommissionen anta rekommendationer för de syften som anges i denna artikel.
5.
När gemenskapen handlar på folkhälsoområdet skall den fullt ut respektera medlemsstaternas ansvar för att organisera och ge hälso- och sjukvård.
Artikel 175
1.
Rådet skall enligt förfarandet i artikel 251 och efter att ha hört Ekonomiska och sociala kommittén och Regionkommittén besluta om vilka åtgärder som skall vidtas av gemenskapen för att uppnå de mål som anges i artikel 174.
Artikel 174
1.
Gemenskapens miljöpolitik skall bidra till att följande mål uppnås:
– Att bevara, skydda och förbättra miljön.
– Att skydda människors hälsa.
– Att utnyttja naturresurserna varsamt och rationellt.
– Att främja åtgärder på internationell nivå för att lösa regionala eller globala miljöproblem.
2.
Gemenskapens miljöpolitik skall syfta till en hög skyddsnivå med beaktande av de olikartade förhållandena inom gemenskapens olika regioner.
Den skall bygga på försiktighetsprincipen och på principerna att förebyggande åtgärder bör vidtas, att miljöförstöring företrädesvis bör hejdas vid källan och att förorenaren skall betala.
I detta sammanhang skall de harmoniseringsåtgärder som motsvarar miljöskyddskraven i förekommande fall innehålla en skyddsklausul som tillåter medlemsstaterna att av icke ‑ekonomiska miljömässiga skäl vidta provisoriska åtgärder, som skall vara föremål för ett kontrollförfarande på gemenskapsnivå.
3.
När gemenskapen utarbetar sin miljöpolitik skall den beakta
– tillgängliga vetenskapliga och tekniska data,
– miljöförhållanden i gemenskapens olika regioner,
– de potentiella fördelar och kostnader som är förenade med att åtgärder vidtas eller inte vidtas,
– den ekonomiska och sociala utvecklingen i gemenskapen som helhet och den balanserade utvecklingen i dess regioner.
4.
Inom sina respektive kompetensområden skall gemenskapen och medlemsstaterna samarbeta med tredje land och med behöriga internationella organisationer.
De närmare villkoren för samarbete från gemenskapens sida kan bli föremål för avtal mellan gemenskapen och berörda tredje parter; avtalen skall förhandlas fram och ingås enligt artikel 300.
Föregående stycke skall inte inverka på medlemsstaternas behörighet att förhandla i internationella organ och att ingå internationella avtal.
Bedömning
I den rättsliga grunden fastställs gemenskapens materiella behörighet.
Enligt motiveringen innehåller förslaget till direktiv följande åtgärder:
· Nationella handlingsplaner som fastställer mål för att minska faror, risker och beroendet av kemisk bekämpning för växtskydd, och som ger utrymme för den flexibilitet som krävs för att anpassa åtgärderna till specifika situationer i medlemsstaterna.
· Berörda parters deltagande i upprättande, genomförande och anpassning av nationella handlingsplaner.
· Ett system för utbildning av och information till distributörer och yrkesmässiga användare av bekämpningsmedel för att säkerställa att de är fullt medvetna om riskerna med användningen.
Bättre information till allmänheten genom upplysningskampanjer och information som lämnas via detaljhandlare och andra lämpliga åtgärder.
· Regelbunden inspektion av spridningsutrustning för att minska negativa effekter av bekämpningsmedel på människors hälsa (särskilt exponering av operatörer) och miljön under spridning.
· Förbud mot flygbesprutning utom i undantagsfall för att begränsa riskerna för betydande negativa hälso- och miljöeffekter, särskilt genom vindavdrift.
· Särskilda åtgärder för att skydda vattenmiljön mot förorening med bekämpningsmedel.
· Fastställande av områden med kraftigt minskad eller ingen användning av bekämpningsmedel i överensstämmelse med åtgärder som vidtagits enligt annan lagstiftning (såsom ramdirektivet om vatten, fågeldirektivet och livsmiljödirektivet) eller för att skydda särskilt känsliga grupper.
· Hantering och lagring av förpackningar och rester av bekämpningsmedel.
· Standarder för integrerat växtskydd på gemenskapsnivå och fastställande av förutsättningar för lantbrukare att tillämpa integrerat växtskydd.
· Lämpliga harmoniserade indikatorer för att mäta framsteg i fråga om riskreduktion.
· Ett system för informationsutbyte för att löpande utarbeta och uppdatera lämplig vägledning, bästa praxis och rekommendationer.
Artikel 152 bör därför betraktas som en lämplig rättslig grund för åtgärder som rör folkhälsa.
Vid utskottssammanträdet den 12 september 2007 antog utskottet för rättsliga frågor enhälligt
Följande ledamöter var närvarande vid slutomröstningen: Giuseppe Gargani (ordförande), Cristian Dumitrescu, Rainer Wieland och Lidia Joanna Geringer de Oedenberg (vice ordförande), Marek Aleksander Czarnecki, Albert Deß, Bert Doorn, Janelly Fourtou, Monica Frassoni, Jean-Paul Gauzès, Othmar Karas, Piia‑Noora K auppi, Barbara Kudrycka, Klaus-Heiner Lehne, Katalin Lévai, Hans-Peter Mayer, Manuel Medina Ortega, Hartmut Nassauer, Michel Rocard, Aloyzas Sakalas, María Sornosa Martínez, Francesco Enrico Speroni, Daniel Strož och Jacques Toubon. följande rekommendation: Den lämpliga rättsliga grunden för Europaparlamentets och rådets direktiv om upprättande av en ram för gemenskapens åtgärder för att uppnå en hållbar användning av bekämpningsmedel bör vara artiklarna 152.4 och 175.1 i EG-fördraget.
Giuseppe Gargani
YTTRANDE från utskottet för industrifrågor, forskning och energi
till utskottet för miljö, folkhälsa och livsmedelssäkerhet
över förslaget till Europaparlamentets och rådets direktiv om upprättande av en ram för gemenskapens åtgärder för att uppnå en hållbar användning av bekämpningsmedel
( KOM(2006)0373 – C6‑0246/2006 – 2006/0132(COD) )
Föredragande:
Dorette Corbey
KORTFATTAD MOTIVERING
För jordbrukare och konsumenter har användningen av bekämpningsmedel eller växtskyddsmedel stora fördelar eftersom det innebär försörjningstrygghet och ett brett urval till ett rimligt pris.
Växtskyddsmedel kan också ha en viktig funktion i vidareutvecklingen och anpassningen av biobränslen, om grödor används i produktionen av biobränslen.
Å andra sidan utvecklas bekämpningsmedel för att bekämpa vissa organismer och de kan därför ha oönskade effekter på folkhälsan och miljön.
För att åstadkomma en ansvarsfull och hållbar användning av bekämpningsmedel infördes redan 1979 en europeisk politik på detta område.
Man måste därför utgå från båda förslagen.
Föredraganden är positiv till kommissionens förslag i följande avseenden:
· Medlemsstaterna skall upprätta nationella handlingsplaner för att identifiera grödor, aktiviteter och områden för vilka riskerna är oroande samt åtgärder för att komma till rätta med dessa problem.
· System skall upprättas för utbildning av distributörer och yrkesmässiga användare av bekämpningsmedel.
· Vid försäljning av bekämpningsmedel skall mer och bättre information ges till allmänheten.
· Regelbunden teknisk inspektion och underhåll av utrustning för spridning skall införas med hjälp av harmoniserade standarder.
· Särskilda åtgärder för att skydda vattenmiljön skall vidtas, t.ex. buffertzoner eller andra lämpliga åtgärder för att begränsa avdrift.
· Förbud mot flygbesprutning måste absolut införas för att begränsa riskerna för vindavdrift och medlemsstaterna måste få möjlighet att göra undantag (dessa skall vara klart angivna).
Med tanke på skillnaderna i medlemsstaternas geografiska läge, deras jordbruk och klimat är föredraganden också positiv till det stora mått av flexibilitet som medlemsstaterna får när det gäller själva genomförandet.
Däremot anser föredraganden att användningen av icke-kemiska bekämpningsmedel skulle kunna främjas mer genom att bästa praxis sprids och genom regelbunden anpassning av integrerade bekämpningsmedel.
ÄNDRINGSFÖRSLAG
Utskottet för industrifrågor, forskning och energi uppmanar utskottet för miljö, folkhälsa och livsmedelssäkerhet att som ansvarigt utskott infoga följande ändringsförslag i sitt betänkande:
Kommissionens förslag
Ännu ej offentliggjort i EUT.
Parlamentets ändringar
Ändringsförslag
1
2.
2.
2
2a.
Medlemsstaterna får bevilja bidrag eller vidta skatteåtgärder för att främja användningen av mindre skadliga växtskyddsmedel.
Motivering
Det måste vara upp till medlemsstaterna att främja en mer hållbar användning av bekämpningsmedel genom skatteåtgärder om de så önskar.
Ändringsförslag
3
(ia) bekämpningsmedel: växtskyddsmedel enligt förordning (EG) nr […] om utsläppande av växtskyddsmedel på marknaden.
Motivering
I texten refererar man ömsom till termen ”bekämpningsmedel”, ömsom till ”växtskyddsmedel”.
För att undvika oklarheter och garantera rättslig säkerhet är det viktigt att definiera termen ”bekämpningsmedel”.
Ändringsförslag
4
1.
Medlemsstaterna skall anta nationella handlingsplaner för att fastställa mål, åtgärder och tidtabeller för minskning av risker, inbegripet faror , och beroendet av bekämpningsmedel.
Motivering
De nationella handlingsplanerna bör först och främst begränsa de risker och faror som uppstår vid användningen av bekämpningsmedel och egentligen inte användningen i sig.
Det är viktigt att de nationella handlingsplanerna även utgår från målsättningarna i ramdirektivet för vatten.
Ändringsförslag
5
De nationella handlingsplanerna skall bland annat omfatta integrerat växtskydd enligt definitionen i artikel 13 och prioriteral växtskyddsåtgärder med icke ‑kemiska metoder.
Motivering
Integrerat växtskydd måste stimuleras.
Ändringsförslag
6
1.
1.
Motivering
Ändringsförslag
7
Artikel 7
Medlemsstaterna skall stödja informationsprogram riktade till allmänheten och underlätta allmänhetens tillgång till information om bekämpningsmedel, särskilt när det gäller hälso- och miljöeffekter och icke-kemiska alternativ.
Medlemsstaterna skall stödja informationsprogram riktade till användare, yrkesmässiga såväl som icke yrkesmässiga och underlätta deras tillgång till information om bekämpningsmedel, särskilt när det gäller effekterna på jordbruk, hälsa och miljö samt icke-kemiska alternativ.
Motivering
Bekämpningsmedel har också sina fördelar, t.ex. bidrar växtskyddsmedel till att öka jordbrukets avkastning, höja kvaliteten på jordbruksvarorna, begränsa jorderosionen, uppfylla växtskyddskraven och möjliggöra internationell handel med jordbruksprodukter.
Ändringsförslag
8
1.
Medlemsstaterna skall, om bekämpningsmedel används i närheten av vatten, i synnerhet vatten som är avsett för mänskligt bruk, se till att företräde ges åt
Motivering
Vatten som är avsett för mänskligt bruk bör skyddas särskilt, i linje med bestämmelserna i artikel 7 i ramdirektivet för vatten.
Ändringsförslag
9
b) Användning av bekämpningsmedel skall förbjudas eller begränsas i särskilda bevarandeområden och andra områden som utsetts i syfte att fastställa nödvändiga bevarandeåtgärder enligt artiklarna 3 och 4 i direktiv 79/409/EEG och artiklarna 6, 10 och 12 i direktiv 92/43/EEG.
Ett förbud eller en begränsning enligt b får grundas på resultaten av relevanta riskbedömningar.
Ett förbud eller en begränsning skall grundas på resultaten av relevanta riskbedömningar.
Motivering
Det är viktigt att man verkligen kontrollerar känsliga områden (med tanke på vilda djur och växter eller känsliga grupper såsom barn) för att se om användningen av bekämpningsmedel måste minskas eller till och med förbjudas.
Man måste bestämma från fall till fall och utifrån en riskbedömning.
Ändringsförslag
10
1.
Medlemsstaterna skall vidta de åtgärder som behövs för att säkerställa att följande arbetsmoment inte medför risk för människors hälsa eller säkerhet eller för miljön:
1.
Medlemsstaterna skall vidta de åtgärder som behövs för att säkerställa att följande arbetsmoment utförda av yrkesmässiga användare inte medför risk för människors hälsa eller säkerhet eller för miljön:
Motivering
Det måste klargöras att kommissionens föreslagna åtgärd är utan betydelse för privat användning.
Ändringsförslag
11
(d) Rengöring av utrustning som använts för spridning.
(d) Förberedning, hantering, rengöring och lagring av utrustning som använts för spridning och eventuella tillbehör, inbegripet spridningsutrustning och kemikalier .
Ändringsförslag
12
1a.
Motivering
Medlemsstaterna skall främja en mer hållbar och miljövänlig användning av bekämpningsmedel.
Det är dessutom viktigt att det finns en tydligare koppling mellan detta direktiv och förordning (EG) nr […] om utsläppande av växtskyddsmedel på marknaden.
Ändringsförslag
13
2.
2.
Medlemsstaterna skall skapa eller stödja skapandet av alla nödvändiga förutsättningar för tillämpning av integrerat växtskydd och för varje gröda beskriva bästa praxis för integrerat växtskydd och ge företräde åt icke-kemiska växtskydd .
Motivering
Bästa praxis när det gäller icke-kemiska växtskyddsmetoder hjälper yrkesmässiga användare att välja ett miljövänligare växtskyddsalternativ.
Ändringsförslag
14
Artikel 15
Kommissionen skall regelbundet lämna en rapport till Europaparlamentet och rådet om framstegen i genomförandet av detta direktiv, vid behov tillsammans med förslag till ändringar.
Kommissionen skall vart tredje år lämna en rapport till Europaparlamentet och rådet om framstegen i genomförandet av detta direktiv och en utvärdering av de nationella handlingsplanerna , vid behov tillsammans med förslag till ändringar.
Ändringsförslag
15
Artikel 15a (ny)
Artikel 15a
Utbyte av information och bästa praxis
Kommissionen skall skapa en plattform för utbyte av information och bästa praxis när det gäller hållbar användning av bekämpningsmedel och integrerat växtskydd.
Motivering
Utbytet av information och bästa praxis mellan medlemsstaterna och andra berörda parter är en viktig del vid främjandet av hållbar användning av bekämpningsmedel och integrerat växtskydd.
På så sätt behöver man inte ständigt etablera en ny praxis.
Existerande initiativ (såsom det europeiska initiativet för att främja hållbar utveckling inom jordbruket) skulle också kunna ingå där.
Ändringsförslag
16
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs.
Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs.
Motivering
Korrekt användning av bekämpningsmedel skall garanteras genom den föregående förordningen.
ÄRENDETS GÅNG
Titel
Ramdirektiv om hållbar användning av bekämpningsmedel
Referensnummer
KOM(2006)0373 – C6-0246/2006 – 2006/0132(COD)
Ansvarigt utskott
ENVI
Yttrande
Tillkännagivande i kammaren
ITRE
5.9.2006
Förstärkt samarbete - tillkännagivande i kammaren
5.9.2006
Föredragande av yttrande
Utnämning
Dorette Corbey
23.11.2006
Behandling i utskott
28.2.2007
3.5.2007
Antagande
3.5.2007
Slutomröstning: resultat
+:
–:
0:
28
14
1
Slutomröstning: närvarande ledamöter
Šarūnas Birutis, Renato Brunetta, Jerzy Buzek, Jorgo Chatzimarkakis, Silvia Ciornei, Pilar del Castillo Vera, Den Dover, Lena Ek, Nicole Fontaine, Adam Gierek, Norbert Glante, Fiona Hall, David Hammerstein, Erna Hennicot-Schoepges, Mary Honeyball, Romana Jordan Cizelj, Romano Maria La Russa, Pia Elda Locatelli, Eugenijus Maldeikis, Angelika Niebler, Reino Paasilinna, Miloslav Ransdorf, Vladimír Remek, Herbert Reul, Mechtild Rothe, Paul Rübig, Andres Tarand, Patrizia Toia, Catherine Trautmann, Claude Turmes, Nikolaos Vakalis, Alejo Vidal-Quadras
Slutomröstning: närvarande suppleanter
YTTRANDE från utskottet för jordbruk och landsbygdens utveckling (*)
till utskottet för miljö, folkhälsa och livsmedelssäkerhet
över förslaget till Europaparlamentets och rådets direktiv om upprättande av en ram för gemenskapens åtgärder för att uppnå en hållbar användning av bekämpningsmedel
( KOM(2006)0373 – C6‑0246/2006 – 2006/0132(COD) )
Föredragande:
Michl Ebner
(*) Förfarande med associerade utskott – artikel 47 i arbetsordningen
KORTFATTAD MOTIVERING
I) Inledning
Det direktiv som lagts fram ingår i den temainriktade strategin för hållbar användning av bekämpningsmedel och därmed i det sjätte miljöhandlingsprogrammet.
Användningen av växtskyddsmedel regleras direkt eller indirekt i många av gemenskapens rättsakter, bland annat följande:
· Direktiv 91/414/EEG (utsläppande av växtskyddsmedel på marknaden), som skall ersättas av förordningen om utsläppande av växtskyddsmedel på marknaden ( KOM(2006)0388 ).
· Direktiv 79/117/EEG (förbud mot växtskyddsprodukter).
· Förordning (EG) nr 396/2005 (gränsvärden för bekämpningsmedelsrester).
· Förordning (EG) nr 882/2004 (offentliga kontroller).
· Förordning (EG) nr 178/2002 (allmänna principer och krav för livsmedelslagstiftning).
· Förordning (EG) nr 852/2004, (EG) nr 853/2004 och (EG) nr 854/2004 (det s.k. hygienpaketet).
· Förordning (EG) nr 1782/2003 (direktstöd inom jordbruket) – föreskriver tillämpning av det s.k. hygienpaketet, direktiv 91/414/EEG och förordning (EG) nr 178/2002 m.m. inom ramen för tvärvillkor.
· Direktiv 79/409/EEG (bevarande av vilda fåglar) och direktiv 79/43/EEG (habitatdirektivet).
· Direktiv 2006/60/EG (ramdirektivet om vatten), medräknat dotterdirektiv och beslut (t.ex. direktiven om grundvatten, dricksvatten och ytvatten, direktivet om miljökvalitetsnormer ( KOM(2006)0937 ), beslutet om prioriterade ämnen m.m.); i alla dessa rättsakter krävs åtgärder mot negativa effekter och utsläpp av växtskyddsmedel.
· Direktiven om skydd av arbetstagarnas hälsa.
· Direktiven om avfall.
Det finns gott om regler.
Ändå finns det tyvärr stora skillnader i fråga om laglig användning av växtskyddsmedel inom den ram som fastställs genom gemenskapsrätten och nationella bestämmelser.
Det har visserligen gjorts tydliga förbättringar under de senaste åren, men trots det hittar man fortfarande oönskade rester av växtskyddsmedel i vatten och livsmedel.
Den föreslagna rättsakten bör bidra till ytterligare harmonisering av bestämmelserna om användning av växtskyddsmedel.
Viktiga instrument som föreslås för detta är följande:
· Upprättande av nationella handlingsplaner.
· Utbildning av användarna.
· Information till allmänheten.
· Kontroll av den utrustning som används.
· Särskilt skydd av vattenmiljön, Natura 2000-områden och områden som används särskilt ofta av allmänheten (parker m.m.).
· Främjande av förfaranden som innefattar ringa användning av bekämpningsmedel, medräknat ett integrerat växtskydd (allmänt och grödspecifikt).
· Utveckling av riskindikatorer.
II) Föreslagna ändringar
Växtskyddsmedlen är en nödvändig del av det moderna jordbruket.
Viktiga aspekter av en miljö‑ och hälsovänlig användning av växtskyddsmedel ingår redan i andra gemenskapsrättsakter.
Därför måste den nationella handlingsplanen utgöra direktivets absoluta kärna.
I den nationella handlingsplanen bör medlemsstaterna med hjälp av olika frivilliga, legislativa och i förekommande fall skattemässiga åtgärder samordna all den verksamhet som krävs för att minska de återstående riskerna och förbättra den ändamålsenliga hanteringen av växtskyddsmedel.
För detta krävs det ovillkorligen bättre utbildning och information, bekämpning av punktkällor, bättre data samt insatser för att genomföra ett integrerat växtskydd i praktiken.
Kontinuerliga insatser är avgörande, eftersom rönen om ett optimalt växtskydd ständigt utvecklas: om insatserna (information, kontroller) avbryts, försämras situationen snabbt.
Med tanke på de omfattande bestämmelser som finns om användningen av växtskyddsmedel bör direktivet begränsas till bestämmelser om vad handlingsplanerna åtminstone skall innehålla.
I annat fall uppstår det, som för Natura 2000, ny gemenskapslagstiftning som klart strider mot de hittillsvarande bestämmelserna.
Ett integrerat växtskydd har också definierats i detalj redan i förslaget till förordning om utsläppande på marknaden, och det är obligatoriskt för samtliga användare från 2014.
Begränsningar för användningen av växtskyddsmedel i avrinningsområden (dricksvatten, grundvatten, vattendrag, besprutningsrestmängder) fastställs även i rättsakter på vattenpolitikens område eller rättsakter om utsläppande av växtskyddsmedel på marknaden.
Liksom för Natura 2000 räcker det i detta sammanhang att medlemsstaterna skall visa särskild uppmärksamhet i handlingsplanerna och uppföljningen av dem.
Bindande bestämmelser bör endast fastställas för områden som hittills inte har behandlats, t.ex. utbildning och fortbildning, information och användning av utrustning.
De nationella handlingsplanernas effektivitet bör förbättras jämfört med kommissionens förslag genom klara bestämmelser om uppdatering och kontroll, måttstockar för uppnåendet av målen och information till allmänheten.
För att förbättra förståelsen har begreppet ”bekämpningsmedel” ersatts med ”växtskyddsmedel”, eftersom direktivet enbart hänför sig till växtskyddsmedel.
ÄNDRINGSFÖRSLAG
Utskottet för jordbruk och landsbygdens utveckling uppmanar utskottet för miljö, folkhälsa och livsmedelssäkerhet att som ansvarigt utskott infoga följande ändringsförslag i sitt betänkande:
Kommissionens förslag
Ännu ej offentliggjort i EUT.
Parlamentets ändringar
Ändringsförslag
1
Titeln
Förslag till Europaparlamentets och rådets direktiv om upprättande av en ram för gemenskapens åtgärder för att uppnå en hållbar användning av bekämpningsmedel
Förslag till Europaparlamentets och rådets direktiv om upprättande av en ram för gemenskapens åtgärder för att uppnå en användning av växtskyddsmedel som följer principen om en hållbar utveckling
Motivering
I direktivet anges inga andra bekämpningsmedel än växtskyddsmedel.
För att tillämpningsområdet skall vara klart bör detta även anges i titeln.
Ändringsförslag
2
Skäl 3
(3) För att underlätta genomförandet av detta direktiv bör medlemsstaterna använda nationella handlingsplaner i syfte att fastställa mål för minskning av risker, inbegripet faror, och beroendet av bekämpningsmedelsanvändning och främja icke-kemiska växtskyddsalternativ.
De nationella handlingsplanerna kan samordnas med genomförandeplaner enligt annan närliggande gemenskapslagstiftning och användas för att gruppera samman mål som skall nås enligt annan gemenskapslagstiftning om bekämpningsmedel.
(3) Kärnan i detta direktiv är medlemsstaternas nationella handlingsplaner som syftar till att minska riskerna med användning av växtskyddsmedel och främja icke-kemiska växtskyddsalternativ.
De nationella handlingsplanerna bör samordnas med genomförandeplaner enligt annan närliggande gemenskapslagstiftning och användas för att gruppera samman mål som skall nås enligt annan gemenskapslagstiftning om bekämpningsmedel.
Ändringsförslag
3
Skäl 3a (nytt)
(3a) Målen med de nationella handlingsplanerna för riskminskning bör definieras så entydigt som möjligt.
Handlingsplanerna bör ses över regelbundet och uppdateras.
Inom ramen för de nationella handlingsplanerna åligger det medlemsstaterna att i enlighet med sina respektive problem och förutsättningar finna den rätta kombinationen av lagstiftningsåtgärder, frivilliga åtgärder och eventuella skatteåtgärder.
Ändringsförslag
4
Skäl 4
(4) Informationsutbytet om de mål och åtgärder som medlemsstaterna fastställer i sina nationella handlingsplaner är en mycket viktig faktor för att nå målen för detta direktiv.
Därför bör medlemsstaterna uppmanas att regelbundet lämna rapporter till kommissionen och övriga medlemsstater, särskilt om genomförandet och resultatet av nationella handlingsplaner och gjorda erfarenheter .
(4) Informationsutbytet och informationen till allmänheten om de mål och åtgärder som medlemsstaterna fastställer i sina nationella handlingsplaner är en mycket viktig faktor för att nå målen för detta direktiv.
Därför bör medlemsstaterna uppmanas att regelbundet lämna rapporter till kommissionen , vilken bör inrätta en databas på Internet som är tillgänglig för allmänheten och som gör det möjligt för allmänheten och de övriga medlemsstaterna att få information om målen med de nationella handlingsplanerna och deras resultat .
Vid utarbetandet av planerna bör åtminstone de aspekter av en hållbar användning av växtskyddsmedel som behandlas i detta direktiv kontrolleras.
Ändringsförslag
5
Skäl 6
(6) Det är önskvärt att medlemsstaterna inrättar system för utbildning av distributörer, rådgivare och yrkesmässiga användare av bekämpningsmedel så att de som använder eller kommer att använda bekämpningsmedel är fullt medvetna om möjliga hälso- och miljörisker och om lämpliga åtgärder för att minska riskerna så mycket som möjligt.
Utbildningar för yrkesmässiga användare kan samordnas med utbildningar som anordnas inom ramen för rådets förordning (EG) nr 1698/2005 av den 20 september 2005 om stöd för landsbygdsutveckling från Europeiska jordbruksfonden för landsbygdsutveckling (EJFLU).
(6) Det är önskvärt att medlemsstaterna inrättar system för kontinuerlig utbildning av distributörer, rådgivare och yrkesmässiga användare av bekämpningsmedel så att de som använder eller kommer att använda bekämpningsmedel är fullt medvetna om möjliga hälso- och miljörisker och om lämpliga åtgärder för att minska riskerna så mycket som möjligt.
Utbildningar för yrkesmässiga användare kan samordnas med utbildningar som anordnas inom ramen för rådets förordning (EG) nr 1698/2005 av den 20 september 2005 om stöd för landsbygdsutveckling från Europeiska jordbruksfonden för landsbygdsutveckling (EJFLU).
Ändringsförslag
6
Skäl 7
(7) Allmänheten bör få bättre kunskaper om de möjliga risker som är förknippade med användning av växtskyddsmedel, liksom om växtskyddsmedlens roll inom jordbruket och livsmedelsproduktionen, genom att den underrättas om fördelar och nackdelar, nytta och risker samt ansvarsfull användning av växtskyddsmedel .
Motivering
Informationskampanjerna till allmänheten bör utöver riskerna med användning av växtskyddsmedel även informera om medlens fördelar och deras betydelse för den nuvarande livsmedelsproduktionen.
Ändringsförslag
7
Skäl 9
(9) I Europaparlamentets och rådets direktiv 2006/42/EG av den 17 maj 2006 om maskiner och om ändring av direktiv 95/16/EG (omarbetning) anges regler för utsläppande av utrustning för spridning av bekämpningsmedel på marknaden som säkerställer att miljökrav uppfylls.
Ändringsförslag
8
Skäl 10
(10) Flygbesprutning av bekämpningsmedel kan ge betydande negativ påverkan på människors hälsa och på miljön, särskilt genom vindavdrift.
(10) Flygbesprutning av bekämpningsmedel kan ge betydande negativ påverkan på människors hälsa och på miljön, särskilt genom vindavdrift.
Det bör därför införas ett generellt anmälnings- eller tillståndsförfarande som avser flygbesprutning, för att säkra att flygbesprutning tillämpas endast om det innebär klara fördelar och ger miljövinster jämfört med andra spridningsmetoder eller om lämpliga alternativ saknas.
Ändringsförslag
9
Skäl 11
(11) Vattenmiljön är särskilt känslig för bekämpningsmedel .
Det är därför nödvändigt att ägna särskild uppmärksamhet åt att undvika förorening av ytvatten och grundvatten genom lämpliga åtgärder , exempelvis att skapa buffertzoner eller plantera häckar längs ytvatten för att minska vattnets exponering för vindavdrift .
Buffertzonernas omfattning bör bland annat avgöras av markförhållanden, klimat, vattendragets storlek och det aktuella områdets jordbruksförhållanden.
Användning av bekämpningsmedel i områden som används som dricksvattentäkt, på eller längs transportleder, t.ex. järnvägslinjer, på hårdgjorda eller mycket genomsläppliga ytor kan leda till högre risker för förorening av vattenmiljön.
I sådana områden bör därför användning av bekämpningsmedel begränsas så långt som möjligt, eller eventuellt undvikas helt.
(11) Vattenmiljön är särskilt känslig för växtskyddsmedel .
Det är därför viktigt att förhindra förorening av ytvatten och grundvatten genom lämpliga bestämmelser och regler för användning som skall fastställas i samband med att växtskyddsmedel godkänns .
Motivering
Vid användning av växtskyddsmedel skall man följa de produktspecifika reglerna för användning och den teknik för att minska skadeverkningarna som fastställts i samband med det officiella godkännandet.
I dessa bestämmelser regleras redan avståndet till vattendrag, så kravet på buffertzoner är onödigt.
Användningen av växtskyddsmedel i skyddsområden för dricksvattentäkter regleras dessutom redan genom nationella förordningar om dricksvatten och behöver därför inte tas upp här.
Ändringsförslag
10
Skäl 12
(12) Användning av bekämpningsmedel kan vara särskilt farlig i mycket känsliga områden, exempelvis Natura 2000-områden som är skyddade enligt rådets direktiv 79/409/EEG av den 2 april 1979 om bevarande av vilda fåglar och rådets direktiv 92/43/EEG av den 21 maj 1992 om bevarande av livsmiljöer samt vilda djur och växter.
På andra platser, exempelvis allmänna parker, sportanläggningar och lekplatser för barn, innebär det stora risker om allmänheten exponeras för bekämpningsmedel.
Användning av bekämpningsmedel i dessa områden bör därför begränsas så långt som möjligt, eller eventuellt undvikas helt .
(12) I mycket känsliga områden, exempelvis Natura 2000-områden som är skyddade enligt rådets direktiv 79/409/EEG av den 2 april 1979 om bevarande av vilda fåglar och rådets direktiv 92/43/EEG av den 21 maj 1992 om bevarande av livsmiljöer samt vilda djur och växter , kan åtgärder för att minska användningen av växtskyddsmedel vara nödvändiga om gemenskapens mål för dessa områden skall kunna uppnås.
Denna aspekt beaktas i de nationella handlingsplanerna och förvaltningsplanerna för särskilt skyddade områden .
På andra platser, exempelvis allmänna parker, sportanläggningar och lekplatser för barn, måste man i samband med godkännandet med hjälp av regler för användningen se till att allmänheten inte utsätts för någon högre risk för exponering för växtskyddsmedel eller att användningen av växtskyddsmedel minimeras .
Motivering
Den minskade användning av tillåtna växtskyddsmedel som eftersträvas är varken vetenskapligt motiverad eller acceptabel.
Genom att begränsa användningen av växtskyddsmedel i så kallade känsliga områden antyder man att användningen av dessa medel innebär en fara, som tack vare stränga statliga regler för godkännande och användning faktiskt inte existerar.
De regler för användning som fastställts i samband med godkännandeförfarandet innebär att ingen fara föreligger för människor och miljö, vilket gör ytterligare bestämmelser överflödiga.
Ändringsförslag
11
Skäl 14
(14) Om alla lantbrukare tillämpar allmänna standarder för integrerat växtskydd skulle det leda till en mer riktad användning av alla tillgängliga bekämpningsmetoder, däribland bekämpningsmedel.
Detta skulle därför bidra till att ytterligare minska riskerna för människors hälsa och för miljön.
Medlemsstaterna bör främja jordbruk med liten användning av bekämpningsmedel, särskilt integrerat växtskydd, och skapa nödvändiga förutsättningar för tillämpning av integrerat växtskydd.
Medlemsstaterna bör också uppmuntra användning av grödspecifika standarder för integrerat växtskydd.
(14) Medlemsstaterna bör inom ramen för de nationella handlingsplanerna främja förutsättningarna för att driva jordbruk med liten användning av bekämpningsmedel, särskilt ekologiskt jordbruk och integrerat växtskydd, i enlighet med definitionen i förordning (EG) nr […] om utsläppande av växtskyddsmedel på marknaden, och skapa nödvändiga förutsättningar för tillämpning av integrerat växtskydd.
Ändringsförslag
12
1.
Detta direktiv skall tillämpas på bekämpningsmedel i form av växtskyddsmedel enligt definitionen i förordning (EG) nr […] om utsläppande av växtskyddsmedel på marknaden.
1.
Detta direktiv skall tillämpas på växtskyddsmedel enligt definitionen i förordning (EG) nr […] om utsläppande av växtskyddsmedel på marknaden.
Ändringsförslag
13
b) yrkesmässig användare: en fysisk eller juridisk person som använder bekämpningsmedel i sin yrkesmässiga verksamhet , inbegripet operatörer, tekniker, arbetsgivare, egenföretagare både inom och utanför jordbrukssektorn .
Till användarna hör även golfbanor, tennisbanor och andra fritidsanläggningar, kommuner och deras parkanläggningar samt infrastrukturområden såsom parkeringsplatser, vägar, järnvägar och liknande.
Motivering
I den engelska texten används uttrycket ”professional user”, vilket betyder yrkesmässig användare.
Den tyska översättningen ”gewerblicher Anwender” är felaktig.
Direktivet bör inte bara rikta sig till jordbrukare utan till alla som använder växtskyddsmedel.
Ändringsförslag
14
d) rådgivare: en fysisk eller juridisk person som ger råd om användningen av bekämpningsmedel, inbegripet privata rådgivningsföretag, handelsagenter, livsmedelsproducenter och detaljhandlare om tillämpligt .
d) rådgivare: en fysisk eller juridisk person som besitter en av medlemsstaterna fastställd utbildningsnivå och som därigenom är behörig att ge råd om användningen av växtskyddsmedel och i det sammanhanget följer de metoder som är godkända i det land där odlingsarealerna finns samt gemenskapens gränsvärden .
Ändringsförslag
15
ia) användningsindikator: en parameter som kan användas för att bedöma intensiteten på och beroendet av användningen av bekämpningsmedel,
Ändringsförslag
16
Nationella handlingsplaner för att minska risker och beroendet av bekämpningsmedel
Nationella handlingsplaner för att minska risker och användningen av bekämpningsmedel
Ändringsförslag
17
1.
Medlemsstaterna skall anta nationella handlingsplaner för att fastställa mål, åtgärder och tidtabeller för minskning av risker , inbegripet faror, och beroendet av bekämpningsmedel .
1.
Medlemsstaterna skall efter samråd med jordbrukarnas representanter, miljöorganisationer, industrin och andra berörda parter anta nationella handlingsplaner för att fastställa mål, åtgärder och tidtabeller för minskning av de risker för hälsan och miljön som är förknippade med användningen av växtskyddsmedel.
Handlingsplanerna skall ta hänsyn till särskilda nationella, regionala och lokala förhållanden .
När medlemsstaterna upprättar och ändrar sina nationella handlingsplaner skall de ta hänsyn till de planerade åtgärdernas sociala, ekonomiska och miljömässiga effekter.
När medlemsstaterna upprättar och ändrar sina nationella handlingsplaner skall de ta hänsyn till de planerade åtgärdernas sociala, ekonomiska och miljömässiga effekter.
Den nationella handlingsplanen kan även bestå av sammanfattningar och på nationell nivå gemensamma regionala planer eller nationella och regionala planer.
Ändringsförslag
18
1a.
De nationella handlingsplanerna skall i nödvändig utsträckning innehålla information om de aspekter som anges i artiklarna 5–13.
I dessa planer bör hänsyn tas till planer som upprättats enligt andra gemenskapsbestämmelser om användning av växtskyddsmedel, t.ex. åtgärdsplaner enligt direktiv 2000/60/EG.
Åtgärderna i de nationella handlingsplanerna kan i synnerhet vara lagstiftningsåtgärder, skatteåtgärder eller frivilliga åtgärder som bör grundas på resultaten av relevanta riskbedömningar.
Motivering
I direktivet bör minimikrav på innehållet anges, eller vilka aspekter som skall kontrolleras då planerna upprättas.
Frågan om när det krävs ytterligare lagstiftning, stödåtgärder, skatteåtgärder eller andra åtgärder bör avgöras av medlemsstaterna.
Ändringsförslag
19
1b.
De nationella handlingsplanerna skall omfatta integrerat växtskydd i den mening som avses i artikel 13 och skall ge prioritet åt icke-kemiska växtskyddsåtgärder samt uppmuntra jordbrukarna att välja icke ‑kemiska växtskyddsmedel.
Ändringsförslag
20
2.
Medlemsstaterna skall inom tre år efter det att detta direktiv har trätt i kraft meddela sina nationella handlingsplaner till kommissionen och övriga medlemsstater .
2.
Medlemsstaterna skall inom tre år efter det att detta direktiv har trätt i kraft meddela sina nationella handlingsplaner till kommissionen.
De nationella handlingsplanerna skall ses över minst vart femte år och alla ändringar av de nationella handlingsplanerna skall utan onödigt dröjsmål rapporteras till kommissionen.
De nationella handlingsplanerna skall ses över minst vart femte år och uppdateras beroende på om målen uppnåtts.
Översynen skall även omfatta en analys av om riskerna har beaktats på lämpligt sätt i handlingsplanen eller om de måste ses över.
Alla ändringar av de nationella handlingsplanerna och de viktigaste resultaten av översynen skall utan onödigt dröjsmål rapporteras till kommissionen.
Motivering
Bestämmelserna om översynen måste preciseras.
Ändringsförslag
21
2a.
Kommissionen skall inrätta en databas på Internet genom vilken allmänheten ges tillgång till de nationella handlingsplanerna, alla ändringar och de viktigaste resultaten av de regelbundna översynerna, särskilt eventuella framsteg eller misslyckanden med att uppnå målen och orsakerna till detta.
Motivering
Involverandet av allmänheten är en viktig del av de nationella handlingsplanerna.
Därför bör dessa planer, ändringar och resultaten av översynen göras tillgängliga för allmänheten i hela Europa via en central databas på Internet.
I och med denna databas bortfaller medlemsstaternas skyldighet att meddela varandra, som ändå är överflödig och som i den form som föreslagits endast omfattade den ursprungliga handlingsplanen men däremot inte några ändringar.
Då information läggs ut på Internet behövs inte längre bestämmelsen om vidarebefordrande av uppgifter till tredjeländer.
Ändringsförslag
22
3.
utgår
Motivering
Ändringsförslag
23
4a.
Utarbetandet och genomförandet av gemenskapsprogram bör kunna få gemenskapsstöd.
Ändringsförslag
24
1.
Medlemsstaterna skall se till att alla yrkesmässiga användare, distributörer och rådgivare har tillgång till lämplig utbildning.
1.
Medlemsstaterna skall se till att alla yrkesmässiga användare, distributörer och rådgivare har tillgång till lämplig och fristående anordnad utbildning eller fortbildning om korrekt användning av växtskyddsmedel som motsvarar de berörda aktörernas ansvarsnivå och specifika roll inom integrerat växtskydd .
Motivering
Det är viktigt att fortbildning anordnas oberoende av vissa aktörers ekonomiska intressen.
Detta utesluter dock inte möjligheten att anlita sakkunniga från industrin eller icke-statliga organisationer.
Medlemsstaterna kan även uppfylla grundkraven enligt detta direktiv genom att erbjuda relevant utbildning.
Ändringsförslag
25
2.
2.
Motivering
Två år är en för kort tid för obligatorisk utbildning av alla lantbrukare.
Ändringsförslag
26
Ändringsförslag
27
1.
1.
Motivering
Eftersom de ramvillkor som anges i lagen och de vetenskapliga rönen om yrkesmässig användning av växtskyddsmedel enligt kommissionens konsekvensbedömning ändras fortlöpande bör intygens giltighetstid begränsas.
Ändringsförslag
28
2.
2.
Ändringsförslag
29
3.
Medlemsstaterna skall ålägga distributörer som släpper ut bekämpningsmedel för icke yrkesmässig användning på marknaden att lämna allmän information om riskerna med bekämpningsmedelsanvändning , särskilt om faror , exponering, korrekt lagring, hantering och spridning samt bortskaffande.
3.
Motivering
Syftet med att producenter och distributörer skall lämna information bör vara en yrkesmässig användning av växtskyddsmedel som i stor utsträckning avvärjer hälso- och miljöfaror.
Informationen bör syfta till att klargöra riskerna med specifika produkter, eftersom dessa kan variera betydligt allt efter medel och användningstyp.
En längre övergångsperiod behövs för att undvika överkapacitet inom utbildningsområdet under de två första åren efter det att utbildningssystemet inrättats.
Ändringsförslag
30
Artikel 7
Medlemsstaterna skall stödja informationsprogram riktade till allmänheten och underlätta allmänhetens tillgång till information om bekämpningsmedel, särskilt när det gäller hälso- och miljöeffekter och icke-kemiska alternativ.
Medlemsstaterna skall stödja informationsprogram riktade till allmänheten och underlätta allmänhetens tillgång till information om fördelar och risker med användning av växtskyddsmedel liksom om möjliga hälso- och miljöeffekter.
Dessutom skall man informera om växtskyddsmedlens roll i jordbruk och livsmedelsproduktion samt om ansvarsfull användning av växtskyddsmedel och icke-kemiska alternativ .
Motivering
Genom ändringsförslaget säkras det att informationsprogram riktade till allmänheten inte bara tar upp riskerna med användning av växtskyddsmedel.
För närvarande är det i första hand riskerna med växtskyddsmedel som tas upp offentligt.
I stället borde man sträva efter att objektivt redogöra för växtskyddsmedelsanvändningens nödvändighet och hållbarhet samt för dess betydelse inom dagens livsmedelsproduktion, såsom det anges i ändringsförslaget.
Ändringsförslag
31
1.
Medlemsstaterna skall se till att utrustning och tillbehör för spridning av bekämpningsmedel i yrkesmässig användning inspekteras med jämna mellanrum.
Medlemsstaterna skall i detta syfte införa system för intyg som gör det möjligt att styrka inspektioner.
1.
Medlemsstaterna skall införa incitamentsystem för att se till att utrustning och tillbehör för spridning av bekämpningsmedel i yrkesmässig användning inspekteras med jämna mellanrum.
Motivering
Incitamentsystem är bättre än tvångsåtgärder för att öka användarnas acceptans för inspektioner av utrustningen.
Ändringsförslag
32
3.
utgår
Motivering
Denna särskilda bestämmelse kan utgå av hänsyn till subsidiaritetsprincipen.
Ändringsförslag
33
4.
Medlemsstaterna skall utse organ med ansvar för att utföra inspektionerna och skall informera kommissionen om detta.
utgår
Motivering
Denna punkt är överflödig.
Ändringsförslag
34
1.
Medlemsstaterna skall förbjuda flygbesprutning , om inte annat följer av punkterna 2–6 .
1.
Medlemsstaterna skall fastställa bestämmelser om flygbesprutning med beaktande av punkt 4 .
Motivering
Ett allmänt förbud mot flygbesprutning är onödigt byråkratiskt och föga motiverat, eftersom det i vissa fall är uppenbart att en annan användning av växtskyddsmedel inte är aktuell (vinodling, skogar).
Medlemsstaterna bör säkra att flygbesprutning endast tillämpas i de fall då det är absolut nödvändigt.
Medlemsstaterna får avgöra om de inför ett tillståndsförfarande eller ett anmälningsförfarande.
Kraven på dokumentation är inte nödvändiga med tanke på bestämmelserna i direktivet om miljöinformation och befintliga nationella bestämmelser.
Ändringsförslag
35
2.
Medlemsstaterna skall fastställa och offentliggöra för vilka grödor och områden, samt på vilka särskilda villkor för spridning, flygbesprutning kan tillåtas genom undantag från punkt 1.
utgår
Motivering
Ändringsförslaget är en följd av de ändringar som görs till punkt 1 och punkt 4.
Ändringsförslag
36
3.
Medlemsstaterna skall utse de myndigheter som är behöriga att medge undantag och skall informera kommissionen om detta.
utgår
Motivering
Denna punkt är överflödig.
Ändringsförslag
37
4.
Undantag får medges endast om följande villkor är uppfyllda:
4.
Flygbesprutning är tillåten endast om följande villkor är uppfyllda:
(a) Det får inte finnas några lämpliga alternativ, eller också skall det innebära klara fördelar i form av minskad påverkan på hälsa och miljö jämfört med markbaserad spridning av bekämpningsmedel.
(a) Det får inte finnas några lämpliga alternativ, eller också skall det innebära klara fördelar i form av minskad påverkan på hälsa och miljö jämfört med markbaserad spridning av bekämpningsmedel.
(b) De bekämpningsmedel som används skall vara uttryckligen tillåtna för flygbesprutning.
(b) De bekämpningsmedel som används skall vara uttryckligen tillåtna för flygbesprutning.
(ca) Det skall säkras att alla nödvändiga åtgärder vidtas för att varna boende och andra närvarande personer i tid och för att skydda miljön i närheten av det besprutade området.
(cb) Flygbesprutningen skall ha förhandsanmälts till eller godkänts av den behöriga myndigheten.
Motivering
Medlemsstaterna får avgöra om de inför ett tillståndsförfarande eller ett anmälningsförfarande.
I vilket fall som helst är flygbesprutning tillåten endast om villkoren i punkt 4 uppfylls.
Kommissionens förslag var dessutom onödigt byråkratiskt.
Ändringsförslag
38
5.
En yrkesmässig användare som vill sprida bekämpningsmedel genom flygbesprutning skall lämna in en begäran till den behöriga myndigheten tillsammans med uppgifter som styrker att de villkor som anges i punkt 4 är uppfyllda.
utgår
Motivering
Ändringsförslaget är en följd av de ändringar som görs till punkt 1 och punkt 4.
Se motiveringen till ändringsförslag 34 och 37.
Ändringsförslag
39
6.
De behöriga myndigheterna skall föra register över de undantag som medges.
utgår
Motivering
Kraven på dokumentation är inte nödvändiga med tanke på bestämmelserna i direktivet om miljöinformation och befintliga nationella bestämmelser.
Ändringsförslag
40
1.
Medlemsstaterna skall, om bekämpningsmedel används i närheten av vatten, se till att företräde ges åt
1.
Då medlemsstaterna utarbetar och genomför de nationella handlingsplanerna skall de , om växtskyddsmedel används i närheten av vatten, vidta åtgärder som på lämpligt sätt ger företräde åt
Motivering
Det är fråga om problem som i första hand skall lösas av medlemsstaterna inom ramen för de nationella handlingsplanerna enligt artikel 4.
Ändringsförslag
41
1a.
Då medlemsstaterna utarbetar och genomför de nationella handlingsplanerna skall de särskilt vidta följande åtgärder för att skydda vattenförekomster:
(b) Vidta lämpliga åtgärder för att begränsa vindavdrift av växtskyddsmedel, åtminstone i högväxande grödor (odlingar av frukt, vin och humle och liknande) i direkt anslutning till ett vattendrag.
(c) Vidta lämpliga åtgärder för att spridning av bekämpningsmedel begränsas så långt som möjligt eller eventuellt undviks helt på och längs vägar, järnvägslinjer, mycket genomsläppliga ytor och annan infrastruktur nära ytvatten eller grundvatten, och på hårdgjorda ytor med hög risk för avrinning till ytvatten eller avloppssystem.
Åtgärder enligt led a skall ingå i varje nationell handlingsplan.
Motivering
Texten i punkt 1a (ny), leden a–c motsvarar i stora drag texten i punkterna 2–4 i kommissionens förslag.
Åtgärderna har samma mål och därför har de sammanfattats i en enda punkt.
Skydds- och buffertzoner för vattendrag och dricksvatten är mycket viktiga beståndsdelar i en nationell handlingsplan.
Som Danmarks exempel visar kan frivilliga åtgärder i detta sammanhang också vara lika effektiva som obligatoriska lagstiftningsförfaranden.
Ändringsförslag
42
2.
utgår
Motivering
Denna punkt ingår nu i punkt 1a (ny), led a, (se ändringsförslag 41).
Ändringsförslag
43
3.
utgår
Motivering
Denna punkt ingår nu i punkt 1a (ny), led b, (se ändringsförslag 41).
Ändringsförslag
44
4.
utgår
Motivering
Denna punkt ingår nu i punkt 1a (ny), led c, (se ändringsförslag 41).
Ändringsförslag
45
Artikel 11, inledningen
Medlemsstaterna skall, med utgångspunkt i resultaten från relevanta riskbedömningar , se till att följande åtgärder vidtas:
Motivering
Ett beslut att minska användningen av växtskyddsmedel i känsliga områden bör baseras på en relevant riskbedömning.
Syftet är inte att förbjuda användningen utan att verka för en försiktig användning av små mängder av ett växtskyddsmedel med hänsyn till det specifika skyddsmålet.
I Natura 2000-förordningarna anges förbud och krav som omfattar samtliga fall, så med hänsyn till subsidiaritetsprincipen behövs ingen ytterligare specifik lagstiftning.
Ändringsförslag
46
(a) Användning av bekämpningsmedel skall begränsas till det absolut nödvändiga eller avskaffas helt i områden som regelbundet används av allmänheten eller av känsliga befolkningsgrupper, åtminstone parker, offentliga trädgårdar, sportanläggningar och lekplatser.
Motivering
Ändringsförslaget syftar till att precisera och förtydliga.
Det som är avgörande är inte själva förbudet, utan att växtskyddsmedel används så litet som möjligt beroende på de särskilda skyddsmålsättningarna för offentliga områden.
Med tanke på att växtskyddsmedel används i liten omfattning i offentliga områden tillämpas denna bestämmelse redan i dag i stor utsträckning i medlemsstaterna.
Ändringsförslag
47
Ett förbud eller en begränsning enligt b får grundas på resultaten av relevanta riskbedömningar.
utgår
Ändringsförslag
48
Begränsningar för användning av växtskyddsmedel i Natura 2000-områden utgör inte något hinder för frivilliga stödåtgärder enligt strukturfondsförordningarna och förordningen om landsbygdsutveckling.
Motivering
Den sista meningen bör tillfogas för att klargöra att begränsningar för användning av växtskyddsmedel i Natura-2000-områden i syfte att uppnå bevarandemålen inte bryter mot frivillighetsprincipen i samband med stödåtgärder.
Hittills har kommissionens enheter inte tillhandahållit entydiga uppgifter om detta, vilket har lett till stor osäkerhet kring rättsläget i medlemsstaterna och försvårar genomförandet av åtgärder till skydd för jordbruksmiljön.
Ändringsförslag
49
1.
Medlemsstaterna skall vidta de åtgärder som behövs för att säkerställa att följande arbetsmoment inte medför risk för människors hälsa eller säkerhet eller för miljön:
1.
Medlemsstaterna skall inom ramen för de nationella handlingsplanerna och på grundval av relevanta riskbedömningar vidta de åtgärder som eventuellt behövs för att säkerställa att följande arbetsmoment inte medför risk för människors hälsa eller säkerhet eller för miljön:
Motivering
De föreslagna åtgärderna bör integreras i de nationella handlingsplanerna.
Det är främst fråga om att de befintliga bestämmelserna verkligen skall genomföras med relevanta insatser.
Det finns gott om föreskrifter i medlemsstaterna.
Ändringsförslag
50
2.
2.
Medlemsstaterna skall inom ramen för de nationella handlingsplanerna och på grundval av relevanta riskbedömningar vidta de åtgärder som eventuellt behövs för att undvika farliga moment i hanteringen av bekämpningsmedel som är tillåtna för icke yrkesmässig användning.
Motivering
Se motiveringen till ändringsförslag 49.
Ändringsförslag
51
3.
3.
Medlemsstaterna skall inom ramen för de nationella handlingsplanerna och på grundval av relevanta riskbedömningar vidta de åtgärder som eventuellt behövs för att säkra att lagringsplatser för bekämpningsmedel utformas på ett sådant sätt att oönskade utsläpp undviks.
Motivering
Se motiveringen till ändringsförslag 49.
Ändringsförslag
52
1.
Medlemsstaterna skall vidta alla åtgärder som behövs för att främja jordbruk med små insatser av bekämpningsmedel, däribland integrerat växtskydd , och för att säkerställa att yrkesmässiga användare av bekämpningsmedel går över till en mer miljövänlig användning av alla tillgängliga växtskyddsåtgärder, företrädesvis lågriskalternativ om sådana kan användas och i annat fall produkter som, av de produkter som är tillgängliga för samma skadegörarproblem, ger minst påverkan på människors hälsa och på miljön .
1.
Medlemsstaterna skall inrätta incitamentsystem för att främja jordbruk med små insatser av bekämpningsmedel, däribland integrerat växtskydd.
Motivering
Incitamentsystem är bättre än tvångsåtgärder för att öka användarnas acceptans för små insatser av växtskyddsmedel eller integrerat växtskydd.
Dessutom bör påpekas att växtskyddsmedlens effekter på människors hälsa och miljön kontrolleras i samband med godkännandeförfarandet.
Man kan utgå från att godkända växtskyddsmedel om de används korrekt bara har effekt på föremålet för behandlingen.
Ändringsförslag
53
2.
utgår
Motivering
Texten har infogats i punkt 1 (se ändringsförslag 52).
Ändringsförslag
54
5.
utgår
Motivering
Punkt 5 regleras redan i artikel 52 i förordningen om utsläppande av växtskyddsmedel på marknaden.
Ändringsförslag
55
6.
utgår
Ändringsförslag
56
7.
7.
För att bistå medlemsstaterna kan kommissionen utarbeta allmänna standarder för integrerad odling som avses i punkt 1 i enlighet med det förfarande som anges i artikel 52 i förordning (EG) nr […].
Detta skall uppmuntra till offentligt deltagande av berörda parter.
Ändringsförslag
57
8.
utgår
Motivering
Införandet av grödspecifika EU-standarder för integrerat växtskydd bör avvisas eftersom gemensamma standarder inte tar hänsyn till skillnaderna i natur- och klimatförhållanden mellan olika odlingsplatser i Europa och strider mot en syn på integrerad odling som innebär att alla åtgärder bör anpassas till lokala förhållanden.
Ändringsförslag
58
8a.
Skyldigheten för mottagare av direktbetalningar enligt artikel 3 och bilaga III till förordning (EG) nr 1782/2003 skall anses vara uppfylld i fråga om användningen av växtskyddsmedel, då styrkta intyg på en utbildnings- eller fortbildningsomgång enligt artiklarna 5 och 6 samt användning av utrustning som uppfyller kraven i artikel 8 har lagts fram.
Motivering
En mycket viktig förutsättning för korrekt användning av växtskyddsmedel är att man har relevanta kunskaper och att utrustningen fungerar som den skall.
Därför förefaller det tillräckligt att lägga fram intyg över utbildning och utrustning som styrker efterlevnaden av tvärvillkoren.
Om man i samband med kontroller av andra bestämmelser (samkörning av uppgifter) ändå fastställer brott mot reglerna, skall påföljder enligt förordning (EG) nr 1782/2003 naturligtvis göras gällande även i fortsättningen.
Ändringsförslag
59
1.
Medlemsstaterna får, fram till dess att indikatorerna har fastställts, fortsätta att använda befintliga nationella indikatorer eller fastställa andra lämpliga indikatorer.
1.
Medlemsstaterna får, fram till dess att indikatorerna har fastställts, fortsätta att använda befintliga nationella indikatorer eller fastställa andra lämpliga indikatorer.
Motivering
Det bör även fastställas indikatorer för användningen av bekämpningsmedel.
Ändringsförslag
60
2.
2.
Motivering
Om statistikförordningen inte antas bör andra statistiska uppgifter användas.
Ändringsförslag
61
a) Beräkning av gemensamma och harmoniserade riskindikatorer på nationell nivå.
a) Beräkning av gemensamma och harmoniserade risk- och användningsindikatorer på nationell nivå.
Motivering
Se ändringsförslag 59.
Ändringsförslag
62
ba) Fastställande av trender för förekomsten av skadegörare och sjukdomar samt utvecklingen av svamp.
Motivering
Man måste även fokusera på ovannämnda frågor eftersom också de påverkar riskindikatorerna för användningen av växtskyddsmedel.
Ändringsförslag
63
ca) Utarbetande, utvärdering och anpassning av de nationella handlingsplanerna.
Ändringsförslag
64
3.
3.
Medlemsstaterna skall meddela kommissionen resultaten av de utvärderingar som gjorts enligt punkt 2.
Motivering
Ändringsförslag
65
4.
4.
Ändringsförslag
66
Motivering
Ändringsförslag
67
5.
5.
Motivering
Se ändringsförslag 59.
Ändringsförslag
68
5a.
När uppgifter samlas in bör man se till att gemenskapens jordbrukare inte belastas med ytterligare dokumentationsskyldigheter och orimliga anmälnings- och rapporteringsskyldigheter.
Motivering
Jordbrukarna omfattas redan av en bred dokumentations- och rapporteringsskyldighet.
Om det i framtiden utarbetas en förordning med statistik för växtskyddsmedel bör man se till att det inte uppstår ytterligare orimliga anmälnings-, rapporterings- och dokumentationsskyldigheter för jordbrukarna.
Det borde räcka med regelbundna stickprov etc. som görs på frivillig basis eller som är resultaten av kontroller som ändå skall genomföras.
Ändringsförslag
69
Artikel 15
Kommissionen skall regelbundet lämna en rapport till Europaparlamentet och rådet om framstegen i genomförandet av detta direktiv, vid behov tillsammans med förslag till ändringar.
Kommissionen skall regelbundet , dock minst vart femte år, lämna en rapport till Europaparlamentet och rådet om framstegen i genomförandet av detta direktiv, vid behov tillsammans med förslag till ändringar.
Motivering
Anpassning av de tidsfrister som även omfattar kontrollen av planerna.
Ändringsförslag
70
Artikel 15a (ny)
Artikel 15a
Kommissionen skall inrätta en europeisk fond för småskalig användning i syfte att uppmuntra forskningsinstitut i medlemsstaterna att samarbeta inom forskning om användning av grödor i småskalig odling.
I anslutning till fonden skall kommissionen inrätta en plattform för utbyte av information och bästa praxis när det gäller växtskyddsmedel i småskalig odling och hållbar användning av växtskyddsmedel.
Ändringsförslag
71
Medlemsstaterna skall fastställa påföljder för överträdelser av de nationella bestämmelser som antas i enlighet med detta direktiv och skall vidta alla åtgärder som behövs för att säkerställa att de tillämpas.
Påföljderna skall vara effektiva, proportionella och avskräckande.
Medlemsstaterna skall fastställa påföljder för överträdelser av de nationella bestämmelser som antas i enlighet med artiklarna 6, 8 och 9 i detta direktiv och skall vidta alla åtgärder som behövs för att säkerställa att de tillämpas.
Påföljderna skall vara effektiva, proportionella och avskräckande.
Motivering
Precisering av bestämmelsen om påföljder.
Ändringsförslag
72
Artikel 16a (ny)
Artikel 16a
Bestämmelserna i direktiv 2004/35/EG skall inte tillämpas när jordbrukare använder växtskyddsmedel i enlighet med godkännandebestämmelserna.
Motivering
Jordbrukare som följer befintliga regler för växtskyddsmedel bör inte hållas ansvariga för miljöskador enligt direktiv 2004/35/EG.
Om godkända växtskyddsmedel används i enlighet med reglerna för användning bör jordbrukaren befrias från ansvar enligt artikel 3.1 i direktiv 2004/35/EG.
Ändringsförslag
73
2.
utgår
Motivering
Korrigering av ett redaktionellt misstag.
Hänvisningen till beslut 1999/468/EG är överflödig, eftersom det inte hänvisas till detta förfarande på något ställe i texten.
Ändringsförslag
74
3.
3.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
Motivering
Ändringsförslag
75
Motivering
Titel
Ramdirektiv om hållbar användning av bekämpningsmedel
Referensnummer
KOM(2006)0373 – C6-0246/2006 – 2006/0132(COD)
Ansvarigt utskott
ENVI
Yttrande
Tillkännagivande i kammaren
AGRI
5.9.2006
Förstärkt samarbete – tillkännagivande i kammaren
5.9.2006
Föredragande av yttrande
Utnämning
Michl Ebner
11.9.2006
Behandling i utskott
21.11.2006
27.2.2007
21.3.2007
12.4.2007
Antagande
12.4.2007
Slutomröstning: resultat
+:
–:
0:
36
2
1
Slutomröstning: närvarande ledamöter
Vincenzo Aita, Katerina Batzeli, Sergio Berlato, Thijs Berman, Niels Busk, Luis Manuel Capoulas Santos, Giuseppe Castiglione, Dumitru Gheorghe Mircea Coşea, Joseph Daul, Albert Deß, Gintaras Didžiokas, Michl Ebner, Carmen Fraga Estévez, Duarte Freitas, Lutz Goepel, Friedrich-Wilhelm Graefe zu Baringdorf, Elisabeth Jeggle, Heinz Kindermann, Diamanto Manolakou, Mairead McGuinness, Rosa Miguélez Ramos, Neil Parish, Radu Podgorean, María Isabel Salinas García, Agnes Schierhuber, Willem Schuth, Czesław Adam Siekierski, Alyn Smith, Marc Tarabella, Jeffrey Titford, Witold Tomczak, Donato Tommaso Veraldi, Janusz Wojciechowski
Slutomröstning: närvarande suppleanter
Herbert Bösch, Bernadette Bourzai, Béla Glattfelder, Christa Klaß, Wiesław Stefan Kuc, Astrid Lulling, Jan Mulder
ÄRENDETS GÅNG
Titel
Ramdirektiv om hållbar användning av bekämpningsmedel
Referensnummer
KOM(2006)0373 – C6-0246/2006 – 2006/0132(COD)
Framläggande för parlamentet
12.7.2006
Ansvarigt utskott
Tillkännagivande i kammaren
ENVI
5.9.2006
Rådgivande utskott
Tillkännagivande i kammaren
ITRE
5.9.2006
AGRI
5.9.2006
Förstärkt samarbete
Tillkännagivande i kammaren
ENVI
29.11.2006
Föredragande
Utnämning
Christa Klaß
3.10.2006
Bestridande av den rättsliga grunden
JURI:s yttrande
JURI
11.9.2007
Behandling i utskott
26.2.2007
5.6.2007
Antagande
26.6.2007
Slutomröstning: resultat
+:
–:
0:
34
11
5
Slutomröstning: närvarande ledamöter
Adamos Adamou, Georgs Andrejevs, Margrete Auken, Pilar Ayuso, Irena Belohorská, Johannes Blokland, Hiltrud Breyer, Dorette Corbey, Chris Davies, Edite Estrela, Jill Evans, Anne Ferreira, Karl-Heinz Florenz, Matthias Groote, Cristina Gutiérrez-Cortines, Satu Hassi, Gyula Hegyi, Jens Holm, Caroline Jackson, Dan Jørgensen, Christa Klaß, Aldis Kušķis, Roberto Musacchio, Riitta Myller, Péter Olajos, Miroslav Ouzký, Vladko Todorov Panayotov, Vittorio Prodi, Guido Sacconi, Richard Seeber, Bogusław Sonik, María Sornosa Martínez, Antonios Trakatellis, Evangelia Tzampazi, Thomas Ulmer, Anja Weisgerber, Åsa Westlund, Anders Wijkman, Glenis Willmott
Slutomröstning: närvarande suppleanter
Jens-Peter Bonde, Christofer Fjellner, Monica Frassoni, Ambroise Guellec, Erna Hennicot-Schoepges, Anne Laperrouze, Kartika Tamara Liotard, David Martin, Renate Sommer, Lambert van Nistelrooij
Slutomröstning: närvarande suppleanter (art.
178.2)
Gabriela Creţu
A6-0415/2007
Föredragande:
Pál Schmitt
PE 390.450v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING..........................................................................................................................12
YTTRANDE från utskottet för sysselsättning och sociala frågor ...15
YTTRANDE från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män 20
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om idrottens roll i utbildningen
( 2007/2086(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av artiklarna 149, 150 och 152 i EG‑fördraget,
– med beaktande av Helsingforsrapporten och Niceförklaringen om idrottens särdrag och sociala funktion i Europa,
– med beaktande av kommissionen vitbok om idrott ( KOM(2007)0391 ),
– med beaktande av kommissionens vitbok om en EU-strategi för hälsofrågor som rör kost, övervikt och fetma ( KOM(2007)0279 ),
– med beaktande av kommissionens utvärdering av Europeiska året för utbildning genom idrott 2004 ( KOM(2005)0680 ),
– med beaktande av Europarådets rekommendation om förbättrad idrottsutbildning och idrott för barn och ungdomar i alla Europas länder (Rec(2003)6),
– med beaktande av kommissionens grönbok ”Främja goda kostvanor och motion: En europeisk dimension i arbetet för att förebygga övervikt, fetma och kroniska sjukdomar” ( KOM(2005)0637 ),
– med beaktande av den studie som har offentliggjorts av Europaparlamentet med titeln ”Current situation and prospects for physical education in the European Union”,
– med beaktande av sin resolution av den 13 juni 1997 om Europeiska unionens roll på idrottens område
EGT C 200, 30.6.1997, s.
244. ,
– med beaktande av sin resolution av den 29 mars 2007 om framtiden för professionell fotboll i Europa
Antagna texter, P6_TA(2007)0100 . ,
– med beaktande av resolutionen av den 14 april 2005 om dopning inom idrotten
EUT C 33, 9.2.2006, s.
497. ,
– med beaktande av artiklarna I–17 och III–282 i fördraget om upprättande av en konstitution för Europa (konstitutionsfördraget),
– med beaktande av artikel 45 i arbetsordningen,
– med beaktande av betänkandet från utskottet för kultur och utbildning och yttrandena från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män och utskottet för sysselsättning och sociala frågor ( A6‑0415/2007 ), och av följande skäl:
A. Idrott är det enda skolämne som syftar till att förbereda barn för en sund livsstil och inriktas på deras totala fysiska och mentala utveckling, samt erbjuder viktiga sociala värden, såsom rättvisa, självdisciplin, solidaritet, laganda, tolerans och rent spel.
B. Övervikt som orsakas av en stillasittande livsstil och felaktig kost och som kan leda till dålig hälsa och psykosociala problem och sjukdomar som medför kostnadskrävande komplikationer, t.ex. högt blodtryck, diabetes och hjärt- och kärlsjukdomar, drabbar en allt större del av EU:s befolkning, varav ungefär en fjärdedel är barn.
C. Skolidrott är ett av de viktigaste redskapen för social integration, men för vissa minoriteter och religiösa samfund, och för funktionshindrade barn, är ett fullt deltagande i skolidrotten i många fall inte säkerställt och är förknippat med problem, som är svåra att lösa.
D. Antalet lektioner som avsätts för idrott har minskat på såväl grundskolenivå som gymnasienivå under det senaste årtiondet, och tillhandahållandet av idrottsanläggningar och utrustning skiljer sig stort mellan medlemsstaterna.
E. Medlemsstaternas utbildningsprogram för idrottslärare skiljer sig mycket åt, och det blir allt vanligare att idrottsundervisningen i skolan ges av lärare med otillräcklig utbildning.
F. Det finns ingen lämplig samordning för att förena idrottsaktiviteter i och utanför skolan och utnyttja befintliga idrottsanläggningar på ett bättre sätt, och kopplingen mellan dem skiljer sig åt mellan olika medlemsstater.
G. Föräldrarna kan spela en avgörande roll i nätverket av partnerskap inom detta område och föräldrars stöd för barnens idrottsaktiviteter är mycket viktigt, eftersom de utgör en förebild för sina barn och det är de som ser till att barnen får tillgång till idrottsanläggningar och program.
H. De rättsliga ramar som styr skolidrott och idrott, och de som styr EU:s finansiering av dessa verksamheter, är båda lika osäkra.
I. Folkhälsa och skydd av minderåriga är prioriterade områden i EU och därför bör särskild vikt läggas vid kampen mot dopning inom idrotten.
Europaparlamentet betonar vikten av att genomföra Amsterdamförklaringen och Niceförklaringen, särskilt när det gäller de särskilda kännetecken för idrott och idrottens sociala funktion i Europa som bör beaktas vid genomförande av den gemensamma politiken.
Europaparlamentet välkomnar de informella arbetsgrupper för idrott som kommissionen och rådet inrättat och föreslår att arbetsgrupperna uttryckligen fäster större uppmärksamhet vid att stärka sambandet mellan hälsa och skolidrott.
Europaparlamentet uppmanar medlemsstaterna att överväga och när så är nödvändigt ändra inriktningen för idrotten som skolämne, med hänsyn till barns hälsomässiga och sociala behov och förväntningar.
Europaparlamentet välkomnar den tidigare omnämnda kommissionens vitbok om en EU‑strategi för hälsofrågor som rör kost, övervikt och fetma, där förebyggande åtgärder prioriteras, huvudsakligen motion och ett ökat antal deltagare i idrott.
Europaparlamentet uppmanar medlemsstaterna att skapa förutsättningar för att det föreskrivna minimiantalet idrottslektioner ska kunna uppfyllas, med tanke på att regelbunden motion bidrar väsentligt till att sänka sjukvårdskostnaderna.
Europaparlamentet uppmanar kommissionen, rådet och medlemsstaterna att, samtidigt som subsidiaritetsprincipen beaktas, inrätta lämpliga rättsliga instrument som kan främja en ökning av investeringarna i ungdomars idrottsaktiviteter och idrottsutrustning.
Europaparlamentet uppmanar alla medlemsstater att intensifiera idrottsprogram och skolidrott för ungdomar från rehabiliteringscentrum för minderåriga, eftersom idrott är medel för socialisering, kommunikation, social integrering och samtidigt lär ut laganda, rättvisa och respekt för regler.
51.
EUT C 68 E, 18.3.2004, s.
605. .
58.
MOTIVERING
Syftet med detta betänkande är främst att behandla skolidrott.
Med skolidrott avses ett lagstadgat ämne i skolans läroplan, som handlar om att utveckla elevernas fysiska kompetens och självförtroende och deras förmåga att använda detta för att lyckas i många olika aktiviteter.
Skolidrott handlar om att lära sig färdigheterna, utveckla mentala förutsättningar och den förståelse som behövs för att delta i fysiska aktiviteter, kännedom om den egna kroppen och dess rörelser och kapacitet till rörelse samt livslånga fysiska aktiviteter som är gynnsamma för hälsan.
”Idrott” har däremot en mycket bredare betydelse och är ett starkt skiftande socialt fenomen som omfattar olika former av fysiska aktiviteter, från tävlingar på hög nivå genom skolan, klubbar eller program som organiseras i samhället till spontan och informell fysisk aktivitet.
Skolan är den perfekta miljön för att främja fysisk aktivitet och en positiv inställning till regelbundna fysiska aktiviteter.
Barn och ungdomar från alla sociala bakgrunder finns regelbundet på plats under minst elva år av sitt liv.
Skolan har även i allmänhet en grundläggande funktion som en plats för lärande.
För närvarande påpekas det dock ofta att skolan inte når upp till sin potential när det gäller att främja fysisk aktivitet.
Den centrala frågan är därför inte om skolidrotten är nyttig eller ej, utan frågan är: vilka förutsättningar är nödvändiga för att skolidrotten ska ge gynnsamma resultat?
Det är denna fråga som behandlas i betänkandet
Se även: Current situation and prospects for physical education in the European Union, studie beställd av Europaparlamentet.
Författare: Ken Hardman, University of Worcester, Bryssel 2007. .
Hälsoproblem
Den allt högre förekomsten av fetma i Europa, särskilt bland ungdomar, är alarmerande och ett stort folkhälsoproblem.
Antalet barn som lider av övervikt och fetma beräknas öka med mer än 400 000 varje år inom EU, utöver de mer än 14 miljoner EU-medborgare som redan är överviktiga (däribland minst 3 miljoner överviktiga barn)
Spanien, Portugal och Italien rapporterar att över 30 procent av barnen mellan 7 och 11 år lider av övervikt och fetma.
Ökningstakten för övervikt och fetma hos barn varierar, och ökningen är kraftigast i Storbritannien och Polen.
Generellt är barn i sämre form än generationerna på 1970- och 1980-talen.
Det finns en stark tendens att övervikten fortsätter att öka från barndomen till medelåldern.
Det är därför viktigt att uppnå en optimal kroppsvikt under hela livet.
Utöver det mänskliga lidande som fetma orsakar är de ekonomiska konsekvenserna av den ökande fetman betydande.
Det beräknas att fetma står för upp till 7 procent av sjukvårdskostnaderna inom EU, och detta belopp kommer att öka ytterligare med tanke på de ökande tendenserna till fetma.
Dessutom har ett antal ”vuxensjukdomar”, exempelvis benskörhet och kranskärlssjukdomar, sitt ursprung i barndomen, och kan delvis mildras genom regelbunden fysisk aktivitet under de tidiga barndomsåren.
Det finns även relativt konsekventa belägg för att regelbunden fysisk aktivitet kan ha en positiv effekt på barns och ungdomars psykologiska välbefinnande, särskilt när det gäller barns självkänsla, och framför allt i missgynnade grupper, bland andra personer med inlärningssvårigheter eller låg självkänsla.
Social kompetens, moralisk utbildning, integration och minskad brottslighet
Idrotten ger med sina bakomliggande begrepp ”rättvisa” och ”frihet” ett rikt sammanhang för att främja den sociomoraliska utvecklingen.
Idrott och skolidrott utgör en effektiv ram för främjandet av personligt och socialt ansvarstagande.
Det har påpekats att det finns ett samband mellan deltagandet i idrott och fysisk aktivitet och sociala relationer och social integration.
I moderna samhällen har ungdomar sämre möjligheter att falla tillbaka på varaktiga sociala band än tidigare.
Detta gör sociala nätverk – däribland skolan och klassen – mycket viktiga.
Uteslutande från gruppen, social isolering, leder till extrem stress.
Integration är däremot bra för självkänslan.
Skolidrott och idrott i allmänhet betraktas som ett viktigt sätt att motverka tendenserna till splittring eftersom idrott ger möjlighet att känna tillhörighet, att uppleva en ”vi‑känsla”, samhällsanda och solidaritet.
Genom idrotten tar man till sig normer, värderingar och färdigheter som kan vara mycket värdefulla i andra sammanhang.
Det finns även starka tecken på att idrott kan bidra till att förebygga brottslighet, inom både rehabilitering och brottsförebyggande.
II.
IDENTIFIERADE PROBLEM
Det finns ett antal problem kring skolidrotten i EU:
Om skolidrotten ska kunna bli ett effektivt instrument för att bekämpa fetma och övervikt bland barn måste aktiviteter i läroplanen som är lockande för alla elevgrupper främjas.
När dataspel blir en allt populärare hobby bland barn växer behovet av att främja en aktiv, sund livsstil bland barn och ungdomar.
För dessa unga befolkningsgrupper har det traditionella innehållet i skolidrotten liten relevans för deras livsstil.
Ø Skolidrotten riskerar att marginaliseras ytterligare inom skoldagen – de senaste åren har den tid som avsätts för skolidrott gradvis minskat inom hela EU.
Sedan 2002 har den avsatta tiden minskat från 121 till 109 minuter per vecka för grundskolan och från 117 till 101 minuter för gymnasiet
Se ”Current situation and prospects for physical education in the European Union”. – forskare rekommenderar att barn och ungdomar ska utföra någon form av fysisk aktivitet i 60 minuter varje dag!
Det finns tecken på att den officiellt redovisade timantalet för skolidrott inte motsvarar verkligheten, eftersom genomförandet inte uppfyller de juridiska kraven eller förväntningarna.
En kontroll av den verkliga situationen är nödvändig!
Ø En närmare granskning av läroplanerna för idrottslärare för att stödja en lärarutbildning av hög kvalitet är nödvändig.
Det måste finnas kompetenta och engagerade lärare som kan utforma idrottslektioner för att motverka hälsoproblem och motivera alla barn att delta.
En effektiv och framgångsrik skolidrott kräver välutbildade idrottslärare med specialkompetens.
Ø Det finns en klyfta mellan skolidrotten och aktiviteter utanför och efter skoltid.
Kopplingen mellan skolan och fritidsaktiviteter skulle kunna stärkas.
Ø Integration : deltagandet i idrottsaktiviteter är särskilt lågt bland etniska minoriteter.
Problemet med deltagande uppstår redan under skoltid – muslimska flickor är en särskilt känslig grupp i detta avseende.
Ett liknande mönster med begränsad tillgång syns bland funktionshindrade ungdomar.
Det är mycket mindre sannolikt att funktionshindrade ungdomar deltar i idrottsaktiviteter utanför läroplanen eller efter skoltid.
Ø Det finns fortfarande en brist på empiriska data på många områden när det gäller idrott, skolidrott och deras effekter på hälsa och sociala trender.
YTTRANDE från utskottet för sysselsättning och sociala frågor
till utskottet för kultur och utbildning
över idrottens roll i utbildningen
( 2007/2086(INI) )
Föredragande:
Evangelia Tzampazi
FÖRSLAG
Utskottet för sysselsättning och sociala frågor uppmanar utskottet för kultur och utbildning att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet erkänner att sport är en sektor som genererar arbetstillfällen och att andra områden, såsom utbildning, medicin, media samt tillverkning och marknadsföring av specialutrustning och specialiserade produkter har ett direkt samband med denna sektor.
Mot bakgrund av Europeiska kommissionens motsedda vitbok om idrott anser Europaparlamentet att det är viktigt att inkludera finansieringsmöjligheter för idrottsrelaterade aktiviteter med koppling till de mål som anges i artikel 149 i EG‑fördraget.
ÄRENDETS GÅNG
Titel
Idrottens roll i utbildningen
Förfarandenummer
2007/2086(INI)
Ansvarigt utskott
CULT
EMPL 24.5.2007
Förstärkt samarbete – tillkännagivande i kammaren
No
Föredragande av yttrande Utnämning
Evangelia Tzampazi 18.1.2006
Tidigare föredragande av yttrande
Behandling i utskott
8.5.2007
14.5.2007
5.6.2007
Antagande
7.6.2007
Slutomröstning: resultat
+:
–:
0:
38
1
Slutomröstning: närvarande ledamöter
Jan Andersson, Alexandru Athanasiu, Emine Bozkurt, Iles Braghetto, Philip Bushill-Matthews, Milan Cabrnoch, Ole Christensen, Derek Roland Clark, Luigi Cocilovo, Proinsias De Rossa, Harlem Désir, Harald Ettl, Richard Falbr, Ilda Figueiredo, Joel Hasse Ferreira, Stephen Hughes, Ona Juknevičienė, Jan Jerzy Kułakowski, Jean Lambert, Raymond Langendries, Elizabeth Lynne, Mary Lou McDonald, Thomas Mann, Ana Mato Adrover, Elisabeth Morin, Csaba Őry, Marie Panayotopoulos-Cassiotou, Kathy Sinnott, Jean Spautz, Gabriele Stauner, Anne Van Lancker, Gabriele Zimmer
Slutomröstning: närvarande suppleanter
Udo Bullmann, Françoise Castex, Monica Maria Iacob-Ridzi, Sepp Kusstatscher, Mario Mantovani, Dimitrios Papadimoulis, Evangelia Tzampazi
Slutomröstning: närvarande suppleanter (art.
178.2)
YTTRANDE från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
till utskottet för kultur och utbildning
över idrottens roll i utbildningen
( 2007/2086(INI) )
Föredragande:
Christa Prets
FÖRSLAG
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män uppmanar utskottet för kultur och utbildning att som ansvarigt utskott införliva följande förslag i sitt resolutionsförslag:
Europaparlamentet vill lyfta fram att ett av idrottens fostrande och sociala värden är dess förmåga att på ett effektivt sätt bekämpa rasism och främlingsfientlighet och dess integrations- och jämlikhetsaspekt i samband med likabehandling och lika möjligheter för kvinnor och män.
Europaparlamentet påminner om sin resolution av den 5 juni 2003 om kvinnor och idrott
EUT C 68E, 18.3.2004, s.
Europaparlamentet begär att medlemsstaterna ägnar särskild uppmärksamhet åt fall då barns talanger exploateras för att de ska lyckas i idrottstävlingar och insisterar på att professionell idrottsaktivitet som inbegriper barn måste ske med respekt för barnens grundläggande rättigheter och att barnens intresse alltid måste komma i första rummet.
Europaparlamentet uppmanar medlemsstaterna och de behöriga myndigheterna att garantera att kvinnor och män representeras jämlikt i de beslutsfattande organen i alla idrottsföreningar och berörda myndigheter samt arbeta för att ge kvinnor ledande ställningar genom positiv särbehandling, med beaktande av de otaliga resolutioner som avgetts om detta ämne.
ÄRENDETS GÅNG
Titel
Idrottens roll i utbildningen
Förfarandenummer
2007/2086(INI)
Ansvarigt utskott
CULT
Yttrande Tillkännagivande i kammaren
FEMM 26.4.2007
Förstärkt samarbete – tillkännagivande i kammaren
Föredragande av yttrande Utnämning
Christa Prets 27.4.2007
Tidigare föredragande av yttrande
Behandling i utskott
4.6.2007
25.6.2007
Antagande
25.6.2007
Slutomröstning: resultat
+:
–:
0:
22
Slutomröstning: närvarande ledamöter
Edit Bauer, Emine Bozkurt, Esther De Lange, Edite Estrela, Věra Flasarová, Esther Herranz García, Urszula Krupa, Pia Elda Locatelli, Marie Panayotopoulos-Cassiotou, Zita Pleštinská, Christa Prets, Raül Romeva i Rueda, Amalia Sartori, Eva-Britt Svensson, Anna Záborská
Slutomröstning: närvarande suppleanter
Gabriela Creţu, Anna Hedh, Mary Honeyball, Elisabeth Jeggle, Maria Petre, Feleknas Uca, Corien Wortmann-Kool
Slutomröstning: närvarande suppleanter (art.
178.2)
Anmärkningar (tillgängliga på ett enda språk)
...
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
10.9.2007
Slutomröstning: resultat
+:
–:
0:
19
1
Slutomröstning: närvarande ledamöter
Ivo Belet, Giovanni Berlinguer, Marie-Hélène Descamps, Milan Gaľa, Ovidiu Victor Ganţ, Vasco Graça Moura, Luis Herrero-Tejedor, Ruth Hieronymi, Manolis Mavrommatis, Ljudmila Novak, Doris Pack, Pál Schmitt, Hannu Takkula, Helga Trüpel, Henri Weber, Thomas Wise, Tomáš Zatloukal
Slutomröstning: närvarande suppleant(er)
Erna Hennicot-Schoepges, Elisabeth Morin, Christel Schaldemose
Slutomröstning: närvarande suppleant(er) (art.
178.2)
A6-0038/2008
***I
BETÄNKANDE
om förslaget till Europaparlamentets och rådets förordning om gemensamma regler för tillträde till den internationella marknaden för godstransporter på väg (omarbetning)
(KOM(2007)0265 – C6‑0146/2007 – 2007/0099(COD))
Utskottet för transport och turism
Föredragande:
Mathieu Grosch
(Omarbetning – artikel 80a i arbetsordningen)
PR_COD_1amRecast
PE 396.395v03-00
Teckenförklaring
* Samrådsförfarandet
majoritet av de avgivna rösterna
**I Samarbetsförfarandet (första behandlingen)
majoritet av de avgivna rösterna
**II Samarbetsförfarandet (andra behandlingen)
majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten
*** Samtyckesförfarandet
majoritet av parlamentets samtliga ledamöter utom i de fall som avses i artiklarna 105, 107, 161 och 300 i EG-fördraget och artikel 7 i EU-fördraget
***I Medbeslutandeförfarandet (första behandlingen)
majoritet av de avgivna rösterna
***II Medbeslutandeförfarandet (andra behandlingen)
majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten
majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
***III Medbeslutandeförfarandet (tredje behandlingen)
majoritet av de avgivna rösterna för att godkänna det gemensamma utkastet
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................22
BILAGA 1: SKRIVELSE FRÅN UTSKOTTET FÖR RÄTTSLIGA FRÅGOR........................24
BILAGA 2: SKRIVELSE FRÅN DE JURIDISKA AVDELNINGARNAS RÅDGIVANDE GRUPP 26
ÄRENDETS GÅNG..................................................................................................................28
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till Europaparlamentets och rådets förordning om gemensamma regler för tillträde till den internationella marknaden för godstransporter på väg (omarbetning)
( KOM(2007)0265 – C6-0146/2007 – 2007/0099(COD) )
(Medbeslutandeförfarandet: första behandlingen – omarbetning)
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2007)0265 ),
EGT C 77, 28.3.2002, s.
1. ,
– med beaktande av skrivelsen från utskottet för rättsliga frågor av den 20 november 2007, i enlighet med artikel 80a.3 i arbetsordningen,
– med beaktande av artiklarna 80a och 51 i arbetsordningen,
2.
3.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
Kommissionens förslag
Parlamentets ändringar
Ändringsförslag
1
Skäl 4a (nytt)
(4a) Ankommande eller avgående transport av gods på väg inom ramen för kombinerad transport enligt bestämmelserna i rådets direktiv 92/106/EEG av den 7 december 1992 om gemensamma regler för vissa former av kombinerad transport av gods mellan medlemsstaterna 1 , och därmed kombinerad järnvägs- och vägtransport och/eller vatten- och vägtransport i båda riktningarna, omfattas inte av definitionen för cabotage.
____________
1 EGT L 368, 17.12.1992, s.
38.
Direktivet senast ändrat genom direktiv 2006/103/EG (EUT L 363, 20.12.2006, s.
344).
Motivering
Gällande praxis i vissa medlemsstater tyder på en annan trend, men det kan eller får inte vara avsikten.
Ändringsförslag
2
Skäl 9
(9) Det bör också skapas ett förartillstånd som gör det möjligt för medlemsstaterna att på ett effektivt sätt kontrollera om förare från tredjeländer har en laglig anställning eller står till förfogande för det transportföretag som ansvarar för en viss transport.
(9) Det bör också skapas ett förartillstånd som gör det möjligt för medlemsstaterna att på ett effektivt sätt kontrollera om förare från tredjeländer har en laglig anställning eller står till förfogande för det transportföretag som ansvarar för en viss transport.
Förartillståndet bör vara förståeligt för alla som utför sådana kontroller.
Motivering
Förtydligande.
Ändringsförslag
25
Skäl 11
(11) Tidigare har sådana nationella transporter varit tillåtna om det har rört sig om trafik av tillfällig karaktär.
I praktiken har det varit svårt att avgöra vilka transporter som är tillåtna.
Det behövs därför tydliga regler för vilka efterlevnaden kan kontrolleras.
(11) Tidigare har sådana nationella transporter varit tillåtna om det har rört sig om trafik av tillfällig karaktär.
I praktiken har det varit svårt att avgöra vilka transporter som är tillåtna.
Det behövs därför tydliga regler för vilka efterlevnaden kan kontrolleras.
På längre sikt kan restriktionerna för cabotage dock inte längre motiveras.
De måste avskaffas fullständigt, eftersom dessa restriktioner inte är förenliga med principerna för en inre marknad utan gränser där fri rörlighet för varor och tjänster garanteras.
Medlemsstaterna måste vidta alla nödvändiga åtgärder för att se till att reglerna tillämpas enhetligt i hela EU.
Motivering
Den fria rörligheten för tjänster och en gemensam transportpolitik ingick redan i fördragen från 1957.
År 1985 inledde Europaparlamentet ett förfarande mot rådet vid domstolen, eftersom rådet misslyckats med att införa en gemensam transportpolitik.
Domstolens dom ledde till de första initiativen för att öppna marknaden för vägtransporter.
Vi får inte nu vrida klockan tillbaka utan måste i stället satsa på att få en helt avreglerad cabotagemarknad 2012.
Ur miljöhänsyn måste transporterna på väg vara så effektiva som möjligt och antalet tomkörningar begränsas så mycket som möjligt.
Ändringsförslag
4
Skäl 12a (nytt)
(12a) Restriktioner i fråga om antalet cabotagetransporter och den tidsperiod inom vilken de får utföras är en nödvändig men endast tillfällig åtgärd som ska uppmuntra medlemsstaterna att i största möjliga utsträckning harmonisera skatte- och arbetsvillkoren.
De restriktioner som fastställs genom denna förordning är därför tillfälliga och bör upphävas från och med den 1 januari 2014.
Motivering
På den inre marknaden bör restriktionerna för cabotagetransporter endast vara tillfälliga.
Därför måste ett specifikt datum anges för att främja harmonisering av skatte- och arbetsvillkoren.
Ändringsförslag
5
Skäl 12b (nytt)
(12b) Vissa angränsande medlemsstater har sedan lång tid tillbaka starka ekonomiska band.
Sådana medlemsstater bör därför kunna tillåta ökat tillträde till cabotage för transportföretag i de berörda angränsande medlemsstaterna.
Motivering
Medlemsstater som gränsar till varandra och har starka ekonomiska band bör kunna ge ökat tillträde till varandras marknader.
Se även det ändringsförslag som syftar till att införa en ny punkt 6b i artikel 8.
Ändringsförslag
6
Skäl 13a (nytt)
(13a) Det bör kunna undvikas att tredjelandstransporter, det vill säga transporter mellan två medlemsstater som ingendera är den medlemsstat där transportföretaget är etablerat, leder till situationer som är så regelbundna, kontinuerliga och systematiska att de kan snedvrida marknaden på grund av att anställnings- och arbetsvillkor tillämpas som är mindre fördelaktiga än de villkor som gäller i de två medlemsstater som tredjelandstransporten utförs emellan.
Motivering
Det måste undvikas att problem uppstår på grund av att transportföretag regelbundet och systematiskt utför transporter och utnyttjar att de sociala villkor och lönevillkor som gäller i de länder där företagen är etablerade är sämre.
Se även det ändringsförslag som syftar till att införa en ny punkt 7a.
Ändringsförslag
7
Skäl 14
(14) De administrativa formaliteterna bör så långt det är möjligt minskas men utan att de kontrollmöjligheter och påföljder avskaffas som säkerställer att denna förordning tillämpas korrekt och att efterlevnaden kontrolleras effektivt.
Därför bör de befintliga reglerna om indragning av gemenskapstillstånd tydliggöras och stärkas.
Reglerna bör anpassas för att även möjliggöra effektiva påföljder för allvarliga överträdelser eller upprepade mindre överträdelser i en annan medlemsstat än den där transportföretaget är etablerat.
Påföljderna bör vara icke-diskriminerande och stå i proportion till hur allvarliga överträdelserna är.
Det bör vara möjligt att överklaga en påföljd .
(14) De administrativa formaliteterna bör så långt det är möjligt minskas men utan att de kontrollmöjligheter och påföljder avskaffas som säkerställer att denna förordning tillämpas korrekt och att efterlevnaden kontrolleras effektivt.
Därför bör de befintliga reglerna om indragning av gemenskapstillstånd tydliggöras och stärkas.
Reglerna bör anpassas för att även möjliggöra effektiva påföljder för allvarliga överträdelser i en annan medlemsstat än den där transportföretaget är etablerat.
Påföljderna bör vara icke-diskriminerande och stå i proportion till hur allvarliga överträdelserna är.
Det bör vara möjligt att överklaga.
Motivering
Om åtgärder ska vidtas vid upprepade mindre överträdelser utanför etableringsmedlemsstaten måste den medlemsstat där överträdelsen skedde anmäla den till etableringsmedlemsstaten.
Detta skulle leda till att en alltför stor del av den administrativa kapaciteten togs i anspråk.
Ändringsförslag
8
Skäl 15
(15) Medlemsstaterna bör i sina nationella register över transportföretag som bedriver godstransporter på väg registrera alla allvarliga överträdelser och upprepade mindre överträdelser som begåtts av transportföretag och för vilka det utmätts påföljder.
(15) Medlemsstaterna bör i sina nationella register över transportföretag som bedriver godstransporter på väg registrera alla allvarliga överträdelser som begåtts av transportföretag och för vilka det utmätts påföljder.
Motivering
Så länge som överträdelser i medlemsstaterna tolkas och åtgärdas på så olika sätt, och det ännu inte finns några konkreta planer på en snabb förbättring, bör bestämmelser om upprepade mindre överträdelser inte ingå i denna förordning.
Ändringsförslag
9
4.
4.
Motivering
Ändringsförslag
10
5.
Denna förordning skall inte tillämpas på följande typer av transporter och resor utan last i samband med sådana transporter:
Ändringsförslag
11
a) Posttrafik som genomförs inom ramen för samhällsomfattande tjänster.
(Berör inte den svenska versionen.)
Motivering
(Berör inte den svenska versionen.)
Ändringsförslag
12
6) cabotage: nationella transporter i yrkesmässig trafik som utförs på tillfällig bas i en värdmedlemsstat,
Motivering
För att andra tolkningar av begreppet ”transporter som utförs på tillfällig bas” ska undvikas, måste det i definitionen av cabotage hänvisas till bestämmelserna i kapitel III.
Ändringsförslag
13
utgår
Motivering
Kravet på gott anseende är oacceptabelt eftersom det innebär ett omotiverat antagande att en yrkesgrupp kan ha gjort sig skyldig till missbruk i moraliskt hänseende.
Ur strikt juridiskt perspektiv är uttrycket olämpligt som grundval för en påföljd.
Vi önskar ändra förslaget till förordning om gemensamma regler beträffande de villkor som ska uppfyllas av personer som yrkesmässigt bedriver transporter på väg (betänkande av Ticau) på samma sätt.
Ändringsförslag
14
7a) tredjelandstransporter: internationella transporter som utförs av ett transportföretag mellan två värdmedlemsstater som ingendera är den medlemsstat där transportföretaget är etablerat.
Motivering
Det måste undvikas att problem uppstår på grund av att transportföretag regelbundet och systematiskt utför transporter och utnyttjar att de sociala villkor och lönevillkor som gäller i de länder där företagen är etablerade är sämre.
Se även det ändringsförslag som syftar till att införa en ny artikel 7a.
Ändringsförslag
15
Artikel 7a (ny)
Artikel 7a
Tredjelandstransporter och utstationering av arbetstagare
När ett godstransportföretag regelbundet, kontinuerligt och/eller systematiskt utför tredjelandstransporter mellan två medlemsstater, kan en värdmedlemsstat kräva att de arbets- och anställningsvillkor som anges i artikel 9 i denna förordning ska tillämpas.
Motivering
Det måste undvikas att problem uppstår på grund av att transportföretag regelbundet och systematiskt utför transporter och utnyttjar att de sociala villkor och lönevillkor som gäller i de länder där företagen är etablerade är sämre.
Se även det ändringsförslag som syftar till att införa ett nytt led 7a.
Ändringsförslag
16
2.
Tranportföretag enligt punkt 1 skall få genomföra upp till tre cabotagetransporter med samma fordon efter en internationell transport, som gått från en annan medlemsstat eller ett tredjeland till värdmedlemsstaten, så snart det gods som transporteras på den ingående resan har levererats.
Den sista lossningen av last inom ramen för en cabotagetransport som genomförs innan fordonet lämnar värdmedlemsstaten skall äga rum inom sju dagar från det att den sista lossningen av den ingående internationella transporten har ägt rum.
2.
Transportföretag enligt punkt 1 skall få genomföra upp till tre cabotagetransporter med samma fordon efter en internationell transport, som gått från en annan medlemsstat eller ett tredjeland till värdmedlemsstaten, så snart det gods som transporteras på den ingående resan har levererats.
Fordonet behöver inte lossas helt och hållet för att dessa cabotagetransporter ska tillåtas.
Den sista lossningen av last inom ramen för en cabotagetransport som genomförs innan fordonet lämnar värdmedlemsstaten skall äga rum inom sju dagar från det att den sista lossningen av den ingående internationella transporten har ägt rum.
Motivering
Cabotage ska tillåtas redan vid den första lossningen av en internationell transport, även om bara en del av lasten lossas.
På så sätt kan man undvika att fordon inte kan köra med full kapacitet och därmed att resor sker med halvtomma fordon.
Ändringsförslag
17
2a.
Cabotagetransporter kan även genomföras i en medlemsstat som ett fordon måste passera igenom efter lossning i en leveransmedlemsstat under en internationell transport, förutsatt att den kortaste vägen tillbaka går genom denna medlemsstat och att återresan efter lossningen i leveranslandet sker inom sju dagar.
Motivering
Cabotage måste tillåtas i länder som passeras på återresan för att resor utan last ska undvikas.
Ändringsförslag
18
2b.
Restriktionerna i fråga om antalet cabotagetransporter och den tidsperiod inom vilken de får utföras ska gradvis upphävas.
Två år efter denna förordnings ikraftträdande ska antalet cabotagetransporter som anges i punkt 2 ökas till sju.
Den 1 januari 2014 ska alla restriktioner i fråga om antalet cabotagetransporter och den tidsperiod inom vilken de får utföras upphävas.
Motivering
På den inre marknaden bör restriktionerna för cabotagetransporter endast vara tillfälliga.
Därför måste ett specifikt datum anges för att främja harmonisering av skatte- och arbetsvillkoren.
Ändringsförslag
19
Bevismaterialet skall som ett minimum innehålla följande uppgifter avseende varje transport:
Bevismaterialet skall innehålla följande uppgifter avseende varje transport:
Motivering
För att minska onödig byråkrati, måste man undvika att medlemsstaterna begär särskilt bevismaterial.
Ändringsförslag
20
3a.
Medlemsstaterna ska inte kräva några ytterligare specifika dokument eller överlappande dokument för att styrka att villkoren i punkt 3 har uppfyllts.
Medlemsstaterna och kommissionen ska se till att bestämmelserna i andra avtal med tredjeländer följer bestämmelserna i denna förordning.
Motivering
Man måste undvika att varje enskild medlemsstat begär särskilda kontrolldokument.
På medellång sikt är en enhetlig och harmoniserad standardfraktsedel för samtliga transporttyper enda sättet att garantera rättssäkerhet, administrativ förenkling, ökad betydelse för transportkontraktet och därmed öppna och rättsligt bindande kommersiella förbindelser.
Ändringsförslag
21
6a.
Bestämmelserna i denna förordning ska inte hindra en medlemsstat från att tillåta godstransportörer från en eller flera medlemsstater att på dess territorium genomföra ett obegränsat antal eller fler cabotagetransporter än vad som avses i punkt 2 inom en för den sista lossningen obegränsad tidsperiod eller en tidsperiod som överstiger den som avses i punkt 2.
Tillstånd som beviljats innan denna förordning träder i kraft ska fortsätta att gälla.
Medlemsstaterna ska underrätta kommissionen om befintliga tillstånd och om tillstånd som de beviljar efter det att denna förordning har trätt i kraft.
Motivering
En anpassning av föredragandens ändringsförslag 14.
Inte enbart grannländer ska kunna komma överens om mer liberala bestämmelser, utan alla medlemsstater som så önskar.
Med andra ord är det inte enbart grannländer som ska kunna enas om mer liberala cabotagebestämmelser.
Ändringsförslag
22
6b.
Ankommande eller avgående transporter av gods på väg inom ramen för kombinerad transport enligt bestämmelserna i direktiv 92/106/EEG omfattas inte av definitionen för cabotage.
Motivering
Gällande praxis i vissa medlemsstater tyder på en annan trend, men det kan eller får inte vara avsikten.
Ändringsförslag
23
ea) Utstationering av arbetstagare enligt direktiv 96/71/EG 1 .
______________
1 EGT L 18, 21.1.1997. s.
1.
Motivering
I skäl 12 förklaras att direktivet om utstationering av arbetstagare gäller för cabotagetransporter.
Detta måste återspeglas även i artiklarna.
Ändringsförslag
24
1.
Om en allvarlig överträdelse av gemenskapens vägtransportlagstiftning begås eller uppdagas i en medlemsstat, skall de behöriga myndigheterna i den medlemsstat där det transportföretag som gjort sig skyldigt till överträdelsen är etablerat utfärda en varning och får, utom annat, utmäta följande administrativa påföljder:
Motivering
Så länge som överträdelser i medlemsstaterna tolkas och åtgärdas på så olika sätt, och det ännu inte finns några konkreta planer på en snabb förbättring, bör bestämmelser om upprepade mindre överträdelser inte ingå i denna förordning.
Ändringsförslag
25
ba) Böter.
Motivering
För att påföljderna också ska ha någon effekt bör även böter uttryckligen införas i förordningen som en möjlig påföljd.
Ändringsförslag
26
Påföljderna skall bestämmas med hänsyn till hur allvarlig överträdelsen är och hur många upprepade mindre överträdelser som innehavaren av gemenskapstillståndet gjort sig skyldig till och hur många bestyrkta kopior av tillståndet han innehar för sin internationella trafik.
Påföljderna skall när ett slutligt beslut har fattats och alla rättsliga möjligheter till ny behandling som står till förfogande för transportföretaget har uttömts bestämmas med hänsyn till hur allvarlig överträdelsen är som innehavaren av gemenskapstillståndet gjort sig skyldig till och hur många bestyrkta kopior av tillståndet han innehar för sin internationella trafik.
Motivering
Så länge som överträdelser i medlemsstaterna tolkas och åtgärdas på så olika sätt, och det ännu inte finns några konkreta planer på en snabb förbättring, bör bestämmelser om upprepade mindre överträdelser inte ingå i denna förordning.
Ändringsförslag
27
2.
2.
Motivering
Så länge som överträdelser i medlemsstaterna tolkas och åtgärdas på så olika sätt, och det ännu inte finns några konkreta planer på en snabb förbättring, bör bestämmelser om upprepade mindre överträdelser inte ingå i denna förordning.
Ändringsförslag
28
ea) Böter.
Motivering
För att påföljderna också ska ha någon effekt bör även böter uttryckligen införas i förordningen som en möjlig påföljd.
Ändringsförslag
29
3.
De skall så snart som möjligt och senast inom tre månader efter det att de fick kännedom om överträdelsen meddela de behöriga myndigheterna i den medlemsstat där överträdelserna uppdagades vilken av påföljderna enligt punkt 1 och 2 i denna artikel som har utmätts.
3.
De skall så snart som möjligt och senast inom tre månader efter det att de fick kännedom om överträdelsen meddela de behöriga myndigheterna i den medlemsstat där överträdelserna uppdagades vilken av påföljderna enligt punkt 1 och 2 i denna artikel som har utmätts.
Motivering
När det är fråga om en allvarlig överträdelse ska en påföljd utmätas.
Ändringsförslag
30
3a.
I beslutet om tillfällig återkallelse av ett dokument (gemenskapstillstånd, förartillstånd, bestyrkt kopia) ska följande anges:
a) Tidsperioden för den tillfälliga återkallelsen.
b) Villkoren för att upphäva den tillfälliga återkallelsen.
c) De fall då gemenskapstillståndet permanent ska återkallas på grund av att de villkor som fastställs i led b inte har uppfyllts inom den tidsperiod som fastställs i led a.
Motivering
Villkoren för att upphäva den tillfälliga återkallelsen måste klart framgå.
Ändringsförslag
31
1.
Om de behöriga myndigheterna i en medlemsstat får kännedom om att ett icke‑hemmahörande transportföretag har begått en allvarlig överträdelse eller upprepade mindre överträdelser mot denna förordning eller mot gemenskapens vägtransportlagstiftning skall den medlemsstat inom vars territorium överträdelsen uppdagades till de behöriga myndigheterna i etableringsmedlemsstaten översända följande information, så snart som möjligt och senast inom en månad efter det att de får kännedom om överträdelsen :
1.
Om de behöriga myndigheterna i en medlemsstat får kännedom om att ett icke hemmahörande transportföretag har begått en allvarlig överträdelse eller upprepade mindre överträdelser mot denna förordning eller mot gemenskapens vägtransportlagstiftning skall den medlemsstat inom vars territorium överträdelsen uppdagades till de behöriga myndigheterna i etableringsmedlemsstaten översända följande information, så snart som möjligt och senast inom en månad från den dag då det slutliga beslutet fattades, efter det att alla rättsliga möjligheter till ny behandling som står till förfogande för det transportföretag som ålagts påföljderna har uttömts :
Motivering
De uppgifter som ska införas i de nationella elektroniska registren måste inhämtas efter det att de slutliga besluten har fattats.
Ändringsförslag
32
1.
Om de behöriga myndigheterna i en medlemsstat får kännedom om att ett icke‑hemmahörande transportföretag har begått en allvarlig överträdelse eller upprepade mindre överträdelser mot denna förordning eller mot gemenskapens vägtransportlagstiftning skall den medlemsstat inom vars territorium överträdelsen uppdagades till de behöriga myndigheterna i etableringsmedlemsstaten översända följande information, så snart som möjligt och senast inom en månad efter det att de får kännedom om överträdelsen:
1.
Om de behöriga myndigheterna i en medlemsstat får kännedom om att ett icke‑hemmahörande transportföretag har begått en allvarlig överträdelse mot denna förordning eller mot gemenskapens vägtransportlagstiftning skall den medlemsstat inom vars territorium överträdelsen uppdagades till de behöriga myndigheterna i etableringsmedlemsstaten översända följande information, så snart som möjligt och senast inom en månad efter det att de får kännedom om överträdelsen:
Motivering
Så länge som överträdelser i medlemsstaterna tolkas och åtgärdas på så olika sätt, och det ännu inte finns några konkreta planer på en snabb förbättring, bör bestämmelser om upprepade mindre överträdelser inte ingå i denna förordning.
Ändringsförslag
33
2.
De skall ålägga sådana påföljder på icke diskriminerande grund.
Påföljderna får exempelvis bestå av en varning eller, i händelse av en allvarlig överträdelse eller upprepade mindre överträdelser , en tidsbegränsad avstängning från cabotage inom den medlemsstats territorium där överträdelsen begicks.
2.
Utan att det påverkar ett eventuellt åtalsförfarande skall de behöriga myndigheterna i värdmedlemsstaten ha rätt att ålägga påföljder mot ett icke hemmahörande transportföretag som har gjort sig skyldigt till överträdelse av denna förordning eller av nationell vägtransportlagstiftning eller av gemenskapens vägtransportlagstiftning i dess territorium vid utförande av cabotage.
De skall ålägga sådana påföljder på icke diskriminerande grund .
Påföljderna får exempelvis bestå av en varning eller, i händelse av en allvarlig överträdelse, en tidsbegränsad avstängning från cabotage inom den medlemsstats territorium där överträdelsen begicks.
Motivering
Så länge som överträdelser i medlemsstaterna tolkas och åtgärdas på så olika sätt, och det ännu inte finns några konkreta planer på en snabb förbättring, bör bestämmelser om upprepade mindre överträdelser inte ingå i denna förordning.
Ändringsförslag
34
Artikel 13
Varje medlemsstat skall se till att uppgifter om allvarliga överträdelser eller upprepade mindre överträdelser av gemenskapens lagstiftning om vägtransport som begåtts av transportföretag som är etablerade på dess territorium och för vilka det i någon medlemsstat utmätts en påföljd registreras i det nationella registret över transportföretag enligt artikel 15 i förordning (EG) nr xx/xxxx [om gemensamma regler beträffande de villkor som skall uppfyllas av personer som yrkesmässigt bedriver transporter på väg] tillsammans med en uppgift om vilken påföljden blev.
Uppgifter om tillfällig eller permanent återkallelse av gemenskapstillstånd skall ligga kvar i databasen under minst två år.
Varje medlemsstat skall se till att uppgifter om allvarliga överträdelser av gemenskapens lagstiftning om vägtransport som begåtts av transportföretag som är etablerade på dess territorium och för vilka det i någon medlemsstat utmätts en påföljd , när ett slutligt beslut har fattats och alla rättsliga möjligheter till ny behandling som står till förfogande för transportföretaget har uttömts, registreras i det nationella registret över transportföretag enligt artikel 15 i förordning (EG) nr xx/xxxx [om gemensamma regler beträffande de villkor som skall uppfyllas av personer som yrkesmässigt bedriver transporter på väg] tillsammans med en uppgift om vilken påföljden blev.
Uppgifter om tillfällig eller permanent återkallelse av gemenskapstillstånd skall ligga kvar i databasen under minst två år.
Motivering
Endast uppgifter om allvarliga överträdelser av gemenskapens lagstiftning bör registreras i de nationella registren.
Ändringsförslag
35
Artikel 18, stycke 2
Den skall tillämpas från och med den [tillämpningsdatum] .
Den skall tillämpas från och med den 1 januari 2009 .
MOTIVERING
Allmän ram
Tillträdet till den internationella marknaden för godstransporter på väg och för cabotage styrs för närvarande av förordningarna (EG) nr 881/92 och (EG) nr 3118/93 samt direktiv 2006/94/EG från 1962.
På den inre marknaden har den internationella transporten mellan medlemsstater helt och hållet avreglerats, medan det för cabotage fortfarande finns ett antal restriktioner.
Bland annat föreslår kommissionen följande:
· Att villkoren för cabotage ska specificeras; cabotage bör enligt definitionen nationella transporter i yrkesmässig trafik som utförs på tillfällig bas i en värdmedlemsstat begränsas till högst tre cabotagetransporter som ska äga rum inom sju dagar.
· Att förenklade och standardiserade modeller ska användas för gemenskapstillstånd, kopior av detta och förartillstånd för att underlätta kontroller.
· Att bestämmelserna om påföljder för överträdelser som begås i andra medlemsstater än den där transportföretaget är etablerat ska skärpas.
Föredragandens ståndpunkt
Föredraganden ser positivt på kommissionens förslag som är tänkt att förenkla och förtydliga de bestämmelser som gäller för godstransporter på väg.
En definition av cabotage medför en mer enhetlig tillämpning av denna princip.
Föredraganden anser dock att kommissionens förslag bör ändras på vissa punkter.
1.
I fråga om cabotage bör den föreslagna regleringen gälla tillfälligt.
På en marknad med mer harmoniserade skatte- och arbetsvillkor skulle det inte längre behövas några restriktioner för cabotage.
Med tanke på detta bör angränsande medlemsstater även i fortsättningen kunna ingå avtal om att ge ökat tillträde till varandras marknader.
Dessutom bör cabotage vara tillåtet i en medlemsstat som ett transportföretag passerar igenom på återresan efter lossning i ett tredje land och efter lossning av en del av den totala lasten.
Man måste se till att det inte finns olika tolkningar i medlemsstaterna av definitionen av cabotage och av de bestämmelser som gäller för det bevismaterial som det transportföretag som utför cabotaget är skyldigt att uppvisa.
2.
Det är viktigt att specificera villkoren för tredjelandstransporter , dvs. transporter mellan två medlemsstater som ingendera är den medlemsstat där transportföretaget är etablerat.
Om sådana transporter utförs regelbundet, kontinuerligt och/eller systematiskt riskerar de att snedvrida den nationella marknaden i en värdmedlemsstat.
En värdmedlemsstat måste således kunna kräva att samma arbets- och anställningsvillkor ska gälla som för dess nationella transportföretag.
3.
I fråga om överträdelser som begås i andra medlemsstater är det viktigt att skilja mellan allvarliga och mindre överträdelser.
För mindre överträdelser vore det tillräckligt att den medlemsstat där överträdelsen har konstaterats meddelar detta till den medlemsstat där transportföretaget är etablerat, vilken i sin tur ska besluta huruvida en påföljd ska utmätas.
För allvarliga överträdelser måste etableringsmedlemsstaten besluta vilken påföljd som ska utmätas och meddela sitt beslut till den medlemsstat där överträdelsen konstaterades.
Vidare måste det anges att en rad mindre överträdelser enligt reglerna om rätten att yrkesmässigt bedriva transporter på väg kan utgöra en allvarlig överträdelse.
Däremot behöver mindre överträdelser inte registreras i det nationella registret förrän de på grund av sitt antal och det antal gånger som de upprepas utgör en allvarlig överträdelse.
BILAGA 1: SKRIVELSE FRÅN UTSKOTTET FÖR RÄTTSLIGA FRÅGOR
COMMITTEE ON LEGAL AFFAIRS
CHAIRMAN
Ref.: D(2008)2164
Mr Paolo COSTA
Chairman of the Committee on Transport and Tourism
LOW T06031
Strasbourg
Subject : Proposal for a recast : Regulation of the European Parliament and of the Council on common rules for access to the international road haulage market ( COM(2007) 265 final -23.5.2007 - 2007/0099 (COD ).
Dear Sir,
The Committee on Legal Affairs, which I am honoured to chair, has examined the proposal referred to above, pursuant to Rule 80a on Recasting, as introduced into the Parliament's Rules of Procedure by its Decision of 10 May 2007.
Paragraph 3 of that Rule reads as follows:
"If the committee responsible for legal affairs considers that the proposal does not entail any substantive changes other than those identified as such in the proposal, it shall inform the committee responsible.
In such a case, over and above the conditions laid down in Rules 150 and 151, amendments shall be admissible within the committee responsible only if they concern those parts of the proposal which contain changes.
However, amendments to the parts which have remained unchanged may be admitted by way of exception and on a case-by-case basis by the chairman of the above committee if he considers that this is necessary for pressing reasons relating to the internal logic of the text or because the amendments are inextricably linked to other admissible amendments.
Such reasons must be stated in a written justification to the amendments".
Following the opinion of the Legal Service, whose representatives participated in the meetings of the Consultative Working Party examining the recast proposal, and in keeping with the recommendations of the draftsperson, the Committee on Legal Affairs considers that the proposal in question does not include any substantive changes other than those identified as such in the proposal and that, as regards the codification of the unchanged provisions of the earlier acts with those changes, the proposal contains a straightforward codification of the existing texts, without any change in their substance.
However, pursuant to Rules 80a(2) and 80(3), the Committee on Legal Affairs considered that the technical adaptations suggested in the opinion of the abovementioned Working Party were necessary in order to ensure that the proposal complied with the codification rules and that they did not involve any substantive change to the proposal.
In conclusion, the Committee on Legal Affairs recommends that your Committee, as the committee responsible, proceed to examine the above proposal in keeping with its suggestions and in accordance with Rule 80a.
Yours faithfully,
Giuseppe GARGANI
BILAGA 2: SKRIVELSE FRÅN DE JURIDISKA AVDELNINGARNAS RÅDGIVANDE GRUPP
Bryssel
YTTRANDE
TILL EUROPAPARLAMENTET
Förslag till Europaparlamentets och rådets förordning om gemensamma regler för tillträde till den internationella marknaden för godstransporter på väg (omarbetning) ( KOM(2007)0265 av den 23 maj 2007 – 2007/0099(COD) )
Vid dessa sammanträden
Gruppen förfogade över alla språkversioner av förslaget och arbetade utifrån den engelska som var textens originalversion. behandlade gruppen förslaget till Europaparlamentets och rådets förordning om omarbetning av rådets förordning (EEG) nr 881/92 av den 26 mars 1992 om tillträde till marknaden för godstransporter på väg inom gemenskapen till eller från en medlemsstats territorium eller genom en eller flera medlemsstaters territorier, rådets förordning (EEG) nr 3118/93 av den 25 oktober 1993 om förutsättningar för transportföretag att utföra inrikes godstransporter på väg i en medlemsstat där de inte är etablerade och Europaparlamentets och rådets direktiv 2006/94/EG av den 12 december 2006 om fastställande av gemensamma regler för vissa godstransporter på väg, och konstaterade enhälligt följande:
1) (Den föreslagna ändringen berör inte den svenska versionen.)
2) I skäl 6 [skäl 5 i den svenska versionen] ska orden ”mellan medlemsstaterna” strykas.
– i artikel 9.1 d: orden ”arbets-” (redan mellan markörer),
– i artikel l1.2 d: ordet ”permanent” (redan mellan markörer),
5) (Den föreslagna ändringen berör inte den svenska versionen.)
6) (Den föreslagna ändringen berör inte den svenska versionen.)
Vid behandlingen kunde den rådgivande gruppen därmed enhälligt konstatera att förslaget inte innehåller några väsentliga ändringar utöver dem som anges i förslaget eller i detta yttrande.
Gruppen konstaterade vidare att förslaget i fråga om kodifieringen av de bibehållna bestämmelserna med de väsentliga ändringarna endast gäller en kodifiering som inte ändrar sakinnehållet i de rättsakter som berörs.
ÄRENDETS GÅNG
Titel
Gemensamma regler för tillträde till den internationella marknaden för godstransporter på väg (omarbetning)
Referensnummer
KOM(2007)0265 – C6-0146/2007 – 2007/0099(COD)
Framläggande för parlamentet
23.5.2007
Ansvarigt utskott
Tillkännagivande i kammaren
TRAN
24.9.2007
Rådgivande utskott
Tillkännagivande i kammaren
JURI
24.9.2007
Inget yttrande avges
Beslut
JURI
18.9.2007
Föredragande
Utnämning
Mathieu Grosch
13.7.2007
Behandling i utskott
9.10.2007
20.11.2007
21.1.2008
Antagande
22.1.2008
Slutomröstning: resultat
+:
–:
0:
32
12
2
Slutomröstning: närvarande ledamöter
Gabriele Albertini, Inés Ayala Sender, Etelka Barsi-Pataky, Paolo Costa, Michael Cramer, Luis de Grandes Pascual, Christine De Veyrac, Petr Duchoň, Saïd El Khadraoui, Robert Evans, Emanuel Jardim Fernandes, Francesco Ferrari, Mathieu Grosch, Georg Jarzembowski, Stanisław Jałowiecki, Timothy Kirkhope, Dieter-Lebrecht Koch, Jaromír Kohlíček, Rodi Kratsa-Tsagaropoulou, Sepp Kusstatscher, Jörg Leichtfried, Bogusław Liberadzki, Eva Lichtenberger, Marian-Jean Marinescu, Erik Meijer, Robert Navarro, Seán Ó Neachtain, Willi Piecyk, Reinhard Rack, Luca Romagnoli, Gilles Savary, Brian Simpson, Renate Sommer, Dirk Sterckx, Ulrich Stockmann, Yannick Vaugrenard, Lars Wohlin, Roberts Zīle
Slutomröstning: närvarande suppleanter
Johannes Blokland, Luigi Cocilovo, Jeanine Hennis-Plasschaert, Lily Jacobs, Anne E. Jensen, Leopold Józef Rutowicz, Ari Vatanen, Corien Wortmann-Kool
A6-0112/2008
BETÄNKANDE
om ansvarsfrihet för genomförandet av budgeten för Europeiska byrån för återuppbyggnad för budgetåret 2006
(C6‑0373/2007 – 2007/2048(DEC))
Budgetkontrollutskottet
Föredragande:
Hans-Peter Martin
PE 396.691v02-00
INNEHÅLL
1.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT.......................................................3
3.
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.............................................7
YTTRANDE från utskottet för utrikesfrågor .................................................15
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................17
1.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
om ansvarsfrihet för genomförandet av budgeten för Europeiska byrån för återuppbyggnad för budgetåret 2006
( C6‑0373/2007 – 2007/2048(DEC) )
Europaparlamentet fattar detta beslut
– med beaktande av den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad för budgetåret 2006
EUT C 261, 31.10.2007, s.
13. ,
– med beaktande av revisionsrättens rapport om den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad för budgetåret 2006, samt byråns svar
EUT C 309, 19.12.2007, s.
40. ,
– med beaktande av rådets rekommendation av den 12 februari 2008 (5843/2008 – C6‑0084/2008 ),
– med beaktande av EG-fördraget, särskilt artikel 276,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1.
Förordningen senast ändrad genom förordning (EG) nr 1525/2007 (EUT L 343, 27.12.2007, s.
9). , särskilt artikel 185,
– med beaktande av rådets förordning (EG) nr 2667/2000 av den 5 december 2000 om Europeiska byrån för återuppbyggnad
EUT L 136, 30.4.2004, s.
7.
Förordningen senast ändrad genom förordning (EG) nr 1756/2006 (EUT L 332, 30.11.2006, s.
18). , särskilt artikel 8,
– med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002
EGT L 357, 31.12.2002, s.
72. , särskilt artikel 94,
– med beaktande av artikel 71 och bilaga V i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för utrikesfrågor ( A6‑0112/2008 ).
2.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
om avslutande av räkenskaperna för Europeiska byrån för återuppbyggnad för budgetåret 2006
( C6‑0373/2007 – 2007/2048(DEC) )
Europaparlamentet fattar detta beslut
– med beaktande av den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad för budgetåret 2006
EUT C 261, 31.10.2007, s.
13. ,
– med beaktande av revisionsrättens rapport om den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad för budgetåret 2006, samt byråns svar
EUT C 309, 19.12.2007, s.
40. ,
– med beaktande av rådets rekommendation av den 12 februari 2008 (5843/2008 – C6‑0084/2008 ),
– med beaktande av EG-fördraget, särskilt artikel 276,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1.
Förordningen senast ändrad genom förordning (EG) nr 1525/2007 (EUT L 343, 27.12.2007, s.
9). , särskilt artikel 185,
– med beaktande av rådets förordning (EG) nr 2667/2000 av den 5 december 2000 om Europeiska byrån för återuppbyggnad
EUT L 136, 30.4.2004, s.
7.
Förordningen senast ändrad genom förordning (EG) nr 1756/2006 (EUT L 332, 30.11.2006, s.
18). , särskilt artikel 8,
– med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002
EGT L 357, 31.12.2002, s.
72. , särskilt artikel 94,
– med beaktande av artikel 71 och bilaga V i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för utrikesfrågor ( A6‑0112/2008 ).
3.
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska byrån för återuppbyggnad för budgetåret 2006
( C6‑0373/2007 – 2007/2048(DEC) )
Europaparlamentet utfärdar denna resolution
– med beaktande av den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad för budgetåret 2006
EUT C 261, 31.10.2007, s.
13. ,
– med beaktande av revisionsrättens rapport om den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad för budgetåret 2006, samt byråns svar
EUT C 309, 19.12.2007, s.
40. ,
– med beaktande av rådets rekommendation av den 12 februari 2008 (5843/2008 – C6‑0084/2008 ),
– med beaktande av EG-fördraget, särskilt artikel 276,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1.
Förordningen senast ändrad genom förordning (EG) nr 1525/2007 (EUT L 343, 27.12.2007, s.
9). , särskilt artikel 185,
– med beaktande av rådets förordning (EG) nr 2667/2000 av den 5 december 2000 om Europeiska byrån för återuppbyggnad
EUT L 136, 30.4.2004, s.
7.
Förordningen senast ändrad genom förordning (EG) nr 1756/2006 (EUT L 332, 30.11.2007, s.
18). , särskilt artikel 8,
– med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002
EGT L 357, 31.12.2002, s.
72. , särskilt artikel 94,
– med beaktande av artikel 71 och bilaga V i arbetsordningen,
A. Revisionsrätten har förklarat att den har uppnått en rimlig säkerhet om att räkenskaperna för budgetåret är tillförlitliga och att de underliggande transaktionerna är lagliga och korrekta.
B. Den 24 april 2007 beviljade Europaparlamentet direktören för Europeiska byrån för återuppbyggnad ansvarsfrihet för genomförandet av detta organs budget för budgetåret 2005
Antagna texter, P6_TA(2007)0136 . , och i sin resolution som åtföljde beslutet om ansvarsfrihet framförde parlamentet bland annat följande synpunkter:
· Europaparlamentet noterade att revisionsrätten i sin rapport för 2004 hade upptäckt, i samband med en genomgång av de verksamheter som överlåtits på UNMIK, att byrån inte utövade vederbörlig finansiell kontroll vid betalningar och att den hade stora svårigheter när den skulle avsluta verksamheterna, främst på grund av att bokföringen för projekten var bristfällig och att utgifterna inte var tillräckligt styrkta.
Allmänna punkter som rör övergripande frågor för de decentraliserade EU-organen och som därmed också är av betydelse för varje enskilt organs ansvarsfrihetsförfarande
Principiella överväganden
Europaparlamentet begär att varje organ ska styras av ett årligt prestationsavtal som formuleras av organet och det ansvariga generaldirektoratet och som ska innehålla de huvudsakliga målsättningarna för det kommande året med en finansieringsram och klara indikatorer för att mäta prestationerna.
Kommissionen uppmanas därför att hitta en snabb lösning för att öka effektiviteten genom att sammanföra de administrativa funktionerna för flera organ så att denna kritiska massa kan uppnås (med beaktande av de nödvändiga ändringarna av de grundförordningar som styr organen och deras budgetmässiga oberoende) eller att omgående utarbeta särskilda regler för organen (i synnerhet genomförandebestämmelser) som gör att de kan uppfylla reglerna helt och hållet.
Europaparlamentet påminner om sitt beslut om ansvarsfrihet för budgetåret 2005 där kommissionen uppmanades att vart femte år genomföra en studie av det mervärde som varje befintligt organ tillför.
Parlamentet begär att kommissionen ska lägga fram åtminstone fem sådana utvärderingar före beslutet om ansvarsfrihet för budgetåret 2007, och då börja med de äldsta organen.
Europaparlamentets resolution innehållande iakttagelser som åtföljer beslutet om ansvarsfrihet för direktören för Europeiska byrån för återuppbyggnad med avseende på genomförandet av byråns budget för budgetåret 2003 (EUT L 196, 27.7.2005, s.
61). där organens direktörer uppmanas att hädanefter låta deras verksamhetsrapporter, som läggs fram tillsammans med ekonomiska och administrativa uppgifter, åtföljas av en revisionsförklaring om transaktionernas laglighet och korrekthet, liknande de förklaringar som undertecknas av kommissionens generaldirektörer.
– en årsrapport, som riktas till en allmän läsekrets, om organets verksamhet, arbete och resultat,
– en ekonomisk årsredovisning och en rapport om genomförandet av budgeten,
– en verksamhetsrapport liknande den som kommissionens generaldirektörer lämnar,
– en revisionsförklaring som undertecknats av organets direktör, med reservationer och iakttagelser som denne anser att den ansvarsfrihetsbeviljande myndigheten lämpligen bör uppmärksamma.
Allmänna iakttagelser från revisionsrätten
EUT C 273, 15.11.2007, s.
1. ) att kommissionens utbetalningar av bidrag från gemenskapsbudgeten inte bygger på tillräckligt motiverade uppskattningar av byråernas behov av likvida medel.
Europaparlamentet noterar att i slutet av 2006 hade 14 byråer ännu inte infört redovisningssystemet ABAC (fotnot till punkt 10.31 i årsrapporten).
Internrevision
22.
23.
Europaparlamentet uppmärksammar följande reservation i internrevisors verksamhetsrapport för 2006:
På grund av personalbrist är kommissionens interrevisor inte i stånd att ordentligt uppfylla den funktion som internrevisor för gemenskapens decentraliserade organ som denne ges i artikel 185 i budgetförordningen.
26.
När det gäller den interna revisionskapaciteten, särskilt i förhållande till mindre organ, noterar Europaparlamentet det förslag som internrevisorn gjorde inför parlamentets ansvariga utskott den 14 september 2006 om att mindre organ ska tillåtas att köpa in interrevisionstjänster från den privata sektorn.
Utvärdering av organ
Rådsdokument DS 605/1/07 Rev1. som förhandlades fram vid medlingen inför Ekofinrådets budgetmöte den 13 juli 2007 där man efterlyser en förteckning på organ som kommissionen avser att utvärdera ii) en förteckning på de organ som redan utvärderats, tillsammans med en sammanfattning av resultaten.
Disciplinära förfaranden
Förslag till interinstitutionellt avtal
I den sammanfattande rapporten om kommissionens förvaltning 2006 (punkt 3.1, KOM(2007)0274 ) sägs att förhandlingarna sedermera avbröts, men att diskussioner om innehållet återupptogs i rådet i slutet av 2006.
Självfinansierade organ
Kontoret för harmonisering inom den inre marknaden har likvida medel på 281 miljoner EUR.
Gemenskapens växtsortsmyndighet har likvida medel på 18 miljoner EUR
Källa: Revisionsrättens särskilda rapport. .
Specifika punkter
Europaparlamentet konstaterar emellertid från byråns räkenskaper att de anslag som överfördes till 2007 uppgick till sammanlagt 678 miljoner EUR.
45.
Europaparlamentet uppmanar kommissionen att informera parlamentets behöriga utskott hur återstoden av outnyttjade anslag vid utgången av byråns mandat skall hanteras.
Europaparlamentet konstaterar att internrevisionsenheten i slutet av 2004 genomförde en granskning av effektiviteten och ändamålsenligheten vid byråns fem arbetsorter och att en serie åtgärder vidtogs under 2006 av byråns ledning för att ta itu med de frågor som internrevisionsenheten tagit upp.
48.
YTTRANDE från utskottet för utrikesfrågor
till budgetkontrollutskottet
över ansvarsfriheten för genomförandet av budgeten för Europeiska byrån för återuppbyggnad för budgetåret 2006
( C6-0373/2007 – 2007/2048(DEC) )
Föredragande: Jelko Kacin
FÖRSLAG
I detta sammanhang upprepar Europaparlamentet sin begäran om att bli regelbundet informerat av kommissionen om överföringen av verksamheten från byrån till delegationerna.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
25.2.2008
Slutomröstning: resultat
+:
–:
0:
27
Slutomröstning: närvarande ledamöter
Angelika Beer, Bastiaan Belder, Colm Burke, Véronique De Keyser, Giorgos Dimitrakopoulos, Michael Gahler, Alfred Gomolka, Klaus Hänsch, Jana Hybášková, Anna Ibrisagic, Jelko Kacin, Metin Kazak, Maria Eleni Koppa, Helmut Kuhne, Vytautas Landsbergis, Johannes Lebech, Francisco José Millán Mon, Philippe Morillon, Annemie Neyts-Uyttebroeck, Baroness Nicholson of Winterbourne, Ioan Mircea Paşcu, Alojz Peterle, Samuli Pohjamo, Libor Rouček, Jacek Saryusz-Wolski, Ari Vatanen
Slutomröstning: närvarande suppleanter
Laima Liucija Andrikienė, Árpád Duka-Zólyomi, Marie Anne Isler Béguin, Inger Segelström
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
25.3.2008
Slutomröstning: resultat
+:
–:
0:
33
4
1
Slutomröstning: närvarande ledamöter
Jean-Pierre Audy, Herbert Bösch, Costas Botopoulos, Mogens Camre, Paulo Casaca, Jorgo Chatzimarkakis, Antonio De Blasio, Esther De Lange, Petr Duchoň, James Elles, Szabolcs Fazakas, Markus Ferber, Christofer Fjellner, Lutz Goepel, Ingeborg Gräßle, Dan Jørgensen, Rodi Kratsa-Tsagaropoulou, Bogusław Liberadzki, Nils Lundgren, Marusya Ivanova Lyubcheva, Hans-Peter Martin, Ashley Mote, Jan Mulder, Bill Newton Dunn, Borut Pahor, Bart Staes, Alexander Stubb, Søren Bo Søndergaard, Jeffrey Titford, Paul van Buitenen, Kyösti Virrankoski
Slutomröstning: närvarande suppleanter
Valdis Dombrovskis, Cătălin-Ioan Nechifor, Dumitru Oprea, Pierre Pribetich, Esko Seppänen, Margarita Starkevičiūtė, Gabriele Stauner, Ralf Walter
A6-0117/2008
BETÄNKANDE
om ansvarsfrihet för genomförandet av budgeten för Europeiska centrumet för förebyggande och kontroll av sjukdomar för budgetåret 2006
(C6‑0386/2007 – 2007/2060(DEC))
Budgetkontrollutskottet
Föredragande:
Hans-Peter Martin
PE 396.703v03-00
INNEHÅLL
1.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT.......................................................3
2.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT.......................................................5
3.
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.............................................7
YTTRANDE från utskottet för miljö, folkhälsa och livsmedelssäkerhets 15
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................17
1.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
om ansvarsfrihet för genomförandet av budgeten för Europeiska centrumet för förebyggande och kontroll av sjukdomar för budgetåret 2006
( C6‑0386/2007 – 2007/2060(DEC) )
Europaparlamentet fattar detta beslut
– med beaktande av den slutliga årsredovisningen för Europeiska centrumet för förebyggande och kontroll av sjukdomar för budgetåret 2006
EUT C 261, 31.10.2007, s.
49. ,
– med beaktande av revisionsrättens rapport om den slutliga årsredovisningen för Europeiska centrumet för förebyggande och kontroll av sjukdomar för budgetåret 2006, samt centrumets svar
EUT C 309, 19.12.2007, s.
99. ,
– med beaktande av rådets rekommendation av den 12 februari 2008 (5843/2008 – C6‑0084/2008 ),
– med beaktande av EG-fördraget, särskilt artikel 276,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1.
Förordningen senast ändrad genom förordning (EG) nr 1525/2007 (EUT L 343, 27.12.2007, s.
9). , särskilt artikel 185,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 851/2004 av den 21 april 2004 om inrättande av ett europeiskt centrum för förebyggande och kontroll av sjukdomar
EUT L 142, 30.4.2004, s.
1. , särskilt artikel 23,
– med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002
EGT L 357, 31.12.2002, s.
72. , särskilt artikel 94,
– med beaktande av artikel 71 och bilaga V i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A6‑0117/2008 ).
2.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
om avslutande av räkenskaperna för Europeiska centrumet för förebyggande och kontroll av sjukdomar för budgetåret 2006
( C6‑0386/2007 – 2007/2060(DEC) )
Europaparlamentet fattar detta beslut
– med beaktande av rådets rekommendation av den 12 februari 2008 (5843/2008 – C6‑0084/2008 ),
– med beaktande av EG-fördraget, särskilt artikel 276,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1.
Förordningen senast ändrad genom förordning (EG) nr 1525/2007 (EUT L 343, 27.12.2007, s.
9). , särskilt artikel 185,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 851/2004 av den 21 april 2004 om inrättande av ett europeiskt centrum för förebyggande och kontroll av sjukdomar
EUT L 142, 30.4.2004, s.
1. , särskilt artikel 23,
– med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002
EGT L 357, 31.12.2002, s.
72. , särskilt artikel 94,
– med beaktande av artikel 71 och bilaga V i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A6‑0117/2008 ).
3.
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska centrumet för förebyggande och kontroll av sjukdomar för budgetåret 2006
( C6‑0386/2007 – 2007/2060(DEC) )
Europaparlamentet utfärdar denna resolution
– med beaktande av den slutliga årsredovisningen för Europeiska centrumet för förebyggande och kontroll av sjukdomar för budgetåret 2006
EUT C 261, 31.10.2007, s.
49. ,
– med beaktande av revisionsrättens rapport om den slutliga årsredovisningen för Europeiska centrumet för förebyggande och kontroll av sjukdomar för budgetåret 2006, samt centrumets svar
EUT C 309, 19.12.2007, s.
99. ,
– med beaktande av rådets rekommendation av den 12 februari 2008 (5843/2008 – C6‑0084/2008 ),
– med beaktande av EG-fördraget, särskilt artikel 276,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1.
9). , särskilt artikel 185,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 851/2004 av den 21 april 2004 om inrättande av ett europeiskt centrum för förebyggande och kontroll av sjukdomar
EUT L 142, 30.4.2004, s.
1. , särskilt artikel 23,
– med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002
EGT L 357, 31.12.2002, s.
72. , särskilt artikel 94,
– med beaktande av artikel 71 och bilaga V i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A6‑0117/2008 ), och av följande skäl:
A. Revisionsrätten har förklarat att den har uppnått en rimlig säkerhet om att räkenskaperna för budgetåret 2006 är tillförlitliga och att de underliggande transaktionerna är lagliga och korrekta.
B. Den 24 april 2007 beviljade Europaparlamentet direktören för Europeiska centrumet för förebyggande och kontroll av sjukdomar ansvarsfrihet för genomförandet av detta organs budget för budgetåret 2005
Antagna texter, P6_TA(2007)0126 . , och i sin resolution som åtföljde beslutet om ansvarsfrihet framförde parlamentet bland annat följande synpunkter:
· Europaparlamentet konstaterade att budgetgenomförandet för 2005 kännetecknades av en låg åtagandegrad (84 procent) och en hög överföringsgrad som generellt sett uppgår till 35 procent och i fråga om driftskostnader till nära 90 procent, men att detta delvis berodde på de inneboende problemen under centrumets inledningsperiod.
· Parlamentet beklagade att det för centrumets kostnader 2005 inte gjordes några budgetåtaganden innan rättsliga åtaganden ingicks och att under samma period verkställdes alla centrumets betalningar av räkenskapsföraren utan betalningsorder från utanordnaren.
· Europaparlamentet noterade att i strid med fastställda bestämmelser i centrums budgetförordning hade det inte tillämpats dubbel bokföring under år 2005, vilket medför risker för fel.
Allmänna punkter som rör övergripande frågor för de decentraliserade EU-organen och som därmed också är av betydelse för varje enskilt organs ansvarsfrihetsförfarande
Europaparlamentet noterar att antalet organ som är föremål för ansvarsfrihetsförfarandet från parlamentets sida har utvecklats enligt följande: Budgetåret 2000: 8, 2001: 10, 2002: 11, 2003: 14, 2004: 14, 2005: 16, 2006: 20 tillsynsmyndigheter och 2 genomförandeorgan (förutom 2 organ som visserligen granskas av revisionsrätten men som blir föremål för ett internt ansvarsfrihetsförfarande).
Principiella överväganden
Europaparlamentet begär att varje organ ska styras av ett årligt prestationsavtal som formuleras av organet och det ansvariga generaldirektoratet och som ska innehålla de huvudsakliga målsättningarna för det kommande året med en finansieringsram och klara indikatorer för att mäta prestationerna.
Europaparlamentet påminner om sitt beslut om ansvarsfrihet för budgetåret 2005 där kommissionen uppmanades att vart femte år genomföra en studie av det mervärde som varje befintligt organ tillför.
Parlamentet begär att kommissionen ska lägga fram åtminstone fem sådana utvärderingar före beslutet om ansvarsfrihet för budgetåret 2007, och då börja med de äldsta organen.
– en årsrapport, som riktas till en allmän läsekrets, om organets verksamhet, arbete och resultat,
– en ekonomisk årsredovisning och en rapport om genomförandet av budgeten,
– en verksamhetsrapport liknande den som kommissionens generaldirektörer lämnar,
– en revisionsförklaring som undertecknats av organets direktör, med reservationer och iakttagelser som denne anser att den ansvarsfrihetsbeviljande myndigheten lämpligen bör uppmärksamma.
Allmänna iakttagelser från revisionsrätten
EUT C 273, 15.11.2007, s.
Europaparlamentet noterar att i slutet av 2006 hade 14 byråer ännu inte infört redovisningssystemet ABAC (fotnot till punkt 10.31 i årsrapporten).
Internrevision
21.
22.
Europaparlamentet uppmärksammar följande reservation i internrevisors verksamhetsrapport för 2006:
På grund av personalbrist är kommissionens interrevisor inte i stånd att ordentligt uppfylla den funktion som internrevisor för gemenskapens decentraliserade organ som denne ges i artikel 185 i budgetförordningen.
25.
När det gäller den interna revisionskapaciteten, särskilt i förhållande till mindre organ, noterar Europaparlamentet det förslag som internrevisorn gjorde inför parlamentets ansvariga utskott den 14 september 2006 om att mindre organ ska tillåtas att köpa in interrevisionstjänster från den privata sektorn.
Utvärdering av organ
Rådsdokument DS 605/1/07 Rev1. som förhandlades fram vid medlingen inför Ekofinrådets budgetmöte den 13 juli 2007 där man efterlyser en förteckning på organ som kommissionen avser att utvärdera ii) en förteckning på de organ som redan utvärderats, tillsammans med en sammanfattning av resultaten.
Disciplinära förfaranden
Förslag till interinstitutionellt avtal
I den sammanfattande rapporten om kommissionens förvaltning 2006 (punkt 3.1, KOM(2007)0274 ) sägs att förhandlingarna sedermera avbröts, men att diskussioner om innehållet återupptogs i rådet i slutet av 2006.
Självfinansierade organ
Kontoret för harmonisering inom den inre marknaden har likvida medel på 281 miljoner EUR.
Gemenskapens växtsortsmyndighet har likvida medel på 18 miljoner EUR
Källa: Revisionsrättens särskilda rapport. .
· Intern kapacitet har avsatts och åtgärder har vidtagits för att hantera de identifierade svagheterna och för att förbättra de interna kontrollsystemen.
Europaparlamentet noterar från centrumets redovisning av det ekonomiska utfallet att det under 2006 uppnådde ett ekonomiskt resultat på 5,3 miljoner EUR på basis av intäkter på 15,8 miljoner EUR, med 7,2 miljoner EUR i likvida medel, och att balansräkningen innehåller en post på 400 000 EUR för förhandsfinansiering som ska betalas tillbaka till kommissionen.
39.
Detta är ett exempel som med fördel skulle kunna följas av alla organ.
3.3.2008
YTTRANDE från utskottet för miljö, folkhälsa och livsmedelssäkerhets
till budgetkontrollutskottet
över ansvarsfrihet för genomförandet av budgeten för Europeiska centrumet för förebyggande och kontroll av sjukdomar för budgetåret 2006
( C6-0386/2007 – 2007/2060(DEC) )
Föredragande: Jutta Haug
FÖRSLAG
Europaparlamentet uttrycker sin tillfredsställelse över det framgångsrika första verksamhetsåret för Europeiska centrumet för förebyggande och kontroll av sjukdomar (ECDC), och det effektiva genomförandet av 2006 års budget både när det gäller åtaganden och betalningar.
Europaparlamentet konstaterar dock att en betydande mängd åtaganden har flyttats över till 2007 på grund av oförutsägbarheten på vissa områden, i synnerhet i fråga om rekrytering.
På grundval av de uppgifter som finns tillgängliga anser Europaparlamentet att direktören för ECDC kan beviljas ansvarsfrihet för genomförandet av centrumets budget för budgetåret 2006.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
26.2.2008
Slutomröstning: resultat
+:
–:
0:
50
1
Slutomröstning: närvarande ledamöter
Adamos Adamou, Margrete Auken, Pilar Ayuso, Johannes Blokland, John Bowis, Magor Imre Csibi, Chris Davies, Avril Doyle, Mojca Drčar Murko, Edite Estrela, Jill Evans, Matthias Groote, Françoise Grossetête, Cristina Gutiérrez-Cortines, Satu Hassi, Gyula Hegyi, Jens Holm, Marie Anne Isler Béguin, Dan Jørgensen, Christa Klaß, Eija-Riitta Korhola, Holger Krahmer, Urszula Krupa, Aldis Kušķis, Peter Liese, Linda McAvan, Roberto Musacchio, Riitta Myller, Miroslav Ouzký, Vladko Todorov Panayotov, Vittorio Prodi, Guido Sacconi, Karin Scheele, Carl Schlyter, Richard Seeber, María Sornosa Martínez, Antonios Trakatellis, Evangelia Tzampazi, Thomas Ulmer, Marcello Vernola, Anja Weisgerber, Åsa Westlund, Anders Wijkman, Glenis Willmott
Slutomröstning: närvarande suppleanter
Kathalijne Maria Buitenweg, Philip Bushill-Matthews, Hélène Goudin, Genowefa Grabowska, Jutta Haug, Johannes Lebech, Lambert van Nistelrooij
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
26.3.2008
Slutomröstning: resultat
+:
–:
0:
27
4
2
Slutomröstning: närvarande ledamöter
Jean-Pierre Audy, Herbert Bösch, Costas Botopoulos, Mogens Camre, Paulo Casaca, Jorgo Chatzimarkakis, Antonio De Blasio, Esther De Lange, Petr Duchoň, James Elles, Szabolcs Fazakas, Markus Ferber, Christofer Fjellner, Ingeborg Gräßle, Dan Jørgensen, Rodi Kratsa-Tsagaropoulou, Bogusław Liberadzki, Nils Lundgren, Marusya Ivanova Lyubcheva, Hans-Peter Martin, Ashley Mote, Jan Mulder, Bill Newton Dunn, Borut Pahor, Bart Staes, Jeffrey Titford, Kyösti Virrankoski, Janusz Wojciechowski
Slutomröstning: närvarande suppleanter
Salvador Garriga Polledo, Edit Herczog, Cătălin-Ioan Nechifor, Dumitru Oprea, Pierre Pribetich, Margarita Starkevičiūtė
A6-0168/2008
BETÄNKANDE
om 2007 års lägesrapport om Turkiet
(2007/2269(INI))
Utskottet för utrikesfrågor
PE 402.879v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
YTTRANDE från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män 13
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................17
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om 2007 års lägesrapport om Turkiet
( 2007/2269(INI) )
Europaparlamentet utfärdar denna resolution,
– med beaktande av kommissionens lägesrapport 2007 om Turkiet ( SEK(2007)1436 ),
– med beaktande av sina tidigare resolutioner av den 27 september 2006 om Turkiets framsteg inför anslutningen
EUT C 306 E, 15.12.2006, s.
284. och den 24 oktober 2007 om förbindelserna mellan EU och Turkiet
Antagna texter, P6_TA(2007)0472 . ,
– med beaktande av de förhandlingsramar för Turkiet som antogs den 3 oktober 2005,
– med beaktande av rådets beslut 2008/158/EG av den 18 februari 2008 om principerna, prioriteringarna och villkoren i partnerskapet för anslutning med Republiken Turkiet
EUT L 51, 26.2.2008, s.
4. (nedan kallat partnerskapet för anslutning), samt rådets föregående beslut om partnerskapet för anslutning 2001, 2003 och 2006,
– med beaktande av artikel 45 i arbetsordningen,
– med beaktande av betänkandet från utskottet för utrikesfrågor och yttrandet från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män ( A6‑0168/2008 ), och av följande skäl:
A. Anslutningsförhandlingarna med Turkiet inleddes den 3 oktober 2005 efter rådets godkännande av förhandlingsramarna och detta utgjorde startpunkten för en lång process vars resultat inte kan garanteras i förväg.
C. En grundförutsättning för anslutning till EU är fortfarande att Köpenhamnskriterierna uppfylls helt och hållet och att EU – som är en gemenskap grundad på gemensamma värderingar – har förmåga att integrera nya medlemsstater i enlighet med slutsatserna från Europeiska rådets möte i december 2006.
D. I sin lägesrapport 2007 konstaterade kommissionen att när det gäller politiska reformer har ”bara begränsade framsteg gjorts under 2007” i Turkiet
Slutsatser om Turkiet, kommissionens lägesrapport 2007 om Turkiet, KOM(2007)0663 , SEK(2007)1436 . .
F. Turkiet har fortfarande inte genomfört de bestämmelser som följer av associeringsavtalet mellan EG och Turkiet och tilläggsprotokollet till detta.
G. Under 2007 öppnades fem förhandlingskapitel.
Reformer för att bygga upp ett demokratiskt och välmående samhälle
Europaparlamentet uppmanar de turkiska myndigheterna att inom ramen för rättsstatsprincipen beslutsamt utreda den kriminella Ergenekon-organisationen, att helt och hållet avslöja dess nätverk som sträcker sig in i de statliga strukturerna och att ställa alla inblandade inför rätta.
Regionala frågor och yttre förbindelser
Europaparlamentet välkomnar inrättandet av ett finansiellt stödinstrument för att främja den ekonomiska utvecklingen i det turkcypriotiska samhället, och uppmanar på nytt kommissionen att särskilt rapportera om tillämpningen av och effektiviteten i detta instrument.
Förbindelserna mellan EU och Turkiet
Europaparlamentet välkomnar nomineringen av Istanbul som 2010 års kulturhuvudstad eftersom detta är en möjlighet att stärka den interkulturella dialogen och det interkulturella samarbetet mellan EU och Turkiet.
Europaparlamentet beklagar att kommissionen inte har följt upp den konsekvensbedömning som lades fram 2004 och kräver att en sådan snarast ska läggas fram för parlamentet.
°
° °
till utskottet för utrikesfrågor
över 2007 års lägesrapport om Turkiet
( 2007/2269(INI) )
Föredragande:
Emine Bozkurt
FÖRSLAG
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män uppmanar utskottet för utrikesfrågor att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
– med beaktande av sina resolutioner av den 6 juli 2005
EUT C 157 E, 6.7.2006, s.
385. och den 13 februari 2007
EUT C 287 E, 29.11.2007, s.
Europaparlamentet framhåller hur viktigt det är att Turkiet bekämpar alla former av diskriminering i överensstämmelse med artikel 13 i EG-fördraget som kräver lika möjligheter för alla oavsett kön, ras, etniskt ursprung, religion eller övertygelse, funktionshinder, ålder eller sexuell läggning.
Europaparlamentet uppmanar den turkiska regeringen att snarast låta den jämställdhetslag som nämns i premiärministerns cirkulär av den 4 juli 2006 träda i kraft.
Europaparlamentet välkomnar den turkiska regeringens initiativ och åtgärder, men framhåller att ytterligare ansträngningar och fler åtgärder krävs för att stoppa alla former av våld mot kvinnor.
Europaparlamentet bekräftar betydelsen av frivilligorganisationer och övriga aktörer i civilsamhället, och uppmanar därför den turkiska regeringen att se till att dialogen med civilsamhället och kvinnoorganisationer stärks, samordnas och institutionaliseras, särskilt vid utarbetandet av den nya konstitutionen, och att se till att civilsamhället kontinuerligt deltar på alla politikområden, även när det gäller socialförsäkringar och förhandlingar med EU.
Europaparlamentet uppmanar de turkiska myndigheterna att fortsätta arbetet för att minska könsskillnaderna i grundskolan och bättre följa upp skolavhoppen särskilt när det gäller flickor.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
14.4.2008
Slutomröstning: resultat
+:
–:
0:
20
1
Slutomröstning: närvarande ledamöter
Emine Bozkurt, Maria Carlshamre, Zita Gurmai, Lívia Járóka, Piia-Noora Kauppi, Astrid Lulling, Siiri Oviir, Doris Pack, Zita Pleštinská, Karin Resetarits, Teresa Riera Madurell, Eva-Britt Svensson, Anne Van Lancker, Anna Záborská
Slutomröstning: närvarande suppleanter
Gabriela Creţu, Lidia Joanna Geringer de Oedenberg, Donata Gottardi, Anna Hedh, Marusya Ivanova Lyubcheva
Slutomröstning: närvarande suppleanter (art.
178.2)
Manolis Mavrommatis, Miroslav Mikolášik
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
21.4.2008
Slutomröstning: resultat
+:
–:
0:
53
2
4
Slutomröstning: närvarande ledamöter
Vittorio Agnoletto, Bastiaan Belder, André Brie, Elmar Brok, Marco Cappato, Philip Claeys, Véronique De Keyser, Giorgos Dimitrakopoulos, Michael Gahler, Georgios Georgiou, Bronisław Geremek, Ana Maria Gomes, Jana Hybášková, Jelko Kacin, Ioannis Kasoulides, Metin Kazak, Maria Eleni Koppa, Johannes Lebech, Willy Meyer Pleite, Francisco José Millán Mon, Philippe Morillon, Pasqualina Napoletano, Annemie Neyts-Uyttebroeck, Baroness Nicholson of Winterbourne, Raimon Obiols i Germà, Ria Oomen-Ruijten, Ioan Mircea Paşcu, Alojz Peterle, Bernd Posselt, Christian Rovsing, José Ignacio Salafranca Sánchez-Neyra, Jacek Saryusz-Wolski, György Schöpflin, Hannes Swoboda, Antonio Tajani, Charles Tannock, Geoffrey Van Orden, Kristian Vigenin, Jan Marinus Wiersma, Josef Zieleniec
Slutomröstning: närvarande suppleanter
Irena Belohorská, Giulietto Chiesa, Andrew Duff, Milan Horáček, Marie Anne Isler Béguin, Evgeni Kirilov, Marios Matsakis, Nickolay Mladenov, Doris Pack, Inger Segelström, Karl von Wogau
Slutomröstning: närvarande suppleanter (art.
178.2)
A6-0248/2008
***I
BETÄNKANDE
om förslaget till Europaparlamentets och rådets förordning om en uppförandekod för datoriserade bokningssystem
(KOM(2007)0709 – C6‑0418/2007 – 2007/0243(COD))
Utskottet för transport och turism
Föredragande:
Timothy Kirkhope
PE 402.929v02-00
Teckenförklaring
* Samrådsförfarandet
majoritet av de avgivna rösterna
**I Samarbetsförfarandet (första behandlingen)
majoritet av de avgivna rösterna
**II Samarbetsförfarandet (andra behandlingen)
*** Samtyckesförfarandet
majoritet av parlamentets samtliga ledamöter utom i de fall som avses i artiklarna 105, 107, 161 och 300 i EG-fördraget och artikel 7 i EU-fördraget
***I Medbeslutandeförfarandet (första behandlingen)
majoritet av de avgivna rösterna
***II Medbeslutandeförfarandet (andra behandlingen)
majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten
majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
***III Medbeslutandeförfarandet (tredje behandlingen)
majoritet av de avgivna rösterna för att godkänna det gemensamma utkastet
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Parlamentets ändringar markeras med fetkursiv stil .
I samband med ändringsakter ska de delar av en återgiven befintlig rättsakt som inte ändrats av kommissionen, men som parlamentet önskar ändra, markeras med fet stil .
Eventuella strykningar ska i sådana fall markeras enligt följande: [...].
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................33
YTTRANDE från utskottet för den inre marknaden och konsumentskydd 38
YTTRANDE från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor 48
ÄRENDETS GÅNG..................................................................................................................53
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till Europaparlamentets och rådets förordning om en uppförandekod för datoriserade bokningssystem
( KOM(2007)0709 – C6‑0418/2007 – 2007/0243(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
– med beaktande av artikel 51 i arbetsordningen,
– med beaktande av betänkandet från utskottet för transport och turism och yttrandena från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor och utskottet för den inre marknaden och konsumentskydd ( A6‑0248/2008 ).
Ändringsförslag
1
Förslag till förordning
Skäl 5a (nytt)
Kommissionens förslag
Ändringsförslag
(5a) Det är nödvändigt att verka för en effektiv konkurrens mellan deltagande transportföretag och moderföretag och att se till att lufttrafikföretag respekterar principen om icke-diskriminering oberoende av om de deltar i datoriserade bokningssystem eller inte.
Motivering
Koden bör utformas så att den främjar konkurrens samtidigt som den förhindrar att datoriserade bokningssystem diskriminerar lufttrafikföretag.
Ändringsförslag
2
Förslag till förordning
Skäl 5b (nytt)
Kommissionens förslag
Ändringsförslag
(5b) För att garantera öppna och jämförbara konkurrensvillkor på marknaden bör särskilda bestämmelser gälla för moderföretag då de investerar i datoriserade bokningssystem.
Motivering
Kompletterande bestämmelser, såsom de i artikel 10, bör gälla för moderföretag, för att förhindra en snedvridning av marknaden.
Ändringsförslag
3
Förslag till förordning
Skäl 5c (nytt)
Kommissionens förslag
Ändringsförslag
(5c) Det ska vara möjligt att hänvisa till EU:s konkurrensbestämmelser och konkurrensförfaranden för att undvika att ett eller flera moderföretag missbrukar sin dominerande ställning.
Motivering
Hänvisningarna till de allmänna konkurrensbestämmelserna bör stramas upp.
Uppförandekoden kompletterar dessa bestämmelser, men ersätter dem inte.
Ändringsförslag
4
Förslag till förordning
Skäl 6
Kommissionens förslag
Ändringsförslag
(6) Systemleverantörer bör göra tydlig åtskillnad mellan de datoriserade bokningssystemen och flygbolagens interna bokningssystem och bör avhålla sig från att låta distributionstjänsterna vara förbehållna moderföretagen, för att undvika att moderföretagen skulle kunna få förmånstillträde till bokningssystemet.
(6) Systemleverantörer bör göra tydlig åtskillnad mellan de datoriserade bokningssystemen och flygbolagens interna bokningssystem eller andra typer av bokningssystem, och bör avhålla sig från att låta distributionstjänsterna vara förbehållna moderföretagen, för att undvika att moderföretagen skulle kunna få förmånstillträde till bokningssystemet.
Ändringsförslag
5
Förslag till förordning
Skäl 7a (nytt)
Kommissionens förslag
Ändringsförslag
(7a) En neutral textbild ökar insynen i de transporttjänster som de deltagande transportföretagen erbjuder och ökar konsumenternas förtroende.
Motivering
Rangordningskriterierna måste vara rättvisa och syfta till att hjälpa resebyrån att erbjuda konsumenten de bästa resealternativen.
Ändringsförslag
6
Förslag till förordning
Skäl 8
Kommissionens förslag
Ändringsförslag
(8) Systemleverantörerna bör säkerställa att ett datoriserat bokningssystems saluföringsuppgifter är tillgängliga för alla deltagande transportföretag utan diskriminering, och transportörerna bör inte kunna använda de uppgifterna för att på ett otillbörligt sätt påverka valet av resebyrå.
(8) Systemleverantörerna bör säkerställa att ett datoriserat bokningssystems saluföringsuppgifter är tillgängliga för alla deltagande transportföretag utan diskriminering, och transportörerna bör inte kunna använda de uppgifterna för att på ett otillbörligt sätt påverka valet av resebyrå eller konsumentens eget val .
Ändringsförslag
7
Förslag till förordning
Skäl 9a (nytt)
Kommissionens förslag
Ändringsförslag
Ändringsförslag
8
Förslag till förordning
Skäl 9b (nytt)
Kommissionens förslag
Ändringsförslag
Denna information kan anges som den genomsnittliga bränsleförbrukningen per person/liter/100km och det genomsnittliga koldioxidutsläppet per person/g/km och kunde jämföras med uppgifter om bästa tåg- och bussförbindelser för resor kortare än 5 timmar.
Ändringsförslag
9
Kommissionens förslag
Ändringsförslag
Denna förordning ska tillämpas på datoriserade bokningssystem, i den mån de omfattar lufttransporttjänster, som tillhandahålls eller används inom gemenskapen.
(Berör inte den svenska versionen.)
Motivering
(Berör inte den svenska versionen.)
Ändringsförslag
10
Förslag till förordning
Kommissionens förslag
Ändringsförslag
Denna förordning ska också tillämpas på järnvägstransporttjänster, som är integrerade jämte lufttransporttjänsterna i den primära textbilden för datoriserade bokningssystem.
Denna förordning ska också tillämpas på järnvägstransporttjänster, som är integrerade jämte lufttransporttjänsterna i den primära textbilden för datoriserade bokningssystem , som tillhandahålls eller används inom gemenskapen .
Motivering
Järnvägstransporttjänster måste behandlas på samma sätt som lufttransporttjänster.
Ändringsförslag
11
Artikel 2 – led d
Kommissionens förslag
Ändringsförslag
d) datoriserat bokningssystem: ett datoriserat system som innehåller information om bland annat tidtabeller, platstillgång , biljettpriser och tjänster i samband med befordran , från mer än ett lufttrafikföretag, med eller utan möjlighet att boka platser eller utfärda biljetter, och där några av eller samtliga dessa tjänster ställs till abonnenternas förfogande.
d) datoriserat bokningssystem: ett datoriserat system som innehåller information om bland annat tidtabeller, platstillgång och biljettpriser, från mer än ett lufttrafikföretag, med eller utan möjlighet att boka platser eller utfärda biljetter, och där några av eller samtliga dessa tjänster ställs till abonnenternas förfogande.
Motivering
Den nuvarande ordalydelsen skapar förvirring om hur ett datoriserat bokningssystem ska definieras och om de tjänster som hör ihop med systemet och som ska ställas till abonnenternas förfogande.
Ändringsförslag
12
Förslag till förordning
Artikel 2 – led g
Kommissionens förslag
Ändringsförslag
g) moderföretag: ett lufttrafikföretag eller järnvägstransportföretag som direkt eller indirekt, ensamt eller tillsammans med andra, äger eller faktiskt kontrollerar en systemleverantör, liksom varje lufttrafikföretag eller järnvägstransportföretag som det äger eller faktiskt kontrollerar.
g) moderföretag: ett lufttrafikföretag eller järnvägstransportföretag som direkt eller indirekt, ensamt eller tillsammans med andra kontrollerar eller deltar i kapitalet eller har lagliga rättigheter och representation i styrelsen, den övervakande styrelsen eller andra ledningsorgan för en systemleverantör, liksom varje lufttrafikföretag eller järnvägstransportföretag som det äger eller faktiskt kontrollerar.
Motivering
Definitionen bör klargöras och utvidgas för att garantera att vederbörlig hänsyn tas till transportföretagens inflytande som en följd av aktieinnehav i systemleverantörer.
Det är berättigat att dra den slutsatsen att de fördelar som flygbolag förväntar sig av att inneha datoriserade bokningssystem har mer att göra med konkurrensfördelar än med kostnader.
Risken för missbruk är särskilt hög då ett dominerande flygbolag är delägare i ett dominerande datoriserat bokningssystem.
Det är svårt att fastställa ett tak för de fall då risken för diskriminering ökar.
Moderföretag bör inte otillbörligt påverka leverantören av datoriserade bokningssystem.
Därför behövs det stängare bestämmelser om moderföretag i syfte att garantera rättvisa och öppenhet.
Ändringsförslag
13
Artikel 2 – led ga (nytt)
Kommissionens förslag
Ändringsförslag
ga) deltagande i en systemleverantörs kapital: en kombination av det rent ekonomiska värdet av ett lufttrafikföretags eller järnvägstransportföretags investering i en systemleverantör och värdet av det berörda företagets äganderätt till systemleverantören.
Motivering
En enda ekonomisk investering i ett datoriserat bokningssystem bör inte medföra att ett flygbolag eller ett järnvägsbolag definieras som ”moderföretag”.
Endast om en sådan investering åtföljs av förvärv av äganderätter ska ett flyg- eller järnvägsbolag betraktas som ”moderföretag” och därmed efterleva kraven i artikel 10.
Detta innebär att hänsyn tas till oavsiktliga investeringar som inte medför någon möjlighet att påverka systemleverantörens verksamhet.
Ändringsförslag
14
Artikel 2 – led h
Kommissionens förslag
Ändringsförslag
h) faktiskt kontroll: ett förhållande som bygger på rättigheter, avtal eller andra medel, som var för sig eller tillsammans , och med hänsyn tagen till faktiska och rättsliga förhållanden, ger möjligheter att direkt eller indirekt utöva ett avgörande inflytande på ett företag, särskilt då det gäller
h) kontroll: ett förhållande som bygger på rättigheter, avtal eller andra medel, som var för sig eller i kombination , och med hänsyn tagen till faktiska och rättsliga förhållanden, ger möjligheter att utöva ett avgörande inflytande på ett företag, särskilt då det gäller
i) rätten att använda alla eller delar av ett företags tillgångar,
i) ägande eller rätten att använda alla eller delar av ett företags tillgångar,
ii) rättigheter eller avtal som ger ett avgörande inflytande på sammansättningen av företagets olika organ och på omröstningar eller beslut i organen , eller som på annat sätt ger ett avgörande inflytande på företagets verksamhet .
ii) rättigheter eller avtal som ger ett avgörande inflytande på sammansättningen av företagets olika organ och på omröstningar eller beslut i organen.
Motivering
Genom ändringsförslaget betonas parallellerna mellan uppförandekoden och konkurrenspolitiken.
Genom att använda samma definitioner som i koncentrationsförordningen kan man också tillämpa samma kriterier för hur kontrollen ska bedömas.
Minoritetsägande, även med mycket små andelar, kan medföra status som ”moderföretag”, om andelarna medför en möjlighet att påverka strategiska beslut inom ett datoriserat bokningssystem.
Detta kommer att vara fallet om ett flygbolag har möjlighet att utöva ett avgörande inflytande på bokningssystemet i det avseendet att flygbolaget kan blockera åtgärder som är avgörande för det datoriserade bokningssystemets strategiska kommersiella agerande.
Ändringsförslag
15
Kommissionens förslag
Ändringsförslag
a) knyta oskäliga villkor till ett avtal med ett deltagande transportföretag eller kräva att tilläggsvillkor godtas, som genom sin karaktär eller enligt kommersiell praxis saknar samband med deltagandet i leverantörens datoriserade bokningssystem,
a) knyta diskriminerande villkor till ett avtal med ett deltagande transportföretag eller kräva att tilläggsvillkor godtas, som genom sin karaktär eller enligt kommersiell praxis saknar samband med deltagandet i leverantörens datoriserade bokningssystem,
Motivering
Ändringsförslaget syftar till att undvika förvirring kring termen ”oskäliga”.
Ändringsförslag
16
Kommissionens förslag
Ändringsförslag
b) ställa som villkor för deltagande i det datoriserade bokningssystemet att ett deltagande transportföretag inte samtidigt deltar i ett annat system.
b) ställa som villkor för deltagande i det datoriserade bokningssystemet att ett deltagande transportföretag inte samtidigt deltar i ett annat system eller att ett deltagande transportföretag inte fritt får använda alternativa bokningssystem, t.ex. sitt eget bokningssystem på Internet eller teletjänstcentraler .
Motivering
Ändringsförslaget syftar till att förhindra att ett datoriserat bokningssystem kan kringgå flygbolagets frihet att förhandla genom att vägra låta flygbolaget delta i systemet om det inte begränsar användningen av andra bokningskanaler.
Ändringsförslag
17
Kommissionens förslag
Ändringsförslag
2a.
Ett lufttrafik- eller järnvägstransportföretags direkta eller indirekta aktieinnehav i en systemleverantör eller en systemleverantörs direkta eller indirekta aktieinnehav i ett lufttrafik- eller järnvägstransportföretag, aktieinnehavets storlek samt den kontroll som ett sådant innehav ger upphov till ska offentliggöras.
Motivering
Denna information bör offentliggöras i syfte att tillämpa bestämmelserna i artiklarna 3 och 10 samt för att få insyn i förhållandena mellan systemleverantörer och lufttrafikföretag.
Ändringsförslag
18
Kommissionens förslag
Ändringsförslag
1.
En systemleverantör får inte reservera någon specifik datainläsningsmetod, databehandlingsmetod eller distributionstjänst – eller några förbättringar av dessa – för ett eller flera av sina moderföretag.
1.
En systemleverantör får inte reservera någon specifik datainläsningsmetod, databehandlingsmetod eller distributionstjänst – eller några förändringar av dessa – för ett eller flera deltagande transportföretag, medräknat sina moderföretag.
Systemleverantören ska tillhandahålla de deltagande transportföretagen information om samtliga förändringar i sina distributionssystem och datainläsnings- eller databehandlingsmetoder.
Motivering
Ändringsförslaget stärker principen om icke-diskriminering mellan flygbolag i fråga om distributionssystem.
Alla flygbolag bör ha tillgång till de senaste tekniska förbättringarna.
För att garantera öppenhet kring de tillgängliga systemen bör de datoriserade bokningssystemen tillhandahålla alla flygbolag information om dem.
Ändringsförslag
19
Kommissionens förslag
Ändringsförslag
1.
Systemleverantören ska via sitt datoriserade bokningssystem tillhandahålla en eller flera primära textbilder för varje enskild transaktion och ska däri inkludera de uppgifter som lämnats in av deltagande transportföretag på ett neutralt och uttömmande sätt som inte är diskriminerande eller partiskt.
Kriterierna för rangordningen av upplysningarna får inte baseras på någon faktor som direkt eller indirekt har samband med transportföretagens identitet och inte tillämpas på ett sätt som diskriminerar något deltagande lufttrafikföretag.
Den eller de primära textbilderna ska vara förenliga med reglerna i bilaga 1.
1.
Systemleverantören ska via sitt datoriserade bokningssystem tillhandahålla en eller flera primära textbilder för varje enskild transaktion och ska däri inkludera de uppgifter som lämnats in av deltagande transportföretag på ett neutralt och uttömmande sätt som inte är diskriminerande , partiskt eller favoriserande .
Kriterierna för rangordningen av upplysningarna får inte baseras på någon faktor som direkt eller indirekt har samband med transportföretagens identitet och inte tillämpas på ett sätt som diskriminerar något deltagande lufttrafikföretag.
Den eller de primära textbilderna får inte avsiktligt vilseleda konsumenter, bör vara lättillgängliga och ska vara förenliga med reglerna i bilaga 1.
Motivering
Det är viktigt att lägga till favorisering som inte ingår i kommissionens ursprungliga formulering.
Den ursprungliga ordalydelsen är inte exakt och kan lämna möjlighet till olika tolkningar.
Ändringsförslag
20
Kommissionens förslag
Ändringsförslag
2.
För de upplysningar som ett datoriserat bokningssystem tillhandahåller ska en abonnent använda en neutral textbild i enlighet med punkt 1, om inte en annan textbild krävs för att tillgodose konsumentens önskemål.
2.
För de upplysningar som ett datoriserat bokningssystem tillhandahåller konsumenten ska en abonnent använda en neutral textbild i enlighet med punkt 1, om inte en annan textbild krävs för att tillgodose konsumentens önskemål.
Motivering
Föredragandens ursprungliga ändringsförslag behöver förtydligas.
Den nya ordalydelsen förhindrar en sådan feltolkning att abonnenten inte skulle få använda information från någon annan källa än det datoriserade bokningssystemets textbild.
Ändringsförslag
21
Kommissionens förslag
Ändringsförslag
2a.
Flygningar som utförs av lufttrafikföretag som förbjudits att bedriva verksamhet enligt förordning (EG) nr 2111/2005 ska klart och specifikt markeras på textbilden.
Motivering
Syftet med detta ändringsförslag är att underlätta tillämpningen av förordning (EG) nr 2111/2005 och att på bästa sätt garantera målen i den.
Ändringsförslag
22
Kommissionens förslag
Ändringsförslag
2b.
Systemleverantören ska införa en särskild symbol i det datoriserade bokningssystemets textbild som användarna ska kunna identifiera för att få information om vilket lufttrafikföretag som utför en viss flygning enligt artikel 11 i förordning (EG) nr 2111/2005.
Motivering
Det är viktigt att de som använder datoriserade bokningssystem (resebyråer eller allmänheten generellt) är medvetna om flygningar som utförs av lufttrafikföretag på EU:s svarta lista, enligt förordning (EG) nr 2111/2005.
Ändringsförslag
23
Kommissionens förslag
Ändringsförslag
3.
Denna artikel ska inte tillämpas på datoriserade bokningssystem som används av ett lufttrafikföretag eller ett järnvägstransportföretag, eller en grupp av lufttrafikföretag eller järnvägstransportföretag, i deras egna klart markerade kontor och försäljningsdiskar.
3.
Denna artikel ska inte tillämpas på datoriserade bokningssystem som används av ett lufttrafikföretag eller ett järnvägstransportföretag, eller en grupp av lufttrafikföretag eller järnvägstransportföretag, i deras egna klart markerade kontor , försäljningsdiskar eller på deras egna webbsidor .
Motivering
Det här är inte rätta forumet för att ta upp frågor som rör företagens egna webbsidor.
Ändringsförslag
24
Kommissionens förslag
Ändringsförslag
1.
En systemleverantör får inte knyta orimliga villkor till ett avtal med en abonnent, t.ex. hindra abonnenten från att abonnera på eller använda ett eller flera andra system, kräva att ytterligare villkor accepteras som inte har samband med deltagandet i dess datoriserade bokningssystem, eller kräva att abonnenten accepterar ett erbjudande om teknisk utrustning eller programvara.
1.
En systemleverantör får inte knyta diskriminerande villkor till ett avtal med en abonnent, t.ex. hindra abonnenten från att abonnera på eller använda ett eller flera andra system, kräva att ytterligare villkor accepteras som inte har samband med deltagandet i dess datoriserade bokningssystem, eller kräva att abonnenten accepterar ett erbjudande om teknisk utrustning eller programvara.
Motivering
Ändringsförslaget syftar till att förhindra förvirring kring termen ”oskäliga”.
Ändringsförslag
25
Förslag till förordning
Artikel 7
Kommissionens förslag
Ändringsförslag
Systemleverantörerna får på följande villkor tillgängliggöra alla saluförings-, boknings- och försäljningsuppgifter :
1.
Systemleverantörerna får tillgängliggöra alla saluförings-, boknings- och försäljningsuppgifter under förutsättning att uppgifterna erbjuds alla deltagande lufttrafikföretag, inklusive moderföretag, inom samma tidsramar och på ett icke-diskriminerande sätt.
Uppgifterna får – och ska på begäran – omfatta alla deltagande transportföretag och abonnenter.
a) Uppgifterna erbjuds alla deltagande lufttrafikföretag, inklusive moderföretag, inom samma tidsramar och på ett icke-diskriminerande sätt.
Uppgifterna får – och ska på begäran – omfatta alla deltagande transportföretag och abonnenter.
2.
Deltagande transportföretag får inte använda sådana uppgifter för att påverka abonnentens val på ett otillbörligt sätt.
b) Om uppgifterna har framkommit då en abonnent med säte i Europeiska unionen använt distributionstjänsterna i ett datoriserat bokningssystem, får de inte innehålla någon identifikation, varken direkt eller indirekt, av abonnenten.
3.
Om uppgifterna har framkommit då en abonnent med säte i gemenskapen använt distributionstjänsterna i ett datoriserat bokningssystem, får de inte innehålla någon identifikation, varken direkt eller indirekt, av abonnenten , om inte abonnenten och systemleverantören har kommit överens om villkoren för lämplig användning av sådana uppgifter .
4.
Alla eventuella avtal mellan abonnenter och systemleverantörer om databand med saluföringsinformation (MIDT) ska offentliggöras.
Motivering
Resebyråerna ska själva få bestämma om deras uppgifter ska tas med i databanden med saluföringsinformation (MIDT).
Därmed skapar artikel 7 b ett monopol för IATA, och de ökade kostnaderna för marknadsuppgifter medför högre priser för konsumenterna.
Ändringsförslag
26
Kommissionens förslag
Ändringsförslag
ba) Avtal mellan abonnenter och systemleverantörer av databand med saluföringsinformation (MIDT) får innehålla ett kompensationssystem som gynnar abonnenterna.
Motivering
I avtal mellan resebyråer och datoriserade bokningssystem om databand med saluföringsinformation ska det finnas möjlighet till kompensation, inklusive ersättning.
Ändringsförslag
27
Kommissionens förslag
Ändringsförslag
Kommissionen ska på begäran av en medlemsstat eller på eget initiativ utreda eventuella fall av diskriminering av EU ‑företag i datoriserade bokningssystem i tredjeländer.
Om det konstateras att diskriminering förekommer ska kommissionen innan den fattar något beslut informera medlemsstaterna och berörda parter och inhämta deras synpunkter, bland annat genom att sammankalla relevanta experter från medlemsstaterna.
Motivering
Utredningen av om lufttrafikföretag i gemenskapen utsätts för diskriminerande eller ojämlik behandling av systemleverantörer utanför EU bör övervakas av kommissionen.
Ändringsförslag
28
Kommissionens förslag
Ändringsförslag
1.
Ett moderföretag får inte, för någon av de lufttransporttjänster som distribueras genom deras eget system, diskriminera ett konkurrerande datoriserat bokningssystem genom att vägra att på begäran och inom samma tidsramar tillhandahålla det senare samma information om tidtabeller, biljettpriser och platstillgång avseende sina egna transporttjänster som det ger de egna datoriserade bokningssystemen, eller genom att distribuera sina egna transporttjänster via ett annat datoriserat bokningssystem eller vägra att inom samma tidsramar godkänna eller bekräfta bokningar som har gjorts via ett konkurrerande system.
Moderföretaget ska bara vara skyldigt att acceptera och bekräfta de bokningar som överensstämmer med dess biljettpriser och villkor.
1.
Ett moderföretag får inte, om det inte är ömsesidigt, för någon av de lufttransporttjänster som distribueras genom deras eget system, diskriminera ett konkurrerande datoriserat bokningssystem genom att vägra att på begäran och inom samma tidsramar tillhandahålla det senare samma information om tidtabeller, biljettpriser och platstillgång avseende sina egna transporttjänster som det ger de egna datoriserade bokningssystemen, eller genom att distribuera sina egna transporttjänster via ett annat datoriserat bokningssystem eller vägra att inom samma tidsramar godkänna eller bekräfta bokningar som har gjorts via ett konkurrerande system.
Moderföretaget ska bara vara skyldigt att acceptera och bekräfta de bokningar som överensstämmer med dess biljettpriser och villkor.
Motivering
Det är önskvärt att införa en ömsesidighetsklausul i förbindelserna mellan de datoriserade bokningssystemen.
Ändringsförslag
29
Kommissionens förslag
Ändringsförslag
1a.
Omvänt kan ett konkurrerande datoriserat bokningssystem inte vägra att på samma villkor som de som beviljas övriga kunder och abonnenter på vilken som helst marknad vara databasvärd för information om tidtabeller, priser och tillgängliga platser vad gäller de transporttjänster som en transportör erbjuder som är knuten till andra datoriserade bokningssystem.
Motivering
Syftet med ändringsförslaget är att klargöra förhållandena mellan konkurrerande datoriserade bokningssystem.
Ändringsförslag
30
Förslag till förordning
2.
Den bokningsavgift som ska betalas till det datoriserade bokningssystemet för en godkänd bokning som gjorts i enlighet med punkt 1, får inte överskrida avgiften för en likvärdig transaktion som ska betalas av andra deltagande lufttrafikföretag till samma datoriserade bokningssystem eller till deras egna datoriserade bokningssystem .
2.
Moderföretaget ska inte vara förpliktat att godta kostnader i samband med detta utom för återgivande av de uppgifter som ska lämnas in och för godkända bokningar.
Den bokningsavgift som ska betalas till det datoriserade bokningssystemet för en godkänd bokning som gjorts i enlighet med punkt 1, ska vara i linje med avgiften för en likvärdig transaktion som ska betalas av andra deltagande lufttrafikföretag till samma datoriserade bokningssystem.
Kommissionen kan när som helst be en systemleverantör att lämna all den information som behövs för att utvärdera om systemleverantören respekterar denna punkt.
Motivering
Det bör klart och tydligt framgå av texten att den avgift som moderföretag betalar bör ligga nära den som andra betalar för samma datoriserade bokningssystem (för likadana transaktioner).
Ändringsförslag
31
Förslag till förordning
3.
3.
Ett moderföretag får inte gynna sitt eget datoriserade bokningssystem genom att , direkt eller indirekt, knyta en abonnents användning av ett visst datoriserat bokningssystem till provision eller någon annan fördel eller nackdel vid försäljningen av företagets transporttjänster.
Motivering
Ett moderföretag får inte förbjudas att förhandla med datoriserade bokningssystem som det inte är knutet till.
Ett moderföretag är, när det gäller dessa datoriserade bokningssystem, i samma situation som andra transportörer.
Förhandlingarna får dock inte gynna det egna datoriserade bokningssystemet.
Ändringsförslag
32
Förslag till förordning
4.
4.
Ett moderföretag får varken direkt eller indirekt gynna sitt eget datoriserade bokningssystem genom att kräva att en abonnent använder ett visst datoriserat bokningssystem för att sälja eller utfärda biljetter för en transporttjänst som företaget självt direkt eller indirekt tillhandahåller.
Motivering
Ett moderföretag får inte förbjudas att förhandla med datoriserade bokningssystem som det inte är knutet till.
Ett moderföretag är, när det gäller dessa datoriserade bokningssystem, i samma situation som andra transportörer.
Förhandlingarna får dock inte gynna det egna datoriserade bokningssystemet.
Ändringsförslag
33
Kommissionens förslag
Ändringsförslag
1.
Personuppgifter ska behandlas av ett datoriserat bokningssystem uteslutande i samband med att bokningar görs eller biljetter utfärdas för transporttjänster.
1.
Personuppgifter som samlats in av ett datoriserat bokningssystem i samband med att bokningar görs eller biljetter utfärdas för transporttjänster ska endast behandlas på ett sätt som är förenligt med dessa ändamål .
Det datoriserade bokningssystemet ska skilja mellan personuppgifter som behövs för passageraruppgifter (PNR-uppgifter) eller kommersiellt bruk enligt principen med blandade uppgifter och all annan eventuell passagerarinformation som finns i systemet.
Sådana personuppgifter får endast göras tillgängliga för andra enheter om personen eller organisationen i fråga uttryckligen har gett sitt skriftliga samtycke.
Motivering
Syftet med detta ändringsförslag är att förbättra den rättsliga klarheten genom att använda den korrekta definitionen (systemleverantör) i stället för det datoriserade bokningssystemet som inte är en rättslig term.
Ändringsförslag
34
Förslag till förordning
3.
3.
När det rör sig om särskilda kategorier av uppgifter i enlighet med artikel 8 i direktiv 95/46/EG, ska sådana uppgifter endast behandlas om den registrerade har gett sitt uttryckliga , informerade medgivande till det.
Motivering
Medgivandet måste grundas på korrekt information.
Ändringsförslag
35
Förslag till förordning
5.
5.
Det ska inte vara möjligt att varken direkt eller indirekt identifiera fysiska personer, eller i tillämpliga fall de organisationer eller företag på vars vägnar de agerar, via de uppgifter om saluföring, bokföring och försäljning som en systemleverantör tillgängliggör.
Motivering
Syftet med detta ändringsförslag är att förbättra den rättsliga klarheten genom att använda den korrekta definitionen (systemleverantör) i stället för det datoriserade bokningssystemet som inte är en rättslig term.
Ändringsförslag
36
Förslag till förordning
7.
7.
Den registrerade ska ha rätt att kostnadsfritt få tillgång till uppgifter om sig själv oberoende av om uppgifterna är lagrade hos systemleverantören eller hos abonnenten.
Motivering
Syftet med detta ändringsförslag är att förbättra den rättsliga klarheten genom att använda den korrekta definitionen (systemleverantör) i stället för det datoriserade bokningssystemet som inte är en rättslig term.
Ändringsförslag
37
Förslag till förordning
8.
8.
De rättigheter som tas upp i denna artikel kompletterar och existerar vid sidan av de rättigheter för registrerade som fastställs i direktiv 95/46/EG , i de nationella bestämmelser som antagits i enlighet därmed och i internationella avtal som EU ingått .
Ändringsförslag
38
Förslag till förordning
9.
Om inte annat anges ska definitionerna i det direktivet gälla.
Denna förordning ska inte påverka bestämmelserna i nämnda direktiv och de nationella bestämmelser som medlemsstaterna antagit i enlighet därmed, om de särskilda bestämmelserna när det gäller bearbetning av personuppgifter i samband med den verksamhet hos ett datoriserat bokningssystem som fastställs i denna artikel inte är tillämpliga.
9.
Bestämmelserna i denna förordning ska precisera och komplettera direktiv 95/46/EG för de ändamål som avses i artikel 1.
Om inte annat anges ska definitionerna i det direktivet gälla.
Denna förordning ska inte påverka bestämmelserna i nämnda direktiv , de nationella bestämmelser som medlemsstaterna antagit i enlighet därmed och internationella avtal som EU ingått , om de särskilda bestämmelserna när det gäller bearbetning av personuppgifter i samband med den verksamhet hos ett datoriserat bokningssystem som fastställs i denna artikel inte är tillämpliga.
Ändringsförslag
39
Kommissionens förslag
Ändringsförslag
9a.
Om en systemleverantör förvaltar databaser i olika egenskaper, t.ex. erbjuder ett datoriserat bokningssystem eller fungerar som databasvärd för flygbolag, ska tekniska och organisatoriska åtgärder vidtas för att förhindra samkörning av databaserna och se till att personuppgifter endast är tillgängliga för de särskilda ändamål som de samlats in för.
Motivering
Ändringsförslaget stärker brandväggen mellan datoriserade bokningssystem och värdtjänster.
Ändringsförslag
40
Förslag till förordning
Artikel 11a (ny)
Kommissionens förslag
Ändringsförslag
Inspektion
1.
Samtliga systemleverantörer, som ett lufttrafikföretag eller ett järnvägstransportföretag investerat kapital i, ska vart tredje år på begäran av kommissionen, lägga fram en oberoende inspektionsrapport med detaljerade uppgifter om ägarstrukturen och förvaltningsmodellen.
Systemleverantören ska stå för kostnaderna för inspektionsrapporten.
2.
Systemleverantören ska säkerställa att en oberoende kontrollant på årsbasis övervakar att dess datoriserade bokningssystem är tekniskt förenligt med artiklarna 4, 7 och 11, samt i tillämpliga fall artikel 10.
Samtliga systemleverantörer ska vart tredje år eller på begäran från kommissionen lämna sin inspektionsrapport till kommissionen.
Systemleverantören ska stå för kostnaderna för inspektionsrapporten.
3.
Samtliga lufttrafikföretag eller järnvägstransportföretag som direkt äger en systemleverantör ska vart tredje år samt på begäran av kommissionen lägga fram en oberoende inspektionsrapport med detaljerade uppgifter om sina anknytningar till systemleverantören och dess förvaltningsmodell.
Lufttrafikföretaget eller järnvägstransportföretaget ska stå för kostnaderna för inspektionsrapporten.
4.
Systemleverantören ska meddela de deltagande transportföretagen och kommissionen namnet på kontrollanten senast tre månader innan utnämningen bekräftas.
Kommissionen ska intyga att kontrollanten är kompetent, såvida inte något av de deltagande företagen inom en månad efter meddelandet ifrågasätter kontrollantens förmåga att utföra sina uppgifter enligt denna artikel.
I sådana fall ska kommissionen inom ytterligare två månader och efter samråd med kontrollanten, systemleverantören och eventuella andra parter som hävdar ett berättigat intresse besluta om kontrollanten ska ersättas.
5.
Kontrollanten ska när som helst beviljas tillträde till de program, metoder, förfaranden och säkerhetskrav som används i de datorer eller datorsystem genom vilka systemleverantören erbjuder sina distributionstjänster.
6.
Kommissionen ska granska de rapporter som avses i punkterna 1, 2 och 3 för att avgöra om den behöver vidta åtgärder enligt artikel 12.
Motivering
Där det fortfarande finns nära förbindelser mellan flygbolag och datoriserade bokningssystem måste insyn ges i dessa företags ägarstruktur och förvaltningsmodell i syfte att bistå kommissionen i dess arbete med att övervaka att konkurrensen är rättvis.
Kontrollanten bör få fullständigt tillträde för att kunna göra en rättvis bedömning.
I texten återinförs bestämmelser om kontroll från den tidigare uppförandekoden som behövs för att få insyn i sektorn.
Ändringsförslag
41
Kommissionens förslag
Ändringsförslag
7.
Kommissionen ska i samråd med berörda parter utarbeta riktlinjer för den inspektionsrapport som avses i punkterna 1, 2 och 3.
Motivering
Där det fortfarande finns nära förbindelser mellan flygbolag och datoriserade bokningssystem måste insyn ges i dessa företags ägarstruktur och förvaltningsmodell i syfte att bistå kommissionen i dess arbete att övervaka att konkurrensen är rättvis.
Ändringsförslag
42
Kommissionens förslag
Ändringsförslag
8.
Kommissionen ska intyga att den kontrollant som det hänvisas till i punkterna 1,2 och 3 är kompetent.
Motivering
Det är kommissionen som ska godkänna kontrollanten.
Ändringsförslag
43
Förslag till förordning
Artikel 12
Kommissionens förslag
Ändringsförslag
Om kommissionen till följd av ett klagomål eller på eget initiativ konstaterar att denna förordning överträds, får den genom beslut ålägga de berörda företagen eller företagssammanslutningarna att se till att överträdelsen upphör.
Om kommissionen till följd av ett klagomål eller på eget initiativ konstaterar att denna förordning överträds, får den genom beslut ålägga de berörda företagen eller företagssammanslutningarna att se till att överträdelsen upphör.
Utredningar av möjliga överträdelser till denna förordning ska till fullo beakta resultaten av en eventuell undersökning enligt artiklarna 81 och 82 i EG-fördraget.
Motivering
Uppförandekoden för datoriserade bokningssystem ersätter inte utan kompletterar bara de gällande konkurrensreglerna, som fortsätter att vara fullt tillämpliga.
Ändringsförslag
44
Förslag till förordning
Artikel 13
Kommissionens förslag
Ändringsförslag
Kommissionen får när den fullgör de uppgifter som den tilldelas genom denna förordning genom en enkel begäran eller genom beslut begära att företag eller företagssammanslutningar överlämnar alla nödvändiga upplysningar.
Kommissionen får när den fullgör de uppgifter som den tilldelas genom denna förordning genom en enkel begäran eller genom beslut begära att företag eller företagssammanslutningar överlämnar alla nödvändiga upplysningar , särskilt i frågor som omfattas av artiklarna 4, 7 och 11, dock med förbehåll för de strängaste kraven för dataskydd som gäller i den berörda medlemsstaten .
Ändringsförslag
45
Förslag till förordning
Artikel 17
Kommissionens förslag
Ändringsförslag
Senast fem år efter det att denna förordning har trätt i kraft ska kommissionen utarbeta en rapport om tillämpningen av denna förordning, där det ska bedömas om det är nödvändigt att bibehålla, ändra eller upphäva förordningen.
Senast tre år efter det att denna förordning har trätt i kraft ska kommissionen utarbeta en rapport om tillämpningen av denna förordning, där det ska bedömas om det är nödvändigt att bibehålla, ändra eller upphäva förordningen.
Motivering
Ändringsförslag
46
Kommissionens förslag
Ändringsförslag
Motivering
Europaparlamentets utskott för transport och turism ska vartannat år regelbundet informeras genom en rapport om hur systemleverantörer som är verksamma i tredjeländer behandlar lufttrafikföretag.
Lufttransportavtal med tredjeländer verkar vara det regelverk som är bäst lämpat för att hantera sådana situationer eller fall.
Ändringsförslag
47
Förslag till förordning
Bilaga I
Kommissionens förslag
Ändringsförslag
1.
När biljettpriserna framgår av den primära textbilden eller när en rangordning görs efter biljettpriserna , ska priserna anges inklusive alla tillämpliga och obligatoriska skatter och avgifter som ska betalas till transportören .
1.
När priserna framgår av den primära textbilden eller när en rangordning görs efter priset , ska priserna anges inklusive biljettpriserna och alla tillämpliga skatter , tillägg och avgifter som ska betalas till lufttrafik- eller järnvägstransportföretaget och som är obligatoriska och förutsebara när de visas i textbilden .
2.
Vad gäller de uppgifter som ska ingå i den primära textbilden får vid sammanställning och val av transporttjänster mellan två givna orter ingen diskriminering ske mellan flygplatser eller järnvägsstationer som betjänar samma ort.
2.
Vad gäller de uppgifter som ska ingå i den primära textbilden får vid sammanställning och val av transporttjänster mellan två givna orter ingen diskriminering ske mellan flygplatser eller järnvägsstationer som betjänar samma ort.
3.
Det ska klart framgå vilken lufttransport som inte är regelbunden.
En konsument ska ha rätt att på begäran få en primär textbild med enbart antingen regelbunden eller icke-regelbunden lufttransport.
3.
Det ska klart framgå vilken lufttransport som inte är regelbunden.
En konsument ska ha rätt att på begäran få en primär textbild med enbart antingen regelbunden eller icke-regelbunden lufttransport.
4.
Det ska klart framgå vilka flygningar som innefattar mellanlandningar.
4.
Det ska klart framgå vilka flygningar som innefattar mellanlandningar.
5.
När en flygning utförs av ett lufttrafikföretag som inte är det lufttrafikföretag som anges i lufttrafikföretagskoden, ska det klart framgå vem som utför flygningen.
Detta krav kommer att gälla vid alla tillfällen, utom vid kortvariga särskilda arrangemang.
5.
När en flygning utförs av ett lufttrafikföretag som inte är det lufttrafikföretag som anges i lufttrafikföretagskoden, ska det klart framgå vem som utför flygningen.
Detta krav kommer att gälla vid alla tillfällen, utom vid kortvariga särskilda arrangemang.
6.
Information om kombinerade tjänster – dvs. en på förhand avtalad kombination av en transport och andra tjänster som inte är bitjänster till transporten, som erbjuds till försäljning till ett totalpris – ska inte visas i den primära textbilden.
6.
Information om kombinerade tjänster – dvs. en på förhand avtalad kombination av en transport och andra tjänster som inte är bitjänster till transporten, som erbjuds till försäljning till ett totalpris – ska inte visas i den primära textbilden.
6a.
Beroende på vad abonnenten väljer ska resealternativen på den primära textbilden rangordnas antingen utifrån biljettpris eller i följande ordning:
(i) alternativ för resa utan uppehåll rangordnade efter avgångstid,
(ii) övriga resealternativ rangordnade efter avverkad restid.
6b.
Med undantag för vad som anges i punkt 6e får inga resealternativ visas mer än en gång i någon primär textbild.
6c.
6d.
När resealternativ som erbjuds via det datoriserade bokningssystemet för två givna orter inkluderar anslutningsflyg eller erbjuds som en kombination av reguljär flyg- och järnvägsförbindelse, ska åtminstone den bästa reguljära flyg- och tågförbindelsen visas på den första sidan av den primära textbilden.
6e.
När olika lufttrafikföretag har flygningar med gemensam linjebeteckning ska de olika enskilda lufttrafikföretagskoderna tydligt anges en gång och det ska framgå vem som utför flygningen.
Motivering
Punkt 1 i bilaga I handlar om biljettpriser.
Detta kan vara förvirrande eftersom definitionen av ”biljettpriser” inte nödvändigtvis omfattar allt som ingår i priset.
För bästa möjliga prisinsyn är det bättre om man hänvisar till priset istället för till biljettpriset.
För kortare avstånd bör även alternativa tågförbindelser visas på den första sidan för att främja mer miljövänliga transportsätt.
När resealternativen för en viss ort erbjuds med anslutningsflyg bör den primära textbilden visa den bästa reguljära flyg- och tågförbindelsen, om det finns någon sådan.
Detta förslag medger ett undantag när det gäller avtal om gemensam linjebeteckning, så att man inte avskräcker från denna typ av avtal som ger framför allt mindre lufttrafikföretag möjlighet att erbjuda sina passagerare ett större flygnät.
Konsumenterna bör tjäna på att få bättre information.
MOTIVERING
Uppförandekoden för datoriserade bokningssystem fastställer hur resebokningar ska hanteras av lufttrafikföretag, järnvägstransportföretag, datoriserade bokningssystem och resebyråer.
Koden gäller i huvudsak flygbokningar, men också järnvägstransporttjänster som är integrerade i lufttransportbokningssystem.
Denna uppförandekod utarbetades under andra marknadsvillkor än de som nu råder.
Det stora flertalet flygbokningar skedde via datoriserade bokningssystem, som till största delen ägdes eller kontrollerades av flygbolag.
Uppförandekoden fastställdes för att främja insyn och förhindra marknadsmissbruk eller en snedvridning av konkurrensen genom tillfälliga bestämmelser.
Denna kod lämpar sig dock allt mindre med tanke på de nya marknadsvillkoren, avregleringen av andra marknader för datoriserade bokningssystem runt om i världen, utvecklingen av alternativa distributionskanaler och flygbolagens ökade delägande i de datoriserade bokningssystemen.
Kommissionens förslag
Huvudsyftet med kommissionens förslag är att göra det möjligt för flygbolag och datoriserade bokningssystem att fritt kunna förhandla om villkoren för tillhandahållandet av lufttjänster.
System ska tävla om priser och kvaliteten på tjänster.
Trots det erkänner man i förslaget att det bör finnas en balans mellan behovet att tillåta större konkurrens och behovet av grundläggande skyddsåtgärder.
Då berörda parter rådfrågades förklarade de att vissa skyddsåtgärder fortfarande behövdes, framför allt för att garantera en rättvis konkurrens i förhållande till ”moderföretag”, för att garantera att textbilderna i de datoriserade bokningssystemen är neutrala och för skydd av personuppgifter.
I kommissionens förslag ändras inte definitionen av moderföretag, vilket innebär att man har kvar det dubbla kriteriet rörande ägarskap och effektiv kontroll.
I kommissionens förslag förenklas reglerna för datoriserade bokningssystem, särskilt reglerna för deras avtalsförhållande med lufttrafikföretag, vilket möjliggör större frihet att förhandla om innehåll och priser.
När det gäller databand med saluföringsinformation (MIDT) föreslår kommissionen dock en ändring till den nuvarande koden.
Genom att ta bort möjligheten att identifiera resebyråer i denna information syftar kommissionen till att förhindra att lufttrafikföretag eventuellt påverkar resebyråer och deras distributionsmetoder.
De viktigaste punkterna i förslaget
Bestämmelser för moderföretag
Under de senaste åren har flygbolag gjort sig av med sitt innehav av datoriserade bokningssystem.
Det finns dock ett undantag: Amadeus.
Amadeus ägs av tre flygbolag med minoritetsandelar, Air France, Iberia och Lufthansa
Flygbolagens ägarandelar i Amadeus: Air France 23 procent, Iberia 11 procent, Lufthansa 11 procent, BC Partners and Cinven 53 procent, (Europeiska kommissionen – DG TREN konsekvensbedömning, SEK(2007)1496 ). .
Det är oklart hur stort strategiskt inflytande detta ägande ger dem, men det är klart att skyddsåtgärder behövs mot eventuellt missbruk.
Databand med saluföringsinformation (MIDT)
Med MIDT avses bokningsuppgifter som ett datoriserat bokningssystem behandlat och sålt till lufttrafikföretag.
Detta kan hjälpa flygbolagen att förstå marknadstrender och konkurrensinformation.
Till följd av alternativa distributionskanaler för bokningar har värdet på dessa uppgifter minskat, eftersom de inte är representativa för hela marknaden.
Medan majoriteten av tillhandahållarna av datoriserade bokningssystem och flygbolagen fortfarande skulle vilja att det skulle vara möjligt att identifiera resebyråer i MIDT kräver resebyråerna att identifieringen ska tas bort från MIDT, eftersom flygbolagen annars kan utöva utpressning mot resebyråerna att minska bokningar med rivaliserande flygbolag.
Textbilden
Textbilden är den bild som resebyråerna använder för att ta fram information från datoriserade bokningssystem.
I vanliga fall är det de datoriserade bokningssystemen som förser resebyråerna med mjukvaran, som en del av affärsavtalet.
Det är viktigt att den information som de datoriserade bokningssystemen ger resebyråerna är neutral och rättvis
Föredragandes kommentarer
Föredraganden ställer sig positiv till kommissionens mål att tillåta flygbolag och datoriserade bokningssystem förhandla om innehåll och priser.
För tillfället leder bristen på konkurrens till högre avgifter inom det datoriserade bokningssystemet.
Efter översynen skulle datoriserade bokningssystem bli tvungna att konkurrera mer aggressivt med varandra om lufttrafikföretag med hjälp av lägre bokningsavgifter och bättre kvalitet på tjänsterna
Förhandlingsfrihet leder i de flesta fall till att lufttrafikföretag ansluter sig till så kallade fullständiga program där de kan erbjuda samtliga priser i de datoriserade bokningssystemen i utbyte mot lägre bokningsavgifter – meddelande från kommissionen, mars 2008. .
Föredraganden är mån om att detta viktiga mål inte rubbas.
I kommissionens förslag ingår också ett ändamålsenligt skydd av personuppgifter, även om de ändringsförslag till kommissionens text som föredraganden föreslår förbättrar rättssäkerheten.
Vissa punkter i kommissionens förslag är dock otillfredsställande.
En undersökning som DG COMP nyligen gjorde visade att Lufthansa inte kan betraktas som ett moderföretag i Amadeus
Air France, Iberia och Lufthansa betraktar sig inte för tillfället som moderföretag.
Inom kort kommer dessa att hävda att de enbart är investerare.
För att svara på den mycket kvistiga frågan om varför flygbolag skulle föredra att vara moderföretag trots de bördor som uppförandekoden medför bör man notera att om flygbolags ekonomiska deltagande i datoriserade bokningssystem i det förgångna kunde motiveras med deras intresse att främja inrättandet av en effektiv kanal för att förmedla uppgifter till marknaden, så kan inte samma motivering användas i dag.
Situationen har ändrats i takt med att de datoriserade bokningssystemen i allt högre grad har blivit självständiga enheter till följd av att ägarandelarna försvunnit.
Det är därför berättigat att dra den slutsatsen att de fördelar som flygbolag förväntar sig av att äga datoriserade bokningssystem har mer att göra med konkurrensfördelar (t.ex. med förmånsvillkor – eller med risken att bli diskriminerad) och strategiska orsaker än enbart med kostnader.
Risken för missbruk är särskilt stor om ett dominerande flygbolag är delägare i ett dominerande datoriserat bokningssystem (t.ex. såsom är fallet med de franska, spanska och tyska marknaderna)
Föredraganden anser att denna punkt ska klargöras och definitionen stramas upp.
Även om man generellt kan säga att ju större ägarandelar man har desto enklare är det att erhålla förmånsvillkor skulle det vara svårt att ange en tröskel för när riskerna för diskriminering ökar
I ett gammalt mål (BAT/Reynolds mot kommissionen – dom av den 17 november 1987, mål 142 och 156/1984) fastställde domstolen följande: ”Även om den omständigheten att ett företag förvärvar aktier i ett konkurrerande företag inte i sig utgör ett konkurrensbegränsande beteende, kan ett sådant förvärv inte desto mindre utgöra ett medel att påverka ifrågavarande företags affärsmässiga uppträdande på ett sådant sätt att konkurrensen begränsas eller snedvrids på [marknaden] (…).
Detta skulle särskilt bli fallet om det investerande företaget genom aktieförvärvet eller genom tilläggsbestämmelser till avtalet erhöll rättslig eller faktisk kontroll över det andra företagets affärsmässiga uppträdande, om avtalet föreskrev att ett affärssamarbete skulle äga rum mellan parterna eller skapade strukturer för att främja ett sådant samarbete” (…)” (punkt 37 – vår fetstil) Se sid.
14 i samma dom. .
I ljuset av detta råder föredraganden utskottet att inte införa ett förbud eller en tröskel för flygbolagens investeringar i datoriserade bokningssystem, utan att i stället införa ett klart och tydligt villkor: Samtliga investeringar som ett flygbolag gör i datoriserade bokningssystem måste vara förenliga med artikel 10.
Detta innebär att moderföretag till datoriserade bokningssystem måste ge andra datoriserade bokningssystem samma prisinformation som sitt eget datoriserade bokningssystem.
Detta innebär att lufttrafikföretag och järnvägstransportföretag utan ägarandelar i datoriserade bokningssystem skyddas mot diskriminering och mot att moderföretag utnyttjar sin dominerande ställning.
Vad gäller MIDT (artikel 7) föreslår föredraganden en kompromiss som skulle göra det möjligt att identifiera resebyråer i MIDT om det finns en överenskommelse om detta mellan resebyrån och det datoriserade bokningssystemet.
Föredraganden föreslår ett kompenseringssystem där resebyrån ersätts för sådan identifiering.
De ovannämnda förslagen ska ses mot bakgrund av det faktum att det rör sig om en sektor med flera inblandade aktörer, i huvudsak lufttrafikföretag och järnvägstransportföretag, datoriserade bokningssystem, resebyråer och konsumenter.
Eftersom kommissionen inte har kommenterat vilka effekter dess konsekvensanalys kan ha på MIDT bör översynen omfatta samtliga element i resedistributionen.
Samtliga beslut att lagstifta om en del av distributionsnätet måste ta i beaktande relevansen för och konsekvenserna på andra områden.
Om identifieringen av resebyråer i MIDT exempelvis begränsas på det sätt som kommissionen föreslår kan det leda till en monopolsituation, eftersom flygbolagen har ett likadant system för datamarknadsföring, t.ex.
Rangordningskriterierna måste vara rättvisa och syfta till att hjälpa resebyrån att erbjuda konsumenten de bästa resealternativen.
Dessa kan ses som ytterligare skyddsåtgärder mot missbruk.
Föredraganden ser detta som en möjlighet för de datoriserade bokningssystemen att utveckla mer användarvänliga och detaljerade sökmöjligheter.
Slutligen har bestämmelser om inspektion av moderföretag införts för att öka insynen i sektorn.
ANNEX
LIST OF STAKEHOLDERS REPRESENTATIVES AND LOBBYSTS
on Code of Conduct Review of Computerised Reservation Systems
The rapporteur would like to make it known that he was contacted during the preparation of his report by the following stakeholder representatives and lobbyists*:
Held meetings with :
Air France
British Airways
Lufthansa
SAS
IATA
Cabinet DN, on behalf Amadeus
APCO, on behalf Sabre Holdings
Travelport
Business Travel Coalition
ECTAA
ITM
Informally involved/written correspondence :
Freshfields
ABTA
BEUC
* Non exhaustive list
YTTRANDE från utskottet för den inre marknaden och konsumentskydd
till utskottet för transport och turism
över förslaget till Europaparlamentets och rådets förordning om en uppförandekod för datoriserade bokningssystem
( KOM(2007)0709 – C6‑0418/2007 – 2007/0243(COD) )
Föredragande:
Wolfgang Bulfon
KORTFATTAD MOTIVERING
Uppförandekoden för datoriserade bokningssystem gäller för researrangörer som bokar flyg- och tågbiljetter via ett datoriserat bokningssystem.
Sedan förordningen trädde i kraft 1989 har den ändrats två gånger, 1993 och 1999.
Den tredje översynen som ska äga rum nu kommer att öka konkurrensen mellan de datoriserade bokningssystemen till följd av att uppförandekoden delvis liberaliserats.
Föredraganden medger att en översyn av den nuvarande uppförandekoden för datoriserade bokningssystem kan leda till större flexibilitet och bättre tjänster.
Den rådande strukturen på den europeiska flygmarknaden, där nationella flygbolag innehar en ledande ställning till följd av den dominans som de har på sina hemmamarknader, har lett till att det dock också råder vissa farhågor för att de dominerande ställningarna på marknaderna kommer att utökas ytterligare.
Genom att flygbolag, datoriserade bokningssystem och resebyråer knyts samman av dominerande marknadsaktörer blir oberoende researrangörer i framtiden tvungna att använda ett visst datoriserat bokningssystem för att få uppgifter om det totala utbudet av priser och tillgång för vissa flygbolag.
Liberaliseringen av uppförandekoden innebär inte enbart ökad konkurrenskraft utan också en ökad splittring av informationen om priser och utbud, som redan nu håller på att utvecklas till följd av att flygbolagen har olika distributionskanaler.
Föredraganden fruktar framför allt att konkurrensen kommer att förvärras för små och medelstora researrangörer, eftersom dessa inte har tillräckligt med resurser för att ingå avtal med flera olika datoriserade bokningssystem, eller att de alternativt måste utnyttja flygbolagens direkta distributionskanaler för att få tillgång till samtliga erbjudanden.
Detta kan leda till att priset för slutkonsumenterna ökar.
Föredraganden stöder de åtgärder som nämns i artikel 10, där det sägs att ett moderföretag måste ge samtliga leverantörer av datoriserade bokningssystem samma information om priser och tillgång (”fullt utbud”), också de leverantörer med vilka de inte ingått något avtal.
Föredraganden stöder helhjärtat kommissionens förslag om att stryka möjligheten att identifiera researrangören i databanden med saluföringsinformation med hjälp av dess IATA‑nummer.
Det är inte tillåtet att i efterhand lägga på avgifter för en bokning via ett datoriserat bokningssystem.
Vad gäller definitionen av de s.k. ”moderföretagen” kräver föredraganden att ett flygbolags eller ett järnvägsföretags direkta eller indirekta deltagande i ett datoriserat bokningssystem ska leda till att bolaget eller företaget klassificeras som ”moderföretag”.
Föredraganden anser att alla former av ägande i ett datoriserat bokningssystem innebär ett visst inflytande.
För att skapa en rättvis konkurrens bör samtliga flygbolag avstå från att delta i datoriserade bokningssystem.
Samtliga flygbolag och järnvägsföretag, som även i fortsättningen vill delta i datoriserade bokningssystem, måste respektera åtgärderna i artikel 3a.
Vid översynen bör man framför allt undersöka hur effektivt förordningen förhindrar diskriminering, hur rättvis konkurrensen är på marknaden för datoriserade bokningssystemstjänster samt effekterna av detta på konsumenternas intressen.
ÄNDRINGSFÖRSLAG
Utskottet för den inre marknaden och konsumentskydd uppmanar utskottet för transport och turism att som ansvarigt utskott infoga följande ändringsförslag i sitt betänkande:
Ändringsförslag
1
Förslag till förordning
Skäl 9a (nytt)
Kommissionens förslag
Ändringsförslag
(9a) Enligt [förordning (…) om gemensamma regler för tillhandahållande av lufttrafiktjänster i gemenskapen] måste lufttrafikföretagen offentliggöra sina priser inklusive alla tillämpliga skatter, avgifter, tilläggsavgifter och avgifter som är oundvikliga och förutsägbara.
De datoriserade bokningssystemens textbilder bör ge information om totalpriser i samma priskategorier för att garantera att resebyråer kan förmedla denna information till sina kunder.
Motivering
Konsumenterna måste få exakta uppgifter om biljettpriserna.
Samtliga aktörer (lufttrafikföretag, innehavare av datoriserade bokningssystem och resebyråer) måste därför öppet redogöra för vad som ingår i biljettpriserna.
Denna bestämmelse är i linje med den pågående omarbetningen av förordningen om gemensamma regler för tillhandahållande av lufttrafiktjänster i gemenskapen.
Ändringsförslag
2
Förslag till förordning
Skäl 11a (nytt)
Kommissionens förslag
Ändringsförslag
(11a) Kommissionen bör regelbundet övervaka hur denna förordning tillämpas, särskilt hur effektivt den förhindrar konkurrenshämmande och diskriminerande praxis på marknaden för distribution av resetjänster via de datoriserade bokningssystemen, särskilt när det finns transportföretag med nära kopplingar till systemleverantörer.
Motivering
Utan att ifrågasätta resultaten från undersökningen om effekterna på moderföretagen bör kommissionen vara uppmärksam och övervaka att konkurrenshämmande praxis förhindras.
Ändringsförslag
3
Förslag till förordning
Skäl 12
Kommissionens förslag
Ändringsförslag
(12) Denna förordning påverkar inte tillämpningen av artiklarna 81 och 82 i fördraget.
(12) Denna förordning påverkar inte tillämpningen av artiklarna 81 och 82 i fördraget.
Denna förordning kompletterar allmänna konkurrensregler som fortfarande är fullt ut tillämpliga på konkurrensbegränsningar såsom överträdelser av kartellagstiftningen eller missbruk av dominerande ställning.
Motivering
Syftet med denna uppförandekod är att bidra till att lufttrafikföretagen åtnjuter rättvisa och neutrala villkor i flygsystemet i de datoriserade bokningssystemen.
Detta är dock inte en isolerad text, utan den kompletterar bestämmelserna i artiklarna 81 och 82.
Ändringsförslag
4
Artikel 2 – led g
Kommissionens förslag
Ändringsförslag
g) moderföretag: ett lufttrafikföretag eller järnvägstransportföretag som direkt eller indirekt, ensamt eller tillsammans med andra, äger eller faktiskt kontrollerar en systemleverantör, liksom varje lufttrafikföretag eller järnvägstransportföretag som det äger eller faktiskt kontrollerar.
g) moderföretag: ett lufttrafikföretag eller järnvägstransportföretag som direkt eller indirekt, ensamt eller tillsammans med andra
– innehar kapitalandelar eller har laglig rätt att nominera personer i företagsledningen, styrelseledamöter, ledamöter i den övervakande styrelsen eller andra ledningsorgan för systemleverantören och
– som erkänts av kommissionen som ett företag som faktiskt kontrollerar en systemleverantör, liksom varje lufttrafikföretag eller järnvägstransportföretag som det äger eller faktiskt kontrollerar.
Kommissionen kan när som helst be ett lufttrafikföretag eller ett järnvägstransportföretag som innehar kapitalandelar i en systemleverantör att lämna kommissionen all information som behövs för att utvärdera dennes eventuella ställning som moderföretag.
Motivering
Kommissionens definition bör preciseras.
Det har inte fastställts någon tröskel för när ett datoriserat bokningssystems deltagande i kapitalet klart och tydligt påverkar datoriserade bokningssystems handelspolitik.
Man bör därför rikta in sig på samtliga företag som innehar kapitalandelar i ett datoriserat bokningssystem och ge kommissionens konkurrensmyndigheter i uppdrag att undersöka vilka företag som effektivt kontrollerar det datoriserade bokningssystemet.
Andra delen av ändringsförslaget innehåller skyldigheter som rör insynen.
Ändringsförslag
5
Kommissionens förslag
Ändringsförslag
1.
Systemleverantören ska via sitt datoriserade bokningssystem tillhandahålla en eller flera primära textbilder för varje enskild transaktion och ska däri inkludera de uppgifter som lämnats in av deltagande transportföretag på ett neutralt och uttömmande sätt som inte är diskriminerande eller partiskt.
Kriterierna för rangordningen av upplysningarna får inte baseras på någon faktor som direkt eller indirekt har samband med transportföretagens identitet och inte tillämpas på ett sätt som diskriminerar något deltagande lufttrafikföretag.
Den eller de primära textbilderna ska vara förenliga med reglerna i bilaga 1.
1.
Systemleverantören ska via sitt datoriserade bokningssystem tillhandahålla en eller flera primära textbilder för varje enskild transaktion och ska däri inkludera de uppgifter som lämnats in av deltagande transportföretag på ett neutralt , öppet och uttömmande sätt som inte är diskriminerande eller partiskt.
Kriterierna för rangordningen av upplysningarna får inte baseras på någon faktor som direkt eller indirekt har samband med transportföretagens identitet och inte tillämpas på ett sätt som diskriminerar något deltagande transportföretag.
Den eller de primära textbilderna ska vara förenliga med reglerna i bilaga 1.
Ändringsförslag
6
Kommissionens förslag
Ändringsförslag
3a.
Då abonnenter tillhandahåller konsumenter information från ett datoriserat bokningssystem ska de informera dem om det slutgiltiga priset för transporttjänsten, inklusive alla tilläggskostnader och serviceavgifter.
Motivering
Åtgärden ökar konsumentens insyn i priset.
Detta gäller för researrangörer på nätet, men även för andra.
Den kompletterar kraven på prisinsyn i den förordning som nyligen antogs om gemensamma regler för tillhandahållande av luftfartstjänster i gemenskapen (det omarbetade tredje paketet) som kräver samma sak av flygbolagen.
Ändringsförslag
7
Artikel 7 − led b
Kommissionens förslag
Ändringsförslag
b) Om uppgifterna har framkommit då en abonnent med säte i Europeiska unionen använt distributionstjänsterna i ett datoriserat bokningssystem, får de inte innehålla någon identifikation, varken direkt eller indirekt, av abonnenten .
b) Deltagande transportföretag ska inte använda uppgifterna för att på ett otillbörligt sätt påverka valet av resebyrå .
Ändringsförslag
8
Förslag till förordning
Artikel 12
Kommissionens förslag
Ändringsförslag
Om kommissionen till följd av ett klagomål eller på eget initiativ konstaterar att denna förordning överträds, får den genom beslut ålägga de berörda företagen eller företagssammanslutningarna att se till att överträdelsen upphör.
Om kommissionen till följd av ett klagomål eller på eget initiativ konstaterar att denna förordning överträds, får den genom beslut ålägga de berörda företagen eller företagssammanslutningarna att se till att överträdelsen upphör.
Utredningar av möjliga överträdelser av denna förordning ska till fullo beakta resultaten av en eventuell undersökning enligt artiklarna 81 och 82 i fördraget.
Motivering
Uppförandekoden för datoriserade bokningssystem ersätter inte utan kompletterar bara de gällande konkurrensreglerna, som fortsätter att vara fullt tillämpliga.
Ändringsförslag
9
Förslag till förordning
Artikel 13
Kommissionens förslag
Ändringsförslag
Kommissionen får när den fullgör de uppgifter som den tilldelas genom denna förordning genom en enkel begäran eller genom beslut begära att företag eller företagssammanslutningar överlämnar alla nödvändiga upplysningar.
Kommissionen får när den fullgör de uppgifter som den tilldelas genom denna förordning genom en enkel begäran eller genom beslut begära att företag eller företagssammanslutningar överlämnar alla nödvändiga upplysningar , inklusive särskilda revisioner, i synnerhet när det gäller frågor som omfattas av artiklarna 4, 7 och 11 i denna förordning .
Motivering
Kommissionen bör ha omfattande befogenheter för att övervaka att uppförandekoden tillämpas på ett bra sätt.
Ändringsförslag
10
Artikel 17 − stycke -1 (nytt)
Kommissionens förslag
Ändringsförslag
Kommissionen ska regelbundet övervaka tillämpningen av denna förordning, vid behov med stöd av särskilda revisioner enligt artikel 13.
Kommissionen ska särskilt undersöka hur effektivt förordningen kan garantera icke ‑diskriminering och rättvis konkurrens på marknaden för datoriserade bokningssystemstjänster.
Ändringsförslag
11
Förslag till förordning
Bilaga I − punkt -1 (ny)
Kommissionens förslag
Ändringsförslag
-1.
Beroende på vad abonnenten väljer ska resealternativen på den primära textbilden rangordnas antingen utifrån biljettpris eller i följande ordning:
a) de direkta resealternativen, rangordnade enligt avgångstid,
b) samtliga övriga resealternativ, rangordnade enligt den totala restiden.
Motivering
Abonnenten bör kunna välja mellan olika alternativ.
Ändringsförslag
12
Förslag till förordning
Bilaga I − punkt 4
Kommissionens förslag
Ändringsförslag
4.
Det ska klart framgå vilka flygningar som innefattar mellanlandningar.
4.
Det ska klart framgå vilka flygningar som innefattar mellanlandningar , och mellanlandningarnas längd måste visas .
Motivering
Konsumenten ska kunna göra det bästa valet som motsvarar hans eller hennes intressen.
ÄRENDETS GÅNG
Titel
Uppförandekod för datoriserade bokningssystem
Referensnummer
KOM(2007)0709 – C6-0418/2007 – 2007/0243(COD)
Ansvarigt utskott
TRAN
Yttrande
Tillkännagivande i kammaren
IMCO
29.11.2007
Föredragande av yttrande
Utnämning
Wolfgang Bulfon
31.1.2008
Behandling i utskott
26.3.2008
6.5.2008
Antagande
27.5.2008
Slutomröstning: resultat
+:
–:
0:
36
1
Slutomröstning: närvarande ledamöter
Cristian Silviu Buşoi, Charlotte Cederschiöld, Gabriela Creţu, Mia De Vits, Janelly Fourtou, Evelyne Gebhardt, Martí Grau i Segú, Małgorzata Handzlik, Malcolm Harbour, Iliana Malinova Iotova, Pierre Jonckheer, Graf Alexander Lambsdorff, Kurt Lechner, Toine Manders, Nickolay Mladenov, Catherine Neris, Zita Pleštinská, Zuzana Roithová, Heide Rühle, Leopold Józef Rutowicz, Salvador Domingo Sanz Palacio, Christel Schaldemose, Andreas Schwab, Marianne Thyssen, Bernadette Vergnaud, Barbara Weiler
Slutomröstning: närvarande suppleanter
Emmanouil Angelakas, Wolfgang Bulfon, Colm Burke, Giovanna Corda, Jan Cremers, Wolf Klinz, Manuel Medina Ortega, Gary Titley
Slutomröstning: närvarande suppleanter (art.
178.2)
YTTRANDE från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
till utskottet för transport och turism
över förslaget till Europaparlamentets och rådets förordning om en uppförandekod för datoriserade bokningssystem
( KOM(2007)0709 – C6‑0418/2007 – 2007/0243(COD) )
Föredragande:
Philip Bradbourn
ÄNDRINGSFÖRSLAG
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor uppmanar utskottet för transport och turism att som ansvarigt utskott infoga följande ändringsförslag i sitt betänkande:
Ändringsförslag
1
Förslag till förordning
Skäl 13b (nytt)
Kommissionens förslag
Ändringsförslag
(13b) Personuppgifter bör endast behandlas i ett datoriserat bokningssystem i samband med bokningar eller utfärdande av biljetter för transporttjänster.
Medlemsstaternas eller tredjelands polismyndigheter bör inte ha rätt till tillgång till personuppgifter i bokningssystemet.
Ändringsförslag
2
Artikel 7 – led b
Kommissionens förslag
Ändringsförslag
b) Om uppgifterna har framkommit då en abonnent med säte i Europeiska unionen använt distributionstjänsterna i ett datoriserat bokningssystem, får de inte innehålla någon identifikation, varken direkt eller indirekt, av abonnenten.
b) Om uppgifterna har framkommit då en abonnent med säte i Europeiska unionen använt distributionstjänsterna i ett datoriserat bokningssystem, får de inte innehålla någon identifikation, varken direkt eller indirekt, av abonnenten , i enlighet med relevant lagstiftning om uppgiftsskydd i medlemsstaterna och EU .
Ändringsförslag
3
Kommissionens förslag
Ändringsförslag
3.
När det rör sig om särskilda kategorier av uppgifter i enlighet med artikel 8 i direktiv 95/46/EG, ska sådana uppgifter endast behandlas om den registrerade har givit sitt uttryckliga medgivande till det.
3.
När det rör sig om särskilda kategorier av uppgifter i enlighet med artikel 8 i direktiv 95/46/EG, ska sådana uppgifter endast behandlas om den registrerade har gett sitt uttryckliga och informerade medgivande till det.
Ändringsförslag
4
Kommissionens förslag
Ändringsförslag
4.
Information som kontrolleras av systemleverantören och som rör identifierbara enskilda bokningar ska lagras offline inom 72 timmar efter det att den sista delen av den enskilda bokningen har avslutats, och den ska förstöras inom tre år.
Det ska endast vara tillåtet att tillgå sådana uppgifter vid faktureringstvister.
4.
Information som kontrolleras av systemleverantören och som rör identifierbara enskilda bokningar ska lagras offline inom 72 timmar efter det att den resa som den enskilda bokningen gäller har avslutats, och den ska förstöras inom tre år.
Det ska endast vara tillåtet att tillgå sådana uppgifter vid faktureringstvister.
Ändringsförslag
5
Kommissionens förslag
Ändringsförslag
5.
Det ska inte vara möjligt att varken direkt eller indirekt identifiera fysiska personer, eller i tillämpliga fall de organisationer eller företag på vars vägnar de agerar, via de uppgifter om saluföring, bokföring och försäljning som ett datoriserat bokningssystem tillgängliggör.
utgår
Ändringsförslag
6
Kommissionens förslag
Ändringsförslag
9a.
Motivering
Det datoriserade bokningssystemet kan fungera som ett globalt gränssnitt för flygbolagen, men också för företag som levererar tjänster till ett visst flygbolag.
Man bör därför anta särskilda säkerhetsbestämmelser för att tydligt skilja på uppgifterna utifrån deras olika funktion.
Ändringsförslag
7
Förslag till förordning
Artikel 13
Kommissionens förslag
Ändringsförslag
Kommissionen får när den fullgör de uppgifter som den tilldelas genom denna förordning genom en enkel begäran eller genom beslut begära att företag eller företagssammanslutningar överlämnar alla nödvändiga upplysningar , särskilt i frågor som omfattas av artiklarna 4, 7 och 11, dock med förbehåll för de strängaste kraven för dataskydd som gäller i den berörda medlemsstaten .
ÄRENDETS GÅNG
Titel
Uppförandekod för datoriserade bokningssystem
Referensnummer
KOM(2007)0709 – C6-0418/2007 – 2007/0243(COD)
Ansvarigt utskott
TRAN
Yttrande
Tillkännagivande i kammaren
LIBE
13.3.2008
Föredragande av yttrande
Utnämning
Philip Bradbourn
27.2.2008
Behandling i utskott
27.3.2008
8.4.2008
6.5.2008
Antagande
6.5.2008
Slutomröstning: resultat
+:
–:
0:
41
Slutomröstning: närvarande ledamöter
Alexander Alvaro, Philip Bradbourn, Mihael Brejc, Kathalijne Maria Buitenweg, Michael Cashman, Giusto Catania, Jean-Marie Cavada, Elly de Groen-Kouwenhoven, Panayiotis Demetriou, Gérard Deprez, Agustín Díaz de Mera García Consuegra, Armando França, Urszula Gacek, Kinga Gál, Roland Gewalt, Jeanine Hennis-Plasschaert, Lívia Járóka, Ewa Klamt, Magda Kósáné Kovács, Stavros Lambrinidis, Henrik Lax, Viktória Mohácsi, Claude Moraes, Martine Roure, Inger Segelström, Csaba Sógor, Vladimir Urutchev, Ioannis Varvitsiotis, Manfred Weber, Tatjana Ždanoka
Slutomröstning: närvarande suppleanter
Edit Bauer, Simon Busuttil, Iliana Malinova Iotova, Sylvia-Yvonne Kaufmann, Marianne Mikko, Bill Newton Dunn, Nicolae Vlad Popa, Rainer Wieland, Stefano Zappalà
Slutomröstning: närvarande suppleanter (art.
178.2)
Emine Bozkurt, Jas Gawronski
ÄRENDETS GÅNG
Titel
Uppförandekod för datoriserade bokningssystem
Referensnummer
KOM(2007)0709 – C6-0418/2007 – 2007/0243(COD)
Framläggande för parlamentet
15.11.2007
Ansvarigt utskott
Tillkännagivande i kammaren
TRAN
29.11.2007
Rådgivande utskott
Tillkännagivande i kammaren
IMCO
29.11.2007
LIBE
13.3.2008
Föredragande
Utnämning
Timothy Kirkhope
9.1.2008
Behandling i utskott
27.2.2008
8.4.2008
28.5.2008
Antagande
29.5.2008
Slutomröstning: resultat
+:
–:
0:
34
1
2
Slutomröstning: närvarande ledamöter
Inés Ayala Sender, Paolo Costa, Arūnas Degutis, Petr Duchoň, Saïd El Khadraoui, Robert Evans, Emanuel Jardim Fernandes, Francesco Ferrari, Brigitte Fouré, Mathieu Grosch, Georg Jarzembowski, Timothy Kirkhope, Sepp Kusstatscher, Jörg Leichtfried, Marian-Jean Marinescu, Erik Meijer, Seán Ó Neachtain, Willi Piecyk, Paweł Bartłomiej Piskorski, Luís Queiró, Reinhard Rack, Brian Simpson
Slutomröstning: närvarande suppleanter
Markus Ferber, Nathalie Griesbeck, Jeanine Hennis-Plasschaert, Aldis Kušķis, Leopold Józef Rutowicz
Slutomröstning: närvarande suppleanter (art.
178.2)
A6-0288/2008
***I
BETÄNKANDE
om förslaget till Europaparlamentets och rådets direktiv om förande av statistik över gods- och passagerarbefordran till sjöss (omarbetning)
(KOM(2007)0859 – C6‑0001/2008 – 2007/0288(COD))
Utskottet för rättsliga frågor
Föredragande:
József Szájer
(Omarbetning – artikel 80a i arbetsordningen)
PE 407.765v02-00
Teckenförklaring
* Samrådsförfarandet
majoritet av de avgivna rösterna
**I Samarbetsförfarandet (första behandlingen)
majoritet av de avgivna rösterna
**II Samarbetsförfarandet (andra behandlingen)
*** Samtyckesförfarandet
majoritet av parlamentets samtliga ledamöter utom i de fall som avses i artiklarna 105, 107, 161 och 300 i EG-fördraget och artikel 7 i EU-fördraget
***I Medbeslutandeförfarandet (första behandlingen)
majoritet av de avgivna rösterna
***II Medbeslutandeförfarandet (andra behandlingen)
majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten
majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
***III Medbeslutandeförfarandet (tredje behandlingen)
majoritet av de avgivna rösterna för att godkänna det gemensamma utkastet
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Parlamentets ändringar markeras med fetkursiv stil .
I samband med ändringsakter ska de delar av en återgiven befintlig rättsakt som inte ändrats av kommissionen, men som parlamentet önskar ändra, markeras med fet stil .
Eventuella strykningar ska i sådana fall markeras enligt följande: [...].
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING............................................................................................................................8
SKRIVELSE FRÅN UTSKOTTET FÖR TRANSPORT OCH TURISM...................................9
BILAGA: YTTRANDE FRÅN DEN RÅDGIVANDE GRUPPEN, SAMMANSATT AV DE JURIDISKA AVDELNINGARNA VID EUROPAPARLAMENTET, RÅDET OCH KOMMISSIONEN 11
ÄRENDETS GÅNG..................................................................................................................13
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till Europaparlamentets och rådets direktiv om förande av statistik över gods- och passagerarbefordran till sjöss (omarbetning)
( KOM(2007)0859 – C6‑0001/2008 – 2007/0288(COD) )
(Medbeslutandeförfarandet – omarbetning)
Europaparlamentet utfärdar denna resolution
– med beaktande av det interinstitutionella avtalet av den 28 november 2001 om en mer strukturerad användning av omarbetningstekniken för rättsakter
EGT C 77, 28.3.2002, s.
1. ,
– med beaktande av artiklarna 80a och 51 i arbetsordningen,
– med beaktande av betänkandet från utskottet för rättsliga frågor och yttrandet från utskottet för transport och turism ( A6‑0288/2008 ), och av följande skäl.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om kommissionen har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
Ändringsförslag
1
Kommissionens förslag
Ändringsförslag
3a.
Kommissionen ska anpassa uppgiftsinsamlingens karakteristika och innehållet i bilagorna I ‑VIII till den ekonomiska och tekniska utvecklingen, om inte en sådan anpassning medför en väsentlig ökning av kostnaderna för medlemsstaterna och/eller en ökning av uppgiftslämnarnas åligganden.
Motivering
Upprepningen av de flesta av dessa delegeringar i artikel 10, särskilt dess inledande mening (”åtgärder som krävs för [direktivets] anpassning till den ekonomiska och tekniska utvecklingen”) kan vara förvirrande och bör därför undvikas.
För att låta förfarandet för ändring av artikel 3 och bilagorna kvarstå inges detta ändringsförslag.
Ändringsförslag
2
Förslag till förordning
Artikel 10
Kommissionens förslag
Ändringsförslag
Artikel 10
utgår
Närmare föreskrifter för genomförandet av detta direktiv, inbegripet åtgärder som krävs för dess anpassning till den ekonomiska och tekniska utvecklingen, skall fastställas, särskilt vad gäller:
a) anpassning av karakteristika för uppgifter som skall insamlas (artikel 3) och för innehållet i bilagorna I-VIII, om inte en sådan anpassning medför en väsentlig ökning av kostnaderna för medlemsstaterna och/eller uppgiftslämnarnas åligganden,
b) den förteckning över hamnar, kodade och indelade efter länder och havskustområden som regelbundet revideras av kommissionen (artikel 4),
c) kraven på noggrannhet (artikel 5),
d) beskrivningen av uppläggningen av uppgiftsinsamlingen och koder för överlämnande av resultat till kommissionen (Eurostat) (artikel 7),
e) sättet för offentliggörande eller spridning av uppgifterna (artikel 9).
Motivering
Upprepningen av de flesta av dessa delegeringar i artikel 10, särskilt dess inledande mening (”åtgärder som krävs för [direktivets] anpassning till den ekonomiska och tekniska utvecklingen”) kan vara förvirrande och bör därför undvikas.
Med tanke på föregående ändringsförslag kan artikel 10 utgå.
MOTIVERING
Rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter
EGT C 203, 17.7.1999, s.
1. ändrades genom rådets beslut 2006/512/EG av den 17 juli 2006
EUT L 200, 22.7.2006, s.
11. .
Genom artikel 5a i det ändrade beslutet 1999/468/EG införs det nya föreskrivande förfarandet med kontroll, som ska tillämpas vid antagande av åtgärder vilka är avsedda att ändra icke väsentliga delar av en grundläggande rättsakt som antagits i enlighet med medbeslutandeförfarandet, inbegripet genom strykning av vissa av dessa delar eller komplettering genom tillägg av nya icke väsentliga delar.
Till följd av en genomgång av befintlig lagstiftning och pågående förfaranden
KOM(2007)0740 . har Europeiska kommissionen lagt fram bland annat detta förslag, som har övergått från att vara en kodifiering till att vara ett förslag till omarbetning så att de ändringar kan införas som krävs för en anpassning till det föreskrivande förfarandet med kontroll.
I sitt beslut av den 12 december 2007 utsåg talmanskonferensen utskottet för rättsliga frågor till ansvarigt utskott, och de specialiserade utskotten till rådgivande utskott, när det gäller denna anpassning till kommittéförfarandet.
Utskottsordförandekonferensen enades den 15 januari 2008 om formerna för samarbetet mellan rättsutskottet och andra berörda utskott.
Med tanke på den föreslagna anpassningen till det föreskrivande förfarandet med kontroll, och efter att ha samrått med det specialiserade utskottet, lägger utskottet för rättsliga frågor fram två ändringsförslag som syftar till att förtydliga kommittébestämmelserna.
När det gäller omarbetningstekniken rekommenderas att man även tar med de tekniska anpassningar som föreslagits av de juridiska avdelningarnas rådgivande grupp.
SKRIVELSE FRÅN UTSKOTTET FÖR TRANSPORT OCH TURISM
Giuseppe Gargani TRAN/D/2008/33600
Ordförande för utskottet för rättsliga frågor
ASP 09E206
Bryssel
Ärende : Förslaget till Europaparlamentets och rådets direktiv om förande av statistik över gods- och passagerarbefordran till sjöss (omarbetning) – ( KOM(2007)0859 - 2007/0288(COD) )
Bäste herr Gargani,
Den 20 maj 2008 behandlade utskottet för transport och turism det ovan nämnda förslaget med anledning av talmanskonferensens beslut av den 12 december 2007 att utse utskottet för rättsliga frågor till ansvarigt utskott för översyn av befintliga rättsakter som ska anpassas till det nya föreskrivande förfarandet med kontroll och för att se till att de specialiserade utskotten associeras och får avge yttranden.
Utskottet för transport och turism rekommenderar enhälligt ert utskott att som ansvarigt utskott godkänna anpassningen med de ändringar (ändringsförslag) som föreslås i bilagan.
Med vänlig hälsning,
Paolo Costa
Bilaga: Sammanställning
Cc: Jarzembowski, föredragande TRAN
Szájer, föredragande JURI
BILAGA
JURI:s kommentarer till kommissionens förslag
Förslag till Europaparlamentets ståndpunkt
Art.
7.2: Inget behov av det föreskrivande förfarandet med kontroll , då ”de tekniska detaljerna beträffande överlämnandet” är av en sådan teknisk karaktär att detta inte kan anses komplettera grundrättsakten.
Art.
9: Inget behov av det föreskrivande förfarandet med kontroll , då ”sättet för offentliggörande eller spridning av statistiska uppgifter” är av en sådan teknisk karaktär att detta inte kan anses komplettera grundrättsakten.
Art.
10, punkterna d och e är överflödiga och bör utgå.
BILAGA: YTTRANDE FRÅN DEN RÅDGIVANDE GRUPPEN, SAMMANSATT AV DE JURIDISKA AVDELNINGARNA VID EUROPAPARLAMENTET, RÅDET OCH KOMMISSIONEN
YTTRANDE
TILL EUROPAPARLAMENTET
RÅDET
KOMMISSIONEN
I enlighet med det interinstitutionella avtalet av den 28 november 2001 om en mer strukturerad användning av omarbetningstekniken för rättsakter, särskilt artikel 9, sammanträdde den rådgivande gruppen, sammansatt av de juridiska avdelningarna vid Europaparlamentet, rådet och kommissionen, den 8 januari 2008 för att bland annat granska det nämnda förslaget som lagts fram av kommissionen.
Vid detta sammanträde
Gruppen förfogade över de engelska, franska och tyska språkversionerna av förslaget och arbetade utifrån den engelska, som var textens originalversion. behandlade gruppen förslaget till Europaparlamentets och rådets direktiv om omarbetning av rådets direktiv 95/46/EG av den 8 december 1995 om förande av statistik över gods- och passagerarbefordran till sjöss och konstaterade enhälligt att de två följande rättelserna hade införts i den befintliga ordalydelsen i de tekniska bilagorna:
1) I bilaga VI hade asterisken efter ordet ” Fiske ” (punkt 41) tagits bort.
2) I bilaga VIII, under uppsättningen uppgifter C1, har man i fotnotens första rad lagt till uppgiften ” 5X ” mellan siffrorna ” 34 ” och ” 51 ”.
Vid behandlingen kunde den rådgivande gruppen därmed enhälligt konstatera att förslaget inte innehåller några betydande ändringar utöver dem som anges.
Gruppen konstaterade vidare att förslaget i fråga om kodifieringen av de bibehållna bestämmelserna med de väsentliga ändringarna endast gäller en kodifiering som inte ändrar sakinnehållet i den text som berörs.
Juridisk rådgivare Juridisk rådgivare Generaldirektör
ÄRENDETS GÅNG
Titel
Förande av statistik över gods- och passagerarbefordran till sjöss (omarbetad version)
Referensnummer
KOM(2007)0859 – C6-0001/2008 – 2007/0288(COD)
Framläggande för parlamentet
21.12.2007
Ansvarigt utskott
Tillkännagivande i kammaren
JURI
19.2.2008
Rådgivande utskott
Tillkännagivande i kammaren
TRAN
19.2.2008
Inget yttrande avges
Beslut
TRAN
22.1.2008
Föredragande
Utnämning
József Szájer
19.12.2007
Antagande
26.6.2008
Slutomröstning: resultat
+:
–:
0:
24
Slutomröstning: närvarande ledamöter
Carlo Casini, Titus Corlăţean, Bert Doorn, Monica Frassoni, Giuseppe Gargani, Neena Gill, Othmar Karas, Piia-Noora Kauppi, Klaus-Heiner Lehne, Hans-Peter Mayer, Manuel Medina Ortega, Hartmut Nassauer, Aloyzas Sakalas, Francesco Enrico Speroni, Diana Wallis, Rainer Wieland, Jaroslav Zvěřina, Tadeusz Zwiefka
Slutomröstning: närvarande suppleanter
A6-0302/2008
BETÄNKANDE
om Bolognaprocessen och studentrörligheten
(2008/2070(INI))
Utskottet för kultur och utbildning
Föredragande:
Doris Pack
PE 404.721v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING............................................................................................................................9
YTTRANDE från budgetutskottet ............................................................................11
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................14
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om Bolognaprocessen och studentrörligheten
( 2008/2070(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av artiklarna 149 och 150 i EG‑fördraget,
– med beaktande av kommissionens meddelande ”Att förverkliga moderniseringsagendan för universiteten – Utbildning, forskning och innovation” ( KOM(2006)0208 ),
– med beaktande av kommissionens meddelande ”Att mobilisera Europas intellektuella resurser: skapa möjligheter för universiteten att lämna sitt fulla bidrag till Lissabonstrategin” ( KOM(2005)0152 ),
– med beaktande av Eurobarometerundersökningen om synen på reformerna av den högre utbildningen, ”Perceptions of Higher Education Reforms”, Europeiska kommissionen, mars 2007,
– med beaktande av sin ståndpunkt vid första behandlingen den 25 september 2007 om förslaget till Europaparlamentets och rådets förordning om framställning och utveckling av statistik om utbildning och livslångt lärande
Antagna texter, P6_TA(2007)0400 . ,
– med beaktande av rådets resolution av den 23 November 2007 om modernisering av universiteten för Europas konkurrenskraft i en global kunskapsekonomi,
– med beaktande av Europeiska rådets slutsatser av den 13–14 mars 2008,
– med beaktande av artikel 45 i arbetsordningen,
– med beaktande av betänkandet från utskottet för kultur och utbildning och yttrandet från budgetutskottet ( A6‑0302/2008 ), och av följande skäl:
A. Bolognaprocessens mål är att skapa ett europeiskt område för högre utbildning senast 2010, vilket inbegriper reformer på området för högre utbildning, avlägsnande av återstående hinder för studenters och lärares rörlighet samt förbättring av den högre utbildningens kvalitet, attraktionskraft och konkurrenskraft i Europa.
B. Studenternas rörlighet och utbildningens kvalitet måste fortsätta att tillhöra de viktigaste aspekterna i Bolognaprocessen.
C. Studentrörligheten ger upphov till nya kulturella, sociala och akademiska värderingar och skapar möjligheter till personlig utveckling, högre akademiska standarder och förbättrad anställbarhet på nationell och internationell nivå.
D. Rörlighet är fortfarande ouppnåeligt för många studenter, forskare och annan personal, i synnerhet i de nya medlemsstaterna och främst på grund av bristen på finansiering, samtidigt som hindren är välkända och har påpekats upprepade gånger av de många berörda parter som har deltagit i diskussionen.
E. Man bör särskilt beakta lämplig finansiering av studenternas lärande, levnadskostnader och rörlighet.
G. Det krävs tillförlitliga statistiska uppgifter om studentrörligheten för att man ska kunna observera, jämföra och utvärdera samt utveckla lämpliga strategier och åtgärder.
H. Erkännandet av informellt och icke‑formellt lärande är hörnstenen i en strategi för livslångt lärande, och vuxenutbildningen är viktig i denna process.
I. Valet att åka utomlands bör inte hindras av administrativa, ekonomiska eller språkliga barriärer.
J. Rörlighet främjar inlärning av främmande språk och förbättrar kommunikationsförmågan generellt.
K. Det är viktigt att snarast reformera och modernisera universiteten med avseende på kvalitet, kursstruktur, innovation och flexibilitet.
M. Olika nationella system för erkännande är ett stort hinder för likabehandling av studenter och för framsteg inom det europeiska området för högre utbildning och på den europeiska arbetsmarknaden.
N. Rörligheten kan försvåras både av att genomgångna kurser inte erkänns fullt ut eller på rätt sätt och av bristande överensstämmelse mellan betyg.
O. Det är brådskande att genomföra, samordna och främja en sammanhållen metod för alla länder som har undertecknat Bolognaprocessen.
Europaparlamentet anser att ökad studentrörlighet och de olika utbildningssystemens kvalitet bör vara en prioritet i samband med fastställandet av Bolognaprocessens viktigaste mål efter 2010.
Europaparlamentet påpekar att man vid genomförandet av Bolognaprocessen särskilt bör eftersträva ett nära och intensivt samarbete och samordning med Europeiska området för forskningsverksamhet.
Studentrörlighet: kvalitet och effektivitet
Reformering av den högre utbildningen och modernisering av universitet en : kvalitet, innovation och flexibilitet
Europaparlamentet upprepar på nytt behovet av ökad dialog över gränserna och utbyte av information och erfarenheter för att underlätta samordning av lärarutbildningen, även för låg- och mellanstadielärare, samt en effektiv och fortlöpande yrkesmässig utveckling.
Finansiering av och investeringar i studentrörlighet och den sociala dimensionen
Kvalitet hos och fullständigt erkännande av examensbevis
Genomförandet av Bolognaprocessen i alla berörda länder
o
o o
MOTIVERING
1.
Bakgrund
Bolognaprocessen, som inleddes 1999, är ett mellanstatligt initiativ som syftar till att senast 2010 skapa ett europeiskt område för högre utbildning.
Grundtanken är att göra det lättare för studenter att välja mellan en mängd olika högkvalitativa kurser och att göra dessa kurser allmänt erkända.
För att kunna uppnå dessa mål finns det i Bolognaprocessen tre prioriterade åtgärdsområden: införandet av ”trestegssystemet” (kandidat, magister och doktor), kvalitetssäkring samt erkännande av kvalifikationer och studieperioder.
Framstegen när det gäller uppnåendet av målen diskuterades vid den offentliga utfrågningen om Bolognaprocessen, som hölls av CULT‑utskottet den 4 oktober 2007.
Den 6 mars 2008 anordnade dessutom PPE‑DE‑gruppen ytterligare en utfrågning om detta ämne (”Higher education: from the Bologna process to educational governance in the EU?"), med Europaparlamentets ledamot Doris Pack som ordförande.
Vid detta tillfälle diskuterades många intressanta slutsatser om Bolognaprocessens effekter på studentrörligheten.
Man tog också upp olika nyckelfrågor, t.ex. vikten av en effektiv ledning av universiteten, den centrala betydelsen av lärarkvalitet och innovativa kursplaner samt de många gemensamma inre och yttre utmaningar som den europeiska högre utbildningen fortfarande måste ta itu med för att förbli konkurrenskraftig och framgångsrik i en alltmer globaliserad värld på 2000‑talet.
Bolognaprocessen drivs framåt genom ett arbetsprogram som får sina riktlinjer från ministerkonferenser som äger rum vartannat år: Prag 2001, Berlin 2003, Bergen 2005, London 2007 och Leuven/Louvaine‑la‑Neuve 2009.
Dessa konferenser organiseras av en uppföljningsgrupp för Bolognaprocessen
Nyckeln till framgång för Bolognasamarbetet är den underliggande partnerskapsmetoden, både när det gäller ledning och genomförande.
I dag förenar processen 46 länder, som alla deltar i det europeiska kulturkonventet och som samarbetar på ett flexibelt sätt och även engagerar internationella organisationer och europeiska föreningar som företräder institutioner för högre utbildning, studenter, personal och arbetsgivare.
Bolognaprocessen är ett bra exempel på europeiskt samarbete, både inom och utanför EU:s ram.
Vi känner alla till att högre utbildning är en grundläggande del i den personliga utvecklingen.
Den stärker den sociala, kulturella och ekonomiska tillväxten, det aktiva medborgarskapet och de etiska värderingarna.
När det gäller EU har emellertid Europeiska kommissionen inget ansvar för den högre utbildningen: det är fortfarande i hög grad en nationell fråga och behörigheten för studiernas innehåll och organisation ligger fortfarande på nationell nivå.
Enligt artikel 149 i Nicefördraget ska dock ”gemenskapen […] bidra till utvecklingen av en utbildning av god kvalitet genom att främja samarbetet mellan medlemsstaterna …”, genom en mängd olika åtgärder som t.ex. främjande av medborgarnas rörlighet, utformande av gemensamma studieprogram, upprättande av nätverk, utbyte av information eller utbildning i EU:s språk.
2.
Föredragandens inställning
Man bör inte glömma bort att rörligheten är ett av de sex främsta målen i Bolognaförklaringen vars signatärer har för avsikt att främja den genom att övervinna hinder mot ett effektivt utövande av den fria rörligheten , då man inte bara tar hänsyn till studenter utan även till lärare, forskare och administrativ personal.
Rörligheten är därför en hörnsten i samband med upprättandet av det europeiska området för högre utbildning, såväl som en av de prioriterade frågorna på dagordningen för 2007–2009.
Föredraganden stöder kommissionens framåtsträvande inställning och dess pågående arbete.
Medlemsstaterna bör stödjas i sina ansträngningar att modernisera och innovativt reformera sina respektive system för högre utbildning, vilket tveklöst krävs om man ska kunna ta itu med globaliseringens utmaningar.
Föredraganden är dock oroad över det tidigare och framtida genomförandet av Bolognaprocessen, eftersom en del av den aktuella utvecklingen i vissa medlemsstater inte går som man hade avsett eller önskat.
Föredraganden anser att det nu, nästan ett decennium efter lanseringen av Bolognaprocessen, är dags för eftertanke och en diskussion om vad man har uppnått och misslyckats med.
Vi bör försöka fastställa hur utbildningssystemen har förändrats som ett resultat av Bolognaprocessen i EU, och även hur denna utveckling och förändring har påverkat kvaliteten på den högre utbildningen i Europa.
Föredraganden vill först och främst understryka att tillgång till högkvalitativ utbildning måste vara möjlig för alla EU‑medborgare, oaktat deras medborgarskap, hemland eller födelseort.
Rörligheten har många positiva effekter, inte bara för den rörliga individen utan även för lärosätena och för samhället som helhet.
Man får inte heller glömma bort dess sociala dimension: rörligheten ger ovärderliga erfarenheter när det gäller akademisk, kulturell och social mångfald.
Den underlättar slutligen nätverkande och samarbete mellan institutionerna för högre utbildning, vilket är helt nödvändigt för en kvalitativ utveckling av den högre utbildningen i Europa och för forskningen.
Föredraganden vill betona och rikta särskild uppmärksamhet mot följande:
1.
Studentrörligheten: kvalitet och effektivitet.
2.
Reformering av den högre utbildningen och modernisering av universiteten: kvalitet, innovation och flexibilitet.
3.
Finansiering av och investeringar i studentrörligheten och den sociala dimensionen.
4.
Examensbevisens kvalitet och fullständiga erkännande.
5.
Genomförande av Bolognaprocessen i alla berörda länder.
Föredraganden erkänner detta mellanstatliga initiativs stora betydelse men betonar att genomförandet är mycket splittrat på nationell nivå.
YTTRANDE från budgetutskottet
till utskottet för kultur och utbildning
över Bolognaprocessen och studentrörligheten
( 2008/2070(INI) )
FÖRSLAG
Budgetutskottet uppmanar utskottet för kultur och utbildning att som ansvarigt utskott införliva följande förslag i sitt förslag till resolution:
Med tanke på det begränsade manöverutrymmet till följd av de små marginaler som återstår i rubrik 1a konstaterar Europaparlamentet att de insatser medlemsstaterna gör inom ramen för det mellanstatliga samarbetet för att förbättra utbildningens kvalitet och konkurrenskraft inom EU, i synnerhet genom att främja rörlighet samt garantera erkännande av kvalifikationer och kvalitetssäkring, är särskilt välkomna.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
6.5.2008
Slutomröstning: resultat
+:
–:
0:
23
Slutomröstning: närvarande ledamöter
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
24.6.2008
Slutomröstning: resultat
+:
–:
0:
30
1
Slutomröstning: närvarande ledamöter
Maria Badia i Cutchet, Katerina Batzeli, Ivo Belet, Giovanni Berlinguer, Nicodim Bulzesc, Marie-Hélène Descamps, Milan Gaľa, Claire Gibault, Vasco Graça Moura, Luis Herrero-Tejedor, Ruth Hieronymi, Mikel Irujo Amezaga, Ramona Nicole Mănescu, Manolis Mavrommatis, Dumitru Oprea, Doris Pack, Zdzisław Zbigniew Podkański, Mihaela Popa, Christa Prets, Pál Schmitt, Hannu Takkula, Helga Trüpel, Thomas Wise, Tomáš Zatloukal
Slutomröstning: närvarande suppleanter
Victor Boştinaru, Mary Honeyball, Ewa Tomaszewska, Cornelis Visser, Jaroslav Zvěřina
A6-0441/2008
***I
BETÄNKANDE
om förslaget till Europaparlamentets och rådets direktiv om leksakers säkerhet
(KOM(2008)0009 – C6‑0039/2008 – 2008/0018(COD))
Utskottet för den inre marknaden och konsumentskydd
Föredragande:
Marianne Thyssen
PE 407.804v02-00
Teckenförklaring
* Samrådsförfarandet
majoritet av de avgivna rösterna
**I Samarbetsförfarandet (första behandlingen)
majoritet av de avgivna rösterna
**II Samarbetsförfarandet (andra behandlingen)
majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten
majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
*** Samtyckesförfarandet
majoritet av parlamentets samtliga ledamöter utom i de fall som avses i artiklarna 105, 107, 161 och 300 i EG-fördraget och artikel 7 i EU-fördraget
***I Medbeslutandeförfarandet (första behandlingen)
majoritet av de avgivna rösterna
***II Medbeslutandeförfarandet (andra behandlingen)
majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten
majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
***III Medbeslutandeförfarandet (tredje behandlingen)
majoritet av de avgivna rösterna för att godkänna det gemensamma utkastet
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Parlamentets ändringar markeras med fetkursiv stil .
I samband med ändringsakter ska de delar av en återgiven befintlig rättsakt som inte ändrats av kommissionen, men som parlamentet önskar ändra, markeras med fet stil .
Eventuella strykningar ska i sådana fall markeras enligt följande: [...].
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................79
YTTRANDE från utskottet för miljö, folkhälsa och livsmedelssäkerhet 83
YTTRANDE från utskottet för industrifrågor, forskning och energi 144
ÄRENDETS GÅNG................................................................................................................163
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till Europaparlamentets och rådets direktiv om leksakers säkerhet
( KOM(2008)0009 – C6‑0039/2008 – 2008/0018(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2008)0009 ),
– med beaktande av artikel 51 i arbetsordningen,
– med beaktande av betänkandet från utskottet för den inre marknaden och konsumentskydd och yttrandena från utskottet för miljö, folkhälsa och livsmedelssäkerhet och utskottet för industrifrågor, forskning och energi ( A6‑0441/2008 ).
Ändringsförslag
1
Förslag till direktiv
Skäl 2
Kommissionens förslag
Ändringsförslag
(2) Direktiv 88/378/EEG bygger på de principer som anges i rådets resolution av den 7 maj 1985 om en ny metod för teknisk harmonisering och standarder.
Där fastställs således endast grundläggande säkerhetskrav för leksaker medan de tekniska detaljerna antas av Europeiska standardiseringsorganisationen (CEN) och Europeiska organisationen för standardisering inom elområdet (Cenelec) i enlighet med Europaparlamentets och rådets direktiv 98/34/EG av den 22 juni 1998 om ett informationsförfarande beträffande tekniska standarder och föreskrifter.
Leksaker som överensstämmer med sådana harmoniserade standarder, till vilka hänvisningar har offentliggjorts i Europeiska unionens officiella tidning, ska förutsättas överensstämma med kraven i direktiv 88/378/EEG.
Dessa grundläggande principer fungerar bra i leksaksbranschen och bör behållas.
(2) Direktiv 88/378/EEG bygger på de principer som anges i rådets resolution av den 7 maj 1985 om en ny metod för teknisk harmonisering och standarder.
Där fastställs således grundläggande säkerhetskrav för leksaker , inklusive särskilda säkerhetskrav för leksakers kemiska, fysikaliska, mekaniska, elektriska och hygieniska egenskaper eller dess brandfarlighet och radioaktivitet .
De tekniska detaljerna antas av Europeiska standardiseringsorganisationen (CEN) och Europeiska organisationen för standardisering inom elområdet (Cenelec) i enlighet med Europaparlamentets och rådets direktiv 98/34/EG av den 22 juni 1998 om ett informationsförfarande beträffande tekniska standarder och föreskrifter.
Leksaker som överensstämmer med sådana harmoniserade standarder, till vilka hänvisningar har offentliggjorts i Europeiska unionens officiella tidning, ska förutsättas överensstämma med kraven i direktiv 88/378/EEG.
Motivering
De grundläggande säkerhetskraven innehåller inte endast de krav som anges i artikel 9 i direktivet, utan även de särskilda säkerhetskrav som anges i bilaga II.
Dessutom är det svårt att låtsas som om saker och ting har fungerat bra i leksaksbranschen, med tanke på de säkerhetsproblem som man nyligen har haft med leksaker.
Ändringsförslag
2
Förslag till direktiv
Skäl 3a (nytt)
Kommissionens förslag
Ändringsförslag
(3a) En annan viktig målsättning med det nya system som inrättas genom detta direktiv är att stimulera och i vissa fall se till att farliga ämnen och material som används i leksaker ersätts med mindre farliga ämnen eller tekniker om det finns lämpliga alternativ som är ekonomiskt och tekniskt genomförbara.
Motivering
Detta ändringsförslag är en anpassning till Reachförordningen (skäl 12).
Ändringsförslag
3
Förslag till direktiv
Skäl 3b (nytt)
Kommissionens förslag
Ändringsförslag
(3b) Försiktighetsprincipen är en princip inom gemenskapslagstiftningen som åter speglas i EG-domstolens avgöranden och är definierad i kommissionens meddelande av den 2 f ebruar i 2000 om försiktighetsprincipen ( KOM(2000)0001 ).
Ändringsförslag
4
Förslag till direktiv
Skäl 8
Kommissionens förslag
Ändringsförslag
(8) Alla ekonomiska aktörer som ingår i leverans- och distributionskedjan bör vidta åtgärder för att se till att de endast tillhandahåller sådana leksaker på marknaden som överensstämmer med den tillämpliga lagstiftningen.
I detta direktiv görs en tydlig och proportionell fördelning av skyldigheterna som svarar mot varje aktörs roll i leverans- och distributionsprocessen.
(8) Alla ekonomiska aktörer som ingår i leverans- och distributionskedjan bör agera så ansvarsfullt och försiktigt som är nödvändigt för att garantera att de leksaker som de släpper ut på marknaden inte har några farliga effekter på barns säkerhet och hälsa vid normal användning och under omständigheter vid användning en som rimligen kan förutses.
De ekonomiska aktörerna bör vidta åtgärder för att se till att de endast tillhandahåller sådana leksaker på marknaden som överensstämmer med den tillämpliga lagstiftningen.
I detta direktiv görs en tydlig och proportionell fördelning av skyldigheterna som svarar mot varje aktörs roll i leverans- och distributionsprocessen.
Motivering
Det räcker inte att påminna de ekonomiska aktörerna om att vidta lämpliga åtgärder, det är också bra att påminna dem om att de är ansvariga.
De måste alltså vara vaksamma så att barns säkerhet och hälsa garanteras.
Hänsyn måste tas till olika typer av användningar.
Ändringsförslag
5
Förslag till direktiv
Skäl 16
Kommissionens förslag
Ändringsförslag
(16) För att barnen ska skyddas mot nyupptäckta risker måste nya grundläggande säkerhetskrav också antas.
Det är särskilt nödvändigt att komplettera och uppdatera bestämmelserna om kemikalier i leksaker.
Dessa bestämmelser bör ange att leksaker bör överensstämma med den allmänna kemikalielagstiftningen, särskilt Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 om registrering, utvärdering, godkännande och begränsning av kemikalier (Reach), inrättande av en europeisk kemikaliemyndighet, ändring av direktiv 1999/45/EG och upphävande av rådets förordning (EEG) nr 793/93 och kommissionens förordning (EG) nr 1488/94 samt rådets direktiv 76/769/EEG och kommissionens direktiv 91/155/EEG, 93/67/EEG, 93/105/EG och 2000/21/EG.
Bestämmelserna bör emellertid också anpassas till barns särskilda behov eftersom de är sårbara konsumenter.
De specifika gränsvärden som anges i direktiv 88/378/EEG för vissa ämnen bör uppdateras mot bakgrund av nya vetenskapliga rön.
(16) För att garantera en hög skyddsnivå för barnen och miljön mot risker , bör ämnen som inger mycket stora betänkligheter, särskilt CMR-ämnen, samt allergiframkallande ämnen och beståndsdelar han teras med yttersta försiktighet .
Nya grundläggande säkerhetskrav måste också antas.
Det är särskilt nödvändigt att komplettera och uppdatera bestämmelserna om kemikalier i leksaker.
Dessa bestämmelser bör ange att leksaker bör överensstämma med den allmänna kemikalielagstiftningen, särskilt Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 om registrering, utvärdering, godkännande och begränsning av kemikalier (Reach), inrättande av en europeisk kemikaliemyndighet, ändring av direktiv 1999/45/EG och upphävande av rådets förordning (EEG) nr 793/93 och kommissionens förordning (EG) nr 1488/94 samt rådets direktiv 76/769/EEG och kommissionens direktiv 91/155/EEG, 93/67/EEG, 93/105/EG och 2000/21/EG.
Bestämmelserna bör emellertid också anpassas till barns särskilda behov eftersom de är sårbara konsumenter.
De specifika gränsvärden som anges i direktiv 88/378/EEG för vissa ämnen bör uppdateras mot bakgrund av nya vetenskapliga rön.
Motivering
Detta ändringsförslag uppmärksammar betydelsen av att ta upp ämnen med särskilt farliga egenskaper.
Detta ändringsförslag är en anpassning till Reachförordningen (skäl 69).
Ändringsförslag
6
Förslag till direktiv
Skäl 17
Kommissionens förslag
Ändringsförslag
(17) De allmänna och särskilda kemikaliekraven i detta direktiv bör syfta till att skydda barns hälsa från farliga ämnen i leksaker, medan miljöproblemen behandlas i övergripande miljölagstiftning som också gäller leksaker, särskilt Europaparlamentets och rådets direktiv 2006/12/EG av den 5 april 2006 om avfall, Europaparlamentets och rådets direktiv 2002/95/EG av den 27 januari 2003 om begränsning av användningen av vissa farliga ämnen i elektriska och elektroniska produkter , Europaparlamentets och rådets direktiv 2002/96/EG av den 27 januari 2003 om avfall som utgörs av eller innehåller elektriska och elektroniska produkter , Europaparlamentets och rådets direktiv 94/62/EG av den 20 december 1994 om förpackningar och förpackningsavfall samt i Europaparlamentets och rådets direktiv 2006/66/EG av den 6 september 2006 om batterier och ackumulatorer och förbrukade batterier och ackumulatorer och om upphävande av direktiv 91/157/EEG.
(17) De allmänna och särskilda kemikaliekraven i detta direktiv bör syfta till att skydda barns hälsa från farliga ämnen i leksaker, medan miljöproblemen behandlas i miljölagstiftning som gäller elektriska och elektroniska leksaker, nämligen Europaparlamentets och rådets direktiv 2002/95/EG av den 27 januari 2003 om begränsning av användningen av vissa farliga ämnen i elektriska och elektroniska produkter och Europaparlamentets och rådets direktiv 2002/96/EG av den 27 januari 2003 om avfall som utgörs av eller innehåller elektriska och elektroniska produkter.
Dessutom regleras miljöfrågor som rör avfall av Europaparlamentets och rådets direktiv 2006/12/EG av den 5 april 2006 om avfall, medan de miljöfrågor som rör förpackningar regleras av Europaparlamentets och rådets direktiv 94/62/EG av den 20 december 1994 om förpackningar och förpackningsavfall, och de miljöfrågor som rör batterier och ackumulatorer regleras av Europaparlamentets och rådets direktiv 2006/66/EG av den 6 september 2006 om batterier och ackumulatorer och förbrukade batterier och ackumulatorer och om upphävande av direktiv 91/157/EEG.
Motivering
Texten ger intrycket av att miljöhänsyn uttryckligen gäller alla leksaker, medan det endast berör elektriska och elektroniska leksaker.
Övergripande lagstiftning är inte uttryckligen tillämplig på leksaker och bör inte klumpas ihop med direktivet om elektriska och elektroniska produkter samt direktivet om avfall som utgörs av eller innehåller elektriska och elektroniska produkter.
Ändringsförslag
7
Förslag till direktiv
Skäl 17a (nytt)
Kommissionens förslag
Ändringsförslag
(17a) Leksaker eller deras delar och förpackningar som rimligen kan förväntas komma i kontakt med livsmedel bör uppfylla kraven i förordning EG) nr 1935/2004 om material och produkter avsedda att komma i kontakt med livsmedel.
Motivering
Bestämmelsen behövs eftersom det hittills inte har varit uppenbart i vissa EU-länder.
Ändringsförslag
8
Förslag till direktiv
Skäl 19
Kommissionens förslag
Ändringsförslag
(19) Eftersom det kan finnas eller komma nya leksaker som medför faror som inte omfattas av särskilda säkerhetskrav i detta direktiv är det nödvändigt att fastställa ett allmänt säkerhetskrav som rättslig grund ör åtgärder mot sådana leksaker.
Leksakernas säkerhet bör då bestämmas utifrån hur de är avsedda att användas eller kan förutses användas med tanke på barns beteende, eftersom de i regel inte är lika försiktiga som vuxna.
(19) Eftersom det kan finnas eller komma nya leksaker som medför faror som inte omfattas av särskilda säkerhetskrav i detta direktiv är det nödvändigt att fastställa ett allmänt säkerhetskrav som rättslig grund för åtgärder mot sådana leksaker.
Leksakernas säkerhet bör då bestämmas utifrån hur de är avsedda att användas eller kan förutses användas med tanke på barns beteende, eftersom de i regel inte är lika försiktiga som vuxna.
Om tillgänglig vetenskaplig bevisning inte medger en sådan bedömning bör medlemsstaterna, särskilt via sina behöriga myndigheter, tillämpa försiktighetsprincipen
Motivering
Det är nödvändigt att tänka på det när leksaken bedöms, så att man tar hänsyn till de olika sätt på vilka barn kan använda en leksak, samtidigt som man utesluter sådana händelser som barn i en viss ålder inte skulle kunna utföra på grund av barnets utvecklingsnivå, fysiska eller intellektuella nivå, etc.
Ändringsförslag
9
Förslag till direktiv
Skäl 21
Kommissionens förslag
Ändringsförslag
(21) CE-märkningen visar att en leksak överensstämmer med kraven och är det synliga resultatet av en hel process av bedömning av överensstämmelse i vid bemärkelse.
Därför bör det i detta direktiv fastställas allmänna principer för hur CE ‑ märkningen ska utformas och användas .
(21) CE-märkningen visar att en leksak överensstämmer med kraven och är det synliga resultatet av en hel process av bedömning av överensstämmelse i vid bemärkelse.
Därför bör det i detta direktiv fastställas hur märkningen ska utformas och anbringas på leksakerna .
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
10
Förslag till direktiv
Skäl 22
Kommissionens förslag
Ändringsförslag
(22) Det är mycket viktigt att klargöra både för tillverkarna och användarna att tillverkaren genom att CE-märka leksaken försäkrar att den överensstämmer med alla tillämpliga krav och tar på sig det fulla ansvaret för detta.
(22) Det är mycket viktigt att klargöra för tillverkarna att tillverkaren genom att CE‑märka leksaken försäkrar att den överensstämmer med alla tillämpliga krav och tar på sig det fulla ansvaret för detta.
Motivering
Endast tillverkaren kan CE-märka.
Tillverkaren måste vara medveten om att användningen av CE-märkningen följer strikta regler, att han är ansvarig och att missbruk är straffbart.
Ändringsförslag
11
Förslag till direktiv
Skäl 34
Kommissionens förslag
Ändringsförslag
(34) Eftersom målen för den föreslagna åtgärden , dvs. att garantera såväl en hög säkerhetsnivå för leksaker som en väl fungerande inre marknad genom att fastställa harmoniserade säkerhetskrav för leksaker och minimikrav för marknadsövervakning, inte i tillräcklig utsträckning kan uppnås av de enskilda medlemsstaterna och de därför, på grund av åtgärdens omfattning och verkningar, bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget.
I enlighet med proportionalitetsprincipen i denna artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå dessa mål.
(34) Eftersom målen för detta direktiv , dvs. att garantera såväl en hög säkerhetsnivå för leksaker för att garantera barns hälsa och säkerhet , som en väl fungerande inre marknad genom att fastställa harmoniserade säkerhetskrav för leksaker och minimikrav för marknadsövervakning, inte i tillräcklig utsträckning kan uppnås av de enskilda medlemsstaterna och de därför, på grund av åtgärdens omfattning och verkningar, bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget.
I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå dessa mål.
Motivering
Man bör påminna om direktivets första målsättning.
Ändringsförslag
12
Förslag till direktiv
Skäl 34a (nytt)
Kommissionens förslag
Ändringsförslag
(34a) För att ge leksakstillverkare och andra ekonomiska aktörer tillräckligt med tid att anpassa sig till de nya kraven är det nödvändigt med en övergångsperiod på två år efter att detta direktiv har trätt i kraft ; en period då leksaker som överensstämmer med direktiv 88/373/EEG kan släppas ut på marknaden.
När det gäller kemiska krav bör denna period vara fyra år , så att det blir möjligt att utveckla de harmoniserade standarder som krävs för efterlevnaden av dessa krav .
Kommissionens förslag
Ändringsförslag
1a.
Detta direktiv baserar sig på principen att tillverkaren är skyldig att se till att leksaker och de eventuella kemikalier som de innehåller varken är skadliga för barns hälsa eller giftiga, i enlighet med bestämmelserna i detta direktiv.
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
1) tillhandahållande på marknaden: varje leverans av en leksak för distribution, förbrukning eller användning på gemenskapsmarknaden i samband med kommersiell verksamhet, mot betalning eller gratis,
1) tillhandahållande på marknaden: varje leverans av en leksak för distribution, förbrukning eller användning på gemenskapsmarknaden i samband med kommersiell verksamhet, mot betalning , utan vinstsyfte eller gratis,
Motivering
Föreningars utdelande av leksaker utan vinstsyfte måste också täckas av detta direktiv.
Ändringsförslag
15
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
(3) tillverkare : varje fysisk eller juridisk person som konstruerar eller tillverkar en leksak eller som låter konstruera eller tillverka en leksak, i eget namn eller under eget varumärke,
(3) tillverkare : varje fysisk eller juridisk person som tillverkar en leksak eller som låter konstruera eller tillverka en leksak och saluför denna leksak , i eget namn eller under eget varumärke,
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
16
Artikel 2 – led 3a (nytt)
Kommissionens förslag
Ändringsförslag
(3a) tillverkarens representant: varje fysisk eller juridisk person som är etablerad i gem enskapen och har tillverkarens skriftliga uppdrag att i dennes ställe utföra vissa uppgifter,
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
17
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
(4) distributör : varje fysisk eller juridisk person i leveranskedjan som tillhandahåller en leksak på marknaden,
(4) distributör : varje fysisk eller juridisk person i leveranskedjan utom tillverkaren eller importören som tillhandahåller en leksak på marknaden,
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
18
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
(7) harmoniserad standard : en standard som i enlighet med artikel 6 i Europaparlamentets och rådets direktiv 98/34/EG antagits av ett europeiskt standardiseringsorgan som upptas i bilaga I till direktiv 98/34/EG ,
(7) harmoniserad standard : en standard som i enlighet med artikel 6 i direktiv 98/34/EG antagits av ett europeiskt standardiseringsorgan som upptas i bilaga I till det direktivet på grundval av en begäran från kommissionen ,
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
19
Artikel 2 – led 7a (nytt)
Kommissionens förslag
Ändringsförslag
(7a) gemenskapslagstiftningen om harmonisering: all gemenskapslagstiftning som harmoniserar villkoren för saluföring av produkter,
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
20
Artikel 2 – led 10a (nytt)
Kommissionens förslag
Ändringsförslag
(10a) organ för bedömning av överensstämmelse: ett organ som bedriver verksamhet inom bedömning av överensstämmelse, bland annat kalibrering, provning, certifiering och inspektion,
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
21
Artikel 2 – led 10b (nytt)
Kommissionens förslag
Ändringsförslag
_____________
1 EUT L 218, 13.8.2008, s.30.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
22
Artikel 2 – led 11a (nytt)
Kommissionens förslag
Ändringsförslag
(11a) doftspel: ett spel vars syfte det är att lära sig känna igen olika dofter eller smaker ,
Ändringsförslag
23
Artikel 2 – led 11b (nytt)
Kommissionens förslag
Ändringsförslag
(11b) kosmetiklåda: en leksak vars syfte det är att hjälpa barn lära sig att tillverka produkter som t.ex. dofter, tvålar, krämer, scha m po , badsalt, läppglans, läppstift, make-up, tandkräm och hårbalsam , som kan innehålla doftämnen eller eteriska oljor,
Ändringsförslag
24
Artikel 2 – led 11c (nytt)
Kommissionens förslag
Ändringsförslag
(11c) smakspel: ett spel där livsmedel kan ingå, t.ex. sötningsmedel, vätskor, pulver eller aromämnen, och som gör det möjligt för barn att tillverka godis eller andra produkter efter recept,
Ändringsförslag
25
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
(13) skada: kroppsskada eller hälsoskada,
(13) skada: kroppsskada eller annan hälsoskada inbegripet långvariga skador ,
Motivering
Denna formulering förtydligar att ”hälsoskada” inbegriper långvariga skador, såsom cancerframkallande effekter och endokrina störningar.
Ändringsförslag
26
Artikel 2 – led 15a (nytt)
Kommissionens förslag
Ändringsförslag
(15a) avsedda för: en förälder eller den som har uppsikt över barnet kan rimligen anta att leksaken är avsedd för barn i den fastställda åldersgruppen.
Varningsmärkning av en produkt som visar att den inte är lämplig för en viss åldersgrupp betraktas inte som ett sätt att få produkten att uppfylla detta direktivs säkerhetskrav.
Motivering
Studier visar att varningstexter på leksaker inte utgör någon effektiv garanti för att grundläggande säkerhetskrav uppfylls.
Framför allt bör en leksak som rimligen kan antas vara avsedd för ett litet barn uppfylla kraven, t.ex. smådelsprovet.
Användningen av formuleringar såsom ”uppenbarligen avsedda för barn under x månader” i detta direktiv bör därför definieras för att förhindra missbruk.
Ändringsförslag
27
Kommissionens förslag
Ändringsförslag
1.
Tillverkarna ska se till att deras leksaker konstrueras och tillverkas i enlighet med de grundläggande säkerhetskraven i artikel 9 och bilaga II.
1.
När tillverkarna släpper ut sina leksaker på marknaden ska de se till att leksakerna har konstruerats och tillverkats i enlighet med de grundläggande säkerhetskraven i artikel 9 och bilaga II.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
28
Kommissionens förslag
Ändringsförslag
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
29
Kommissionens förslag
Ändringsförslag
4.
Tillverkarna ska se till att det finns rutiner som garanterar att serietillverkningen fortsätter att överensstämma med kraven.
Det ska också tas hänsyn till ändringar i produktens konstruktion eller egenskaper och ändringar i de harmoniserade standarder som det hänvisas till vid försäkran om överensstämmelse för en leksak.
4.
Tillverkarna ska se till att det finns rutiner som garanterar att serietillverkningen fortsätter att överensstämma med kraven.
Det ska också tas hänsyn till ändringar i produktens konstruktion eller egenskaper och ändringar i de harmoniserade standarder som det hänvisas till vid försäkran om överensstämmelse för en leksak.
Tillverkarna ska i alla tillämpliga fall utföra slumpvis provning av saluförda leksaker, granska och vid behov registerföra inkomna klagomål samt informera distributörerna om denna övervakning.
När det anses lämpligt med tanke på de risker som en leksak utgör ska tillverkarna, för att skydda konsumenternas hälsa och säkerhet, utföra slumpvis provning av saluförda leksaker, granska och vid behov registerföra inkomna klagomål , leksaker som inte överensstämmer med kraven och återkallanden av leksaker samt informera distributörerna om all sådan övervakning.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
30
Kommissionens förslag
Ändringsförslag
6.
Tillverkarnas ska ange namn och en kontaktadress på leksaken eller, om detta inte är möjligt på grund av leksakens storlek eller art , på förpackningen eller i ett medföljande dokument.
6.
Tillverkarna ska ange namn , sin registrerade handelsbeteckning eller sitt registrerade varumärke och en kontaktadress på leksaken eller, om detta inte är möjligt, på förpackningen eller i ett medföljande dokument.
Den angivna adressen ska ange en enda kontaktpunkt genom vilken tillverkaren kan kontaktas .
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
31
Kommissionens förslag
Ändringsförslag
6a.
Tillverkarna ska se till att leksaken åtföljs av bruksanvisningar och säkerhetsföreskrifter på ett språk som lätt kan förstås av konsumenterna och andra slutanvändare och som bestämts av den berörda medlemsstaten.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
32
Kommissionens förslag
Ändringsförslag
7.
Tillverkare som anser eller har skäl att tro att en leksak som de har släppt ut på marknaden inte överensstämmer med den tillämpliga gemenskapslagstiftningen ska antingen vidta de korrigerande åtgärder som krävs för att få leksaken att överensstämma med kraven eller i förekommande fall dra tillbaka leksaken från marknaden och återkalla den från slutanvändarna .
De ska omedelbart underrätta de nationella myndigheterna i de medlemsstater där de har tillhandahållit leksaken, och lämna detaljerade uppgifter om i synnerhet den bristande överensstämmelsen och de korrigerande åtgärder som vidtagits.
7.
Tillverkare som anser eller har skäl att tro att en leksak som de har släppt ut på marknaden inte överensstämmer med den tillämpliga gemenskapslagstiftningen om harmonisering ska omedelbart vidta de korrigerande åtgärder som krävs för att få leksaken att överensstämma med kraven eller i förekommande fall dra tillbaka leksaken eller återkalla den.
Om leksaken utgör en risk ska tillverkarna dessutom omedelbart underrätta de behöriga nationella myndigheterna i de medlemsstater där de har tillhandahållit leksaken, och lämna detaljerade uppgifter om i synnerhet den bristande överensstämmelsen och de eventuella korrigerande åtgärder som vidtagits.
Tillverkarna ska omedelbart upphöra att släppa ut leksaken på marknaden tills den motsvarar kraven i den tillämpliga gemenskapslagstiftningen .
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
33
Kommissionens förslag
Ändringsförslag
8.
Tillverkarna ska på begäran ge de behöriga nationella myndigheterna all information och dokumentation som behövs för att visa att leksaken överensstämmer med kraven.
De ska på begäran samarbeta med de behöriga myndigheterna i de åtgärder som vidtas för att undvika riskerna med de leksaker som de har släppt ut på marknaden.
8.
Tillverkarna ska på motiverad begäran ge en behörig nationell myndighet all information och dokumentation som behövs för att visa att leksaken överensstämmer med kraven , på ett språk som lätt kan förstås av denna myndighet.
De ska på begäran samarbeta med denna myndighet i de åtgärder som vidtas för att undanröja riskerna med de leksaker som de har släppt ut på marknaden.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
34
Kommissionens förslag
Ändringsförslag
Tillverkarens representant
Skyldigheter för tillverkarens representant
1.
Tillverkarna får genom skriftlig fullmakt utse en fysisk eller juridisk person som är etablerad i gemenskapen (nedan kallad tillverkarens representant) att i deras ställe utföra specificerade uppgifter som följer av tillverkarnas skyldigheter enligt detta direktiv .
1.
Motivering
För att titeln ska överensstämma med artiklarna 3 och 5.
En definition av begreppet ”tillverkarens representant” har lagts till i artikel 2.
Ändringsförslag
35
Kommissionens förslag
Ändringsförslag
2.
2.
Ändringsförslag
36
Kommissionens förslag
Ändringsförslag
3.
Om en tillverkare har utsett en representant ska denne åtminstone
3.
Tillverkarens representant ska utföra de uppgifter som anges i fullmakten från tillverkaren.
Enligt fullmakten ska representanten åtminstone
(a) kunna uppvisa EG-försäkran om överensstämmelse och den tekniska dokumentationen för de nationella myndigheterna under en period på tio år,
(a) kunna uppvisa EG-försäkran om överensstämmelse och den tekniska dokumentationen för de nationella myndigheterna under en period på tio år,
(b) på begäran ge de nationella behöriga myndigheterna all information och dokumentation som behövs för att visa att leksaken överensstämmer med kraven,
(b) på motiverad begäran från en behörig nationell myndighet ge denna myndighet all information och dokumentation som behövs för att visa att en leksak överensstämmer med kraven,
(c) på begäran samarbeta med de behöriga myndigheterna i de åtgärder som vidtas för att undvika riskerna med de leksaker som omfattas av fullmakten.
(c) på begäran samarbeta med de behöriga nationella myndigheterna i de åtgärder som vidtas för att undanröja riskerna med de leksaker som omfattas av fullmakten.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
37
Kommissionens förslag
Ändringsförslag
1.
När importörerna släpper ut en leksak på marknaden ska de iaktta vederbörlig omsorg för att se till att de tillämpliga kraven uppfylls .
1.
Importörerna får endast släppa ut sådana leksaker på gemenskapsmarknaden som uppfyller kraven.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
38
Kommissionens förslag
Ändringsförslag
2.
Innan importörerna släpper ut en leksak på marknaden ska de kontrollera att tillverkaren har utfört bedömningen av överensstämmelse.
2.
Innan importörerna släpper ut en leksak på marknaden ska de se till att tillverkaren har utfört bedömningen av överensstämmelse.
Om en importör anser eller har skäl att tro att en leksak inte överensstämmer med de grundläggande säkerhetskraven i artikel 9 och bilaga II får han eller hon inte släppa ut produkten på marknaden förrän den överensstämmer.
Om leksaken utgör en risk ska importören dessutom underrätta tillverkaren och myndigheterna för marknads kontroll om detta.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
39
Kommissionens förslag
Ändringsförslag
3.
Importörerna ska ange namn och en kontaktadress på leksaken eller, om detta inte är möjligt på grund av leksakens storlek eller art , på förpackningen eller i ett medföljande dokument.
3.
Importörerna ska ange namn , sin registrerade handelsbeteckning eller sitt registrerade varumärke och en kontaktadress på leksaken eller, om detta inte är möjligt, på förpackningen eller i ett medföljande dokument.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
40
Kommissionens förslag
Ändringsförslag
3a.
Importörerna ska se till att leksaken åtföljs av bruksanvisningar och säkerhetsföreskrifter på ett språk som lätt kan förstås av konsumenterna och andra slutanvändare och som bestämts av den berörda medlemsstaten.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
41
Kommissionens förslag
Ändringsförslag
4a.
När det anses lämpligt med tanke på de risker som en leksak utgör ska importörerna, för att skydda konsumenternas hälsa och säkerhet, utföra slumpvis provning av saluförda leksaker, granska och vid behov registerföra inkomna klagomål, leksaker som inte överensstämmer med kraven och återkallanden av leksaker samt informera distributörerna om all sådan övervakning.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
42
Kommissionens förslag
Ändringsförslag
5.
Importörer som anser eller har skäl att tro att en leksak som de har släppt ut på marknaden inte överensstämmer med den tillämpliga gemenskapslagstiftningen ska antingen vidta de korrigerande åtgärder som krävs för att få leksaken att överensstämma med kraven eller i förekommande fall dra tillbaka leksaken från marknaden och återkalla den från slutanvändarna .
De ska omedelbart underrätta de nationella myndigheterna i de medlemsstater där de har tillhandahållit leksaken, och lämna detaljerade uppgifter om i synnerhet den bristande överensstämmelsen och de korrigerande åtgärder som vidtagits.
5.
Importörer som anser eller har skäl att tro att en leksak som de har släppt ut på marknaden inte överensstämmer med den tillämpliga gemenskapslagstiftningen om harmonisering ska omedelbart antingen vidta de korrigerande åtgärder som krävs för att få leksaken att överensstämma med kraven eller i förekommande fall dra tillbaka leksaken eller återkalla den.
Om produkten utgör en risk ska importörerna dessutom omedelbart underrätta de behöriga nationella myndigheterna i de medlemsstater där de har tillhandahållit leksaken, och lämna detaljerade uppgifter om i synnerhet den bristande överensstämmelsen och de eventuella korrigerande åtgärder som vidtagits.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
43
Kommissionens förslag
Ändringsförslag
7.
Importörerna ska på begäran ge de behöriga myndigheterna all information och dokumentation som behövs för att visa att leksaken överensstämmer med kraven.
De ska på begäran samarbeta med de behöriga myndigheterna i de åtgärder som vidtas för att undvika riskerna med de leksaker som de har släppt ut på marknaden.
7.
Importörerna ska på motiverad begäran ge en behörig nationell myndighet all information och dokumentation som behövs för att visa att leksaken överensstämmer med kraven , på ett språk som lätt kan förstås av denna myndighet .
De ska på begäran samarbeta med denna myndighet i de åtgärder som vidtas för att undanröja riskerna med de leksaker som de har släppt ut på marknaden.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
44
Kommissionens förslag
Ändringsförslag
2.
2.
Distributören ska informera tillverkaren eller importören om detta.
Om en distributör anser eller har anledning att tro att leksaken inte överensstämmer med de grundläggande säkerhetskraven i artikel 9 och bilaga II får han eller hon inte tillhandahålla produkten på marknaden förrän den överensstämmer med dessa krav.
Om produkten dessutom innebär en risk ska distributören informera tillverkaren eller importören samt myndigheten för marknadskontroll om detta.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
45
Kommissionens förslag
Ändringsförslag
4.
Distributörer som anser eller har skäl att tro att en leksak som de har tillhandahållit på marknaden inte överensstämmer med den tillämpliga gemenskapslagstiftningen ska antingen vidta de korrigerande åtgärder som krävs för att få leksaken att överensstämma med kraven eller i förekommande fall dra tillbaka leksaken från marknaden och återkalla den från slutanvändarna .
De ska omedelbart underrätta de nationella myndigheterna i de medlemsstater där de har tillhandahållit leksaken, och lämna detaljerade uppgifter om i synnerhet den bristande överensstämmelsen och de korrigerande åtgärder som vidtagits.
4.
Distributörer som anser eller har skäl att tro att en leksak som de har släppt ut på marknaden inte överensstämmer med den tillämpliga gemenskapslagstiftningen om harmonisering ska antingen se till att de korrigerande åtgärder vidtas som krävs för att få leksaken att överensstämma med kraven eller i förekommande fall dra tillbaka leksaken eller återkalla den.
Om leksaken utgör en risk ska distributörerna dessutom omedelbart underrätta de behöriga nationella myndigheterna i de medlemsstater där de har tillhandahållit leksaken, och lämna detaljerade uppgifter om i synnerhet den bristande överensstämmelsen och de eventuella korrigerande åtgärder som vidtagits.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
46
Kommissionens förslag
Ändringsförslag
5.
Distributörerna ska på begäran ge de nationella behöriga myndigheterna den information och dokumentation som behövs för att visa att leksaken överensstämmer med kraven.
De ska på begäran samarbeta med de behöriga myndigheterna när det gäller de åtgärder som vidtas för att undvika riskerna med de leksaker som de tillhandahållit på marknaden.
5.
Distributörerna ska på motiverad begäran från en behörig nationell myndighet ge denna myndighet den information och dokumentation som behövs för att visa att en leksak överensstämmer med kraven, De ska på begäran samarbeta med denna myndighet när det gäller de åtgärder som vidtas för att undanröja riskerna med de leksaker som de har släppt ut på marknaden.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
47
Förslag till direktiv
Artikel 7
Kommissionens förslag
Ändringsförslag
En importör eller distributör som släpper ut en leksak på marknaden i eget namn eller under eget varumärke ska ha samma skyldigheter som tillverkaren har enligt artikel 3.
I detta direktiv ska en importör eller distributör anses som tillverkare och ha samma skyldigheter som tillverkaren har enligt artikel 3 när denne släpper ut en leksak på marknaden i eget namn eller under eget varumärke eller ändrar en leksak på ett sådant sätt att det kan påverka överensstämmelsen med de tillämpliga kraven .
En importör eller distributör som ändrar en leksak på ett sådant sätt att det kan påverka överensstämmelsen med de grundläggande säkerhetskraven i artikel 9 och bilaga II, ska ha samma skyldigheter som tillverkaren har enligt artikel 3 när det gäller dessa ändringar.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
48
Förslag till direktiv
Artikel 8
Kommissionens förslag
Ändringsförslag
De ekonomiska aktörerna ska kunna ange
De ekonomiska aktörerna ska på begäran kunna lämna information till myndigheterna för marknads kontroll under en period på tio år om
(a) alla ekonomiska aktörer som har levererat en leksak till dem,
(a) alla ekonomiska aktörer som har levererat en leksak till dem,
(b) alla ekonomiska aktörer som de har levererat en leksak till.
(b) alla ekonomiska aktörer som de har levererat en leksak till.
I detta syfte ska de ha system och förfaranden för att på begäran kunna lämna denna information till myndigheterna för marknadsövervakning under en period på tio år.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
49
Kommissionens förslag
Ändringsförslag
Hänsyn ska tas till barnets förmåga, och i förekommande fall förmågan hos den som har uppsikt över barnet, att hantera leksaken, särskilt när det gäller leksaker som på grund av sin funktion, storlek och särskilda egenskaper är avsedda för barn under 36 månader.
Hänsyn ska tas till barnets förmåga, och i förekommande fall förmågan hos den som har uppsikt över barnet, att hantera leksaken, särskilt när det gäller leksaker som på grund av sin funktion, storlek och särskilda egenskaper är avsedda för barn under 36 månader.
För särskilda leksakskategorier kan andra åldersgränser fastställas i enlighet med säkerhetskraven i de harmoniserade standarder som avses i artikel 12.
Motivering
Ändringsförslag
50
Kommissionens förslag
Ändringsförslag
Märkningen på leksaken eller förpackningen samt medföljande bruksanvisning ska varna barnet, eller den som har uppsikt över barnet, för faror och skaderisker som leksaken kan medföra vid användning och upplysa om hur dessa risker kan undvikas.
Märkningen på leksaken och/eller förpackningen samt medföljande bruksanvisning ska varna barnet, eller den som har uppsikt över barnet, för faror och relaterade risker som leksaken kan medföra vid användning och upplysa om hur dessa risker kan undvikas.
Motivering
Det är ibland förvirrande för konsumenten med en varningstext om vilken del av leksaken som kan orsaka skada eller om att leksaken innehåller en särskild kemikalie.
Det är inte självklart för konsumenten att varningen ”små bollar” betyder att leksaken kan orsaka kvävning.
Varningstexter bör därför ge användare tydlig information om både faror och relaterade risker som leksaken kan medföra.
Ändringsförslag
51
Kommissionens förslag
Ändringsförslag
3a.
När de behöriga myndigheterna i medlemsstaterna vidtar sådana åtgärder som föreskrivs i detta direktiv, särskilt åtgärderna i artikel 37, ska de ta vederbörlig hänsyn till försiktighetsprincipen.
Ändringsförslag
52
Kommissionens förslag
Ändringsförslag
De varning stexter som avses i del B punkt 1 i bilaga V ska inte användas för leksaker som på grund av funktion, storlek eller utmärkande drag är avsedda för barn under 36 månader.
Ändringsförslag
53
Kommissionens förslag
Ändringsförslag
För de kategorier av leksaker som förtecknas i del B i bilaga V ska de varningstexter som anges där användas.
För de kategorier av leksaker som förtecknas i del B punkterna 2–5 i bilaga V ska de varningstexter som anges där användas med identisk ordalydelse .
Ändringsförslag
54
Kommissionens förslag
Ändringsförslag
2.
Tillverkaren ska på lämpligt sätt förse leksakerna med väl synliga och lättlästa varningstexter , antingen direkt på leksaken, på en etikett på leksaken eller på förpackningen och i tillämpliga fall på den bruksanvisning som medföljer leksaken.
Tillverkaren ska förse leksakerna med väl synliga , korrekta och lättlästa varningstexter direkt på leksaken, på en etikett på leksaken eller på konsumentförpackningen och i tillämpliga fall på den bruksanvisning som medföljer leksaken.
Varningstexterna ska vara på ett språk som konsumenten förstår.
För små leksaker som säljs utan förpackning ska lämpliga varningstexter finnas på själva leksaken.
Varningstexterna ska föregås av ordet ”varning” respektive ”varningar” beroende på omständigheterna .
Ändringsförslag
55
Artikel 10 – punkt 2 - stycke 2
Varningstexter som anger en leksaks säkerhet i samband med den avsedda användaren enligt artikel 10.1 andra stycket, och som är avgörande för köpbeslutet , måste finnas på förpackningen.
Om leksaken köps via Internet ska varningstexten finnas på webbsidan på ett iögonfallande sätt.
Ändringsförslag
56
Kommissionens förslag
Ändringsförslag
1.
När en medlemsstat eller kommissionen anser att en harmoniserad standard inte helt uppfyller de krav som den omfattar och som fastställs i artikel 9 och bilaga II, ska kommissionen eller den berörda medlemsstaten ta upp frågan i den kommitté som inrättats genom artikel 5 i direktiv 98/34/EG (nedan kallad kommittén) och redovisa sina skäl för detta.
Kommittén ska yttra sig utan dröjsmål.
1.
När en medlemsstat eller kommissionen anser att en harmoniserad standard inte helt uppfyller de krav som den omfattar och som fastställs i artikel 9 och bilaga II, ska kommissionen eller den berörda medlemsstaten ta upp frågan i den kommitté som inrättats genom artikel 5 i direktiv 98/34/EG och redovisa sina skäl för detta.
Kommittén ska efter samråd med de berörda europeiska standardiseringsorganen yttra sig utan dröjsmål.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
57
Förslag till direktiv
2.
EG-försäkran om överensstämmelse ska utformas i enlighet med mallen i bilaga III .
2.
Den ska översättas till det eller de språk som begärs av den medlemsstat på vars marknad produkten släpps ut eller görs tillgänglig.
________________
1 EUT L 218, 13.8.2008, s.82.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
58
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
Allmänna principer för CE-märkning
CE-märkning
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
59
Förslag till direktiv
2.
2.
Genom att CE-märka eller låta CE-märka en leksak ska tillverkaren ta ansvar för att den överensstämmer med kraven i detta direktiv.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
60
Kommissionens förslag
Ändringsförslag
4.
CE-märkningen ska vara den enda märkning som intygar att leksaken överensstämmer med de tillämpliga kraven.
utgår
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
61
Kommissionens förslag
Ändringsförslag
5.
Medlemsstaterna får inte införa, eller ska dra tillbaka, hänvisningar i sina nationella bestämmelser till någon annan märkning om överensstämmelse än CE ‑märkningen när det gäller överensstämmelse med bestämmelserna i detta direktiv.
utgår
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
62
Kommissionens förslag
Ändringsförslag
6.
Det ska vara förbjudet att förse leksaker med märkning, symboler och inskriptioner som troligen kan vilseleda tredje part i fråga om CE-märkningens innebörd eller utformning.
Leksakerna får förses med annan märkning, förutsatt att den inte försämrar CE-märkningens synlighet eller läsbarhet eller ändrar dess innebörd.
utgår
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
63
Kommissionens förslag
Ändringsförslag
7.
Icke CE-märkta leksaker som inte överensstämmer med kraven i detta direktiv får visas på handelsmässor och utställningar, förutsatt att det finns en tydlig angivelse om att leksakerna inte uppfyller kraven i detta direktiv och därför varken får säljas eller delas ut gratis.
7.
Icke CE-märkta leksaker eller leksaker som på annat sätt inte överensstämmer med kraven i detta direktiv får visas på handelsmässor och utställningar, förutsatt att det finns en tydlig angivelse om att leksakerna inte uppfyller kraven i detta direktiv och därför varken får säljas eller delas ut gratis.
Motivering
Leksaker på mässor anses inte som utsläppta på den inre marknaden, och inga åtgärder får vidtas mot dem, även om de är farliga.
En skylt måste visa bl.a. importörer och distributörer på mässan att de inte får säljas på marknaden.
De flesta leksaker på mässor är dock EG-märkta.
Den nuvarande formuleringen gör att det är svårt för marknadsövervakare att tvinga utställare att sätta upp en sådan skylt, eftersom leksaker som inte uppfyller kraven och som är EG-märkta inte omfattas.
Ändringsförslag
64
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
Regler och villkor för utformning och placering av CE-märkning
Regler och villkor för utformning och placering av CE-märkning på leksaker
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
65
Kommissionens förslag
Ändringsförslag
1.
CE-märkningen ska bestå av bokstäverna ”CE” i följande utformning:
utgår
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
66
Förslag till direktiv
2.
utgår
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
67
Kommissionens förslag
Ändringsförslag
3.
Om det inte i någon rättsakt föreskrivs särskilda mått ska CE-märkningen vara minst 5 mm hög.
utgår
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
68
Förslag till direktiv
Artikel 17
Kommissionens förslag
Ändringsförslag
Innan tillverkarna släpper ut en leksak på marknaden ska de analysera eventuella faror som beror på leksakens kemiska, fysikaliska, mekaniska, elektriska och hygieniska egenskaper eller dess brandfarlighet och radioaktivitet samt bedöma den möjliga exponeringen för dessa faror.
Innan tillverkarna släpper ut en leksak på marknaden ska de analysera eventuella faror som beror på leksakens kemiska, fysikaliska, mekaniska, elektriska och hygieniska egenskaper eller dess brandfarlighet och radioaktivitet samt bedöma den möjliga exponeringen för dessa faror.
Att det inte finns några uppgifter om tidigare olyckor får inte automatiskt tas till intäkt för en låg risk.
Ändringsförslag
69
Kommissionens förslag
Ändringsförslag
2.
Medlemsstaterna får bestämma att den bedömning och kontroll som avses i punkt 1 ska utföras av deras nationella ackrediteringsorgan i den betydelse som anges i och i enlighet med förordning (EG) nr […].
2.
Medlemsstaterna får bestämma att den bedömning och kontroll som avses i punkt 1 ska utföras av ett nationellt ackrediteringsorgan i den betydelse som anges i och i enlighet med förordning (EG) nr […].
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
70
Kommissionens förslag
Ändringsförslag
3.
Om den anmälande myndigheten delegerar, anlitar en underentreprenör eller på annat sätt överlåter den bedömning, anmälan eller kontroll som avses i punkt 1 till ett organ som inte är offentligt, ska det organ till vilket uppgiften har delegerats, lagts ut på underentreprenad eller på annat sätt överlåtits vara en juridisk person och ha vidtagit åtgärder för att kunna hantera ansvarsskyldighet som kan uppstå i samband med dess verksamhet.
3.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
71
Kommissionens förslag
Ändringsförslag
3a.
Den anmälande myndigheten ska ta det fulla ansvaret för uppgifter som utförs av det organ som avses i punkt 3.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
72
Kommissionens förslag
Ändringsförslag
3b.
Den anmälande myndigheten ska etablera rapporterings ställen för säkerhetsanmälningar dit konsumenter och människor som arbetar med barn kan anmäla leksaker som inte följer bestämmelserna eller olyckor som är relaterade till användningen av en leksak.
Motivering
Genom att sätta upp ställen för säkerhetsanmälningar i medlemsstaterna skulle man ge konsumenterna inflytande och underlätta direkt kommunikation med tillverkare och producenter ifall det finns problem med en särskild produkt.
Tillverkare och producenter skulle då kunna reagera mer direkt på konsumenternas krav.
Ändringsförslag
73
Kommissionens förslag
Ändringsförslag
1.
Den anmälande myndigheten ska uppfylla kraven i punkterna 2–7.
utgår
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
74
Kommissionens förslag
Ändringsförslag
5.
Den anmälande myndigheten får inte erbjuda eller utföra sådan verksamhet som utförs av organet för bedömning av överensstämmelse och får heller inte erbjuda eller utföra konsultverksamhet.
5.
Den anmälande myndigheten får inte erbjuda eller utföra sådan verksamhet som utförs av organet för bedömning av överensstämmelse och får heller inte erbjuda eller utföra konsultverksamhet på kommersiell eller konkurrensmässig grund .
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
75
Kommissionens förslag
Ändringsförslag
6.
Den anmälande myndigheten ska ha rutiner som säkerställer att den information som erhållits behandlas konfidentiellt.
6.
Den anmälande myndigheten ska säkerställa att den information som den erhåller behandlas konfidentiellt.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
76
Kommissionens förslag
Ändringsförslag
Medlemsstaterna ska informera kommissionen och de andra medlemsstaterna om sina nationella förfaranden för bedömning och anmälan av organ för bedömning av överensstämmelse och för kontroll av anmälda organ samt om eventuella ändringar.
Medlemsstaterna ska informera kommissionen om sina förfaranden för bedömning och anmälan av organ för bedömning av överensstämmelse och för kontroll av anmälda organ samt om eventuella ändringar.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
77
Kommissionens förslag
Ändringsförslag
3.
Organet för bedömning av överensstämmelse ska vara oberoende av den organisation eller produkt som den bedömer.
3.
Organet för bedömning av överensstämmelse ska vara oberoende av den organisation eller produkt som den bedömer.
Ett organ som tillhör en företags- eller branschsammanslutning där företag ingår som deltar i konstruktion, tillverkning, leverans, montering, användning eller underhåll av de leksaker som det bedömer kan, under förutsättning att dess oberoende och frånvaro av varje intressekonflikt visas, betraktas som ett sådant organ.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
78
Kommissionens förslag
Ändringsförslag
4.
Organet för bedömning av överensstämmelse, dess högsta ledning och den personal som ansvarar för att bedömningen av överensstämmelse görs får inte utgöras av den som konstruerar, tillverkar, levererar, installerar, köper, äger, använder eller underhåller de produkter som bedöms och inte heller av den som företräder någon av dessa parter.
De får varken delta direkt i konstruktion, tillverkning, marknadsföring, installation, användning eller underhåll av dessa produkter eller företräda parter som bedriver sådan verksamhet.
4.
Organet för bedömning av överensstämmelse, dess högsta ledning och den personal som ansvarar för att bedömningen av överensstämmelse görs får inte utgöras av den som konstruerar, tillverkar, levererar, installerar, köper, äger, använder eller underhåller de leksaker som bedöms och inte heller av den som företräder någon av dessa parter.
Detta får inte utesluta sådan användning av bedömda leksaker som krävs för det arbete som utförs av organet för bedömning av överensstämmelse, eller produkternas användning för personliga ändamål.
Organet för bedömning av överensstämmelse, dess högsta ledning och den personal som ansvarar för att bedömningen av överensstämmelse görs får inte delta direkt i konstruktion, tillverkning, marknadsföring, installation, användning eller underhåll av dessa leksaker eller företräda parter som bedriver sådan verksamhet.
De får inte delta i någon verksamhet som kan påverka deras objektivitet och integritet i samband med den bedömning av överensstämmelse för vilken de har anmälts.
Detta ska särskilt gälla för konsultverksamhet.
De får inte utföra konsultverksamhet som har anknytning till den bedömning av överensstämmelse för vilken de har anmälts eller till de produkter som ska släppas ut på gemenskapsmarknaden .
Detta ska inte utesluta utbyte av teknisk information mellan tillverkaren och organet för bedömning av överensstämmelse eller användning av bedömda produkter som är nödvändiga för organets arbete.
Organet för bedömning av överensstämmelse ska se till att dess dotterbolags eller underentreprenörers verksamhet inte påverkar sekretessen, objektiviteten och opartiskheten i dess bedömningar av överensstämmelse.
Organet för bedömning av överensstämmelse ska se till att dess dotterbolags eller underentreprenörers verksamhet inte påverkar sekretessen, objektiviteten eller opartiskheten i dess bedömningar av överensstämmelse.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
79
Kommissionens förslag
Ändringsförslag
6.
Organet för bedömning av överensstämmelse ska kunna utföra alla de uppgifter avseende bedömning av överensstämmelse som fastställs i artikel 19 för ett sådant organ och för vilka det har anmälts, oavsett om dessa uppgifter utförs av organet för bedömning av överensstämmelse eller för dess räkning och under dess ansvar.
6.
Organet för bedömning av överensstämmelse ska kunna utföra alla de uppgifter avseende bedömning av överensstämmelse som fastställs i artikel 19 för organet och för vilka det har anmälts, oavsett om dessa uppgifter utförs av organet för bedömning av överensstämmelse eller för dess räkning och under dess ansvar.
Vid alla tidpunkter, vid varje bedömning av överensstämmelse och för varje typ eller kategori av produkter för vilka det har anmälts ska organet för bedömning av överensstämmelse ha erforderlig personal med teknisk kunskap och tillräcklig erfarenhet för att utföra bedömningen av överensstämmelse.
Det ska ha de nödvändiga medlen för att korrekt kunna utföra de tekniska och administrativa uppgifterna i samband med bedömningen av överensstämmelse och det ska ha tillgång till den utrustning och de faciliteter som är nödvändiga.
Vid alla tidpunkter, vid varje bedömning av överensstämmelse och för varje typ eller kategori av produkter för vilka det har anmälts ska organet för bedömning av överensstämmelse ha erforderlig
a) personal med teknisk kunskap och tillräcklig erfarenhet för att utföra bedömningen av överensstämmelse ,
c) förfaranden som gör det möjligt för organet att utöva sin verksamhet med hänsyn till företagens storlek, bransch och struktur, den berörda produktteknikens komplexitet och produktionsprocessens seriemässiga karaktär.
Det ska ha de nödvändiga medlen för att korrekt kunna utföra de tekniska och administrativa uppgifterna i samband med bedömningen av överensstämmelse och det ska ha tillgång till den utrustning och de faciliteter som är nödvändiga.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
80
Kommissionens förslag
Ändringsförslag
(c) kännedom och insikt om de grundläggande kraven, de tillämpliga harmoniserade standarderna och de relevanta bestämmelserna i gemenskapslagstiftningen och de relevanta tillämpningsföreskrifterna,
(c) kännedom och insikt om de grundläggande kraven, de tillämpliga harmoniserade standarderna och de relevanta bestämmelserna i gemenskapslagstiftningen om harmonisering och tillämpningsföreskrifterna,
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
81
Kommissionens förslag
Ändringsförslag
11.
Organet för bedömning av överensstämmelse ska delta i, eller se till att dess bedömningspersonal känner till, det relevanta standardiseringsarbetet och det arbete som utförs i samordningsgruppen för anmälda organ, som inrättats i enlighet med artikel 36 , och det ska som generella riktlinjer använda de administrativa beslut och dokument gruppens arbete har resulterat i.
11.
Organet för bedömning av överensstämmelse ska delta i, eller se till att dess bedömningspersonal känner till, det relevanta standardiseringsarbetet och det arbete som utförs i samordningsgruppen för anmälda organ, som inrättats i enlighet med den relevanta gemenskapslagstiftningen om harmonisering , och det ska som generella riktlinjer använda de administrativa beslut och dokument gruppens arbete har resulterat i.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
82
Förslag till direktiv
Artikel 26
Kommissionens förslag
Ändringsförslag
Ett organ för bedömning av överensstämmelse som kan visa att det uppfyller kriterierna i de harmoniserade standarderna, till vilka hänvisningar har offentliggjorts i Europeiska unionens officiella tidning, ska förutsättas uppfylla kraven i artikel 25.
Ett organ för bedömning av överensstämmelse som visar att det uppfyller kriterierna i de relevanta harmoniserade standarderna eller delar av dessa , till vilka hänvisningar har offentliggjorts i Europeiska unionens officiella tidning, ska förutsättas uppfylla kraven i artikel 25 i den utsträckning som de tillämpliga harmoniserade standarderna täcker dessa krav .
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
83
Förslag till direktiv
Artikel 26a (ny)
Kommissionens förslag
Ändringsförslag
Artikel 26a
Formell invändning mot en harmoniserad standard
Om en medlemsstat eller kommissionen har en formell invändning mot de harmoniserade standarder som avses i artikel 26 ska bestämmelserna i artikel 13 gälla.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
84
Kommissionens förslag
Ändringsförslag
1.
Om organet för bedömning av överensstämmelse lägger ut specifika uppgifter med anknytning till bedömningen av överensstämmelse på underentreprenad eller anlitar ett dotterbolag, ska det se till att underentreprenören eller dotterbolaget uppfyller kraven i artikel 25.
1.
Om det anmälda organet lägger ut specifika uppgifter med anknytning till bedömningen av överensstämmelse på underentreprenad eller anlitar ett dotterbolag, ska det se till att underentreprenören eller dotterbolaget uppfyller kraven i artikel 25 och informera den anmälande myndigheten i enlighet härmed .
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
85
Kommissionens förslag
Ändringsförslag
2.
Organet för bedömning av överensstämmelse ska ta det fulla ansvaret för underentreprenörernas eller dotterbolagens uppgifter, oavsett var de är etablerade.
2.
Det anmälda organet ska ta det fulla ansvaret för underentreprenörernas eller dotterbolagens uppgifter, oavsett var de är etablerade.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
86
Kommissionens förslag
Ändringsförslag
4.
Organet för bedömning av överensstämmelse ska se till att de nationella myndigheterna har tillgång till de relevanta dokumenten rörande bedömningen av underentreprenörens eller dotterbolagets kvalifikationer och det arbete som underentreprenören eller dotterbolaget har utfört i enlighet med artikel 19.
4.
Det anmälda organet ska se till att den anmälande myndigheten har tillgång till de relevanta dokumenten rörande bedömningen av underentreprenörens eller dotterbolagets kvalifikationer och det arbete som dessa har utfört i enlighet med artikel 19.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
87
Kommissionens förslag
Ändringsförslag
4.
4.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
88
Kommissionens förslag
Ändringsförslag
5.
Det berörda organet får fungera som anmält organ endast om kommissionen och de andra medlemsstaterna inte har rest invändningar inom två månader efter anmälan.
5.
Det berörda organet får fungera som anmält organ endast om kommissionen eller de andra medlemsstaterna inte har rest invändningar inom två veckor efter en anmälan, om ett ackrediteringsintyg används, och inom två månader efter en anmälan , om ackreditering inte används .
Endast ett sådant organ ska anses vara ett anmält organ i enlighet med detta direktiv.
Endast ett sådant organ ska anses vara ett anmält organ i enlighet med detta direktiv.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
89
Kommissionens förslag
Ändringsförslag
1.
Om en anmälande myndighet har konstaterat eller har informerats om att ett anmält organ inte längre uppfyller de krav som avses i artikel 25 eller att det underlåter att fullgöra sina skyldigheter, ska myndigheten i förekommande fall belägga anmälan med restriktioner eller återkalla den tillfälligt eller slutgiltigt.
Den ska omedelbart underrätta kommissionen och de andra medlemsstaterna om detta.
1.
Om en anmälande myndighet har konstaterat eller har informerats om att ett anmält organ inte längre uppfyller de krav som fastställs i artikel 25 eller att det underlåter att fullgöra sina skyldigheter, ska myndigheten i förekommande fall belägga anmälan med restriktioner eller återkalla den tillfälligt eller slutgiltigt , där åtgärdens omfattning beror på hur allvarlig underlåtenheten att uppfylla dessa krav eller fullgöra dessa skyldigheter är .
Den ska omedelbart underrätta kommissionen och de andra medlemsstaterna om detta.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
90
Kommissionens förslag
Ändringsförslag
3.
Kommissionen ska se till att all information som erhållits i samband med undersökningarna behandlas konfidentiellt.
3.
Kommissionen ska se till att all känslig information som erhållits i samband med undersökningarna behandlas konfidentiellt.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
91
Kommissionens förslag
Ändringsförslag
2.
Bedömningarna av överensstämmelse ska vara proportionella så att de ekonomiska aktörerna inte belastas i onödan , och man ska särskilt ta hänsyn till företagens storlek och till hur komplex produkttekniken är .
2.
Bedömningarna av överensstämmelse ska vara proportionella så att de ekonomiska aktörerna inte belastas i onödan .
Organen för bedömning av överensstämmelse ska utöva sin verksamhet med hänsyn till företagens storlek , bransch och struktur, den berörda produktteknikens komplexitet och produktionsprocessens seriemässiga karaktär .
Samtidigt ska de dock respektera den noggrannhet och den skyddsnivå som krävs för att leksaken ska överensstämma med bestämmelserna i detta direktiv.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
92
Kommissionens förslag
Ändringsförslag
(c) Begäran om information från myndigheterna för marknadsövervakning .
(c) Begäran om information om bedömningar av överensstämmelse från myndigheterna för marknads kontroll .
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
93
Kommissionens förslag
Ändringsförslag
Medlemsstaterna ska se till att de organ som de har anmält deltar i gruppens arbete.
Medlemsstaterna ska se till att de organ som de har anmält deltar i gruppens eller gruppernas arbete , direkt eller genom ombud .
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
94
Förslag till direktiv
Artikel 37
Kommissionens förslag
Ändringsförslag
Medlemsstaterna ska organisera och genomföra övervakning av leksaker som släpps ut på marknaden i enlighet med artiklarna 6, 8 och 9 i direktiv 2001/95/EG .
Förutom de bestämmelserna gäller artiklarna 38, 39 och 40 i det här direktivet.
Medlemsstaterna ska organisera och genomföra övervakning av leksaker som släpps ut på marknaden i enlighet med artiklarna 15 till 29 i förordning (EG) nr 765/2008 .
Förutom de bestämmelserna gäller artikel 39 i det här direktivet.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
95
Förslag till direktiv
Artikel 38
Kommissionens förslag
Ändringsförslag
Artikel 38
utgår
Marknadsövervakningsmyndigheternas befogenhet
1.
Marknadsövervakningsmyndigheterna får av de berörda ekonomiska aktörerna begära all information som de bedömer nödvändig för en effektiv marknadsövervakning, inklusive den tekniska dokumentation som avses i artikel 20.
2.
Marknadsövervakningsmyndigheterna får be ett anmält organ att tillhandahålla information om alla EG-typintyg som det organet har utfärdat eller återkallat samt information om avslag på ansökan om EG-typintyg, inklusive provningsrapporterna och den tekniska dokumentationen.
3.
Marknadsövervakningsmyndigheterna ska ha tillträde till de berörda ekonomiska aktörernas lokaler om det är nödvändigt för att kunna övervaka leksakerna i enlighet med artikel 37.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
96
Artikel 39 – punkt -1a (ny)
Kommissionens förslag
Ändringsförslag
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
97
Förslag till direktiv
Artikel 40
Kommissionens förslag
Ändringsförslag
Artikel 40
utgår
Samarbete om marknadsövervakning
1.
Medlemsstaterna ska säkerställa effektivt samarbete och informationsutbyte i alla frågor som gäller leksaker som utgör en risk, dels mellan sina marknadsövervakningsmyndigheter och myndigheterna i andra medlemsstater, dels mellan sina egna myndigheter och kommissionen och berörda gemenskapsorgan.
2.
För de syften som avses i punkt 1 ska marknadsövervakningsmyndigheterna i en medlemsstat på begäran bistå motsvarande myndigheter i en annan medlemsstat genom att tillhandhålla information eller dokumentation, utföra lämpliga undersökningar eller åtgärder eller delta i undersökningar som inletts i en annan medlemsstat.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
98
Kommissionens förslag
Ändringsförslag
1.
Om en medlemsstats myndigheter för marknadsövervakning har vidtagit åtgärder enligt artikel 12 i direktiv 2001/95/EG eller om de har tillräckliga skäl att anta att en leksak som omfattas av det här direktivet utgör en risk för människors hälsa eller säkerhet, ska de tillsammans med de berörda ekonomiska aktörerna utvärdera leksaken med avseende på alla de krav som fastställs i det här direktivet.
1.
Om en medlemsstats myndigheter för marknads kontroll har vidtagit åtgärder enligt artikel 20 i förordning (EG) nr 756/2008 , eller om de har tillräckliga skäl att anta att en leksak som omfattas av det här direktivet utgör en risk för människors hälsa eller säkerhet eller andra aspekter av skydd i allmänhetens intresse som omfattas av detta direktiv , ska de utvärdera leksaken med avseende på alla de krav som fastställs i det här direktivet.
De berörda ekonomiska aktörerna ska samarbeta i den utsträckning som behövs med myndigheterna för marknads kontroll .
Om myndigheterna för marknadsövervakning vid utvärderingen konstaterar att en leksak inte uppfyller kraven i detta direktiv ska de ålägga de berörda ekonomiska aktörerna att vidta lämpliga korrigerande åtgärder för att leksaken ska uppfylla dessa krav eller dra tillbaka leksaken från marknaden eller återkalla den inom en rimlig tid som de fastställer i förhållande till typen av risk.
Om myndigheterna för marknads kontroll vid utvärderingen konstaterar att en leksak inte uppfyller kraven i detta direktiv ska de utan dröjsmål ålägga de berörda ekonomiska aktörerna att vidta lämpliga korrigerande åtgärder för att leksaken ska uppfylla dessa krav eller dra tillbaka leksaken från marknaden eller återkalla den inom en rimlig tid som de fastställer i förhållande till typen av risk.
Myndigheterna för marknads kontroll ska informera det relevanta anmälda organet om detta.
Artikel 21 i förordning (EG) nr 765/2008 ska gälla för de åtgärder som avses i andra stycke t i denna punkt .
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
99
Kommissionens förslag
Ändringsförslag
3.
De ekonomiska aktörerna ska se till att det vidtas korrigerande åtgärder i fråga om alla berörda leksaker som de har tillhandahållit på gemenskapsmarknaden.
3.
De ekonomiska aktörerna ska se till att alla lämpliga korrigerande åtgärder vidtas i fråga om alla berörda leksaker som de har tillhandahållit på gemenskapsmarknaden.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
100
Kommissionens förslag
Ändringsförslag
5.
I den information som avses i punkt 4 ska alla tillgängliga uppgifter ingå, särskilt de uppgifter som krävs för att kunna identifiera den leksak som inte uppfyller kraven, dess ursprung, den risk leksaken utgör, vilken typ av nationell åtgärd som vidtagits och dess giltighetstid.
Myndigheterna för marknadsövervakning ska särskilt ange om den bristande överensstämmelsen beror på
5.
I den information som avses i punkt 4 ska alla tillgängliga uppgifter ingå, särskilt de uppgifter som krävs för att kunna identifiera den leksak som inte uppfyller kraven, dess ursprung, typ av påstådd bristande överensstämmelse och den risk leksaken utgör, vilken typ av nationell a åtgärd er som vidtagits och de ra s giltighetstid samt de argument som framförts av den berörda ekonomiska aktören .
Myndigheterna för marknads kontroll ska särskilt ange om den bristande överensstämmelsen beror på
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
101
Kommissionens förslag
Ändringsförslag
7a.
Medlemsstaterna ska se till att lämpliga restriktiva åtgärder vidtas i fråga om den berörda leksaken, till exempel att leksaken utan dröjsmål återkallas från marknaden.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
102
Kommissionens förslag
Ändringsförslag
3.
3.
Kommittén ska efter samråd med det berörda europeiska standardiseringsorganet eller de berörda europeiska standardiseringsorganen yttra sig utan dröjsmål.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
103
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
104
Kommissionens förslag
Ändringsförslag
da) Den tekniska dokumentationen är antingen inte tillgänglig eller ofullständig.
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
105
Kommissionens förslag
Ändringsförslag
1.
Kommissionen kan ändra följande bestämmelser i syfte att anpassa dem till den tekniska och vetenskapliga utvecklingen:
1.
Kommissionen kan ändra följande bestämmelser i syfte att anpassa dem till den tekniska , vetenskapliga och praktiska utvecklingen:
-a) Bilaga I:
(a) Punkterna 7 och 8 i del III i bilaga II.
(a) Punkterna 7 och 8 i del III i bilaga II.
(b) Bilaga V.
(b) Bilaga V.
Motivering
Denna artikel berör doftämnen och tungmetaller (samt varningstexter).
Ändringsförslag
106
Kommissionens förslag
Ändringsförslag
(Berör inte den svenska versionen.)
Ändringsförslag
107
Kommissionens förslag
Ändringsförslag
2.
Kommissionen får besluta att ämnen eller preparat som enligt bilaga I till direktiv 67/548/EEG klassificerats som cancerframkallande, mutagena eller reproduktionstoxiska i kategori 1, 2 eller 3 får användas i leksaker.
2.
Kommissionen får besluta att ämnen eller preparat som enligt bilaga I till direktiv 67/548/EEG klassificerats som cancerframkallande, mutagena eller reproduktionstoxiska i kategori 1, 2 eller 3 får ingå i leksaker.
Motivering
Byter ut ”användas” till ”ingå”.
Direktivet blir på så sätt tydligare.
Det blir också tydligare att det är själva utsläppandet av en leksak på marknaden som regleras (oavsett var leksaken tillverkas) och inte tillverkningen av leksaken.
Genom den andra ändringen klargörs endast den vetenskapliga kommitténs deltagande i direktivet, på samma sätt som i bilagan om kemikalier.
Ändringsförslag
108
Förslag till direktiv
Artikel 52
Kommissionens förslag
Ändringsförslag
Medlemsstaterna får inte förhindra att leksaker som överensstämmer med direktiv 88/378/EEG och som släpptes ut på marknaden innan det här direktivet trädde i kraft eller under de första två åren efter ikraftträdandet görs tillgängliga på marknaden.
2.
Med avvikelse från punkt 1 får medlemsstaterna inte hindra att leksaker som uppfyller kraven i detta direktiv görs tillgängliga på marknaden, med undantag av kraven i del III i bilaga II, under förutsättning att de leksaker som inte uppfyller kraven i del III i bilaga II i detta direktiv uppfyller kraven i del II avsnitt 3 i bilaga II till d ire k tiv 88/378/EE G och släpptes ut på marknaden inom fyra år efter att det direktivet trädde i kraft .
Motivering
Syftet med ändringsförslaget är att klargöra dels att det nya direktivet inte har retroaktiv effekt, dels att den minsta övergångsperioden på två år måste respekteras vid införlivandet av direktivet.
Ändringsförslag
109
Kommissionens förslag
Ändringsförslag
Ändringsförslag
110
Förslag till direktiv
Bilaga I – punkt 4
Kommissionens förslag
Ändringsförslag
4.
Cyklar, sparkcyklar och andra transportmedel avsedda för idrottsutövning eller framförande på allmän väg eller allmän gång- och cykelväg.
4.
Sparkcyklar och andra transportmedel avsedda för idrottsutövning eller framförande på allmän väg eller allmän gång- och cykelväg.
Cyklar med en högsta sadelhöjd på mer än 435 mm, mätt som det vertikala avståndet från marken till sadelns ovansida, med sadeln i horisontellt läge och sadelstolpen placerad i högsta tillåtna läge.
Motivering
De nuvarande europeiska normerna för barncyklar är otydliga och skiljer mellan cyklar med en maximal sadelhöjd på mindre än 435 mm (EN 71-1), cyklar med en maximal sadelhöjd på mer än 435 mm men mindre än 635 mm (EN 14765) och cyklar med en sadelhöjd på över 635 mm (EN 14764).
Den första typen av cykel är inte avsedd att användas på allmän väg och betraktas i vissa länder som cykel och i andra länder inte som cykel, beroende på medlemsstatens lagstiftning.
Denna inkonsekvens leder till oklarhet både för marknadskontrollen och tillverkarna .
Ändringsförslag
111
Förslag till direktiv
Bilaga I – punkt 17a (ny)
Kommissionens förslag
Ändringsförslag
17a.
Barn b öcker som är utformade för eller tydligt avsedda att användas av barn och som endast är tillverkade av papp eller papper och endast innehåller sådana delar som är tillverkade av papp eller papper .
Ändringsförslag
112
Förslag till direktiv
Bilaga II – avsnitt I – punkt 4 – stycke 1
Kommissionens förslag
Ändringsförslag
4.
Leksaker och deras delar får inte medföra risk för strypning eller kvävning .
4.
Leksaker och deras delar får inte medföra risk för strypning
Motivering
Vissa leksakers form har förorsakat flera allvarliga olyckor och har nu förbjudits enligt standarden.
Samma regler bör gälla för förpackningar eftersom barn ofta leker även med dessa.
De flesta tillverkarna av försäljningsautomater och de största tillverkarna av överraskningsägg har redan vidtagit åtgärder och ersatt dessa kapslar med kapslar av ett säkrare slag.
Detta välkomnas men samtliga förpackningar bör uppfylla dessa strängare normer.
För att förebygga att mindre ansvarskännande tillverkare återinför den gamla sortens kapslar krävs det lagstiftning.
Ändringsförslag
113
Förslag till direktiv
Bilaga II – avsnitt I – punkt 4 – stycke 2
Kommissionens förslag
Ändringsförslag
Förpackningarna i vilka leksakerna saluförs i detaljhandeln får inte medföra risk för strypning eller kvävning genom att på yttre väg täppa till luftvägarna till munnen och näsan.
Förpackningarna i vilka leksakerna saluförs i detaljhandeln får inte medföra risk för strypning eller stopp i lufttillförseln genom att på yttre väg täppa till luftvägarna till munnen och näsan.
Sfäriska, äggformade eller ellipsformade förpackningar får inte vara av ett sådant format att de kan fastna i munnen eller i svalget och därigenom täppa till de nedre luftvägarna.
Motivering
Vissa leksakers form har förorsakat flera allvarliga olyckor och har nu förbjudits enligt standarden.
Samma regler bör gälla för förpackningar eftersom barn ofta leker även med dessa.
De flesta tillverkarna av försäljningsautomater och de största tillverkarna av överraskningsägg har redan vidtagit åtgärder och ersatt dessa kapslar med kapslar av ett säkrare slag.
Detta välkomnas men samtliga förpackningar bör uppfylla dessa strängare normer.
För att förebygga att mindre ansvarskännande tillverkare återinför den gamla sortens kapslar krävs det lagstiftning.
Ändringsförslag
114
Förslag till direktiv
Bilaga II – avsnitt I – punkt 4 – stycke 2a (nytt)
Kommissionens förslag
Ändringsförslag
Leksaker och deras delar får inte medföra risk för s topp i lufttillförseln genom att på yttre väg täppa till luftvägarna till munnen och näsan.
Motivering
Vissa leksakers form har förorsakat flera allvarliga olyckor och har nu förbjudits enligt standarden.
Samma regler bör gälla för förpackningar eftersom barn ofta leker även med dessa.
De flesta tillverkarna av försäljningsautomater och de största tillverkarna av överraskningsägg har redan vidtagit åtgärder och ersatt dessa kapslar med kapslar av ett säkrare slag.
Detta välkomnas men samtliga förpackningar bör uppfylla dessa strängare normer.
För att förebygga att mindre ansvarskännande tillverkare återinför den gamla sortens kapslar krävs det lagstiftning.
Ändringsförslag
115
Förslag till direktiv
Bilaga II – del I – punkt 4 – stycke 3
Kommissionens förslag
Ändringsförslag
Leksaker som uppenbarligen är avsedda för barn under 36 månader, deras beståndsdelar och delar som kan tas loss från leksakerna ska ha sådana dimensioner att de inte kan sväljas eller inandas.
Detta gäller också andra leksaker som är avsedda att stoppas i munnen, deras beståndsdelar och alla delar som kan tas loss från dem .
Leksaker som på grund av funktion, storlek eller utmärkande drag uppenbarligen är avsedda för barn under 36 månader samt leksakernas beståndsdelar och delar som kan tas loss från dem ska ha sådana dimensioner att de inte kan sväljas eller inandas.
Detta gäller också munstycken från andra leksaker som på grund av funktion, storlek eller utmärkande drag är avsedda att stoppas i munnen, deras beståndsdelar och alla delar som kan tas loss från munstycken, oavsett viken åldersgrupp som leksaken är avsedd för .
Motivering
Den nuvarande formuleringen är alltför restriktiv, eftersom en leksak för äldre barn, avsedd att stoppa i munnen, inte får bestå av några smådelar.
Ändringsförslag
116
Förslag till direktiv
Bilaga II – avsnitt I – punkt 4 – stycke 4
Kommissionens förslag
Ändringsförslag
Leksaker i livsmedel eller livsmedelsförpackningar måste ha sin egen förpackning.
Denna förpackning ska, i det skick den levereras, ha sådana dimensioner att den inte kan sväljas eller inandas.
Leksaker i livsmedel eller livsmedelsförpackningar måste ha sin egen förpackning.
Denna förpackning ska, i det skick den levereras, ha sådana dimensioner att den inte kan sväljas eller inandas och måste uppfylla övriga krav för förpackning av leksaker som fastställs i stycke 2 i denna punkt .
Cylinderformade inneremballage med avrundade ändar och som kan delas upp i två enskilda delar får inte vara utformade på ett sådant sätt att de kan täppa till de nedre luftvägarna.
Motivering
Vissa leksakers form har förorsakat flera allvarliga olyckor och har nu förbjudits enligt standarden.
Samma regler bör gälla för förpackningar eftersom barn ofta leker även med dessa.
De flesta tillverkarna av försäljningsautomater och de största tillverkarna av överraskningsägg har redan vidtagit åtgärder och ersatt dessa kapslar med kapslar av ett säkrare slag.
Detta välkomnas men samtliga förpackningar bör uppfylla dessa strängare normer.
För att förebygga att mindre ansvarskännande tillverkare återinför den gamla sortens kapslar krävs det lagstiftning.
Ändringsförslag
117
Förslag till direktiv
Bilaga II – avsnitt I – punkt 4 – stycke 5
Kommissionens förslag
Ändringsförslag
Leksaker som sitter så fast ihop med ett livsmedel att man att man måste konsumera det för att komma åt leksaken ska förbjudas.
Leksaker som sitter så fast ihop med ett livsmedel att man att man måste konsumera det för att komma åt leksaken ska förbjudas.
Delar av leksaker som annars direkt sitter ihop med ett livsmedel ska up pfylla de krav som fastställs i stycke 2 a i denna punkt .
Motivering
Vissa leksakers form har förorsakat flera allvarliga olyckor och har nu förbjudits enligt standarden.
Samma regler bör gälla för förpackningar eftersom barn ofta leker även med dessa.
De flesta tillverkarna av försäljningsautomater och de största tillverkarna av överraskningsägg har redan vidtagit åtgärder och ersatt dessa kapslar med kapslar av ett säkrare slag.
Detta välkomnas men samtliga förpackningar bör uppfylla dessa strängare normer.
För att förebygga att mindre ansvarskännande tillverkare återinför den gamla sortens kapslar krävs det lagstiftning.
Ändringsförslag
118
Förslag till direktiv
Bilaga II – avsnitt I – punkt 10
Kommissionens förslag
Ändringsförslag
10.
Ljudleksaker ska vara utformade och konstruerade så att ljudet inte skadar barnens hörsel.
10.
Ljudleksaker ska vara utformade och konstruerade så att ljudet inte skadar barnens hörsel.
Detta ska gälla alla leksaker, oavsett vilken åldersgrupp de är avsedda för.
Motivering
Studier pekar på att långvarig exponering för ljud över 80 dB kan orsaka hörselskador.
Barn är särskilt sårbara då deras öron är mer känsliga för höga decibelnivåer än vuxnas, vilket återspeglas i senare års ökning av barnhörselskador.
Decibelnivån för särskilt skadliga leksaker, s.k. impulsljudleksaker, bör av den anledningen sättas vid 115 dB.
Ändringsförslag
119
Förslag till direktiv
Bilaga II – del III – punkt 1
Kommissionens förslag
Ändringsförslag
1.
1.
Motivering
Se ändringsförslag 3.
Ändringsförslag
120
Förslag till direktiv
Bilaga II – avsnitt III – punkt 3
Kommissionens förslag
Ändringsförslag
3.
3.
Ändringsförslag
121
Förslag till direktiv
Bilaga II – del III – punkt 4
Kommissionens förslag
Ändringsförslag
4.
Ämnen eller preparat som klassificeras som CMR-ämnen i kategori 1 och 2 enligt direktiv 67/548/EEG får användas i leksaker om följande villkor är uppfyllda:
4.
Ämnen eller preparat som klassificeras som CMR-ämnen i kategori 1 och 2 enligt direktiv 67/548/EEG får användas i leksaker om följande villkor är uppfyllda:
4.1 Användningen av ämnet har utvärderats av behörig vetenskaplig kommitté och funnits vara säker, särskilt med tanke på exponeringen, och ett beslut enligt artikel 45.2 har antagits.
4.2.
Det finns inga lämpliga ersättningsämnen, vilket framgår av en analys av möjliga alternativ.
b) Det finns inga lämpliga ersättningsämnen eller preparat , vilket framgår av en analys av möjliga alternativ.
c) De är inte förbjudna att användas i konsumentvaror enligt förordning (EG) nr 1907/2006 (Reach).
Följande användning av ämnen eller preparat ska vara undantagna från förbudet i punkt 3:
[lägg till förteckning]
Ändringsförslag
122
Förslag till direktiv
Bilaga II – del III – punkt 5
Kommissionens förslag
Ändringsförslag
5.
5.
Ämnen eller preparat som klassificeras som CMR-ämnen i kategori 3 enligt direktiv 67/548/EEG ska vara förbjudna att använda i leksaker , om inte
a) användningen av ämnet har utvärderats av den behöriga vetenskapliga kommittén och funnits vara säker, särskilt med tanke på exponeringen,
c) de inte är förbjudna i konsumentvaror enligt förordning (EG) nr 1907/2006 (Reach).
Ändringsförslag
123
Förslag till direktiv
Bilaga II – avsnitt III – punkt 5a (ny)
Kommissionens förslag
Ändringsförslag
Ändringsförslag
124
Förslag till direktiv
Bilaga II – del III – led 5b (ny)
Kommissionens förslag
Ändringsförslag
Motivering
Användningen av farliga ämnen i leksaker är inte begränsad till CMR-ämnen, doftämnen eller ämnen som innehåller vissa beståndsdelar.
Alla farliga ämnen bör regelbundet utvärderas av kommissionen.
Skulle det vid denna utvärdering avslöjas en oacceptabel risk, bör kommissionen ges befogenhet att vidta lämpliga åtgärder inom ramen för kommittéförfarandet.
Ändringsförslag
125
Förslag till direktiv
Bilaga II – del III – led 5c (ny)
Kommissionens förslag
Ändringsförslag
Programmet ska ta hänsyn till rapporter från marknads kontrollerande organ och till synpunkter som medlemsstater och intressenter ger uttryck för.
Kommissionen ska besluta, med ledning av den behöriga vetenskapliga kommitténs åsikt, att vidta lämpliga restriktiva åtgärder, om nödvändigt.
Motivering
Användningen av farliga ämnen i leksaker är inte begränsad till CMR-ämnen, doftämnen eller ämnen som innehåller vissa beståndsdelar.
Alla farliga ämnen bör regelbundet utvärderas av kommissionen.
Skulle det vid denna utvärdering avslöjas en oacceptabel risk, bör kommissionen ges befogenhet att vidta lämpliga åtgärder inom ramen för kommittéförfarandet.
Ändringsförslag
126
Förslag till direktiv
Bilaga II – del III – punkt 6a (ny)
Kommissionens förslag
Ändringsförslag
6a.
Leksaker som är avsedda att komma i frekvent kontakt med huden, t.ex. fingerfärg eller modellera, ska uppfylla kraven på sammansättning och märkning i direktiv 76/768/EEG.
Motivering
Det finns inga skäl att i leksaksdirektivet ha mindre stränga krav för leksaker som kommer i frekvent kontakt med huden, än de normer som återfinns i kosmetikadirektivet.
Ändringsförslag
127
Förslag till direktiv
Bilaga II – avsnitt III – punkt 7
Kommissionens förslag
Ändringsförslag
7.
7.
Leksaker får inte innehålla följande allergiframkallande doftämnen:
(1) Ålandsrot (Inula helenium)
(2) Allylisotiocyanat
(4) 4-Tert-butylfenol
(5) Chenopodiumolja
(6) Cyklamenalkohol
(7) Dietylmaleat
(8) Dihydrokumarin
(9) 2,4-Dihydroxi-3-metylbensaldehyd
(10) 3,7-Dimetyl-2-okten-1-ol (6,7-dihydrogeraniol)
(12) Dimetylcitrakonat
(13) 7,11-Dimetyl-4,6,10-dodekatrien-3-on
(14) 6,10-Dimetyl-3,5,9-undekatrien-2-on
(15) Difenylamin
(16) Etylakrylat
(18) Trans-2-heptenal
(19) Trans-2-hexenaldietylacetal
(20) Trans-2-hexenaldimetylacetal
(22) 4-Etoxifenol
(23) 6-lsopropyl-2-dekahydronaftalenol
(25) 4-Metoxifenol
(26) 4-(p-Metoxifenyl)-3-buten-2-on
(27) 1-(p-Metoxifenyl)-1-penten-3-on
(28) Metyl-trans-2-butenoat
(29) 6-Metylkumarin
(30) 7-Metylkumarin
(31) 5-Metyl-2,3-hexanedion
(33) 7-Etoxi-4-metylkumarin
(34) Hexahydrokumarin
(35) Perubalsam (Myroxylon pereirae Klotzsch)
(36) 2-Pentyliden-cyklohexanon
(37) 3,6,10-Trimetyl-3,5,9-undekatrien-2-on
(38) Citronverbenaolja (Lippia citriodora Kunth).
(39) Ambrettmysk
(40) 4-fenyl-3-buten-2-on
(41) Amylkanelaldehyd
(42) Amylkanelalkohol
(43) Bensylalkohol
(44) Bensylsalicylat
(45) Kanelalkohol
(46) Kanelaldehyd
(47) Citral
(48) Kumarin
(49) Eugenol
(50) Geraniol
(51) Hydroxicitronellal
(52) Hydroxymethylpentylcyclohe
(53) Isoeugenol
(54) Ekmosseextrakt
(55) Trämosseextrakt
Spår av dessa ämnen ska dock tillåtas förutsatt att förekomsten är tekniskt oundviklig med god tillverkningssed.
Spår av dessa ämnen ska dock tillåtas förutsatt att förekomsten är tekniskt oundviklig med god tillverkningssed och inte överskrider 10 ppm .
Dessutom ska följande allergiframkallande doftämnen anges om de används i leksaker i koncentrationer över 0,01 viktprocent.
(1) Anisylalkohol
(2) Amylkanelalkohol
(3) Anisylalkohol
(4) Bensylalkohol
(5) Bensylbensoat
(6) Bensylcinnamat
(7) Bensylsalicylat
(8) Kanelaldehyd
(9) Kanelalkohol
(10) Citral
(11) Citronellol
(12) Kumarin
(13) Eugenol
(14) Farnesol
(15) Geraniol
(16) Hexylkanelaldehyd
(17) Hydroxicitronellal
(18) Hydroxi-metylpentylcyklohexenkarboxaldehyd
(19) Isoeugenol
(21) d-Limonen
(22) Linalol
(23) Metylheptinkarbonat
(24) 3-Metyl-4-(2,6,6-trimetyl-2-cyklohexen-1-yl)-3-buten-2-on
(25) Ekmosseextrakt
(26) Trämosseextrakt
Ändringsförslag
128
Förslag till direktiv
Bilaga III – del III – punkt 7a (ny)
Kommissionens förslag
Ändringsförslag
7a.
Användningen av de doftämnen som anges i punkterna 41–55 i förteckningen under punkt 7.1 och de doftämnen som anges i punkterna 1–11 i förteckningen under punkt 7.3 ska vara tillåtna i doftspel, kosmetiklådor och smakspel under förutsättning att
i) dessa doftämnen tydligt anges på förpackningen och förpackningen innehåller varningstexten ”innehåller allergiframkallande doftämnen”,
ii) de produkter som barnet tillverkar i enlighet med anvisningarna måste överensstämma med kraven i direktiv 76/768/EEG [ Kosmetikadirektivet ] och,
iii) i förekommande fall, att dessa doftämnen överensstämmer med den relevanta livsmedelslagstiftningen.
Barn under 36 månader ska inte tillåtas använda sådana doftspel, kosmetiklådor och smakspel, och dessa leksaker ska uppfylla bestämmelserna i del B avsnitt 1 i bilaga V.
Ändringsförslag
129
Förslag till direktiv
Bilaga II – avsnitt III – punkt 8 - tabell
Kommissionens förslag
Ändringsförslag
Grundämne
mg/kg
i vätske-formigt eller klibbigt leksaks-material
Grundämne
mg/kg
Aluminium
5625
1406
Aluminium
5625
1406
Antimon
45
11,3
Antimon
45
11,3
Arsenik
7,5
1,9
Barium
4500
1125
Barium
4500
1125
Bor
1200
300
Bor
1200
300
Kadmium
3,8
0,9
Krom (III)
37,5
9,4
Krom (III)
37,5
9,4
Krom (VI)
0,04
0,01
Kobolt
10,5
2,6
Kobolt
10,5
2,6
Koppar
622,5
156
Koppar
622,5
156
Bly
27
6,8
Mangan
1200
300
Mangan
1200
300
Kvicksilver
15
3,8
Nickel
75
18,8
Nickel
75
18,8
Selen
37,5
9,4
Selen
37,5
9,4
Strontium
4500
1125
Strontium
4500
1125
Tenn
15000
3750
Tenn
15000
3750
Organiskt tenn
1,9
0,5
Zink
3750
938
Zink
3750
938
Motivering
Arsenik, kadmium, bly, krom (VI), kvicksilver och organiskt tenn är mycket toxiska och bör totalförbjudas i leksaker.
Kadmium, bly, krom (VI) och kvicksilver är redan förbjudna i bilar och elektriska och elektroniska apparater.
Krom (VI) i cement behöver reduceras till en oskadlig form genom tillsats av järnsulfat.
Arsenik är förbjudet i färg och för behandling av trä (med vissa undantag).
Organiska tennföreningar är förbjudna som biocider.
Dessa ämnen bör helt klart inte ingå i leksaker.
Ändringsförslag
130
Förslag till direktiv
Bilaga II – del III – punkt 8a (ny)
Kommissionens förslag
Ändringsförslag
8a.
Det är förbjudet att använda arsenik, kadmium, krom (VI) bly, kvicks i lver och organiskt tenn i leksaker.
Spår av dessa ämnen kan tillåtas såvida det inte kan undvikas tekniskt, i enlighet med god tillverkningssed.
Denna punkt ska gälla utan hinder av punkterna 3–5.
Ändringsförslag
131
Förslag till direktiv
Bilaga II – del V – punkt 2
Kommissionens förslag
Ändringsförslag
2.
Tygleksaker för barn under 36 månader ska gå att tvätta och ska uppfylla säkerhetskraven även efter tvätt.
2.
Tygleksaker för barn under 36 månader ska gå att tvätta och ska uppfylla kraven på funktionsduglighet och säkerhet även efter tvätt.
Motivering
En hög nivå på hygienen ska vara förenlig med garantin för leksakernas funktionsduglighet och säkerhet.
Ändringsförslag
132
Förslag till direktiv
Bilaga III – punkt 2
Kommissionens förslag
Ändringsförslag
2.
(Berör inte den svenska versionen.)
Motivering
(Berör inte den svenska versionen.)
Ändringsförslag
133
Förslag till direktiv
Bilaga III – punkt 4
Kommissionens förslag
Ändringsförslag
4.
Föremål för försäkran (identifiera leksaken så att den kan spåras):
4.
Föremål för försäkran (identifiera leksaken så att den kan spåras .
Om det är lämpligt kan ett fotografi bifogas. ):
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
134
Förslag till direktiv
Bilaga III – punkt 7
Kommissionens förslag
Ändringsförslag
7.
Det anmälda organet … (namn, nummer) har utfört ... (beskrivning av åtgärden) och utfärdat intyg: …
7.
Det anmälda organet … (namn, nummer) har utfört ... (beskrivning av åtgärden) och utfärdat intyg: …
Motivering
Teknisk anpassning till åtgärdspaketet för den inre marknaden för varor.
Ändringsförslag
135
Förslag till direktiv
Bilaga V – del A – stycke 1a (nytt)
Kommissionens förslag
Ändringsförslag
Alla varningar i form av varningstext eller varningssymbol ska föregås av or det ”varning”.
Motivering
Alla varningar ska börja med ordet ”varning” för att klargöra för konsumenterna att texten avser säkerhetsfrågor och för att uppmärksamma dem på varningen.
Detta gäller särskilt varningar i form av varningssymbol.
Ändringsförslag
136
Förslag till direktiv
Bilaga V – del B – punkt 1
Kommissionens förslag
Ändringsförslag
1.
Leksaker som inte är avsedda för barn under 36 månader
1.
[Varningssymbol]
[Varningssymbol]
Varningstexterna ska kompletteras med en kortfattad upplysning, som kan finnas i bruksanvisningen, om vilka specifika faror som ligger till grund för åldersgränsen.
Varningstexterna ska kompletteras med en kortfattad upplysning, som kan finnas i bruksanvisningen, om vilka specifika faror som ligger till grund för åldersgränsen.
Dessa varningstexter får inte användas för leksaker som är utformade för eller, som på grund av funktion, storlek eller utmärkande drag, är avsedda för barn under 36 månader.
Denna bestämmelse gäller inte leksaker som på grund av funktion, storlek, utmärkande drag, egenskaper eller andra viktigare omständigheter uppenbarligen inte är avsedda för barn under 36 månader.
Denna bestämmelse gäller inte leksaker som på grund av funktion, storlek, utmärkande drag, egenskaper eller andra viktigare omständigheter uppenbarligen inte är avsedda för barn under 36 månader.
Motivering
Mjukt stoppade leksaker som nallar och mjuka dockor bör aldrig innehålla små lösa delar eftersom barn sannolikt kommer att leka med dem oavsett vad tillverkaren tänkt sig.
Ändringsförslag 1
37
Förslag till direktiv
Bilaga V – del B – punkt 7
Kommissionens förslag
Ändringsförslag
Leksaker i livsmedel och livsmedelsförpackningar ska vara försedda med texten:
Leksaker i livsmedel och livsmedelsförpackningar ska vara försedda med texten:
”Tillsyn av en vuxen rekommenderas”
” Leksak i förpackningen.
Ändringsförslag
138
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
7a.
Skyddsmasker och skyddshjälmar i form av leksaker
Denna leksak ger inte något skydd”.
Motivering
Varningarna ska inte kräva någon närmare förklaring utan man bör kunna vara säker på att konsumenten förstår deras innebörd och vidtar erforderliga åtgärder.
Ändringsförslag
139
Förslag till direktiv
Bilaga V – del B – punkt 7b (ny)
Kommissionens förslag
Ändringsförslag
7b.
Leksaker som är avsedda att fästas tvärs över en vagga, barnsäng eller barnvagn med hjälp av snoddar, band, resårband eller remmar ska ha följande varningstext dels på förpackningen, dels permanent anbringad på själva leksaken:
”För att förhindra eventuell skada genom att barnet trasslar in sig, avlägsna denna leksak så snart barnet börjar kunna resa sig på händer och knän.”
MOTIVERING
1.
Bakgrund och nya element i förslaget
Kommissionens förslag syftar till att till upphäva direktiv 88/378/EEG av den 3 maj 1988 om leksakers säkerhet och ersätta det med ett nytt direktiv.
Direktiv 88/378/EEG var det första direktiv som infördes enligt den s.k. nya metoden, där de grundläggande säkerhetskraven infördes i själva lagstiftningen och man hänvisade till harmoniserade normer när det gällde de tekniska specifikationerna.
Det föreslagna nya direktivet baserar sig på samma principer.
Även om direktivet från 1988 har levt upp till förväntningarna och redan garanterar en hög säkerhetsnivå för leksaker i Europeiska unionen, är det efter 20 år redo för en modernisering.
Man måste också tänka på nya säkerhetsrisker som kan uppkomma genom utveckling och marknadsföring av nya typer av leksaker, eventuellt tillverkade av nya material.
Huvuddragen i översynen är enligt kommissionen följande:
En effektivare och mer konsekvent användning av direktivet.
Anpassning till den allmänna lagstiftningen om saluföring av produkter.
Det föreslagna direktivet handlar bara om leksakers (fysiska) säkerhet och innehåller inga bestämmelser rörande med pedagogiskt värde eller moraliska aspekter.
2.
Anpassning av förslaget till de godkända nya bestämmelserna i åtgärdspaketet för den inre marknaden för varor
De rättsliga ramarna för saluföring av produkter kommer snart att ändras.
– En ny förordning för saluföring av produkter.
Denna förordning innehåller bestämmelser om ackreditering och marknadsövervakning.
Det nya direktivet måste anpassas till denna nya rättsliga ram.
Kommissionens förslag stämmer överens med det förslag till förordning och beslut som kommissionen från början lade fram, med inte med den text som Europaparlamentet antog den 21 februari 2008, och som kanske kommer att godkännas av rådet.
Kommissionen har förklarat att man inte kommer att utforma ett ändrat förslag till leksaksdirektiv för att anpassa det till det nya åtgärdspaketet för den inre marknaden för varor.
För att komma vidare med det föreslagna direktivet föreslår föredraganden att Europaparlamentet för in de tekniska anpassningarna i texten till det föreslagna direktivet i den av Europaparlamentet nyligen godkända ramtexten (åtgärdspaketet för den inre marknaden för varor).
Det gäller anpassningar avseende
- definitioner
- allmänna villkor för de ekonomiska aktörerna
- presumtion om överensstämmelse
- formell invändning mot harmoniserade standarder
- bestämmelser för CE-märkning
- krav avseende organ för bedömning av överensstämmelse
- anmälningsförfaranden
- förfaranden för produkter som medför risker
Ändringsförslagen 1–79 avser dessa tekniska anpassningar till den nya ramlagstiftningen.
De ligger i linje med Europaparlamentets val och beslut i samband med denna allmänna ram.
3.
Bedömning
– allmänt
Föredraganden anser att barn, som är de mest utsatta konsumenterna, måste skyddas så fullständigt som möjligt och att deras föräldrar och ledsagare måste kunna lita på att de leksaker som erbjuds på europamarknaden uppfyller stränga säkerhetskrav.
Därför instämmer parlamentet i de av kommissionen uppställda målen: Modernisering, förtydligande och skärpning av direktivets säkerhetskrav och dess genomförandebestämmelser.
Parlamentet instämmer också i stora drag i de av kommissionen gjorda tilläggen till och ändringarna av bestämmelserna i det gällande direktivet 88/378/EEG.
Närmare upplysningar om föredragandens ändringsförslag
– kemiska egenskaper
Det finns ingen anledning att göra någon skillnad mellan ämnen i kategorierna 1 och 2 å ena sidan och kategori 3 å andra sidan
Föredraganden föreslår att villkoret för att undantagsvis tillåta dess ämnen ska vara lika för de tre kategorierna, nämligen att den vetenskapliga kommittén har bedömt användningen av ämnet i leksaker och kommit fram till att det är acceptabelt, och att det dessutom inte finns något lämpligt alternativt ämne.
Föredraganden föreslår också att man helt ska förbjuda användningen av allergiframkallande doftämnen.
– mekaniska egenskaper
Även om föredraganden är bekymrad över de risker som kan uppkomma vid användning av små men mycket kraftiga magneter i leksaker anser hon att det inte är nödvändigt att i direktivet infoga en särskild bestämmelse för magneter.
En särskild norm för magnetiska leksaker förbereds av CEN, och kommissionen har vidtagit interimsåtgärder (krav på en varning om att det kan vara farligt att svälja mer än en magnet).
– hantverksmässigt tillverkade eller icke serietillverkade leksaker
Föredraganden är medveten om att det för små eller medelstora företag som tillverkar leksaker på hantverksmässigt sätt, eller i varje fall inte seriemässigt, inte är lätt att uppfylla de strängare kraven i direktivet.
Hon arbetar på en lösning, men har ännu inte funnit något juridiskt hållbart koncept.
Hon vill gärna få reda på kollegornas uppfattning i denna fråga.
– leksaker som uttryckligen är avsedda för barn i en bestämd åldersgrupp
Alltför ofta förses leksaker som är avsedda för spädbarn och mycket små barn med en varning om att leksaken inte är lämplig för barn under 36 månader.
Tillverkarna försöker på detta sätt att kringgå strängare säkerhetsföreskrifter för att undgå eventuellt juridiskt ansvar.
Detta är oförsvarligt och måste förbjudas.
Dessutom är dessa felaktiga åldersangivelser mycket förvirrande för köparna och befrämjar inte det förtroende som konsumenten borde ha för leksakers säkerhet.
De relevanta bestämmelserna i direktivets artikel 10 måste förtydligas.
– leksaker som kommer i kontakt med munnen eller huden
Leksaker som är avsedda att ofta stoppas i munnen (t.ex. leksaksinstrument, bitringar, etc.) måste, oavsett åldern på de barn för vilka de är avsedda, uppfylla samma stränga gränsvärden för migration som återfinns i direktiv 1935/2004/EG.
Leksaker som är avsedda att ofta komma i kontakt med barns hud måste, oavsett åldern på barnen, uppfylla etiketterings- och sammansättningsbestämmelserna i kosmetikadirektivet.
– rapporteringscentrum för leksakers säkerhet
I vissa medlemsstater eller regioner har man inrättat rapporteringscentrum för farliga leksaker, dit professionella barnskötare men också konsumenter/föräldrar kan anmäla egenskaper som gör att leksaker inte är säkra samt olyckor eller tillbud i samband med leksaker.
Utan att förespråka att sådana rapporteringscentrum ska inrättas i varje medlemsstat, anser föredraganden att det skulle kunna vara lämpligt att undersöka huruvida konsumenterna vet att de, när de kommer i kontakt med farliga leksaker, kan anmäla detta hos en instans som kan ha nytta av dessa upplysningar.
– språk
Det är grundläggande att de varningar som krävs enligt direktivet, och även bruksanvisningarna, skrivs på ett språk som är begripligt för konsumenterna.
YTTRANDE från utskottet för miljö, folkhälsa och livsmedelssäkerhet
till utskottet för den inre marknaden och konsumentskydd
över förslaget till Europaparlamentets och rådets direktiv om leksakers säkerhet
( KOM(2008)0009 – C6‑0039/2008 – 2008/0018(COD) )
Föredragande:
Anne Ferreira
KORTFATTAD MOTIVERING
Leksakers säkerhet omfattas av ett direktiv som antogs 1988 och ändrades 1993.
Texten har gjort det möjligt att harmonisera de befintliga bestämmelserna i medlemsstaterna och att ge barn ett bättre skydd.
Men direktivet måste anpassas till det ekonomiska sammanhang som vi lever i, till de nya vetenskapliga rön vi har, samtidigt som det måste ta hänsyn till statistik över riskerna och de nya samhälleliga kraven.
Nya uppgifter att beakta
Det ekonomiska sammanhanget
Det allt större kommersiella utbytet har bidragit till att i stor utsträckning ändra den ekonomiska leksakssektorn.
Ungefär 80 procent av de leksaker som saluförs i EU är importerade och man bör påminna om att under 2007 återkallades miljontals leksaker från Kina på grund av att de inte uppfyllde EU:s standarder.
Varuhandeln gör att man måste se över bestämmelserna för utsläppandet på marknaden och för kontrollen av att standarderna följs.
Nya vetenskapliga rön
Leksakerna innehåller alltmer kemiska ämnen vilket gör att man måste anpassa lagstiftningen till de risker som finns med de ämnenas närvaro och till det särskilda sätt som barn kan använda leksaker på (suga, kasta etc.).
Statistik och riskhantering
De olyckor som anmäls i samband med leksaker är i huvudsak allvarliga olyckor.
Man bör beakta samtliga olyckor för att bättre förstå farorna och riskerna i samband med att leksaker används.
I syfte att bättre förebygga olyckor som orsakas av att leksaker används bör vi stödja oss på de vetenskapliga bedömningar och riskbedömningar som finns tillgängliga.
Försiktighetsprincipen bör tillämpas inte bara för en särskild produktkategori utan allmänt.
Nya samhälleliga krav
Leksaker återspeglar vårt samhälle och de blir därmed allt fler och mer varierande.
De följer barnen i deras känslomässiga och intellektuella utveckling och ingår i barnens värld både i hemmet och i samband med inlärning.
Slutkonsumenterna har rätt att vänta sig och att kräva att de produkter de köper är av god kvalitet och att de inte kan vara farliga för vare sig barnen eller de som har barnen i uppsikt.
Slutkonsumenterna är miljömedvetna och kräver också att produkterna ska vara miljövänliga.
Detta krav gäller produktens livscykel, dess förpackning samt leksakernas livslängd.
Undersökningar visar att många av de leksaker som släpps på marknaden inte är tillräckligt tåliga och att de fort blir till avfall.
Kommissionens förslag innehåller framsteg men det krävs preciseringar.
Ändringsförslagen har avfattats i det syftet, särskilt beträffande:
Vikten av varningstexten och de föreskrifter som åtföljer produkten
De begrepp som används bör vara en definition som alla förstår och de ska följa EU:s nomenklatur, till exempel vad avser risken för kvävning.
Handlingarna bör dessutom vara lättlästa.
Det är även mycket viktigt att de skrivs på det officiella språket eller de officiella språken i de medlemsstater där de saluförs.
Bestämmelserna för tidsfristen för svar på frågor och information bör anges i detalj.
Det gäller även bestämmelserna för avhjälpande åtgärder, tillbakadragning och återkallelse av leksaker som inte uppfyller standarderna.
Produktkvalitén och risker i samband med innehåll av kemiska ämnen
Faktum är att organen inte är fullt utvecklade förrän efter en viss ålder och att CMR-ämnen utgör ett hinder för barns utveckling och deras hälsa på sikt.
Man måste alltså se till även annan lagstiftning (förpackningar för livsmedel, kosmetika etc.) där man satt gränsvärden för ämnesinnehåll eller ämnens överföring, och bedöma dessa med avseende på hur barnet kan använda produkten (suga, hudkontakt etc.)
Föredraganden uppskattar att bestämmelserna om kemiska ämnen även bör omfatta PBT‑ämnen etc.
I kommissionens förslag prioriteras den fria rörligheten framför leksakers säkerhet.
I detta sammanhang måste bevisbördan vara omvänd i likhet med Reach.
Även de ekonomiska aktörerna bör visa att deras leksaker är säkra och att de uppfyller kraven för barns hälsa.
Till följd av många utlokaliseringar importeras 80 procent av de leksaker som saluförs i EU, i huvudsak från Kina, där arbetsvillkoren är dåliga och miljöstandarderna låga.
Det är alltså många som delar på ansvaret för leksakernas säkerhet.
Men de stora västerländska märkena och beställarna dominerar fortfarande leksaksmarknaden och det är deras samt importörernas och distributörernas uppgift att se till att produktspecifikationerna, som ska följa gemenskapslagstiftningen, fastställs och efterlevs och sålunda garanterar en hög nivå för våra barns hälsoskydd.
ÄNDRINGSFÖRSLAG
Utskottet för miljö, folkhälsa och livsmedelssäkerhet uppmanar utskottet för den inre marknaden och konsumentskydd att som ansvarigt utskott infoga följande ändringsförslag i sitt betänkande:
Ändringsförslag
1
Förslag till direktiv
Skäl 3a (nytt)
Kommissionens förslag
Ändringsförslag
Motivering
Eftersom det inte finns några uppgifter om de faror och risker som leksaker kan medföra för barns säkerhet och hälsa och eftersom barn tillhör de grupper av befolkningen som är mycket sårbara eller sårbara beroende på ålder, bör försiktighetsprincipen tas med i lagstiftningen om leksakers säkerhet så att både medlemsstaternas behöriga myndigheter och de ekonomiska aktörerna kan vidta åtgärder för att hindra att vissa leksaker kommer ut på marknaden.
Lagstiftningen bör ha en allmän räckvidd.
Ändringsförslag
2
Förslag till direktiv
Skäl 8
Kommissionens förslag
Ändringsförslag
(8) Alla ekonomiska aktörer som ingår i leverans- och distributionskedjan bör vidta åtgärder för att se till att de endast tillhandahåller sådana leksaker på marknaden som överensstämmer med den tillämpliga lagstiftningen.
I detta direktiv görs en tydlig och proportionell fördelning av skyldigheterna som svarar mot varje aktörs roll i leverans- och distributionsprocessen.
(8) Alla ekonomiska aktörer som ingår i leverans- och distributionskedjan bör agera så ansvarsfullt och försiktigt som det krävs för att garantera att de leksaker som de släpper ut på marknaden inte har några farliga effekter på barns säkerhet och hälsa vid normal användning och under användningsomständigheter som rimligen kan förutses.
De ekonomiska aktörerna bör vidta åtgärder för att se till att de endast tillhandahåller sådana leksaker på marknaden som överensstämmer med den tillämpliga lagstiftningen.
I detta direktiv görs en tydlig och proportionell fördelning av skyldigheterna som svarar mot varje aktörs roll i leverans- och distributionsprocessen.
Motivering
Det räcker inte att påminna de ekonomiska operatörerna om att vidta lämpliga åtgärder, det är också bra att påminna dem om att de är ansvariga.
Ändringsförslag
3
Förslag till direktiv
Skäl 16
Kommissionens förslag
Ändringsförslag
(16) För att barnen ska skyddas mot nyupptäckta risker måste nya grundläggande säkerhetskrav också antas .
Det är särskilt nödvändigt att komplettera och uppdatera bestämmelserna om kemikalier i leksaker.
Dessa bestämmelser bör ange att leksaker bör överensstämma med den allmänna kemikalielagstiftningen, särskilt Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 om registrering, utvärdering, godkännande och begränsning av kemikalier (Reach), inrättande av en europeisk kemikaliemyndighet, ändring av direktiv 1999/45/EG och upphävande av rådets förordning (EEG) nr 793/93 och kommissionens förordning (EG) nr 1488/94 samt rådets direktiv 76/769/EEG och kommissionens direktiv 91/155/EEG, 93/67/EEG, 93/105/EG och 2000/21/EG.
Bestämmelserna bör emellertid också anpassas till barns särskilda behov eftersom de är sårbar konsumenter.
De specifika gränsvärden som anges i direktiv 88/378/EEG för vissa ämnen bör uppdateras mot bakgrund av nya vetenskapliga rön.
(16) För att garantera en hög skydds- och hälsonivå för barn och miljön mot olika slags risker , bör man vara särskilt vaksam mot farliga och mycket farliga ämnen .
Det är också nödvändigt att anta grundläggande säkerhetskrav.
Det är särskilt nödvändigt att komplettera och uppdatera bestämmelserna om kemikalier i leksaker.
Dessa bestämmelser bör ange att leksaker bör överensstämma med den allmänna kemikalielagstiftningen, särskilt Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 om registrering, utvärdering, godkännande och begränsning av kemikalier (Reach), inrättande av en europeisk kemikaliemyndighet, ändring av direktiv 1999/45/EG och upphävande av rådets förordning (EEG) nr 793/93 och kommissionens förordning (EG) nr 1488/94 samt rådets direktiv 76/769/EEG och kommissionens direktiv 91/155/EEG, 93/67/EEG, 93/105/EG och 2000/21/EG.
Bestämmelserna bör emellertid också anpassas till barns särskilda behov eftersom de är sårbara konsumenter.
De specifika gränsvärden som anges i direktiv 88/378/EEG för vissa ämnen bör uppdateras mot bakgrund av nya vetenskapliga rön.
Motivering
I fördragen och den relevanta gemenskapslagstiftningen hänvisas det hela tiden till målsättningen med en hög hälsoskyddsnivå för de berörda personerna och miljön.
Man bör ta samma hänsyn vid översynen av lagstiftningen om leksakers säkerhet.
Eftersom detta skäl gäller kemiska ämnen är det absolut nödvändigt att hänvisa till farliga och mycket farliga ämnen.
Ändringsförslag
4
Förslag till direktiv
Skäl 16a (nytt)
Kommissionens förslag
Ändringsförslag
(16a) De ekonomiska aktörer som begär ett undantag för att använda ett mycket farligt ämne i leksaker bör bevisa att det inte finns något säkrare alternativ.
Motivering
Man bör generellt undvika att använda mycket farliga ämnen på grund av de eventuella risker som de kan ha på barns hälsa under en kortare eller längre tid.
Det kan emellertid vara möjligt att använda sådana ämnen, men då måste tillverkarna visa att det inte finns något ersättningsämne som är säkrare.
Ändringsförslag
5
Förslag till direktiv
Skäl 16b (nytt)
Kommissionens förslag
Ändringsförslag
(16b) Ansvaret för riskerna i samband med leksaker, särskilt de som är knutna till användandet av kemiska ämnen i leksaker, bör ligga på de fysiska eller juridiska personer som tillverkar, importerar eller släpper ut leksakerna på marknaden.
Motivering
De ekonomiska aktörerna i leksakssektorn bör även vara helt medvetna om de eventuellt farliga effekterna av att använda vissa kemiska ämnen eller blandningar på barns hälsa.
De bör alltså ta med problematiken kring kemiska ämnen när de hanterar riskerna i samband med användning av leksaker.
Ändringsförslag
6
Förslag till direktiv
Skäl 17
Kommissionens förslag
Ändringsförslag
(17) De allmänna och särskilda kemikaliekraven i detta direktiv bör syfta till att skydda barns hälsa från farliga ämnen i leksaker, medan miljöproblemen behandlas i övergripande miljölagstiftning som också gäller leksaker, särskilt Europaparlamentets och rådets direktiv 2006/12/EG av den 5 april 2006 om avfall, Europaparlamentets och rådets direktiv 2002/95/EG av den 27 januari 2003 om begränsning av användningen av vissa farliga ämnen i elektriska och elektroniska produkter, Europaparlamentets och rådets direktiv 2002/96/EG av den 27 januari 2003 om avfall som utgörs av eller innehåller elektriska och elektroniska produkter, Europaparlamentets och rådets direktiv 94/62/EG av den 20 december 1994 om förpackningar och förpackningsavfall samt i Europaparlamentets och rådets direktiv 2006/66/EG av den 6 september 2006 om batterier och ackumulatorer och förbrukade batterier och ackumulatorer och om upphävande av direktiv 91/157/EEG 5 .
(17) De allmänna och särskilda kemikaliekraven i detta direktiv bör syfta till att skydda barns hälsa från farliga ämnen i leksaker, medan miljöproblemen behandlas i den miljölagstiftning som gäller elektriska och elektroniska leksaker, nämligen Europaparlamentets och rådets direktiv 2002/95/EG av den 27 januari 2003 om begränsning av användningen av vissa farliga ämnen i elektriska och elektroniska produkter samt Europaparlamentets och rådets direktiv 2002/96/EG av den 27 januari 2003 om avfall som utgörs av eller innehåller elektriska och elektroniska produkter.
Dessutom regleras miljöfrågor som rör avfall av Europaparlamentets och rådets direktiv 2006/12/EG av den 5 april 2006 om avfall, medan de miljöfrågor som rör förpackningar regleras av Europaparlamentets och rådets direktiv 94/62/EG av den 20 december 1994 om förpackningar och förpackningsavfall , och de miljöfrågor som rör batterier och ackumulatorer regleras i Europaparlamentets och rådets direktiv 2006/66/EG av den 6 september 2006 om batterier och ackumulatorer och förbrukade batterier och ackumulatorer och om upphävande av direktiv 91/157/EEG.
Motivering
Kommissionens text ger intrycket av att miljöhänsyn uttryckligen gäller alla leksaker, medan det endast berör elektriska och elektroniska leksaker.
Övergripande lagstiftning är inte uttryckligen tillämplig på leksaker och bör inte klumpas ihop med direktivet om elektriska och elektroniska produkter samt direktivet om avfall som utgörs av eller innehåller elektriska och elektroniska produkter.
Ändringsförslag
7
Förslag till direktiv
Skäl 18
Kommissionens förslag
Ändringsförslag
(18) I enlighet med försiktighetsprincipen bör det fastställas särskilda säkerhetskrav för att förebygga den särskilda fara som leksaker i livsmedel kan innebära, eftersom kombinationen leksak och mat skulle kunna medföra en annan typ av kvävningsrisk än den som leksaken ensam medför och som alltså inte omfattas av några specifika gemenskapsåtgärder.
(18) Det bör fastställas särskilda säkerhetskrav för att förebygga den särskilda fara som leksaker i livsmedel kan innebära, eftersom kombinationen leksak och mat skulle kunna medföra en annan typ av kvävningsrisk än den som leksaken ensam medför och som alltså inte omfattas av några specifika gemenskapsåtgärder.
Motivering
Försiktighetsprincipen bör tillämpas allmänt inom ramen för detta omarbetade direktiv.
Detta ändringsförslag har även samband med ändringsförslag 1 avseende skäl 3a.
Ändringsförslag
8
Förslag till direktiv
Skäl 19
Kommissionens förslag
Ändringsförslag
(19) Eftersom det kan finnas eller komma nya leksaker som medför faror som inte omfattas av särskilda säkerhetskrav i detta direktiv är det nödvändigt att fastställa ett allmänt säkerhetskrav som rättslig grund för åtgärder mot sådana leksaker.
Leksakernas säkerhet bör då bestämmas utifrån hur de är avsedda att användas eller kan förutses användas med tanke på barns normala beteende, eftersom de i regel inte är lika försiktiga som vuxna.
(19) Eftersom det kan finnas eller komma nya leksaker som medför faror som inte omfattas av särskilda säkerhetskrav i detta direktiv är det nödvändigt att fastställa ett allmänt säkerhetskrav som rättslig grund för åtgärder mot sådana leksaker.
Leksakernas säkerhet bör då bestämmas utifrån hur de är avsedda att användas eller rimligen kan förutses användas med tanke på barns normala beteende, eftersom de i regel inte är lika försiktiga som vuxna.
Motivering
Man måste ange de olika typerna av förutsebara användningar som ska bedömas.
Det är nödvändigt att tänka på det när leksaken bedöms så att man tar hänsyn till de olika sätt på vilka barn kan använda en leksak samtidigt som man utesluter sådana händelser som barn i en viss ålder inte skulle kunna utföra på grund av barnets utvecklingsnivå, fysiska eller intellektuella nivå, etc.
Ändringsförslag
9
Förslag till direktiv
Skäl 21
Kommissionens förslag
Ändringsförslag
(21) CE-märkningen visar att en leksak överensstämmer med kraven och är det synliga resultatet av en hel process av bedömning av överensstämmelse i vid bemärkelse.
Därför bör det i detta direktiv fastställas allmänna principer för hur CE‑märkningen ska utformas och användas.
(Berör inte den svenska versionen.)
Motivering
(Berör inte den svenska versionen.)
Ändringsförslag
10
Förslag till direktiv
Skäl 22
Kommissionens förslag
Ändringsförslag
(22) Det är mycket viktigt att klargöra både för tillverkarna och användarna att tillverkaren genom att CE-märka leksaken försäkrar att den överensstämmer med alla tillämpliga krav och tar på sig det fulla ansvaret för detta.
(22) Det är mycket viktigt att klargöra för tillverkarna att tillverkaren genom att CE‑märka leksaken försäkrar att den överensstämmer med alla tillämpliga krav och tar på sig det fulla ansvaret för detta.
Motivering
Har samband med ändringsförslag 8.
Ändringsförslag
11
Förslag till direktiv
Skäl 32
Kommissionens förslag
Ändringsförslag
(32) Kommissionen bör särskilt få befogenhet att i vissa väl definierade fall anpassa kemikaliekraven och i vissa fall bevilja undantag från förbudet mot CMR‑ämnen samt anpassa ordalydelsen i varningstexterna för vissa kategorier av leksaker.
Eftersom detta är åtgärder med allmän räckvidd som avser att ändra icke väsentliga delar av detta direktiv, eller att komplettera det genom tillägg av nya icke väsentliga delar, ska de antas enligt det föreskrivande förfarandet med kontroll i artikel 5a i beslut 1999/468/EG.
(32) Kommissionen bör särskilt få befogenhet att i vissa väl definierade fall anpassa kemikaliekraven och i vissa fall bevilja undantag från förbudet mot mycket farliga ämnen och CMR-ämnen samt anpassa ordalydelsen i varningstexterna för vissa kategorier av leksaker.
Eftersom detta är åtgärder med allmän räckvidd som avser att ändra icke väsentliga delar av detta direktiv, eller att komplettera det genom tillägg av nya icke väsentliga delar, ska de antas enligt det föreskrivande förfarandet med kontroll i artikel 5a i beslut 1999/468/EG.
Motivering
Ändringsförslaget har samband med ändringsförslagen till skälen 16, artikel 47 och bilaga II, del III.
Ändringsförslag
12
Förslag till direktiv
Skäl 34
Kommissionens förslag
Ändringsförslag
(34) Eftersom målen för den föreslagna åtgärden, dvs. att garantera såväl en hög säkerhetsnivå för leksaker som en väl fungerande inre marknad genom att fastställa harmoniserade säkerhetskrav för leksaker och minimikrav för marknadsövervakning, inte i tillräcklig utsträckning kan uppnås av de enskilda medlemsstaterna och de därför, på grund av åtgärdens omfattning och verkningar, bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget.
I enlighet med proportionalitetsprincipen i denna artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå dessa mål.
(34) Eftersom målen för den föreslagna åtgärden, dvs. att garantera såväl en hög säkerhetsnivå för leksaker för att säkerställa barns säkerhet och hälsa, som en väl fungerande inre marknad genom att fastställa harmoniserade säkerhetskrav för leksaker och minimikrav för marknadsövervakning, inte i tillräcklig utsträckning kan uppnås av de enskilda medlemsstaterna och de därför, på grund av åtgärdens omfattning och verkningar, bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget.
I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå dessa mål.
Motivering
Man bör påminna om direktivets första målsättning.
Ändringsförslag
13
Kommissionens förslag
Ändringsförslag
1a.
Detta direktiv grundar sig på principen om att tillverkarna, importörerna och de övriga ekonomiska aktörerna intygar att tillverkningen av leksaker eller utsläppandet på marknaden av leksaker, och särskilt de kemiska ämnen som leksakerna innehåller, inte har några skadliga eller giftiga effekter på barns hälsa eller miljön.
Åtgärderna grundar sig på försiktighetsprincipen.
Motivering
I fördragen och den relevanta gemenskapslagstiftningen hänvisas det hela tiden till målsättningen med en hög hälsoskyddsnivå för de berörda personerna och miljön.
Man bör ta samma hänsyn vid översynen av lagstiftningen om leksakers säkerhet inklusive de kemiska ämnen som används för tillverkning av leksaker.
Där är nödvändigt att man därvid påminner om att försiktighetsprincipen bör tas med i lagstiftningen om leksakers säkerhet.
Ändringsförslag
14
Artikel 2 – led 8a (nytt)
Kommissionens förslag
Ändringsförslag
(8a) varningstext: särskild information till slutanvändaren eller den person som har uppsikt över barnet, om säkerhetsaspekterna av villkoren för användning eller montering av en leksak,
Motivering
Det är nödvändigt att definiera begreppet ”varningstext” för att undvika att det blandas ihop med märkningen.
Ändringsförslag
15
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
(9) tillbakadragande: varje åtgärd för att förhindra att en leksak i leveranskedjan tillhandahålls på marknaden,
(9) tillbakadragande: varje åtgärd för att förhindra att en leksak i leveranskedjan tillhandahålls , distribueras, erbjuds eller visas på marknaden,
Motivering
Man måste absolut precisera vilka åtgärder tillbakadragandet täcker exakt.
Ändringsförslag
16
Artikel 2 – led 11a (nytt)
Kommissionens förslag
Ändringsförslag
(11a) asfyxi: blockering av mycket viktiga eller livsviktiga organ på grund av syrebrist, av följande fem olika orsaker: ett föremål i halsen, drunkning, kvävning, strypning eller krossning,
Motivering
Man bör definiera begreppet asfyxi eftersom det står för olika slags fenomen orsakade av syrebrist.
Asfyxi är följden av en av de händelser som framkallar syrebrist och utgör en allvarlig eller livsfarlig risk för barns hälsa.
Ändringsförslag
17
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
(13) skada: kroppsskada eller hälsoskada,
(13) skada: kroppsskada eller annan hälsoskada , inbegripet långvariga skador ,
Motivering
Det är lämpligt att precisera denna definition och ta med de andra skador än fysiska skador som en leksak kan orsaka, samt långvariga skador i samband med användningen av vissa ämnen.
Ändringsförslag
18
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
(14) fara: möjlig källa till skada,
(14) fara: möjlig källa till skada på människors hälsa eller välbefinnande ,
Motivering
Det är nödvändigt att precisera vad som kan skadas.
Ändringsförslag
19
Artikel 2 – led 15 a (nytt)
Kommissionens förslag
Ändringsförslag
15a) ”utformad eller ämnad uttryckligen för barn i åldersgruppen x”: ett begrepp, som betyder, att barnet måste förfoga över sådan händighet och intellektuell förmåga, som motsvarar den avsedda åldersgruppens.
Motivering
Det måste säkerställas att tillverkaren mot bättre vetande inte på etiketten anger en fiktiv åldersgrupp, för att undandra sig vissa bestämda skyldigheter och ansvar.
Ändringsförslag
20
Kommissionens förslag
Ändringsförslag
8.
Tillverkarna ska på begäran ge de behöriga nationella myndigheterna all information och dokumentation som behövs för att visa att leksaken överensstämmer med kraven.
De ska på begäran samarbeta med de behöriga myndigheterna när det gäller de åtgärder som vidtas för att undvika riskerna med de leksaker som de har släppt ut på marknaden.
8.
Tillverkarna ska på begäran , och inom två veckor, ge de behöriga nationella myndigheterna all information och dokumentation som behövs för att visa att leksaken överensstämmer med kraven.
De ska på begäran samarbeta med de behöriga myndigheterna i de åtgärder som vidtas för att undvika riskerna med de leksaker som de har släppt ut på marknaden.
Motivering
Tidsfristerna för tillhandahållande av alla dokument och all information bör anges.
Därmed förbättras tillämpningen av säkerhetsåtgärderna och barnens hälsa säkerställs.
Ändringsförslag
21
Artikel 4 – punkt 1a (ny)
Kommissionens förslag
Ändringsförslag
1a.
Tillverkarna ska informera de nationella behöriga myndigheterna om utnämnanden av representanter på de marknader där leksakerna saluförs senast fyra veckor efter datumet för utnämnandet.
Motivering
Det är nödvändigt att de behöriga nationella myndigheterna får denna information.
Informationen ska ges inom en viss tid.
Ändringsförslag
22
Kommissionens förslag
Ändringsförslag
1b.
Informationen i samband med utnämnandet av en representant ska åtminstone innehålla uppgifter om representanten (namn, adress, telefonnummer, e-postadress och Internetadress), de leksaker för vilka representanten är underställd skyldigheterna i punkt 3 samt leksakernas identifieringsnummer.
Motivering
Ändringsförslag
23
Kommissionens förslag
Ändringsförslag
(b) på begäran ge de nationella behöriga myndigheterna all information och dokumentation som behövs för att visa att leksaken överensstämmer med kraven,
(b) på begäran , och inom två veckor, ge de behöriga nationella myndigheterna all information och dokumentation som behövs för att visa att leksaken överensstämmer med kraven.
Motivering
Tidsfristerna för tillhandahållande av alla dokument och all information bör anges.
Därmed ökas tillämpningen av säkerhetsåtgärderna och barnens hälsa säkerställs.
Ändringsförslag
24
Kommissionens förslag
Ändringsförslag
1.
När importörerna släpper ut en leksak på marknaden ska de iaktta vederbörlig omsorg för att se till att de tillämpliga kraven uppfylls .
1.
Motivering
Det är absolut nödvändigt att ange att även importörerna har en del av ansvaret för att detta direktiv tillämpas och att målsättningarna med omarbetningen av detta direktiv efterlevs.
Ändringsförslag
25
Kommissionens förslag
Ändringsförslag
2.
Innan importörerna släpper ut en leksak på marknaden ska de kontrollera att tillverkaren har utfört bedömningen av överensstämmelse.
2.
Innan importörerna släpper ut en leksak på marknaden ska de kontrollera att tillverkaren har utfört bedömningen av överensstämmelse i enlighet med artiklarna 18 och 19 .
Om en importör upptäcker att leksaken inte överensstämmer med de grundläggande säkerhetskraven i artikel 9 och bilaga II får han eller hon inte släppa ut produkten på marknaden förrän den överensstämmer med dessa krav.
Motivering
Det är nödvändigt att påminna om de relevanta bestämmelser i detta direktiv som de olika punkterna hänvisar till.
Ändringsförslag
26
Kommissionens förslag
Ändringsförslag
3.
Importörerna ska ange namn och en kontaktadress på leksaken eller, om detta inte är möjligt på grund av leksakens storlek eller art, på förpackningen eller i ett medföljande dokument.
3.
Importörerna ska klart och tydligt ange namn samt den adress, det telefonnummer och den e-postadress där de kan nås på leksaken eller, om detta inte är möjligt på grund av leksakens storlek eller art, på förpackningen eller i ett medföljande dokument , på ett sådant sätt att det är tydligt och skilt från beskrivningen av leksaken .
Motivering
De uppgifter som inledningsvis föreslagits bör kompletteras och de bör vara lätt- och snabbtillgängliga.
Ändringsförslag
27
Kommissionens förslag
Ändringsförslag
7.
Importörerna ska på begäran ge de behöriga myndigheterna all information och dokumentation som behövs för att visa att leksaken överensstämmer med kraven.
De ska på begäran samarbeta med de behöriga myndigheterna i de åtgärder som vidtas för att undvika riskerna med de leksaker som de har släppt ut på marknaden.
7.
De ska på begäran samarbeta med de behöriga myndigheterna i de åtgärder som vidtas för att undvika riskerna med de leksaker som de har släppt ut på marknaden.
Motivering
Se ändringsförslag 26.
Ändringsförslag
28
Kommissionens förslag
Ändringsförslag
1.
När distributörerna tillhandahåller en leksak på marknaden ska de iaktta vederbörlig omsorg för att se till att de tillämpliga kraven uppfylls .
1.
Motivering
Se ändringsförslag 27.
Ändringsförslag
29
Kommissionens förslag
Ändringsförslag
5.
Distributörerna ska på begäran ge de nationella behöriga myndigheterna den information och dokumentation som behövs för att visa att leksaken överensstämmer med kraven.
De ska på begäran samarbeta med de behöriga myndigheterna när det gäller de åtgärder som vidtas för att undvika riskerna med de leksaker som de tillhandahållit på marknaden.
5.
De ska på begäran samarbeta med de behöriga myndigheterna i de åtgärder som vidtas för att undvika riskerna med de leksaker som de har släppt ut på marknaden.
Motivering
Se ändringsförslag 26.
Ändringsförslag
30
Förslag till direktiv
Artikel 7a (ny)
Kommissionens förslag
Ändringsförslag
Artikel 7a
Register
De ekonomiska aktörerna i leksakssektorn, enligt definitionen i artikel 1, ska föra ett register över avhjälpande åtgärder, tillbakadraganden från marknaden, återkallelser, reklamationer och klagomål som erhållits från övriga ekonomiska aktörer och slutanvändare samt uppföljningen av de ovan nämnda åtgärderna.
Registret ska behållas i tio år.
Aktörerna ska tillhandahålla de behöriga myndigheterna registren på begäran.
Motivering
Därför är det viktigt att precisera de villkor som tillämpas för förandet av det nämnda registret i detta direktiv.
Ändringsförslag
31
Artikel 8 – stycke 2
Kommissionens förslag
Ändringsförslag
I detta syfte ska de ha system och förfaranden för att på begäran kunna lämna denna information till myndigheterna för marknadsövervakning under en period på tio år.
I detta syfte ska de ha system och förfaranden för att på begäran , och inom två veckor, kunna lämna denna information till myndigheterna för marknadsövervakning under en period på tio år.
Motivering
Se ändringsförslag 23.
Ändringsförslag
32
Artikel 9 – punkt -1 (ny)
Kommissionens förslag
Ändringsförslag
-1.
Det ska erinras om att barn tillhör kategorin sårbara personer eftersom deras hälsa är mer ömtålig och reagerar starkare biologiskt mot vissa ämnens närvaro.
Dessutom är riskerna vid utsatthet för kemiska ämnen större än för vuxna eftersom barn fortfarande utvecklas.
Motivering
Det är tvunget att i denna artikel med mycket viktiga säkerhetskrav påminna om att barn tillhör den befolkningsgrupp som är sårbar eller mycket sårbar beroende på deras ålder.
Det är också nödvändigt att man tar hänsyn till säkerhetskraven och hälsoskyddet för de barn som använder leksakerna, särskilt vad beträffar kemiska ämnen.
Ändringsförslag
33
Kommissionens förslag
Ändringsförslag
Medlemsstaterna ska följa försiktighetsprincipen.
Motivering
Se ändringsförslag 1.
Ändringsförslag
34
Kommissionens förslag
Ändringsförslag
2.
Leksaker får inte innebära en risk för användarens eller någon annan persons säkerhet och hälsa när de används på avsett eller förutsebart sätt med tanke på barns normala beteende.
2.
Hänsyn ska tas till barnets förmåga , och i förekommande fall förmågan hos den som har uppsikt över barnet, att hantera leksaken, särskilt när det gäller leksaker som på grund av sin funktion, storlek och särskilda egenskaper är avsedda för barn under 36 månader.
Hänsyn ska tas till barnets förmåga att hantera leksaken, särskilt när det gäller leksaker som på grund av sin funktion, storlek och särskilda egenskaper är avsedda för barn under 36 månader.
Märkningen på leksaken eller förpackningen samt medföljande bruksanvisning ska varna barnet, eller den som har uppsikt över barnet, för faror och skaderisker som leksaken kan medföra vid användning och upplysa om hur dessa risker kan undvikas.
Motivering
Se ändringsförslag 7 för den första delen av ändringsförslaget.
Vid bedömningen av de mycket viktiga säkerhetskraven kan man inte ta hänsyn till en person som har uppsikt över barnet eftersom det är leksakernas säkerhet i sig som ska bedömas.
Man bör ha uppsikt över barnen, men detta kan inte ske jämt, eftersom barn bör kunna och behöver leka ensamma för att utvecklas och bli självständiga.
Ändringsförslag
35
Kommissionens förslag
Ändringsförslag
3.
Leksaker som släpps ut på marknaden ska uppfylla de grundläggande säkerhetskraven under hela den tid som de normalt sett förväntas användas.
3.
Motivering
Se ändringsförslag 2.
Ändringsförslag
36
Kommissionens förslag
Ändringsförslag
Varningstexterna i del B punkt 1 i bilaga V får inte användas för leksaker som med hänsyn till funktion, mått eller andra egenskaper än vikten, är avsedda för barn under 36 månader.
Motivering
Leksaker för barn under tre år är ofta märkta med ”ej för barn under tre år” även om de är avsedda för den ålderskategorin.
Vissa tillverkare försöker på så sätt komma undan sitt ansvar eller friskriva sig från rättsliga påföljder.
Eftersom det i bilaga V inte uttryckligen står att det är förbjudet att märka leksaker med denna text är det mycket lättare i marknadsövervakningshänseende att se till att lagstiftningen följs genom att denna bestämmelse tas med i direktivet.
Ändringsförslag
37
Kommissionens förslag
Ändringsförslag
För de kategorier av leksaker som förtecknas i del B i bilaga V ska de varningstexter som anges där användas.
Motivering
I överensstämmelse med ändringsförslag 102.
Det är även lämpligt att ange bestämmelsens räckvidd.
Ändringsförslag
38
Förslag till direktiv
2.
För små leksaker som säljs utan förpackning ska lämpliga varningstexter finnas på själva leksaken.
2.
Varningstexter ska vara avfattade på ett exakt, synligt, tydligt och lättläst sätt samt vara begripliga för användarna eller de personer som övervakar användarna.
De ska fästas på leksaken eller, om detta inte är tekniskt möjligt , på en etikett fäst vid leksaken eller på konsumentförpackningen .
Varningstexter ska upprepas i den bruksanvisning som medföljer leksaken.
För små leksaker som säljs utan förpackning ska lämpliga varningstexter finnas på själva leksaken.
Varningstexter som anger användarnas lägsta eller högsta tillåtna ålder ska vara synliga och lättlästa och placerade på ett iögonfallande sätt på försäljningsstället.
Varningstexter som anger användarnas lägsta eller högsta tillåtna ålder ska vara synliga , tydliga, lättlästa och exakta samt placerade på ett iögonfallande sätt på leksaksförpackningen och på försäljningsstället.
Tillverkarens representant, importörer och distributörer ska informeras om dessa varningstexter, så att man placerar de varningstexter som anger användarnas lägsta och högsta tillåtna ålder på ett korrekt sätt på försäljningsstället.
Varningstexter ska alterneras på ett sådant sätt att de förekommer regelbundet.
Varningstexten ska tryckas på styckförpackningens mest synliga yta och på alla yttre omslag som förekommer vid detaljförsäljning av varan, med undantag av genomskinliga ytteromslag.
Medlemsstaterna får bestämma var på dessa ytor varningstexten ska placeras med tanke på de krav som språken ställer.
För att kunna beakta de krav som språken ställer ska medlemsstaterna ha rätt att bestämma storleken på typsnittet, förutsatt att den typsnittsstorlek som fastställs i deras lagstiftning gör varningstexten mycket lättläst och tydlig.
Varningstexten ska tryckas på det/de officiella språket/språken i den medlemsstat där leksaken släpps ut på marknaden.
Ändringsförslag
39
Kommissionens förslag
Ändringsförslag
3.
Medlemsstaterna får kräva att varningstexter eller säkerhetsanvisningar, eller en del av dem , finns på deras officiella språk när leksakerna släpps ut på marknaden på deras territorium.
3.
Varningstexter , i enlighet med vad som anges i denna artikel och i bilaga V, och säkerhetsanvisningar ska finnas på den berörda medlemsstatens officiella språk när leksakerna släpps ut på marknaden på statens territorium.
Motivering
Avfattandet av varningstexter och säkerhetsanvisningar på det eller de officiella språk som finns i medlemsstaten där leksakerna släpps ut på marknaden är en viktig del för barns säkerhet och hälsa.
Ändringsförslag
40
Förslag till direktiv
Artikel 10b (ny)
Kommissionens förslag
Ändringsförslag
Artikel 10b
Gemensamma bestämmelser för ekonomiska aktörer om åtgärder för tillbakadragande av leksaker med bristande överensstämmelse eller förmodad bristande överensstämmelse
1.
I enlighet med artiklarna 3, 5 och 6 ska de ekonomiska operatörer som har problem med leksaker med bristande överensstämmelse eller förmodad bristande överensstämmelse med bestämmelserna om säkra leksaker omedelbart vidta åtgärder för tillbakadraganden av leksakerna.
2.
De ekonomiska operatörer som har problem med leksaker med bristande överensstämmelse eller förmodad bristande överensstämmelse med bestämmelserna om säkra leksaker ska omedelbart informera de andra ekonomiska aktörerna, konsumentorganisationerna och de nationella myndigheterna i de medlemsstater de har tillhandahållit leksaken och ge en detaljerad beskrivning av i synnerhet problemet med bristande överensstämmelse och de åtgärder för tillbakadragande som vidtagits.
3.
Åtgärderna för tillbakadragande ska vidtas omedelbart och utföras så fort som möjligt, senast inom två veckor efter att den bristande överensstämmelsen har konstaterats.
Om åtgärder inte kan vidtas inom ovannämnda tidsfrist, ska de ekonomiska aktörer som har problem med bristande överensstämmelse omedelbart informera de andra berörda ekonomiska aktörerna och de ansvariga nationella myndigheterna.
De ansvariga nationella myndigheterna ska så fort som möjligt besluta om en begäran om ytterligare en tidsfrist och omedelbart informera de berörda ekonomiska aktörerna om beslutet, i synnerhet om den eventuella tidsfrist som krävs för åtgärdande av bristande överensstämmelse för berörda leksaker.
4.
Saluföringen av leksakerna till slutanvändarna ska avbrytas på obestämd tid.
Efter att den bristande överensstämmelsen åtgärdats för de leksaker som dragits tillbaka från marknaden, ska dessa leksaker anses som nya, och de ska stämma överens med alla bestämmelser i detta direktiv när de på nytt tillhandahålls slutanvändarna.
Motivering
Det är nödvändigt att precisera bestämmelserna om åtgärderna för tillbakadragande som nämns i artiklarna 3, 5 och 6 i detta direktiv.
Dessa preciseringar går hand i hand med förstärkningen av bestämmelserna om säkra leksaker och barns hälsa.
De närmare bestämmelserna för tillbakadragande ska vara kraftfullare än de korrigerande åtgärderna eftersom leksakernas säkerhet och barnens hälsa kan påverkas på ett allvarligare sätt.
Ändringsförslag
41
Artikel 17 – stycke 1a (nytt)
Kommissionens förslag
Ändringsförslag
Vid bedömningen av leksakernas säkerhet ska man ta hänsyn till alla relevanta aspekter, i synnerhet de barn eller barngrupper som är särskilt sårbara eller som har en ovanlig åkomma, till exempel barn med särskilda behov.
Motivering
Förutom att det handlar om att återkalla det föremål som är viktigt för bedömningen, är det också nödvändigt att precisera kompletterande aspekter av denna, särskilt att även beakta barn med olika funktionsnedsättningar.
Ändringsförslag
42
Artikel 17 – stycke 1b (nytt)
Kommissionens förslag
Ändringsförslag
Det är nödvändigt att beakta samtliga olyckor, även små och mindre allvarliga, som barn råkar ut för, när risk- och farlighetsnivåerna för leksakerna fastställs.
Motivering
Detta ändringsförslag syftar till att olyckor med inte alltför allvarlig utgång och framför allt småolyckor i större omfattning beaktas, så att olycksbenägenheten i samband med leksaker återges på ett korrektare sätt.
Ändringsförslag
43
Kommissionens förslag
Ändringsförslag
3.
När ett organ för bedömning av överensstämmelse som anmälts enligt artikel 21 (nedan kallat anmält organ) utför EG-typkontrollen ska den vid behov och tillsammans med tillverkaren utvärdera tillverkarens analys enligt artikel 17 av de faror som leksaken kan medföra.
3.
När ett organ för bedömning av överensstämmelse som anmälts enligt artikel 21 (nedan kallat anmält organ) utför EG-typkontrollen ska den tillsammans med tillverkaren utvärdera tillverkarens analys enligt artikel 17 av de faror som leksaken kan medföra.
Motivering
Denna bedömning kan inte vara frivillig med tanke på syftet att förstärka leksakernas säkerhet.
Ändringsförslag
44
Kommissionens förslag
Ändringsförslag
Intyget ska ses över när det anses nödvändigt, särskilt när leksakens tillverkningsprocess, utgångsmaterial eller ingående delar ändras, men i alla händelser vart femte år.
Motivering
Tidsfristen måste minskas med tanke på syftet att förstärka leksakernas säkerhet.
Ändringsförslag
45
Artikel 20 – punkt -1 (ny)
Kommissionens förslag
Ändringsförslag
-1.
Motivering
Det finns anledning att precisera i denna artikel att den tekniska dokumentationen måste finnas tillgänglig för all inspektion eller kontroll hos leksakstillverkaren.
Ändringsförslag
46
Kommissionens förslag
Ändringsförslag
Om en myndighet för marknadsövervakning begär att få den tekniska dokumentationen eller en översättning av delar av den från en tillverkare kan den fastställa en tidsfrist för detta som ska vara 30 dagar, såvida inte en kortare tidsfrist är berättigad på grund av en allvarlig eller omedelbar risk.
På begäran av behöriga nationella myndigheter ska tillverkaren eller dennes representant tillhandahålla den tekniska dokumentationen eller en översättning av delar av den inom en tidsfrist på högst 14 dagar, såvida inte en kortare tidsfrist är berättigad på grund av en allvarlig eller omedelbar risk.
Motivering
Det är nödvändigt att vara mer precis och omgående fastställa tidsfristen för överlämnandet av dokumentationen.
Detta förstärker leksakernas säkerhet och gör det möjligt att bättre garantera barnens säkerhet och hälsa vilket är målet med denna omarbetning.
Ändringsförslag
47
Kommissionens förslag
Ändringsförslag
4.
Om tillverkaren inte uppfyller sina skyldigheter enligt punkterna 1, 2 och 3 får myndigheten för marknadsövervakning begära att tillverkaren på egen bekostnad låter ett anmält organ utföra en provning av leksaken inom en viss föreskriven tid för att kontrollera att den uppfyller de harmoniserade standarderna och grundläggande säkerhetskraven.
4.
Ändringsförslag
48
Kommissionens förslag
Ändringsförslag
4a.
Om tillverkaren inte uppfyller sina skyldigheter enligt punkt 4 ska myndigheten för marknadsövervakning vidta de åtgärder som man anser nödvändiga för att tillse att leksakerna inte tillhandahålls på marknaden och i distributionsnätet på det territorium som myndigheten övervakar.
Motivering
Den föreliggande artikeln är ofullständig.
Om tillverkaren inte respekterar de skyldigheter som åligger denne, ska behöriga nationella myndigheter vidta åtgärder som gör det möjligt att garantera barnens säkerhet och hälsa.
Ändringsförslag
49
Kommissionens förslag
Ändringsförslag
3a.
Den anmälande myndigheten ska sätta upp ställen för säkerhetsanmälningar dit konsumenter och människor som arbetar med barn kan rapportera in leksaker som inte följer bestämmelserna eller olyckor som är relaterade till användningen av en leksak.
Motivering
Genom att sätta upp ställen för säkerhetsanmälningar i medlemsstaterna skulle man ge konsumenterna inflytande och underlätta direkt kommunikation med tillverkare och producenter ifall det finns problem med en särskild produkt.
Tillverkare och producenter skulle då kunna reagera mer direkt på konsumenternas krav.
Ändringsförslag
50
Kommissionens förslag
Ändringsförslag
(a) fullgod teknisk och yrkesinriktad utbildning som täcker all slags bedömning av överensstämmelse på det område inom vilket organet för bedömning av överensstämmelse har anmälts,
(a) fullgod teknisk och yrkesinriktad utbildning , som ska bevisas genom, bland annat, formella meriter, yrkeserfarenhet eller intyg, som täcker all slags bedömning av överensstämmelse på det område inom vilket organet för bedömning av överensstämmelse har anmälts,
Motivering
Det är nödvändigt att intyga den tekniska och yrkesinriktade utbildningen hos personalen i de anmälda organen.
Ändringsförslag
51
Kommissionens förslag
Ändringsförslag
11a.
Organet för bedömning av överensstämmelse ska ha som mål att bli certifierad enligt ISO 9001, version 2000.
Motivering
Denna certifiering är en extra garanti för bedömningens kvalitet och respekten för standarderna när denna genomförs.
Ändringsförslag
52
Kommissionens förslag
Ändringsförslag
4a.
Dotterbolagen och underentreprenörerna ska vara certifierade enligt ISO 9001, version 2000.
Motivering
Denna certifiering är en extra garanti för kvaliteten på tillverkningsprocesserna samt den regelbundna bedömningen och kontrollerna av dessa.
Ändringsförslag
53
Kommissionens förslag
Ändringsförslag
3a.
För övervakning av leksaker som släpps ut på marknaden i enlighet med artikel 37 får myndigheterna för marknadsövervakning, eller något annat anmält organ till vilket myndigheterna ger uppdraget, utföra icke planerade kontroller i de ekonomiska aktörernas lokaler en gång om året om det är möjligt och minst vartannat år.
Motivering
Ändringsförslag
54
Kommissionens förslag
Ändringsförslag
1.
Om en medlemsstats myndigheter för marknadsövervakning har vidtagit åtgärder enligt artikel 12 i direktiv 2001/95/EG eller om de har tillräckliga skäl att anta att en leksak som omfattas av det här direktivet utgör en risk för människors hälsa eller säkerhet, ska de tillsammans med de berörda ekonomiska aktörerna utvärdera leksaken med avseende på alla de krav som fastställs i det här direktivet.
1.
Om en medlemsstats myndigheter för marknadsövervakning har vidtagit åtgärder enligt artikel 12 i direktiv 2001/95/EG eller om de misstänker att en leksak som omfattas av det här direktivet kan utgöra en risk för människors hälsa eller säkerhet, ska de omedelbart utföra alla nödvändiga bedömningar av leksaken med avseende på alla de krav som fastställs i det här direktivet.
De ekonomiska aktörerna ska inom två veckor tillhandahålla myndigheterna all information eller alla handlingar de ber om.
Om myndigheterna för marknadsövervakning vid utvärderingen konstaterar att en leksak inte uppfyller kraven i detta direktiv ska de ålägga de berörda ekonomiska aktörerna att vidta lämpliga korrigerande åtgärder för att leksaken ska uppfylla dessa krav eller dra tillbaka leksaken från marknaden eller återkalla den inom en rimlig tid som de fastställer i förhållande till typen av risk .
Om myndigheterna för marknadsövervakning vid utvärderingen konstaterar att en leksak inte uppfyller kraven i detta direktiv ska de ålägga de berörda ekonomiska aktörerna att vidta lämpliga korrigerande åtgärder för att leksaken ska uppfylla dessa krav eller dra tillbaka leksaken från marknaden eller återkalla den inom den tidsfrist som anges i artiklarna 10a, 10b och 10c .
Motivering
Alla problem med överensstämmelse skall omedelbart bedömas.
De ekonomiska aktörernas medverkan ska begränsas till att de tillhandahåller information för bedömningen av leksaken i fråga.
Om överensstämmelsen inte har respekterats, ska lämpliga korrigerande åtgärder i förhållande till det konstaterade problemet genomföras inom utsatt tid.
Ändringsförslag
55
Kommissionens förslag
Ändringsförslag
Om myndigheterna för marknadsövervakning vid utvärderingen konstaterar att en leksak inte uppfyller kraven i detta direktiv ska de ålägga de berörda ekonomiska aktörerna att vidta lämpliga korrigerande åtgärder för att leksaken ska uppfylla dessa krav eller dra tillbaka leksaken från marknaden eller återkalla den inom en rimlig tid som de fastställer i förhållande till typen av risk
Om myndigheterna för marknadsövervakning vid utvärderingen konstaterar att en leksak inte uppfyller kraven i detta direktiv ska de, samtidigt som ett meddelande går ut till konsumenterna, ålägga de berörda ekonomiska aktörerna att vidta lämpliga korrigerande åtgärder för att leksaken ska uppfylla dessa krav eller dra tillbaka leksaken från marknaden eller återkalla den inom en rimlig tid som de fastställer i förhållande till typen av risk
Motivering
Den direkta informationen till konsumenterna utgör en avgörande förutsättning för att säkerställa att en fara undviks.
Ändringsförslag
56
Kommissionens förslag
Ändringsförslag
2.
Om myndigheterna för marknadsövervakning anser att den bristande överensstämmelsen inte bara gäller det nationella territoriet, ska de informera kommissionen och de andra medlemsstaterna om utvärderingsresultaten och om de åtgärder som de har ålagt de ekonomiska aktörerna att vidta
2.
Om myndigheterna för marknadsövervakning anser att den bristande överensstämmelsen inte bara gäller det nationella territoriet, ska de informera kommissionen och de andra medlemsstaterna om utvärderingsresultaten och om de åtgärder som de har ålagt de ekonomiska aktörerna att vidta.
De ska officiellt informera medlemsstaterna och kommissionen om det svar och den vilja att åtgärda den bristande överensstämmelsen eller att inte göra det som den ekonomiske aktören har meddelat.
Motivering
Inom ramarna för öppenhet och full upplysning av allmänheten, ska en ekonomisk aktör vara tvungen att svara och svaret ska komma medlemsstaterna och kommissionen tillhanda.
Ändringsförslag
57
Kommissionens förslag
Ändringsförslag
3.
De ekonomiska aktörerna ska se till att det vidtas korrigerande åtgärder i fråga om alla berörda leksaker som de har tillhandahållit på gemenskapsmarknaden.
3.
Den berörda ekonomiska aktören eller de berörda ekonomiska aktörerna ska se till att det vidtas korrigerande åtgärder , tillbakadragande eller återkallelse i fråga om alla berörda leksaker som de har tillhandahållit på gemenskapsmarknaden.
Motivering
Det finns anledning att vara precis och alltså inkludera alla ekonomiska aktörer och alla verksamheter som berörs av de åtgärder som ska vidtas om överensstämmelse med regelverket inte föreligger.
Ändringsförslag
58
Kommissionens förslag
Ändringsförslag
4.
4.
Motivering
Se ändringsförslag 64.
Ändringsförslag
59
Kommissionens förslag
Ändringsförslag
7.
Åtgärden ska anses vara motiverad om ingen medlemsstat eller kommissionen har rest invändningar inom tre månader efter mottagandet av den information som avses i punkt 4 mot en provisorisk åtgärd som vidtagits av en medlemsstat med avseende på den berörda leksaken.
7.
Åtgärden ska anses vara motiverad om ingen medlemsstat eller kommissionen har rest invändningar inom fyra veckor efter mottagandet av den information som avses i punkt 4 mot en provisorisk åtgärd som vidtagits av en medlemsstat med avseende på den berörda leksaken.
Motivering
De åtgärder som föreslagits av behöriga nationella myndigheter ska behandlas av andra myndigheter och kommissionen inom en rimlig tidsfrist i syfte att fatta beslut om de åtgärder i samband med bristande överensstämmelse som den behöriga nationella myndigheten begärt att de ekonomiska aktörer som berörs av leksaken i fråga ska vidta.
Ändringsförslag
60
Kommissionens förslag
Ändringsförslag
2.
Om den nationella åtgärden anses vara motiverad ska alla medlemsstater vidta de åtgärder som krävs för att säkerställa att den leksak som inte uppfyller kraven dras tillbaka från deras marknader.
Medlemsstaterna ska underrätta kommissionen om detta.
2.
Om den nationella åtgärden anses vara motiverad ska alla medlemsstater vidta de åtgärder som krävs för att säkerställa att den leksak som inte uppfyller kraven dras tillbaka eller återkallas från deras marknader.
Medlemsstaterna skall underrätta kommissionen om detta.
Motivering
Se ändringsförslag 64.
Ändringsförslag
61
Kommissionens förslag
Ändringsförslag
3.
3.
Motivering
Bristerna när det gäller en harmoniserad standard avseende leksakernas överensstämmelse och säkerhet ska korrigeras så snabbt som möjligt.
Ändringsförslag
62
Kommissionens förslag
Ändringsförslag
2.
Om det fortfarande råder sådan bristande överensstämmelse som avses i punkt 1 ska medlemsstaten vidta lämpliga åtgärder för att begränsa eller förbjuda tillhandahållandet av leksaken på marknaden eller se till att den återkallas eller dras tillbaka från marknaden.
2.
Om det fortfarande råder sådan bristande överensstämmelse som avses i punkt 1 ska medlemsstaten omedelbart vidta lämpliga åtgärder för att begränsa eller förbjuda tillhandahållandet av leksaken på marknaden eller se till att den återkallas eller dras tillbaka från marknaden.
Motivering
Man bör så snabbt som möjligt garantera leksakernas säkerhet och barnens hälsa.
Ändringsförslag
63
Kommissionens förslag
Ändringsförslag
1.
Kommissionen kan ändra följande bestämmelser i syfte att anpassa dem till den tekniska och vetenskapliga utvecklingen:
1.
Kommissionen ska ändra följande bestämmelser i syfte att anpassa dem till den tekniska och vetenskapliga utvecklingen så fort som man får in nya uppgifter :
(-a) Bilaga I.
(a) Punkterna 7 och 8 i del III i bilaga II.
(a) Del III i bilaga II , med undantag för punkterna 1 och 2 .
(b) Bilaga V.
(b) Bilaga V.
Motivering
Det beslutade kommittéförfarandet kan bara tillämpas för dessa punkter.
Det bör utvidgas till att omfatta andra frågor eftersom standardiserings- eller harmoniseringsförfarandet är för långsamt för brådskande ändringar, vilket visas av de faror och risker som magneter utgör för barns hälsa.
Ändringsförslag
64
Kommissionens förslag
Ändringsförslag
Motivering
(Berör inte den svenska versionen.)
Ändringsförslag
65
Kommissionens förslag
Ändringsförslag
1a.
– fastställa gränsvärden eller andra restriktioner för ämnen eller preparat som utgör en fara för hälsan utöver de som listas i leden 7 och 8 i del III i bilaga II,
– införa eller anpassa gränsvärden för buller och hastigheter.
Motivering
Kommissionen bör ges befogenhet att införa nya restriktioner för nya ämnen eller bullergränsvärden inom ramarna för kommittéförfarandet.
Ändringsförslag
66
Förslag till direktiv
Artikel 47
Kommissionens förslag
Ändringsförslag
Rapporten ska innehålla en utvärdering av dels situationen när det gäller leksakers säkerhet, dels hur verkningsfullt detta direktiv är samt en beskrivning av marknadsövervakningen i medlemsstaten.
Rapporten ska innehålla en utvärdering av dels situationen när det gäller leksakers säkerhet, dels hur verkningsfullt detta direktiv är samt en beskrivning av marknadsövervakningen i medlemsstaten.
Kommissionen ska utarbeta och offentliggöra en sammanfattning av de nationella rapporterna .
Kommissionen ska utarbeta och offentliggöra en rapport så fort som möjligt med, i tillämpliga fall, förslag till ändring eller omarbetning av detta direktiv .
Kommissionen ska överlämna rapporten till Europaparlamentet och rådet.
Kommissionen ska omedelbart offentliggöra åtminstone en sammanfattning och slutsatserna i rapporten på sin webbplats på Europeiska unionens samtliga officiella språk.
Motivering
Kommissionen ska utarbeta en rapport om utvärderingsrapporterna om tillämpningen av detta direktiv i medlemsstaterna.
Kommissionen ska utan dröjsmål överlämna den till de två lagstiftningsorganen och offentliggöra rapporten i sin helhet, eller åtminstone en sammanfattning och slutsatserna, på sin webbplats.
I detta ändringsförslag begärs alltså att minimiåtgärderna när det gäller insyn tillämpas.
Ändringsförslag
67
Artikel 50 – stycke 1
Kommissionens förslag
Ändringsförslag
Medlemsstaterna ska fastställa regler för påföljder, även straffrättsliga påföljder för allvarliga överträdelser, vid överträdelser av de nationella bestämmelser som antas i enlighet med detta direktiv och de ska vidta alla åtgärder som krävs för att säkerställa att påföljderna verkställs.
Påföljderna ska vara effektiva, proportionella och avskräckande.
Motivering
Det är nödvändigt men otillräckligt att medlemsstaterna fastställer påföljderna för överträdelser av bestämmelserna i detta direktiv.
De måste också kunna tillämpa dem för att förverkliga dessa påföljder.
Ändringsförslag
68
Förslag till direktiv
Artikel 52
Kommissionens förslag
Ändringsförslag
Medlemsstaterna får inte förhindra att leksaker som överensstämmer med direktiv 88/378/EEG och som släpptes ut på marknaden innan det här direktivet trädde i kraft eller senast två år efter ikraftträdandet släpps ut på marknaden
Medlemsstaterna får inte förhindra att leksaker som överensstämmer med direktiv 88/378/EEG och som släpptes ut på marknaden innan det här direktivet trädde i kraft eller senast tre år efter ikraftträdandet släpps ut på marknaden.
Ändringsförslag
69
Förslag till direktiv
Artikel 54a (ny)
Kommissionens förslag
Ändringsförslag
Artikel 54a
Översyn
Kommissionen ska vart åttonde år se över detta direktiv, baserat på den behöriga vetenskapliga kommitténs bedömningar och expertgruppens utlåtande.
Motivering
En revidering av direktivet, åtminstone vart åttonde år eller tidigare om nödvändigt på grund av nya upptäckter eller olyckor, behövs för att säkerställa att säkerhetskrav i direktivet är tillräckliga för att täcka de risker som kan uppstå genom t.ex. nya leksaker och ny teknik, men även genom nya vetenskapliga rön.
Ändringsförslag
70
Förslag till direktiv
Bilaga II – del I – punkt 2
Kommissionens förslag
Ändringsförslag
2.
Åtkomliga kanter, utskjutande partier, rep, snören, kablar och fästanordningar ska vara utformade och konstruerade på ett sådant sätt att risken för kroppsskada vid kontakt minimeras.
2.
Åtkomliga kanter, utskjutande partier, rep, snören, kablar och fästanordningar ska vara utformade och konstruerade på ett sådant sätt att risken för kroppsskada vid kontakt minimeras så mycket som möjligt .
Motivering
Det är nödvändigt att minska riskerna i detta sammanhang så långt som möjligt för att förbättra leksakernas säkerhet och garantera barnens integritet och hälsa.
Ändringsförslag
71
Förslag till direktiv
Bilaga II – del I – led 4 – stycke 2
Kommissionens förslag
Ändringsförslag
Ändringsförslag
72
Förslag till direktiv
Bilaga II – del I – punkt 5
Kommissionens förslag
Ändringsförslag
5.
Leksaker avsedda att användas på grunt vatten och till att hålla barn över vatten eller stödja dem ska vara utformade och konstruerade så att risken för sämre flytkraft eller stöd för barnet begränsas så långt möjligt med hänsyn till rekommenderat användningssätt.
5.
Leksaker avsedda att användas på grunt vatten och till att hålla barn över vatten eller stödja dem ska vara utformade och konstruerade så att risken för sämre flytkraft eller stöd för barnet begränsas maximalt med hänsyn till ett rekommenderat och i möjligaste mån förutsägbart användningssätt.
Motivering
Se ändringsförslag 74 respektive 2.
Ändringsförslag
73
Förslag till direktiv
Bilaga II – del I – punkt 7 – stycke 1
Kommissionens förslag
Ändringsförslag
7.
Leksaker med vars hjälp användaren kan förflytta sig ska så långt möjligt vara försedda med broms, anpassad till typ av leksak och till den rörelseenergi som leksaken utvecklar.
Bromssystemet ska vara enkelt att använda utan risk för att användaren kastas ur leksaken eller att denne eller andra personer skadas.
7.
Leksaker med vars hjälp användaren kan förflytta sig ska vara försedda med broms, anpassad till typ av leksak och till den rörelseenergi som leksaken utvecklar.
Bromssystemet ska vara enkelt att använda utan risk för att användaren kastas ur leksaken eller att denne eller andra personer skadas.
Motivering
Avsaknad av bromssystem eller ett otillräckligt sådant gäller en betydande del av de leksaker som är försedda med hjul.
Det finns därför anledning att vara striktare för att förbättra säkerheten när det gäller barns användning av denna typ av leksaker.
Ändringsförslag
74
Förslag till direktiv
Bilaga II – del I – led 10
Kommissionens förslag
Ändringsförslag
10) Ljudleksaker ska vara utformade och konstruerade så att ljudet inte skadar barnens hörsel.
Detta ska gälla alla leksaker oavsett vilken åldersgrupp de är avsedda för.
Gränser för ihållande buller ska sättas baserat på örats känslighet för ett litet barn som är under 36 månader gammalt.
Motivering
Nuvarande normer för bullergränser hanterar inte på ett betryggande sätt möjligheterna att barns hörsel skadas.
För det första gäller normerna inte för alla leksaker (normen för ”nära örat-leksaker” gäller exempelvis endast barn under 10 månaders ålder).
För det andra, behöver en lägre gräns sättas för impulsljud.
Med tanke på den verkliga livssituationen för barn i olika åldrar inom en familj, bör bullernivåer sättas baserat på de mest sårbara, dvs. barn under 36 månaders ålder.
Ändringsförslag
75
Förslag till direktiv
Bilaga II – del I – punkt 11
Kommissionens förslag
Ändringsförslag
11.
Aktivitetsleksaker ska vara utformade så att risken att klämma sig eller fastna med kroppsdelar eller kläder och risken att falla, kollidera eller drunkna minimeras.
11.
Aktivitetsleksaker ska vara utformade så att risken att klämma sig eller fastna med kroppsdelar eller kläder och risken att falla, kollidera eller drunkna minimeras så mycket som möjligt .
Motivering
Se ändringsförslag 74.
Ändringsförslag
76
Förslag till direktiv
Bilaga II – del III – punkt 1
Kommissionens förslag
Ändringsförslag
1.
1.
Motivering
Se ändringsförslag 3.
Ändringsförslag
77
Förslag till direktiv
Bilaga II – del III – punkt 3
Kommissionens förslag
Ändringsförslag
3.
3.
Användningen i leksaker av ämnen som är klassificerade som cancerframkallande, mutagena eller reproduktionstoxiska (CMR) kategori 3 enligt direktiv 67/548/EEG i koncentrationer som var för sig är lika med eller högre än 0,1 procent ska vara förbjuden.
Motivering
Förekomsten av ämnen som är klassificerade som CMR över det uppsatta tröskelvärdet bör förbjudas för att säkra en hög nivå på skyddet av barnens hälsa.
Detta tröskelvärde bör sänkas genom ett kommittéförfarande så fort som möjligt, på grundval av ny information.
Ändringsförslag
78
Förslag till direktiv
Bilaga II – del III – punkt 4
Kommissionens förslag
Ändringsförslag
4.
Ämnen eller preparat som klassificeras som CMR-ämnen i kategori 1 och 2 enligt direktiv 67/548/EEG får användas i leksaker om följande villkor är uppfyllda:
4.
Ämnen eller preparat som klassificeras som CMR-ämnen i kategori 1 , 2 och 3 enligt direktiv 67/548/EEG får användas i leksaker om följande villkor är uppfyllda:
Motivering
Användningen av dessa kan bara motiveras om de villkor som är uppräknade i styckena i punkt 4 är uppfyllda.
Ändringsförslag
79
Förslag till direktiv
Bilaga II – del III – punkt 4.2
Kommissionens förslag
Ändringsförslag
4.2.
Motivering
Det är nödvändigt att precisera det som ersättningen täcker.
Ändringsförslag
80
Förslag till direktiv
Bilaga II – del III – punkt 4.3a (ny)
Kommissionens förslag
Ändringsförslag
4.3a.
Leksaker eller delar av leksaker som är avsedda att stoppas i munnen, måste, oavsett viken åldersgrupp som de är avsedda för, uppfylla de bestämmelser för överföringsgränsvärden som gäller för livsmedelsförpackningar i Europaparlamentets och rådets förordning (EG) nr 1935/2004 av den 27 oktober 2004 om material och produkter avsedda att komma i kontakt med livsmedel.
Ändringsförslag
81
Förslag till direktiv
Motivering
En ny bedömning av dessa ämnen eller preparat ska äga rum oftare.
Ändringsförslag
82
Förslag till direktiv
Bilaga II – del III – punkt 4a (ny)
Kommissionens förslag
Ändringsförslag
4a.
Ämnen som klassificeras som farliga för det endokrina systemet och som står med på EU:s lista över prioriterade ämnen är förbjudna att användas i leksaker och leksakernas beståndsdelar förutom om tillverkaren bevisar att det inte finns några ersättningsämnen som är säkrare eller mindre skadliga för hälsan.
Motivering
Ämnen som klassificeras som farliga för det endokrina systemet utgör en allvarlig risk för barns utveckling och deras hälsa i vuxen ålder.
Det finns också anledning att slå fast principen om förbud för dessa samtidigt som man tillåter att de används om det inte finns några ersättningsämnen som är säkrare eller mindre skadliga för hälsan, vilket tillverkaren ska bevisa.
Ändringsförslag
83
Förslag till direktiv
Bilaga II – del III – punkt 4b (ny)
Kommissionens förslag
Ändringsförslag
4b.
Ämnen som klassificeras som persistenta, bioackumulerande eller toxiska (PBT) eller mycket persistenta och mycket bioackumulerande (vPvB) är förbjudna att användas i leksaker och leksakernas beståndsdelar förutom om tillverkaren bevisar att det inte finns några ersättningsämnen som är säkrare eller mindre skadliga för hälsan.
Motivering
Se ändringsförslag 87 när det här gäller ämnen som klassificeras som PBT och vPvB.
Ändringsförslag
84
Förslag till direktiv
Bilaga II – del III – punkt 5
Kommissionens förslag
Ändringsförslag
5.
utgår
Motivering
Ändringsförslag
85
Förslag till direktiv
Bilaga II – del III – led 5a och 5b (nya)
Kommissionens förslag
Ändringsförslag
5a) Leksaker eller delar av leksaker måste, oavsett viken åldersgrupp som de är avsedda för, uppfylla de bestämmelser om utlösning av nitrosaminer och nitroserbara ämnen från nappar av elastomer eller gummi som fastställts i kommissionens direktiv 93/11/EEG av den 15 mars 1993 om utlösning av N-nitrosaminer och N-nitroserbara ämnen från dinappar och tröstnappar av elastomer eller gummi.
Programmet ska ta hänsyn till rapporter från marknadsövervakande organ och till synpunkter som medlemsstater och intressenter ger uttryck för.
Kommissionen ska besluta, med ledning av den behöriga vetenskapliga kommitténs åsikt, att vidta lämpliga restriktiva åtgärder, om nödvändigt.
Motivering
Användningen av farliga ämnen i leksaker är inte begränsad till CMR-ämnen, doftämnen eller ämnen som innehåller vissa beståndsdelar.
Alla farliga ämnen bör regelbundet utvärderas av kommissionen.
Skulle det vid denna utvärdering avslöjas en oacceptabel risk, bör kommissionen ges befogenhet att vidta lämpliga åtgärder inom ramen för kommittéförfarandet.
Ändringsförslag
86
Förslag till direktiv
Bilaga II – del III – punkt 7
Kommissionens förslag
Ändringsförslag
7.
Leksaker får inte innehålla följande allergiframkallande doftämnen:
7.
Leksaker får inte innehålla följande allergiframkallande doftämnen .
1) Ålandsrot (Inula helenium)
1) Ålandsrot (Inula helenium)
2) Allylisotiocyanat
2) Allylisotiocyanat
3) Bensylcyanid
3) Bensylcyanid
4) 4-Tert-butylfenol
4) 4-Tert-butylfenol
5) Chenopodiumolja
5) Chenopodiumolja
6) Cyklamenalkohol
6) Cyklamenalkohol
7) Dietylmaleat
7) Dietylmaleat
8) Dihydrokumarin
8) Dihydrokumarin
9) 2,4-Dihydroxi-3-metylbensaldehyd
9) 2,4-Dihydroxi-3-metylbensaldehyd
10) 3,7-Dimetyl-2-okten-1-ol (6,7‑dihydrogeraniol)
10) 3,7-Dimetyl-2-okten-1-ol (6,7‑dihydrogeraniol)
11) 4,6-Dimetyl-8-tert-butylkumarin
11) 4,6-Dimetyl-8-tert-butylkumarin
12) Dimetylcitrakonat
12) Dimetylcitrakonat
13) 7,11-Dimetyl-4,6,10-dodekatrien-3-on
13) 7,11-Dimetyl-4,6,10-dodekatrien-3-on
14) 6,10-Dimetyl-3,5,9-undekatrien-2-on
14) 6,10-Dimetyl-3,5,9-undekatrien-2-on
15) Difenylamin
15) Difenylamin
16) Etylakrylat
16) Etylakrylat
17) Fikonblad, färska och beredda
17) Fikonblad, färska och beredda
18) Trans-2-heptenal
18) Trans-2-heptenal
19) Trans-2-hexenaldietylacetal
19) Trans-2-hexenaldietylacetal
20) Trans-2-hexenaldimetylacetal
20) Trans-2-hexenaldimetylacetal
21) Hydroabietylalkohol
21) Hydroabietylalkohol
22) 4-Etoxifenol
22) 4-Etoxifenol
23) 6-lsopropyl-2-dekahydronaftalenol
23) 6-lsopropyl-2-dekahydronaftalenol
24) 7-Metoxikumarin
24) 7-Metoxikumarin
25) 4-Metoxifenol
25) 4-Metoxifenol
26) 4-(p-Metoxifenyl)-3-buten-2-on
26) 4-(p-Metoxifenyl)-3-buten-2-on
27) 1-(p-Metoxifenyl)-1-penten-3-on
27) 1-(p-Metoxifenyl)-1-penten-3-on
28) Metyl-trans-2-butenoat
28) Metyl-trans-2-butenoat
29) 6-Metylkumarin
29) 6-Metylkumarin
30) 7-Metylkumarin
30) 7-Metylkumarin
31) 5-Metyl-2,3-hexanedion
31) 5-Metyl-2,3-hexanedion
32) Costusrotolja (Saussurea lappa Clarke)
32) Costusrotolja (Saussurea lappa Clarke)
33) 7-Etoxi-4-metylkumarin
33) 7-Etoxi-4-metylkumarin
34) Hexahydrokumarin
34) Hexahydrokumarin
35) Perubalsam (Myroxylon pereirae Klotzsch)
35) Perubalsam (Myroxylon pereirae Klotzsch)
36) 2-Pentyliden-cyklohexanon
36) 2-Pentyliden-cyklohexanon
37) 3,6,10-Trimetyl-3,5,9-undekatrien-2-on
37) 3,6,10-Trimetyl-3,5,9-undekatrien-2-on
38) Citronverbenaolja (Lippia citriodora Kunth)
38) Citronverbenaolja (Lippia citriodora Kunth)
Spår av dessa ämnen ska dock tillåtas förutsatt att förekomsten är tekniskt oundviklig med god tillverkningssed
Dessutom ska följande allergiframkallande doftämnen anges om de används i leksaker i koncentrationer över 0,01 viktprocent
1) Amylkanelaldehyd
39) Amylkanelaldehyd
2) Amylkanelalkohol
40) Amylkanelalkohol
3) Anisylalkohol
41) Anisylalkohol
4) Bensylalkohol
42) Bensylalkohol
5) Bensylbensoat
43) Bensylbensoat
6) Bensylcinnamat
44) Bensylcinnamat
7) Bensylsalicylat
45) Bensylsalicylat
8) Kanelaldehyd
46) Kanelaldehyd
9) Kanelalkohol
47) Kanelalkohol
10) Citral
48) Citral
11) Citronellol
49) Citronellol
12) Kumarin
50) Kumarin
13) Eugenol
51) Eugenol
14) Farnesol
52) Farnesol
15) Geraniol
53) Geraniol
16) Hexylkanelaldehyd
54) Hexylkanelaldehyd
17) Hydroxicitronellal
55) Hydroxicitronellal
18) Hydroxi-metylpentylcyklohexenkarboxaldehyd
56) Hydroxi-metylpentylcyklohexenkarboxaldehyd
19) Isoeugenol
57) Isoeugenol
20) Lilial (i kosmetikadirektivet upptaget i post 83 som 2-(4-tert-butylbensyl)-propionaldehyd)
58) Lilial (i kosmetikadirektivet upptaget i post 83 som 2-(4-tert-butylbensyl)-propionaldehyd)
21) d-Limonen
59) d-Limonen
22) Linalol
60) Linalol
23) Metylheptinkarbonat
61) Metylheptinkarbonat
24) 3-Metyl-4-(2,6,6-trimetyl-2-cyklohexen-1-yl)-3-buten-2-on
62) 3-Metyl-4-(2,6,6-trimetyl-2-cyklohexen-1-yl)-3-buten-2-on
25) Ekmosseextrakt
63) Ekmosseextrakt
26) Trämosseextrakt
64) Trämosseextrakt
Ändringsförslag
87
Förslag till direktiv
Bilaga II – del III – punkt 7a (ny)
Kommissionens förslag
Ändringsförslag
7a.
Leksaker som är avsedda att ofta komma i kontakt med huden, t.ex. fingerfärg eller modellera, ska uppfylla kraven på sammansättning och märkning i direktiv 76/768/EEG.
Motivering
För leksaker som ofta kommer i kontakt med huden ska samma stränga bestämmelser tillämpas som dem som föreskrivs i direktivet för kosmetikaprodukter.
Ändringsförslag
88
Förslag till direktiv
Bilaga II – del III – punkt 7b (ny)
Kommissionens förslag
Ändringsförslag
7b.
Leksaker som är avsedda att ofta komma i kontakt med huden och som innehåller andra allergiframkallande ämnen än doftämnen som är kända för att framkalla allvarliga eller till och med dödliga reaktioner hos barn (t.ex. dem som framkallar en anafylaktisk chock) ska uppfylla bestämmelserna om märkning i kommissionens direktiv 2006/125/EG av den 5 december 2006 om spannmålsbaserade livsmedel och barnmat för spädbarn och småbarn 1 .
________________
16.
Motivering
Närvaron av andra allergiframkallande ämnen än doftämnen ska alltså bli föremål för märkning.
Ändringsförslag
89
Förslag till direktiv
Bilaga II – del III – punkt 7c (ny)
Kommissionens förslag
Ändringsförslag
7.c Användningen av allergiframkallande doftämnen är tillåten i luktleksaker och vetenskapsleksaker.
Luktleksaker och vetenskapsleksaker måste uppfylla kraven på sammansättning i direktiv 76/768/EEG och bestämmelserna i del III punkt 6 i bilaga II.
Allergiframkallande doftämnen som används i dessa två leksakskategorier måste märkas som allergiframkallande på ett sätt som skiljer dem från andra använda doftämnen och med en exakt, väl synlig och lättläst information, i syfte att upplysa konsumenterna om användningen och förekomsten av allergiframkallande doftämnen.
Kommissionen kan anmoda den behöriga vetenskapliga kommittén att fastställa koncentrationsgränsvärdena för de allergiframkallande doftämnen som används i dessa två leksakskategorier.
Den behöriga vetenskapliga kommittén måste lämna sitt utlåtande inom tre månader.
Flaskor som innehåller doftämnen i dessa två leksakskategorier ska förses med en anordning vid öppningen som kräver att ett särskilt verktyg används för att ta mycket små prover av de flytande ämnena eller pulverämnena/doftämnena och därmed undvika risken att dessa ämnen/doftämnen sväljs i annat än små kvantiteter.
Leksaker som omfattas av denna punkt är förbjudna för barn under sex års ålder.
De leksaker som omfattas av denna punkt definieras enligt följande:
a) en luktleksak är en leksak för att lära sig att känna igen eller urskilja olika lukter eller smaker från basämnen eller parfymextrakt,
b) en vetenskapsleksak är en leksak för att lära sig framställa produkter från basämnen eller parfymextrakt och andra råvaror än parfymämnen.
Ändringsförslag
90
Förslag till direktiv
Bilaga II – del III – punkt 8 – inledningen
Kommissionens förslag
Ändringsförslag
1.
8.
Följande gränsvärden för migration får inte överskridas i någon leksakskomponent .
Motivering
Bestämmelserna för gränser för överföring måste vara striktare i syfte att förverkliga målet att förbättra leksakernas säkerhet och hålla en hög skyddsnivå för barns hälsa.
Ändringsförslag
91
Förslag till direktiv
Bilaga II – del III – punkt 8 – tabellrubrik – kolumn 2
Kommissionens förslag
Ändringsförslag
mg/kg i torrt, sprött, pulverliknande eller böjligt leksaksmaterial
mg/kg i fast, torrt, sprött, pulverliknande eller böjligt leksaksmaterial
Motivering
Det finns anledning att vara precis och täcka alla typer av material som används i leksakstillverkningen i syfte att förverkliga målet att förbättra leksakernas säkerhet och hålla en hög skyddsnivå för barns hälsa.
Ändringsförslag
92
Förslag till direktiv
Bilaga II – del III – punkt 8 – tabellen
Kommissionens förslag
Grundämne
mg/kg i torrt, sprött, pulverliknande eller böjligt leksaksmaterial
mg/kg
i vätskeformigt eller klibbigt leksaksmaterial
Aluminium
5 625
1 406
Antimon
45
11,3
Arsenik
7,5
1,9
Barium
4 500
1 125
Bor
1 200
300
Kadmium
3,8
0,9
Krom (III)
37,5
9,4
Krom (VI)
0,04
0,01
Kobolt
10,5
2,6
Koppar
622,5
156
Bly
27
6,8
Mangan
1 200
300
Kvicksilver
15
3,8
Nickel
75
18,8
Selen
37,5
9,4
Strontium
4 500
1 125
Tenn
15 000
3 750
Organiskt tenn
1,9
0,5
Zink
3 750
938
Ändringsförslag från parlamentet
Grundämne
mg/kg i fast, torrt, sprött, pulverliknande eller böjligt leksaksmaterial
mg/kg
i vätskeformigt eller klibbigt leksaksmaterial
Aluminium
5 625
1 406
Antimon
45
11,3
utgår
utgår
utgår
Barium
4 500
1 125
Bor
1 200
300
utgår
utgår
utgår
Krom (III)
37,5
9,4
utgår
utgår
utgår
Kobolt
10,5
2,6
Koppar
622,5
156
utgår
utgår
utgår
Mangan
1 200
300
utgår
utgår
utgår
Nickel
75
18,8
Selen
37,5
9,4
Strontium
4 500
1 125
Tenn
15 000
3 750
utgår
utgår
utgår
Zink
3 750
938
Motivering
Arsenik, kadmium, bly, krom (VI), kvicksilver och organiskt tenn är mycket toxiska.
Kadmium, bly, krom (VI) och kvicksilver är redan förbjudna i bilar och elektriska och elektroniska apparater.
Krom (VI) i cement behöver reduceras till en oskadlig form genom tillsats av järnsulfat.
Det är uppenbart att ämnen som är baserade på dessa beståndsdelar inte bör användas i leksaker.
Det finns anledning att vara precis och täcka alla typer av material som används i leksakstillverkningen i syfte att förverkliga målet att förbättra leksakernas säkerhet och hålla en hög skyddsnivå för barns hälsa.
Ändringsförslag
93
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
utgår
Motivering
Den sista punkten behöver också utgå eftersom den tillåter alltför stora undantag från CMR-förbudet.
Ändringsförslag
94
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
Användning i leksaker eller i leksakskomponenter av ämnen eller preparat som är baserade på någon av de följande beståndsdelarna ska förbjudas:
1) Arsenik
2) Kadmium
3) Krom (V)
4) Bly
5) Kvicksilver
6) Organiskt tenn
Motivering
Arsenik, kadmium, bly, krom (VI), kvicksilver och organiskt tenn är mycket toxiska.
Kadmium, bly, krom (VI) och kvicksilver är redan förbjudna i bilar och elektriska och elektroniska apparater.
Krom (VI) i cement behöver reduceras till en oskadlig form genom tillsats av järnsulfat.
Det är uppenbart att ämnen som är baserade på dessa beståndsdelar inte bör användas i leksaker.
Ändringsförslag
95
Förslag till direktiv
Bilaga II – del III – punkt 8a (ny)
Kommissionens förslag
Ändringsförslag
8a.
Leksaker eller delar av leksaker som är avsedda att stoppas i munnen, måste, oavsett viken åldersgrupp som de är avsedda för, uppfylla de bestämmelser för överföringsgränsvärden som gäller för livsmedelsförpackningar i Europaparlamentets och rådets förordning (EG) nr 1935/2004 av den 27 oktober 2004 om material och produkter avsedda att komma i kontakt med livsmedel.
Ändringsförslag
96
Förslag till direktiv
Bilaga II – del V
Kommissionens förslag
Ändringsförslag
1.
Leksaker ska vara utformade och tillverkade så att de uppfyller kraven på hygien och renlighet för att undvika infektion, sjukdom och smitta.
1.
Leksaker ska vara utformade och tillverkade så att de uppfyller kraven på hygien och renlighet för att undvika infektion, sjukdom och smitta.
Leksaker ska gå att tvätta, skrubba eller desinficera utan att leksakernas funktionsduglighet eller säkerhet förändras.
2.
Tygleksaker för barn under 36 månader ska gå att tvätta och ska uppfylla säkerhetskraven även efter tvätt.
2.
Tygleksaker för barn under 36 månader ska gå att tvätta och ska uppfylla kraven på funktionsduglighet och säkerhet även efter tvätt.
Motivering
En hög nivå på hygienen ska vara förenlig med garantin för leksakernas funktionsduglighet och säkerhet.
Ändringsförslag
97
Förslag till direktiv
Bilaga IV – led a
Kommissionens förslag
Ändringsförslag
a) Ingående beskrivning av konstruktion och tillverkning, inklusive en lista på delar och material som använts i leksakerna samt kemikalieleverantörens säkerhetsdatablad för de kemikalier som använts;
a) Ingående beskrivning av konstruktion och tillverkning, inklusive en lista på delar , material och råvaror som använts i leksakerna liksom även detaljerad information om de kemikalier som använts i leksakerna och leksakskomponenterna, samt de använda kvantiteterna.
Motivering
Detta är ett tillägg till ändringsförslag 100 av föredraganden för att även inkludera information om råvaror.
Testresultaten gällande kemikalier kan variera avsevärt från parti till parti på grund av användningen av olika råvaror.
Det är därför viktigt att information om råvaror också tillhandahålls.
Ändringsförslag
98
Förslag till direktiv
Bilaga V – del B – punkt 1 – stycke 2
Kommissionens förslag
Ändringsförslag
Varningstexterna ska kompletteras med en kortfattad upplysning , som kan finnas i bruksanvisningen, om vilka specifika faror som ligger till grund för åldersgränsen.
Varningstexterna ska kompletteras med en kortfattad upplysning om de specifika faror som ligger till grund för åldersgränsen.
Upplysningen ska vara lättläst och sitta klart synlig på leksaken eller, om detta är tekniskt omöjligt, på en etikett fäst vid leksaken eller på förpackningen, och i bruksanvisningen .
För små leksaker utan förpackning ska dessa upplysningar finnas på själva leksaken.
Motivering
Förslagets bestämmelser är inte tillräckligt precisa och tvingande.
Ändringsförslaget syftar till att göra de bestämmelser som ändrats här tydligare och lättbegripligare.
Ändringsförslag
99
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
Motivering
Förslagets bestämmelser är inte tillräckligt precisa.
Den föreslagna texten är förenlig med tillämpningsområdet för detta förslag men den varnar inte i tillräcklig grad för en fara eller en risk.
Ändringsförslag
100
Förslag till direktiv
Bilaga V – del B – punkt 2 – stycke 2a (nytt)
Kommissionens förslag
Ändringsförslag
Motivering
Det måste tydligt klargöras att det är nödvändigt att läsa instruktionerna innan man börjar montera eller sätta ihop leksaken, så att personen som utför uppgiften vet hur denne ska agera för att undvika skador.
Ändringsförslag
101
Förslag till direktiv
Kommissionens förslag
Ändringsförslag
”Tillsyn av en vuxen rekommenderas ”
” Innehåller en leksak som endast får användas under tillsyn av en vuxen” .
Motivering
Den föreslagna texten varnar inte i tillräcklig grad för en fara eller en risk.
Den ska tydligt varsko om de åtgärder som ska vidtas.
ÄRENDETS GÅNG
Titel
Leksakers säkerhet
Referensnummer
KOM(2008)0009 – C6-0039/2008 – 2008/0018(COD)
Ansvarigt utskott
IMCO
Yttrande
Tillkännagivande i kammaren
ENVI
11.3.2008
Föredragande av yttrande
Utnämning
Anne Ferreira
7.3.2008
Behandling i utskott
15.7.2008
8.9.2008
Antagande
7.10.2008
Slutomröstning: resultat
+:
–:
0:
45
6
2
Slutomröstning: närvarande ledamöter
Adamos Adamou, Georgs Andrejevs, Margrete Auken, Liam Aylward, Pilar Ayuso, Irena Belohorská, Johannes Blokland, John Bowis, Frieda Brepoels, Hiltrud Breyer, Martin Callanan, Dorette Corbey, Avril Doyle, Mojca Drčar Murko, Jill Evans, Anne Ferreira, Elisabetta Gardini, Matthias Groote, Satu Hassi, Gyula Hegyi, Jens Holm, Marie Anne Isler Béguin, Dan Jørgensen, Christa Klaß, Urszula Krupa, Marie-Noëlle Lienemann, Peter Liese, Jules Maaten, Marios Matsakis, Linda McAvan, Roberto Musacchio, Riitta Myller, Miroslav Ouzký, Vladko Todorov Panayotov, Vittorio Prodi, Frédérique Ries, Guido Sacconi, Daciana Octavia Sârbu, Amalia Sartori, Bogusław Sonik, María Sornosa Martínez, Salvatore Tatarella, Thomas Ulmer, Anja Weisgerber, Åsa Westlund, Glenis Willmott
Slutomröstning: närvarande suppleanter
Iles Braghetto, Antonio De Blasio, Bairbre de Brún, Caroline Lucas, Miroslav Mikolášik
Slutomröstning: närvarande suppleanter (art.
178.2)
Pervenche Berès, Dieter-Lebrecht Koch
till utskottet för den inre marknaden och konsumentskydd
över förslaget till Europaparlamentets och rådets direktiv om leksakers säkerhet
( KOM(2008)0009 – C6‑0039/2008 – 2008/0018(COD) )
Föredragande:
David Hammerstein
KORTFATTAD MOTIVERING
Behovet av särskilda bestämmelser för leksaksindustrin resulterade i direktivet om leksakers säkerhet, vilket antogs i maj 1988.
Direktivet har onekligen varit till stor nytta för industrin sedan det infördes.
Återkallandet av miljoner leksaker från ledande tillverkare 2007 var dock ett tydligt bevis på att bestämmelserna i direktivet från 1988 inte var i fas med den dynamiska och snabba utvecklingen inom leksaksindustrin och att den aktuella lagstiftningen inte kunde hantera de problem som uppstod inom detta område.
Som ett svar på den snabba utvecklingen och den ökande oron bland konsumenter över säkerheten för leksaker som tillverkats i Europa lade kommissionen i januari 2008 fram ett förslag till ett omarbetat direktiv för leksakers säkerhet som syftar till att införa bestämmelser gällande:
Ett förtydligande av direktivets tillämpningsområde och begrepp – beträffande de produkter som inte omfattas av direktivet och en förteckning över de begrepp som förekommer i direktivet.
Föredraganden välkomnar initiativet till den mycket välbehövliga revideringen av direktivet om leksakers säkerhet.
Förslaget går i rätt riktning genom att stärka aktuella åtgärder och introducera nya för alla de områden som blivit kritiserade i syfte att reglera leksakers säkerhet i Europa.
För att garantera den högsta nivån av skydd för barn behöver dock vissa åtgärdskategorier utredas ytterligare utifrån hur ingående de är.
Leksakers kemiska egenskaper: Cancerframkallande ämnen (alla CMR-ämnen i kategori 1, 2 och 3) såväl som farliga ämnen utgör en mycket allvarlig risk för barns hälsa.
Obotliga och negativa hälsoeffekter uppkommer kanske inte alltid över en natt utan snarare efter en längre tids exponering av sådana ämnen.
Det är även allmänt känt att vissa doftämnen orsakar allergier som är relativt svåra att behandla.
Föredraganden anser därför att man ska vidta så strama åtgärder som möjligt för att minska hälsoriskerna genom att införa ett allmänt förbud mot CMR-ämnen i kategori 1 och 2 samt ett förbud mot ämnen i kategori 3 men med möjlighet till undantag för vissa ämnen.
Alla doftämnen samt de farliga ämnena arsenik, kvicksilver, bly, organiskt tenn, kadmium och krom IV ska också förbjudas.
Förfarande för säkerhetsbedömning: Förfarandet för säkerhetsbedömning är ett av de viktigaste momenten för att säkerställa en hög säkerhetsnivå för leksaker på marknaden och bör därför stärkas.
Utan att för den delen belasta industrin måste det införas krav på EG‑typkontroller för åtminstone de farligaste leksakskategorierna och årliga stickprovskontroller inom dessa kategorier för att garantera att det även genomförs regelbundna säkerhetskontroller efter den första prototyptesten.
Flexibla bestämmelser: Leksaksindustrin har visat sig vara ytterst dynamisk och snabb när det gäller att ta fram nya produkter och ny produktdesign och använda sig av nya material osv. De nya bestämmelserna i det reviderade direktivet måste därför formuleras på ett sådant sätt att de snabbt kan anpassas till oförutsedda risker och utvecklingar så att man kan undvika ödesdigra misstag som skulle ha kunnat förhindras genom snabba åtgärder (snarare än en snabb reaktion) från tillverkarnas, lagstiftarnas och de brottsbekämpande myndigheternas sida.
Det föreskrivande förfarandet med kontroll ska följaktligen tillämpas oftare och ha en framträdande roll på följande områden: ändring av gränsvärdena för leksakers fysikaliska egenskaper (hastighet, buller, temperatur), ändring av förteckningen över de produkter som enligt direktivet inte räknas som leksaker och ändring av förteckningen över de leksaker som omfattas av de fyra farligaste leksakskategorierna och som ska genomgå EG-typkontroll.
ÄNDRINGSFÖRSLAG
Utskottet för industrifrågor, forskning och energi uppmanar utskottet för den inre marknaden och konsumentskydd att som ansvarigt utskott infoga följande ändringsförslag i sitt betänkande:
Ändringsförslag
1
Förslag till direktiv
Skäl 3a (nytt)
Kommissionens förslag
Ändringsförslag
(3a) En annan viktig målsättning med det nya system som inrättas genom detta direktiv är att stimulera och i vissa fall se till att farliga ämnen och material som används i leksaker ersätts med mindre farliga ämnen eller tekniker om det finns lämpliga alternativ som är ekonomiskt och tekniskt genomförbara.
Motivering
Detta ändringsförslag är en anpassning till Reach-förordningen (skäl 12).
Ändringsförslag
2
Förslag till direktiv
Skäl 8
Kommissionens förslag
Ändringsförslag
(8) Alla ekonomiska aktörer som ingår i leverans- och distributionskedjan bör vidta åtgärder för att se till att de endast tillhandahåller sådana leksaker på marknaden som överensstämmer med den tillämpliga lagstiftningen.
I detta direktiv görs en tydlig och proportionell fördelning av skyldigheterna som svarar mot varje aktörs roll i leverans- och distributionsprocessen.
(8) Detta direktiv bygger på principen att alla ekonomiska aktörer som ingår i leverans- och distributionskedjan bör tillverka, importera eller släppa ut leksaker på marknaden med det ansvar och den försiktighet som krävs för att garantera att barns säkerhet och hälsa under normala och rimligen förutsebara användningsförhållanden inte påverkas negativt.
De ekonomiska aktörerna bör vidta åtgärder för att se till att de endast tillhandahåller sådana leksaker på marknaden som överensstämmer med den tillämpliga lagstiftningen.
I detta direktiv görs en tydlig och proportionell fördelning av skyldigheterna som svarar mot varje aktörs roll i leverans- och distributionsprocessen.
Motivering
Detta ändringsförslag inför skyldigheten för ekonomiska aktörer att iaktta försiktighet.
Det är en anpassning som inspirerats av bestämmelserna i Reach-förordningen (skäl 16).
Ändringsförslag
3
Förslag till direktiv
Skäl 16
Kommissionens förslag
Ändringsförslag
(16) För att barnen ska skyddas mot nyupptäckta risker måste nya grundläggande säkerhetskrav också antas.
Det är särskilt nödvändigt att komplettera och uppdatera bestämmelserna om kemikalier i leksaker.
Dessa bestämmelser bör ange att leksaker bör överensstämma med den allmänna kemikalielagstiftningen, särskilt Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 om registrering, utvärdering, godkännande och begränsning av kemikalier (Reach), inrättande av en europeisk kemikaliemyndighet, ändring av direktiv 1999/45/EG och upphävande av rådets förordning (EEG) nr 793/93 och kommissionens förordning (EG) nr 1488/94 samt rådets direktiv 76/769/EEG och kommissionens direktiv 91/155/EEG, 93/67/EEG, 93/105/EG och 2000/21/EG.
Bestämmelserna bör emellertid också anpassas till barns särskilda behov eftersom de är sårbar konsumenter.
De specifika gränsvärden som anges i direktiv 88/378/EEG för vissa ämnen bör uppdateras mot bakgrund av nya vetenskapliga rön.
Nya grundläggande säkerhetskrav måste också antas.
Det är särskilt nödvändigt att komplettera och uppdatera bestämmelserna om kemikalier i leksaker.
Dessa bestämmelser bör ange att leksaker bör överensstämma med den allmänna kemikalielagstiftningen, särskilt Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 om registrering, utvärdering, godkännande och begränsning av kemikalier (Reach), inrättande av en europeisk kemikaliemyndighet, ändring av direktiv 1999/45/EG och upphävande av rådets förordning (EEG) nr 793/93 och kommissionens förordning (EG) nr 1488/94 samt rådets direktiv 76/769/EEG och kommissionens direktiv 91/155/EEG, 93/67/EEG, 93/105/EG och 2000/21/EG.
Bestämmelserna bör emellertid också anpassas till barns särskilda behov eftersom de är sårbara konsumenter.
Det bör därför införas nya begränsningar för ämnen som klassificeras som CMR-ämnen enligt direktiv 67/548/EEG av den 27 juni 1967 om tillnärmning av lagar och andra författningar om klassificering, förpackning och märkning av farliga ämnen och doftämnen i leksaker, med tanke på att dessa ämnen kan utgöra en särskild hälsorisk.
De specifika gränsvärden som anges i direktiv 88/378/EEG för vissa ämnen bör uppdateras mot bakgrund av nya vetenskapliga rön.
Motivering
Detta ändringsförslag uppmärksammar betydelsen av att ta upp ämnen med särskilt farliga egenskaper.
Detta ändringsförslag är en anpassning till Reach-förordningen (skäl 69).
Ändringsförslag
4
Förslag till direktiv
Skäl 16a (nytt)
Kommissionens förslag
Ändringsförslag
Motivering
Man måste undvika att olika EU-organ gör samma utvärdering av ett ämne som ska användas i leksaker.
Ändringsförslag
5
Förslag till direktiv
Skäl 16b (nytt)
Kommissionens förslag
Ändringsförslag
Motivering
Enligt förslaget får medlemsstaterna inte förhindra att leksaker som uppfyller kraven i det nuvarande direktivet 88/378/EEG om leksakers säkerhet ”senast två år efter ikraftträdandet” släpps ut på marknaden.
Detta innebär att medlemsstater får besluta att tillämpa de nya bestämmelserna i direktivet efter det att direktivet trätt i kraft.
Av rättssäkerhetsskäl är det viktigt att en sådan situation inte uppstår.
Ändringsförslag
6
Artikel 2 – led 3a (nytt)
Kommissionens förslag
Ändringsförslag
(3a) Tillverkarens representant: varje fysisk eller juridisk person etablerad inom gemenskapen som tillverkaren skriftligen utsett till sin företrädare att i dennes ställe utföra specificerade uppgifter som följer av tillverkarens skyldigheter enligt detta direktiv.
Motivering
En definition av begreppet ”tillverkarens representant” behöver läggas till i artikel 2.
Ändringsförslag
7
Kommissionens förslag
Ändringsförslag
7.
Tillverkare som anser eller har skäl att tro att en leksak som de har släppt ut på marknaden inte överensstämmer med den tillämpliga gemenskapslagstiftningen ska antingen vidta de korrigerande åtgärder som krävs för att få leksaken att överensstämma med kraven eller i förekommande fall dra tillbaka leksaken från marknaden och återkalla den från slutanvändarna.
De ska omedelbart underrätta de nationella myndigheterna i de medlemsstater där de har tillhandahållit leksaken, och lämna detaljerade uppgifter om i synnerhet den bristande överensstämmelsen och de korrigerande åtgärder som vidtagits.
7.
Tillverkare som anser eller har skäl att tro att en leksak som de har släppt ut på marknaden inte överensstämmer med den tillämpliga gemenskapslagstiftningen ska antingen vidta de korrigerande åtgärder som krävs för att få leksaken att överensstämma med kraven eller i förekommande fall dra tillbaka leksaken från marknaden och återkalla den från slutanvändarna.
De ska omedelbart underrätta de nationella myndigheterna i de medlemsstater där de har tillhandahållit leksaken, och lämna detaljerade uppgifter om i synnerhet den bristande överensstämmelsen och de korrigerande åtgärder som vidtagits.
Tillverkare ska omedelbart skjuta upp utsläppandet på marknaden av leksakerna till dess att de uppfyller kraven i den tillämpliga gemenskapslagstiftningen.
Ändringsförslag
8
Kommissionens förslag
Ändringsförslag
Tillverkarens representant
Skyldigheter för tillverkarens representant
1.
Tillverkarna får genom skriftlig fullmakt utse en fysisk eller juridisk person som är etablerad i gemenskapen (nedan kallad tillverkarens representant) att i deras ställe utföra specificerade uppgifter som följer av tillverkarnas skyldigheter enligt detta direktiv .
1.
Motivering
För att titeln ska överensstämma med artiklarna 3 och 5.
En definition av begreppet ”tillverkarens representant” har lagts till i artikel 2.
Ändringsförslag
9
Kommissionens förslag
Ändringsförslag
3.
Medlemsstaterna får kräva att varningstexter eller säkerhetsanvisningar , eller en del av dem, finns på deras officiella språk när leksakerna släpps ut på marknaden på deras territorium.
3.
Medlemsstaterna ska kräva att alla varningstexter eller säkerhetsanvisningar finns på deras officiella språk när leksakerna släpps ut på marknaden på deras territorium.
Motivering
Det är inte tillåtet att ange säkerhetsinformation som är viktig för konsumenten på ett annat språk än det officiella språket på den marknad där produkten släpps ut.
Ändringsförslag
10
Kommissionens förslag
Ändringsförslag
1.
Kommissionen kan ändra följande bestämmelser i syfte att anpassa dem till den tekniska och vetenskapliga utvecklingen:
1.
Kommissionen kan ändra följande bestämmelser i syfte att anpassa dem till den tekniska , vetenskapligt möjliga utvecklingen:
(a) Punkterna 7 och 8 i del III i bilaga II.
(a) Punkterna 7 och 8 i del III i bilaga II.
(b) Bilaga V.
(b) Bilaga V.
Motivering
Den vetenskapliga kommittén måste vara delaktig i översynen av Bilaga II och V för vetenskaplig och teknisk rådgivning mot bakgrund av den vetenskapliga utvecklingen.
Ändringsförslag
11
Kommissionens förslag
Ändringsförslag
2.
Kommissionen får besluta att ämnen eller preparat som enligt bilaga I till direktiv 67/548/EEG klassificerats som cancerframkallande, mutagena eller reproduktionstoxiska i kategori 1, 2 eller 3 får användas i leksaker.
2.
Kommissionen får besluta att ämnen eller preparat som enligt bilaga I till direktiv 67/548/EEG klassificerats som cancerframkallande, mutagena eller reproduktionstoxiska i kategori 1, 2 eller 3 får ingå i leksaker.
Motivering
Den vetenskapliga kommittén måste vara delaktig i översynen av Bilaga II och V för vetenskaplig och teknisk rådgivning mot bakgrund av den vetenskapliga utvecklingen.
Ändringsförslag
12
Förslag till direktiv
Artikel 52
Kommissionens förslag
Ändringsförslag
Medlemsstaterna får inte förhindra att leksaker som överensstämmer med direktiv 88/378/EEG och som släpptes ut på marknaden innan det här direktivet trädde i kraft eller senast två år efter ikraftträdandet släpps ut på marknaden.
Motivering
Det är viktigt att detta direktiv träder i kraft samtidigt i alla medlemsstater.
Ytterligare en period är nödvändig för att centrala organ ska få tid på sig att ta fram nya tester och för att näringslivet ska kunna uppfylla nya tekniska krav på kemikalier.
Ändringsförslag
13
Förslag till direktiv
Bilaga I – punkt 17a (ny)
Kommissionens förslag
Ändringsförslag
17a.
Böcker som inte innehåller andra delar eller föremål (annat än av papper eller papp).
Motivering
Vissa medlemsstater har i samband med genomförandet av direktivet om leksakers säkerhet från 1988 kommit att betrakta barnböcker som leksaker.
I flera medlemsstater har detta resulterat i att de som publicerar barnböcker drabbats av stora problem.
Eftersom böcker är viktiga, framför allt för små barn för att förbättra deras läsförmåga, är det viktigt att man även fortsättningsvis främjar läsandet.
Därför bör man när det gäller detta direktiv inte betrakta böcker som leksaker förutsatt att de inte har en uppenbar funktion som leksak.
Ändringsförslag
14
Förslag till direktiv
Bilaga II – del I – punkt 4 – stycke 2
Kommissionens förslag
Ändringsförslag
Förpackningarna i vilka leksakerna saluförs i detaljhandeln får inte medföra risk för strypning eller kvävning genom att täppa till munnen och näsan.
Förpackningarna i vilka leksakerna saluförs i detaljhandeln får inte medföra risk för strypning eller kvävning genom att på inre och yttre väg täppa till munnen och näsan.
Ändringsförslag
15
Förslag till direktiv
Bilaga II – del III – punkt 3
Kommissionens förslag
Ändringsförslag
3.
3.
Ämnen som klassificeras som cancerframkallande, mutagena eller reproduktionstoxiska i kategorierna 1 eller 2 enligt bilaga 1 i direktiv 67/548/EEG i koncentrationer som var för sig är lika med eller högre än de relevanta koncentrationer som enligt direktiv 1999/45/EG fastställts för klassificeringen av preparat som innehåller ämnena i fråga ska, utan att det påverkar tillämpningen av begränsningarna i punkt 2 första meningen, inte ingå i leksaker, utom om ämnena förekommer i leksakernas beståndsdelar som barn inte kan komma åt i enlighet med standard EN 71 .
Motivering
Om man inte kan komma åt CMR-ämnen i kategori 1 och 2 (dvs. ingen exponering) innebär det inga risker att använda leksakerna.
Säkerheten kommer inte att förbättras för att man utökar begränsningen till delar av leksaker som inte går att komma åt.
För en bättre definiering av begreppet är det viktigt att införa definitionen åtkomst i enlighet med EU‑standarden EN 71.
Ändringsförslag
16
Förslag till direktiv
Bilaga II – del III – punkt 4 – inledningen
Kommissionens förslag
Ändringsförslag
4.
Ämnen eller preparat som klassificeras som CMR-ämnen i kategori 1 och 2 enligt direktiv 67/548/EEG får användas i leksaker om följande villkor är uppfyllda:
4.
Ämnen som klassificeras som CMR‑ämnen i kategori 1 och 2 i bilaga I i direktiv 67/548/EEG får användas i leksaker om följande villkor är uppfyllda:
Motivering
Strykningen av ordet preparat och tillägget av bilaga I behövs för att förtydliga rättsläget.
Ändringsförslag
17
Förslag till direktiv
Bilaga II – del III – punkt 4 – led 4.1
Kommissionens förslag
Ändringsförslag
4.1.
Tillverkare kan i detta syfte, innan den övergångsperiod som avses i artikel 52 löper ut, lämna in begäran till kommissionen om att den behöriga vetenskapliga kommittén ska göra en utvärdering av de risker som ämnen som klassificeras som CMR-ämnen i kategori 1 och 2 enligt bilaga I i direktiv 67/548/EEG utgör.
En sådan begäran ska åtföljas av relevant information, särskilt i fråga om exponering.
När en begäran kommit in ska kommissionen omedelbart ge den vetenskapliga kommittén i uppdrag att avge ett yttrande.
Tillverkarna får, fram till dess att ett beslut antagits, fortsätta att släppa ut leksaker på marknaden som innehåller ämnen som klassificeras som CMR ‑ämnen i kategori 1 och 2 enligt bilaga I i direktiv 67/548/EEG för vilka en begäran har lämnats in.
Motivering
Man vinner inget säkerhetsmässigt på att tillämpa begränsningar på inre delar av leksaker.
Det är i standarden som alla tekniska detaljer om leksakers säkerhet utarbetas, inbegripet sannolikheten för att de ska gå sönder.
Det är därför vi rekommenderar att definitionen av åtkomst är den som fastställs i standarden.
När beståndsdelarna inte exponeras föreligger ingen risk för barns hälsa.
Ändringsförslag
18
Förslag till direktiv
Bilaga II – del III – punkt 4 – led 4.2
Kommissionens förslag
Ändringsförslag
utgår
Motivering
Kravet på att en kemikalie ska ersättas därför att det finns ett alternativ bör strykas för att främja barns säkerhet.
Om riskbedömningen visar att ämnet inte utgör någon risk för barn, finns det ingen anledning att man ska experimentera med nya kemikalier med risk för att det material där det ingår ändras.
Barns säkerhet beror först och främst på hur säkert det material som används för att konstruera en leksak är, t.ex. om plasten kommer att spricka eller gå i bitar.
Säkerheten ökar därför när man använder material som uppfyller kraven i inarbetade tester.
Ändringsförslag
19
Förslag till direktiv
Bilaga II – del III – punkt 5
Kommissionens förslag
Ändringsförslag
5.
5.
Leksaker ska inte innehålla ämnen som klassificeras som cancerframkallande, mutagena eller reproduktionstoxiska i kategori 3 enligt bilaga I i direktiv 67/548/EEG, utan att det påverkar tillämpningen av begränsningarna i punkt 2 första meningen, om
(i) de har förbjudits i konsumentvaror enligt förordning (EG) nr 1907/2006 (Reach) eller
Motivering
Skillnaden mellan CMR-ämnen i kategori 1–2 och CMR-ämnen i kategori 3 är uppenbar.
Med hänvisning till barns hälsa och EU:s åtagande om bättre lagstiftning krävs det en enhetlig strategi för alla konsumentprodukter.
CMR-ämnen i kategori 3 som är förbjudna bör förtecknas i en ny bilaga IIb.
Ändringsförslag
20
Förslag till direktiv
Bilaga II – del III – punkt 5a (ny)
Kommissionens förslag
Ändringsförslag
5a.
Tillverkarna får, fram till dess att ett beslut antagits, fortsätta att släppa ut leksaker på marknaden som innehåller ämnen som klassificeras som CMR ‑ämnen enligt direktiv 67/548/EEG för vilka en begäran har lämnats in.
Ändringsförslag
21
Förslag till direktiv
Bilaga II – del III – punkt 7 – stycke 1 – nya led efter led 38
Kommissionens förslag
Ändringsförslag
(39) Ambrettmysk
(40) 4-fenyl-3-buten-2-on
(41) Amylkanelaldehyd
(42) Amylcinnamylalkohol
(43) Benzylalkohol
(44) Bensylsalicylat
(45) Kanelalkohol
(46) Kanelaldehyd
(47) Citral
(48) Cumarin
(49) Eugenol
(50) Geraniol
(51) Hydroxicitronellal
(52) Hydroximetylpentylcyklohexenkarboxaldehyd
(53) Isoeugenol
Motivering
Scientific reports show that there are 40 forbidden fragrances.
These are contained in the list of banned fragrances in the Proposal on the safety of toys with the exception of 2 substances.
These 2 substances (= musk ambrette and 4 phenyl-3-buten-2-one) which have been considered as allergenic by the SCCNFP in 2003 were not included in the list of the TSD and need to be added.
It is also appropriate to ban13 fragrances that are subject to labelling in the Commission's Porposal because Scientific reports indicated that these 13 fragrance chemicals are most frequently reported as contact allergens.
Ändringsförslag
22
Förslag till direktiv
Bilaga II – del III – punkt 7 – stycke 2
Kommissionens förslag
Ändringsförslag
(1) Amylkanelaldehyd
(2) Amylkanelalkohol
(3) Anisylalkohol
(3) Anisylalkohol
(4) Bensylalkohol
(5) Bensylbensoat
(5) Bensylbensoat
(6) Bensylcinnamat
(6) Bensylcinnamat
(7) Bensylsalicylat
(8) Kanelaldehyd
(9) Kanelalkohol
(10) Citral
(11) Citronellol
(11) Citronellol
(12) Kumarin
(13) Eugenol
(14) Farnesol
(14) Farnesol
(15) Geraniol
(16) Hexylkanelaldehyd
(16) Hexylkanelaldehyd
(17) Hydroxicitronellal
(18)Hydroxi-metylpentylcyklohexenkarboxaldehyd
(19) Isoeugenol
(21) d-Limonen
(21) d-Limonen
(22) Linalol
(22) Linalol
(23) Metylheptinkarbonat
(23) Metylheptinkarbonat
(24) 3-Metyl-4-(2,6,6-trimetyl-2-cyklohexen-1-yl)-3-buten-2-on
(24) 3-Metyl-4-(2,6,6-trimetyl-2-cyklohexen-1-yl)-3-buten-2-on
(25) Ekmosseextrakt
(25) Ekmosseextrakt
(26) Trämosseextrakt
(26) Trämosseextrakt
Motivering
Några viktiga ämnen saknas i kommissionen förteckning över allergiframkallande doftämnen.
Dessa måste läggas till.
Ändringsförslag
23
Förslag till direktiv
Bilaga II – del III – punkt 8 – inledningen och tabellen
Kommissionens förslag
Grundämne
mg/kg i torrt, sprött, pulverliknande eller böjligt leksaksmaterial
mg/kg
i vätskeformigt eller klibbigt leksaksmaterial
Aluminium
5625
1406
Antimon
45
11,3
Arsenik
7,5
1,9
Barium
4500
1125
Bor
1200
300
Kadmium
3,8
0,9
Krom (III)
37,5
9,4
Krom (VI)
0,04
0,01
Kobolt
10,5
2,6
Koppar
622,5
156
Bly
27
6,8
Mangan
1200
300
Kvicksilver
15
3,8
Nickel
75
18,8
Selen
37,5
9,4
Strontium
4500
1125
Tenn
15000
3750
Organiskt tenn
1,9
0,5
Zink
3750
938
Ändringsförslag
För att skydda barns hälsa får dagligen högst följande mängder av nedanstående ämnen vara biologiskt tillgängliga till följd av kontakt med en leksak:
0,2 µg Antimon
0,01 µg Arsenik
0,85 µg Barium
5,0 µg Bor
0,25 µg Kadmium
0,25 µg Krom*(härlett ur Cr III)
0,35 µg Bly
0,2 µg Kvicksilver
1,25 µg Selen
Därutöver får högst följande mängder av organiska tennföreningar vara biologiskt tillgängliga:
0,025 µg Tenn
0,075 µg Summan av de organiska tennföreningarna
Vid oral exponering via en leksak får högst 10 % av det för barn anpassade acceptabla dagliga intaget (ADI) vara biologiskt tillgängligt till följd av kontakt med en leksak.
Motivering
Ämnen som exempelvis strontium, som inte förekommer i leksakstillverkning, bör utgå ur direktivet och i stället bedömas enligt gängse toxikologiska förfaranden.
Vidare är gränsvärdena för andra ämnen på tok för höga och måste därför sänkas.
Framför allt bör ett lägre gränsvärde införas för bly.
Mätvärdet för de uppräknade ämnena bör bygga på det för barn anpassade acceptabla dagliga intaget.
Ändringsförslag
24
Förslag till direktiv
Bilaga V – del B – punkt 7 – stycke 2
Kommissionens förslag
Ändringsförslag
”Tillsyn av en vuxen rekommenderas”
”Tillsyn av en vuxen rekommenderas starkt ”
Motivering
Barns säkerhet skyddas bättre genom denna formulering.
ÄRENDETS GÅNG
Titel
Leksakers säkerhet
Referensnummer
KOM(2008)0009 – C6-0039/2008 – 2008/0018(COD)
Ansvarigt utskott
IMCO
Yttrande
Tillkännagivande i kammaren
David Hammerstein
27.5.2008
Behandling i utskott
27.5.2008
16.7.2008
7.10.2008
Antagande
7.10.2008
Slutomröstning: resultat
+:
–:
0:
29
2
1
Slutomröstning: närvarande ledamöter
Jan Březina, Jerzy Buzek, Jorgo Chatzimarkakis, Giles Chichester, Dragoş Florin David, Pilar del Castillo Vera, Den Dover, Nicole Fontaine, Norbert Glante, András Gyürk, David Hammerstein, Erna Hennicot-Schoepges, Mary Honeyball, Ján Hudacký, Romana Jordan Cizelj, Werner Langen, Pia Elda Locatelli, Eluned Morgan, Angelika Niebler, Reino Paasilinna, Atanas Paparizov, Francisca Pleguezuelos Aguilar, Miloslav Ransdorf, Herbert Reul, Teresa Riera Madurell, Paul Rübig, Britta Thomsen, Patrizia Toia, Claude Turmes, Nikolaos Vakalis, Adina-Ioana Vălean
Slutomröstning: närvarande suppleanter
Gabriele Albertini, Etelka Barsi-Pataky, Manuel António dos Santos, Juan Fraile Cantón, Neena Gill, Pierre Pribetich, Silvia-Adriana Ţicău, Vladimir Urutchev
Slutomröstning: närvarande suppleanter (art.
178.2)
Domenico Antonio Basile, José Javier Pomés Ruiz, Stefano Zappalà
ÄRENDETS GÅNG
Titel
Leksakers säkerhet
Referensnummer
KOM(2008)0009 – C6-0039/2008 – 2008/0018(COD)
Framläggande för parlamentet
25.1.2008
Ansvarigt utskott
Tillkännagivande i kammaren
IMCO
11.3.2008
Rådgivande utskott
Tillkännagivande i kammaren
ENVI
11.3.2008
ITRE
11.3.2008
Föredragande
Utnämning
Marianne Thyssen
28.2.2008
Behandling i utskott
7.4.2008
27.5.2008
23.6.2008
24.6.2008
6.10.2008
Antagande
6.11.2008
Slutomröstning: resultat
+:
–:
0:
40
Slutomröstning: närvarande ledamöter
Mia De Vits, Janelly Fourtou, Evelyne Gebhardt, Martí Grau i Segú, Małgorzata Handzlik, Malcolm Harbour, Anna Hedh, Iliana Malinova Iotova, Pierre Jonckheer, Alexander Graf Lambsdorff, Kurt Lechner, Lasse Lehtinen, Toine Manders, Catiuscia Marini, Arlene McCarthy, Nickolay Mladenov, Zita Pleštinská, Giovanni Rivera, Zuzana Roithová, Heide Rühle, Leopold Józef Rutowicz, Salvador Domingo Sanz Palacio, Christel Schaldemose, Andreas Schwab, Marianne Thyssen, Jacques Toubon, Bernadette Vergnaud, Barbara Weiler, Marian Zlotea
Slutomröstning: närvarande suppleanter
Emmanouil Angelakas, Wolfgang Bulfon, Colm Burke, Joel Hasse Ferreira, Filip Kaczmarek, Guntars Krasts, Marine Le Pen, Andrea Losco, Manuel Medina Ortega, José Javier Pomés Ruiz, Olle Schmidt, Francesco Enrico Speroni, Anja Weisgerber
Slutomröstning: närvarande suppleanter (art.
178.2)
Maddalena Calia, Francesco Ferrari, Mario Mauro, Willem Schuth, Csaba Őry
Ingivande
12.11.2008
A6-0457/2008
***I
BETÄNKANDE
om förslaget till Europaparlamentets och rådets beslut om ändring av rådets beslut 2001/470/EG om inrättande av ett europeiskt rättsligt nätverk på privaträttens område
(KOM(2008)0380 – C6‑0248/2008 – 2008/0122(COD))
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Föredragande:
Ona Juknevičienė
PE 414.369v03-00
Teckenförklaring
* Samrådsförfarandet
majoritet av de avgivna rösterna
**I Samarbetsförfarandet (första behandlingen)
majoritet av de avgivna rösterna
**II Samarbetsförfarandet (andra behandlingen)
majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten
majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
*** Samtyckesförfarandet
majoritet av parlamentets samtliga ledamöter utom i de fall som avses i artiklarna 105, 107, 161 och 300 i EG-fördraget och artikel 7 i EU-fördraget
***I Medbeslutandeförfarandet (första behandlingen)
majoritet av de avgivna rösterna
***II Medbeslutandeförfarandet (andra behandlingen)
majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten
majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
***III Medbeslutandeförfarandet (tredje behandlingen)
majoritet av de avgivna rösterna för att godkänna det gemensamma utkastet
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Parlamentets ändringar markeras med fetkursiv stil .
I samband med ändringsakter ska de delar av en återgiven befintlig rättsakt som inte ändrats av kommissionen, men som parlamentet önskar ändra, markeras med fet stil .
Eventuella strykningar ska i sådana fall markeras enligt följande: [...].
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
FÖRKLARING OM EUROPEISKA GEMENSKAPERNAS DOMSTOL..............................17
YTTRANDE från utskottet för rättsliga frågor ...........................................20
ÄRENDETS GÅNG..................................................................................................................32
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till Europaparlamentets och rådets beslut om ändring av rådets beslut 2001/470/EG om inrättande av ett europeiskt rättsligt nätverk på privaträttens område
( KOM(2008)0380 – C6‑0248/2008 – 2008/0122(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
– med beaktande av artiklarna 61 d och 66 i EG-fördraget,
– med beaktande av yttrandet från utskottet för rättsliga frågor över den föreslagna rättsliga grunden,
– med beaktande av artiklarna 51 och 35 i arbetsordningen,
– med beaktande av betänkandet från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor och yttrandet från utskottet för rättsliga frågor ( A6‑0457/2008 ).
PARLAMENTETS ÄNDRINGSFÖRSLAG
till kommissionens förslag
Förslag till Europaparlamentets och rådets beslut om ändring av rådets beslut 2001/470/EG om inrättande av ett europeiskt rättsligt nätverk på privaträttens område
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA BESLUT
med beaktande av kommissionens förslag,
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande
(Ännu ej offentliggjort i EUT). , och
i enlighet med förfarandet i artikel 251 i fördraget
Europaparlamentets ståndpunkt av den ...
2008. , och
av följande skäl:
(1) Tanken bakom det europeiska rättsliga nätverket på privaträttens område, som inrättades mellan medlemsstaterna genom rådets beslut 2001/470/EG av den 28 maj 2001
25. , var att ett område med frihet, säkerhet och rättvisa förutsätter ett förbättrat, förenklat och påskyndat rättsligt samarbete mellan medlemsstaterna och en verklig möjlighet för medborgarna att få sin sak prövad i domstol i gränsöverskridande tvister.
Beslutet trädde i kraft den 1 december 2002.
I programmet läggs särskild tonvikt vid genomförandet av de rättsakter som Europaparlamentet och rådet antagit på civilrättens område och vid ett stärkt samarbete mellan medlemmar av de juridiska yrkeskårerna i syfte att fastställa bästa metoder.
(3) I enlighet med artikel 19 i beslut 2001/470/EG lade kommissionen den 16 maj 2006 fram en rapport om nätverkets verksamhet
Rapport från kommissionen till rådet, Europaparlamentet och Europeiska ekonomiska och sociala kommittén om tillämpningen av rådets beslut 2001/470/EG om inrättande av ett europeiskt rättsligt nätverk på privaträttens område av den 16 maj 2006, KOM(2006)0203 . .
I rapporten fastställs att målen från 2001 visserligen allmänt sett har uppnåtts, men att nätverket inte på långa vägar uttömt sina möjligheter.
(4) För att uppnå Haagprogrammets mål i fråga om stärkt rättsligt samarbete och medborgarnas tillgång till domstolsprövning och för att nätverket ska kunna axla det större antal arbetsuppgifter som väntas under de kommande åren , bör nätverket ges en ▌rättslig ram som är bättre lämpad att ge nätverket större manöverutrymme.
(5) ▌ Det är mycket viktigt att villkoren förbättras för nätverkets verksamhet i medlemsstaterna genom nationella kontaktpunkter och på så sätt stärka kontaktpunkternas roll både inom nätverket och gentemot domarna ▌och juristkåren .
(6) Medlemsstaterna bör därför göra en bedömning av vilka resurser de måste ställa till kontaktpunkternas förfogande för att de ska kunna utföra sina uppgifter fullständigt.
Den interna behörighetsfördelningen i medlemsstaterna för finansieringen av de nationella nätverksmedlemmarna bör inte påverkas av detta beslut.
(7) För att detta mål ska kunna uppnås måste det i varje medlemsstat finnas en eller flera ▌kontaktpunkter som ▌kan utföra de uppgifter som de anförtrotts .
Om det finns mer än en kontaktpunkt bör medlemsstaten sörja för effektiv samordning dem emellan.
(8) Om det av ett gemenskapsrättsligt instrument eller en internationell konvention följer att en annan medlemsstats lagstiftning är tillämplig , bör kontaktpunkterna medverka när det gäller att informera rättsliga och icke-rättsliga myndigheter i medlemsstaterna om innehållet i den utländska lagstiftningen.
(9) Kontaktpunkternas bör behandla framställningar om rättsligt samarbete tillräckligt snabbt för att det ska vara förenligt med beslutets allmänna mål.
(10) Vid beräkningen av tidsfrister enligt bestämmelserna i detta beslut bör förordning (EEG, Euratom) nr 1182/71 av den 3 juni 1971 om regler för bestämning av perioder, datum och frister
EGT L 124, 8.6.1971, s.
1. gälla.
(11) Syftet med det elektroniska registret är att tillhandahålla information för bedömningen av nätverkets insats och den konkreta tillämpningen av gemenskapsinstrument.
Det bör därför inte omfatta all information som förmedlas mellan kontaktpunkterna.
(12) ▌De inom juristkåren, särskilt advokater, notarier, utmätningsmän solicitors eller barristers, som är direkt involverade i tillämpningen av gemenskapsrättsliga och internationella instrument på civilrättens område , kan bli medlemmar i nätverket genom sina nationella organisationer för att tillsammans med nätverket kunna bidra till en del av nätverkets särskilda uppgifter och verksamhet .
(13) För att ytterligare kunna utveckla nätverkets uppgifter när det gäller möjligheten till rättslig prövning, bör kontaktpunkterna i medlemsstaterna bidra till information till allmänheten med den tekniska utrustning som är lämpligast och åtminstone genom att på justitieministeriets webbplats i medlemsstaterna ha länkar till det europeiska rättsliga nätverket och de myndigheter som ansvarar för instrumentens faktiska tillämpning.
Detta beslut bör inte tolkas som en skyldighet för medlemsstaterna att göra kontaktpunkterna direkt åtkomliga för allmänheten.
(14) Vid tillämpningen av detta beslut bör hänsyn tas till ett successivt införande av det europeiska e-juridiksystemet som särskilt är tänkt att underlätta det rättsliga samarbetet och medborgarnas möjlighet till rättslig prövning.
(15) För att öka förtroendet mellan domarna i EU och förbättra synergierna mellan de berörda europeiska nätverken , bör nätverket ▌upprätthålla förbindelser med andra europeiska nätverk som har samma mål, särskilt nätverk av rättsliga organ och nätverk av domare.
(16) För att främja det internationella rättsliga samarbetet bör nätverket utveckla kontakter med andra nätverk för rättsligt samarbete i världen samt med internationella organisationer som främjar internationellt samarbete i rättsfrågor.
(17) För att möjliggöra en regelbunden uppföljning av arbetet med att uppnå beslutets mål bör kommissionen lägga fram rapporter om nätverkets verksamhet för Europaparlamentet och rådet.
(18) Rådets beslut 2001/470/EG bör ändras i enlighet med detta.
(19) Eftersom målen för detta beslut ▌inte i tillräcklig utsträckning kan uppnås av medlemsstaterna och de därför på grund av detta besluts omfattning och verkningar bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget.
I enlighet med proportionalitetsprincipen i samma artikel går detta beslut inte utöver vad som är nödvändigt för att uppnå dessa mål.
(20) ║Förenade kungariket och Irland har i enlighet med artikel 3 i protokollet om Förenade kungarikets och Irlands ställning, som är fogat till fördraget om Europeiska unionen och fördraget om upprättandet av Europeiska gemenskapen, meddelat att de önskar delta i antagandet och tillämpningen av detta beslut.║
(21) I enlighet med artiklarna 1 och 2 i protokollet om Danmarks ställning, som är fogat till fördraget om Europeiska unionen och fördraget om upprättandet av Europeiska gemenskapen, deltar Danmark inte i antagandet av detta beslut, som därför varken är bindande för eller tillämpligt i Danmark.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Beslut 2001/470/EG ska ändras på följande sätt:
1) Artikel 2 ska ändras på följande sätt:
(a) Punkt 1 ska ändras på följande sätt:
(i) I led c ska ”samarbete på privaträttens område” ersättas med ”rättsligt samarbete på privaträttens område”. ii) Följande led ska läggas till som led e:
(ii) Följande led e ska läggas till:
” e) Yrkessammanslutningar som på nationell nivå i medlemsstaterna företräder personer med rättsliga yrken som är direkt involverade i tillämpning av gemenskapsrättsliga eller internationella instrument rörande rättsligt samarbete på privaträttens område. ”
(b) I punkt 2 ska följande stycke läggas till:
▌
Om den kontaktpunkt som utses i enlighet med denna punkt inte är en domare ska den berörda medlemsstaten föreskriva om förbindelser med de nationella domstolarna .
För att underlätta detta får medlemsstaterna utse en domare för att stödja detta arbete .
Denna domare ska vara ▌medlem av nätverket.”
(c) Följande punkt 2a ska införas:
” 2a.
Medlemsstaterna ska garantera kontaktpunkten tillräckliga och lämpliga medel vad beträffar personal, resurser och modern kommunikationsutrustning för att korrekt kunna utföra uppgiften som kontaktpunkt. ”
(d) Följande punkt ska införas som punkt 4a:
” 4a.
I detta syfte ska de inhämta de berörda yrkessammanslutningarnas samtycke till att delta i nätverket. ”
När det i en medlemsstat finns flera yrkessammanslutningar som på nationell nivå företräder ett juridiskt yrke, ska medlemsstaten sörja för att yrket i fråga företräds på lämpligt sätt i nätverket. ”
” e) Punkt 5 ska ändras på följande sätt :
i) Första meningen skall ersättas med följande:
” Medlemsstaterna ska till kommissionen översända uppgifter, i enlighet med artikel 20, om namn och fullständig adress för de myndigheter som avses i punkterna 1 och 2, med uppgift om ”
ii) Led c skall ersättas med följande:
” c) när så är lämpligt, deras särskilda funktioner i nätverket samt, om det finns mer än en kontaktpunkt, kontaktpunkternas särskilda ansvarsområden. ”
2) Artikel 3 ska ändras på följande sätt:
(a) I punkt 1 ska led b ersättas med följande:
”b) förbättra allmänhetens faktiska möjlighet till rättslig prövning , ▌ genom att tillhandahålla information om hur de gemenskapsrättsliga och internationella instrument som rör rättsligt samarbete på privaträttens område fungerar.”
b) ║Punkt 2 ║ ändras på följande sätt :
i) Led b ska ersättas med följande:
” b) Att gemenskapsrättsliga instrument eller gällande konventioner mellan två eller flera medlemsstater tillämpas ändamålsenligt i praktiken, framför allt ▌ när en annan medlemsstats lagstiftning är tillämplig, att berörda domstolar eller myndigheter får vända sig till nätverket för att få information om innehållet i denna lagstiftning.”
ii) Led c ska ersättas med följande:
” c) Att inrätta, underhålla och främja ett informationssystem för allmänheten om det rättsliga samarbetet på privaträttens område inom Europeiska unionen, om relevanta gemenskapsrättsliga och internationella instrument samt om medlemsstaternas nationella lagstiftning, särskilt när det gäller möjligheten till rättslig prövning.
Den viktigaste informationskällan ska vara nätverkets webbplats, som ska innehålla uppdaterad information på samtliga officiella språk vid EU:s institutioner. ”
a) Följande led -a ska införas:
(b) Följande led ska införas som led aa:
(c) Följande led ska införas som led ca:
” c a) bidra till att på nätverkets webbplats allmänt informera allmänheten om det rättsliga samarbetet på privaträttens område i Europeiska unionen ▌ och om de relevanta gemenskapsinstrumenten och internationella instrumenten samt om den nationella rätten i medlemsstaterna , särskilt med avseende på möjligheten till rättslig prövning ,”
(d) Följande led ska läggas till som led f – g :
” f) sörja för samordningen mellan medlemmarna i nätverket på nationell nivå, ”
” g) vartannat år utarbeta en rapport om sin verksamhet , inbegripet i lämpliga fall bästa praxis i nätverket, ▌lägga fram den vid ett möte med nätverkets medlemmar och ta särskild hänsyn till möjligheterna att förbättra nätverket . ”
4) Följande artikel ska införas som artikel 5a:
” Artikel 5a
Yrkessammanslutningar
1.
2.
De kontakter som avses i punkt 1 får omfatta i synnerhet följande verksamhet:
a) Utbyte av erfarenheter och information avseende ändamålsenlig tillämpning av gemenskapsrättsliga och internationella instrument.
b) Samarbete vid utformning och uppdatering av de faktablad som avses i artikel 15.
3.
Yrkessammanslutningarna får inte begära information om enskilda ärenden hos kontaktpunkterna.
” Varje medlemsstat ska i detta syfte , i enlighet med de närmare bestämmelser som den själv ska fastställa, se till att kontaktpunkten eller kontaktpunkterna och de behöriga myndigheterna förfogar över tillräckliga medel för att kunna sammanträda regelbundet .”
7) Artikel 8 ska ersättas med följande:
”Artikel 8
▌Behandling av framställningar om rättsligt samarbete
1.
Kontaktpunkterna ska besvara alla framställningar utan dröjsmål och senast femton dagar efter det att de mottagits.
Om en kontaktpunkt inte är i stånd att besvara en framställning inom femton dagar från och med mottagandet , ska den kortfattat informera den framställande parten om detta och ange hur lång tid den anser sig behöva för att besvara framställningen, men denna tid ska normalt sett inte överstiga 30 dagar .
2.
För att så effektivt och så snabbt som möjligt kunna besvara framställningar enligt punkt 1 ska kontaktpunkterna använda den bäst lämpade tekniska utrustningen, som ska ställas till deras förfogande av medlemsstaterna.
3.
4.
Kommissionen ska minst en gång var sjätte månad förse kontaktpunkterna med statistik över de framställningar om rättsligt samarbete och de svar som avses i punkt 3.”
8) ▌Artikel 9 ska ändras på följande sätt :
a) Punkt 1 ska ersättas med följande:
” 1.
Kontaktpunkterna i nätverket ska mötas minst en gång var sjätte månad i enlighet med artikel 12.
(b) Punkt 2 ska ersättas med följande:
”2.
Vid mötena ska varje medlemsstat företrädas av en eller flera kontaktpunkter som kan åtföljas av andra medlemmar i nätverket, dock högst sex företrädare per medlemsstat .”
(c) Punkt 3 ska utgå.
9) Följande artikel ska införas som artikel 11a:
”Artikel 11a
Deltagande av observatörer i nätverkets möten
1.
2.
Anslutningsländer och kandidatländer får inbjudas att delta i dessa möten som observatörer.
Även sådana tredjeländer som är parter i internationella avtal om rättsligt samarbete på privaträttens område ▌ som Europeiska gemenskapen ingått får ▌ inbjudas att delta som observatörer vid vissa möten i nätverket .
3.
Varje stat som är observatör får vid dessa möten låta sig företrädas av en eller flera personer, som dock inte under några omständigheter får vara fler än tre per stat.”
10) Följande artikel ska införas som artikel 12a i slutet av avdelning II :
”Artikel 12a
Förbindelser med andra nätverk och internationella organisationer
1.
Nätverket ska upprätthålla förbindelser och utbyta erfarenheter och bästa praxis med de övriga europeiska nätverk som har samma mål, till exempel det europeiska rättsliga nätverket på straffrättens område ▌.
Nätverket ska även upprätthålla sådana förbindelser med det europeiska nätverket för utbildning av domare för att i lämpliga fall och utan att påverka nationell praxis främja kurser i rättsligt samarbete på privaträttens område som riktar sig till de lokala rättsliga myndigheterna i sin medlemsstat.
2.
Nätverket ska ha förbindelser med ECC-nätverket (European Consumer Centres Network) .
Kontaktpunkterna i det europeiska rättsliga nätverket på privaträttens område ska i synnerhet bistå medlemmarna i nätverket av europeiska konsumentcentrum med all sådan allmän information om hur gemenskapsinstrument och internationella instrument fungerar som förbättrar konsumenternas möjlighet till rättslig prövning .
3.
För att kunna fullgöra de uppgifter som avses i artikel 3 när det gäller internationella instrument rörande rättsligt samarbete på privaträttens område , ska nätverket upprätthålla kontakter och utbyta erfarenheter med andra nätverk för rättsligt samarbete som inrättats mellan tredjeländer samt med internationella organisationer som främjar internationellt rättsligt samarbete ▌.
4.
Kommissionen ska vara ansvarig för att i nära samarbete med rådets ordförandeskap och medlemsstaterna genomföra bestämmelserna i denna artikel.”
11) Rubriken till avdelning III skall ersättas med följande:
”AVDELNING III
TILLGÄNGLIG INFORMATION INOM NÄTVERKET OCH INFORMATION TILL ALLMÄNHETEN”
”(c) den information som avses i artikel 8 .”
13) Följande artikel ska införas som artikel 13a:
”Artikel 13a
Allmän information till allmänheten ▌
▌Nätverket ▌ska bidra till att förse allmänheten med allmän information genom den bäst lämpade tekniska utrustningen för att ge upplysningar om innehållet i och tillämpningen av de gemenskapsrättsliga eller internationella instrument som rör det rättsliga samarbetet på privaträttens område.
”b) ▌sörja för att information om de relevanta aspekterna i gemenskapsrätten och gemenskapens förfaranden, däribland gemenskapens rättspraxis, de allmänna sidorna i informationssystemet och de faktablad som avses i artikel 15, översätts till unionens officiella språk och görs tillgängliga på nätverkets webbplats.
16) Artikel 19 ska ersättas med följande:
”Artikel 19
Utvärdering
Rapporten ska vid behov åtföljas av förslag till anpassning och ska omfatta nätverkets verksamhet för att förbättra den europeiska e-juridikens utformning, utveckling och genomförande, särskilt med avseende på att underlätta för medborgarna att få möjlighet till rättslig prövning .”
17) Artikel 20 ska ersättas med följande:
”Artikel 20
Underrättelse
Artikel 2
Ikraftträdande
Detta beslut träder i kraft den […].
Det ska tillämpas från och med den […], med undantag av artiklarna 2 och 20 som ska tillämpas från och med den dag då beslutet delges de medlemsstater som det riktar sig till.
Detta beslut riktar sig till medlemsstaterna i enlighet med fördraget om upprättandet av Europeiska gemenskapen.
Utfärdat ║ den ...
På Europaparlamentets vägnar På rådets vägnar
Ordförande Ordförande
FÖRKLARING OM EUROPEISKA GEMENSKAPERNAS DOMSTOL
Europaparlamentet och rådet uppmanar kommissionen att be representanter för domstolen, att på en nivå och på ett sätt som domstolen anser vara lämpligt, närvara vid de sammanträden som hålls av det europeiska rättsliga nätverket på privaträttens område.
YTTRANDE FRÅN UTSKOTTET FÖR RÄTTSLIGA FRÅGOR ÖVER DEN RÄTTSLIGA GRUNDEN
Gérard Deprez
Ordförande
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
BRYSSEL
Artikel 61 d:
d) besluta om lämpliga åtgärder för att främja och stärka administrativt samarbete, i enlighet med vad som föreskrivs i artikel 66,
och artikel 66:
Rådet skall enligt förfarandet i artikel 67 vidta åtgärder för att säkerställa samarbete mellan de relevanta enheterna i medlemsstaternas förvaltningar inom de områden som omfattas av denna avdelning samt mellan dessa enheter och kommissionen.
Detta tillägg tycks mest vara en korrigering eftersom rådets förslag återger exakt den rättsliga grund som tas upp i det ursprungliga beslutet 2001/470/EG, som ändras genom det beslut som nu är under behandling.
Även om artikel 66 fortfarande omfattas av samrådsförfarandet, och inte medbeslutandeförfarandet, ansåg utskottet att dessa tillägg inte påverkar innehållet och därför kan godkännas.
Slutsats
Vid utskottssammanträdet den 17 november 2008 antog utskottet för rättsliga frågor därför enhälligt
Med vänlig hälsning
Giuseppe Gargani
till utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
över förslaget till Europaparlamentets och rådets beslut om ändring av rådets beslut 2001/470/EG om inrättande av ett europeiskt rättsligt nätverk på privaträttens område
( KOM(2008)0380 – C6‑0248/2008 – 2008/0122(COD) )
Föredragande:
Diana Wallis
ÄNDRINGSFÖRSLAG
Utskottet för rättsliga frågor uppmanar utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor att som ansvarigt utskott infoga följande ändringsförslag i sitt betänkande:
Ändringsförslag
1
Förslag till beslut – ändringsakt
Skäl 4
Kommissionens förslag
Ändringsförslag
(4) För att uppnå Haagprogrammets mål i fråga om stärkt rättsligt samarbete och medborgarnas tillgång till domstolsprövning och för att nätverket ska kunna axla det större antal arbetsuppgifter som väntas under de kommande åren behövs en ny rättslig ram som ger nätverket större manöverutrymme.
(4) För att uppnå Haagprogrammets mål i fråga om stärkt rättsligt samarbete och för att nätverket ska kunna axla det större antal arbetsuppgifter som väntas under de kommande åren behövs en ny rättslig ram som ger nätverket större manöverutrymme.
Ändringsförslag
2
Förslag till beslut – ändringsakt
Skäl 5
Kommissionens förslag
Ändringsförslag
(5) Först och främst är det mycket viktigt att bättre strukturera nätverkens verksamhet i medlemsstaterna kring en nationell kontaktpunkt och med utgångspunkt därifrån stärka kontaktpunktens roll inom nätverket gentemot domare , rättstillämpare och det civila samhället .
(5) Först och främst är det mycket viktigt att bättre strukturera nätverkens verksamhet i medlemsstaterna kring en eller flera nationella kontaktpunkter och med utgångspunkt därifrån stärka kontaktpunkternas roll inom nätverket gentemot domare och vissa yrkesorganisationer .
Ändringsförslag
3
Förslag till beslut – ändringsakt
Skäl 6
Kommissionens förslag
Ändringsförslag
(6) För att detta mål ska uppnås bör varje medlemsstat utse en huvudsaklig kontaktpunkt som uteslutande bör ägna sig åt nätverkets uppgifter och på så vis till fullo utöva de befogenheter som fastställs i beslut 2001/470/EG.
(6) För att detta mål ska uppnås bör varje medlemsstat utse en eller flera huvudsakliga kontaktpunkter som endast ägnar sig åt nätverkets uppgifter och därmed är fullt kapabla att utöva de befogenheter som tilldelats kontaktpunkterna enligt beslut 2001/470/EG.
Ändringsförslag
4
Förslag till beslut – ändringsakt
Skäl 6a (nytt)
Kommissionens förslag
Ändringsförslag
(6a) En särskild kontaktpunkt bör inrättas vid EG-domstolen med uppgift att ta sig an frågor av allmän karaktär, särskilt frågor som rör fastställande av referensramarna för förhandsavgöranden.
Ändringsförslag
5
Förslag till beslut – ändringsakt
Skäl 7
Kommissionens förslag
Ändringsförslag
(7) Om det av ett gemenskapsrättsligt instrument eller en internationell konvention följer att en annan medlemsstats lagstiftning är tillämplig bör kontaktpunkterna spela en viktig roll när det gäller att informera rättsliga och icke-rättsliga myndigheter i medlemsstaterna om innehållet i den utländska lagstiftningen.
(7) Om det av ett gemenskapsrättsligt instrument eller en internationell konvention följer att en annan medlemsstats lagstiftning är tillämplig bör kontaktpunkterna vara beredda att spela en viktig roll när det gäller att informera rättsliga och icke-rättsliga myndigheter i medlemsstaterna om innehållet i den lagstiftningen.
Ändringsförslag
6
Förslag till beslut – ändringsakt
Skäl 8
Kommissionens förslag
Ändringsförslag
(8) Kontaktpunkternas behandling av framställningarna om samarbete bör vara så snabb att den är förenlig med beslutets allmänna mål.
(8) Kontaktpunkternas behandling av framställningarna om samarbete bör vara så effektiv och snabb som möjligt så att den är förenlig med beslutets allmänna mål.
Ändringsförslag
7
Förslag till beslut – ändringsakt
Skäl 9
Kommissionens förslag
Ändringsförslag
(9) För att uppnå målen med beslut 2001/470/EG i fråga om bättre rättsligt samarbete i unionen och bättre tillgång till domstolsprövning för medborgarna bör de juridiska yrkeskårer som är direkt involverade i tillämpningen av gemenskapsrättsliga och internationella instrument på civilrättens område bli medlemmar i nätverket genom sina nationella organisationer .
(9) För att uppnå målen med beslut 2001/470/EG i fråga om bättre rättsligt samarbete i unionen och bättre tillgång till domstolsprövning för medborgarna kan de av medlemsstaterna utsedda yrkesorganisationer som är direkt involverade i tillämpningen av gemenskapsrättsliga och internationella instrument på civilrättens område bli medlemmar i nätverket.
Ändringsförslag
8
Förslag till beslut – ändringsakt
Skäl 10
Kommissionens förslag
Ändringsförslag
(10) För att ytterligare utveckla nätverkets uppgifter när det gäller tillgång till domstolsprövning bör kontaktpunkterna i medlemsstaterna dessutom stegvis göras tillgängliga för allmänheten genom moderna kommunikationsmedel .
(10) För att ytterligare främja tillgången till domstolsprövning bör kontaktpunkterna i medlemsstaterna uppmuntras att ta aktiv del i utvecklingen av europeisk e-juridik genom att bidra till utformningen av framtida webbplatser, inbegripet medborgarnas webbplats för e-juridik, som led i gemenskapens politik på området för e-juridik vars främsta syfte är att ge medborgarna direkt tillgång till rättsväsendet.
Som ett första steg bör de nationella justitieministeriernas webbplatser förses med länkar till det europeiska rättsliga nätverkets webbplats .
Ändringsförslag
9
Förslag till beslut – ändringsakt
Skäl 11
Kommissionens förslag
Ändringsförslag
(11) För att öka förtroendet mellan domarna i EU och förbättra synergierna mellan de berörda europeiska nätverken bör nätverket kunna upprätthålla förbindelser med andra europeiska nätverk som har samma mål, särskilt nätverk av rättsliga organ och nätverk av domare.
(11) För att öka förtroendet mellan domarna eller andra jurister i EU och förbättra synergierna mellan de berörda europeiska nätverken bör nätverket kunna upprätthålla förbindelser med andra europeiska nätverk som har samma mål, särskilt nätverk av rättsliga organ , domare och jurister .
Motivering
Det bör tydliggöras att samarbetet med andra officiella nätverk, inbegripet juristnätverk, bör utvidgas.
Ändringsförslag
10
Förslag till beslut – ändringsakt
Beslut 2001/470/EG
Kommissionens förslag
Ändringsförslag
ia) Följande led da ska läggas till:
” da) En särskild kontaktpunkt vid EG ‑domstolen med uppgift att ta sig an frågor av allmän karaktär om mål hos denna institution, särskilt frågor som rör fastställande av referensramarna för förhandsavgöranden. ”
Ändringsförslag
11
Förslag till beslut – ändringsakt
Beslut 2001/470/EG
Kommissionens förslag
Ändringsförslag
e) Yrkesorganisationer som på nationell nivå i medlemsstaterna företräder advokater, notarier, utmätningsmän och andra juridiska yrkeskårer som är direkt involverade i tillämpning av gemenskapsrättsliga eller internationella instrument rörande rättsligt samarbete på privaträttens område.
e) Yrkesorganisationer som på nationell nivå i medlemsstaterna företräder advokater, notarier enligt romersk rätt , utmätningsmän och andra juridiska yrkeskårer som är direkt involverade i tillämpning av gemenskapsrättsliga eller internationella instrument rörande rättsligt samarbete på privaträttens område och som medlemsstaterna kan utse, med deras samtycke, i syfte att ge omdömen om hur det civilrättsliga systemet fungerar på europeisk nivå, samt ge befogenhet att ställa allmänna frågor .
Ändringsförslag
12
Förslag till beslut – ändringsakt
Kommissionens förslag
Ändringsförslag
Om en medlemsstat utser flera kontaktpunkter ska den bland dem utse en huvudsaklig kontaktpunkt och se till att lämpliga samordningsmekanismer tillämpas kontaktpunkterna emellan.
Om en medlemsstat utser flera kontaktpunkter ska den bland dem utse en eller flera huvudsakliga kontaktpunkter och se till att lämpliga samordningsmekanismer tillämpas kontaktpunkterna emellan.
Ändringsförslag
13
Förslag till beslut – ändringsakt
Kommissionens förslag
Ändringsförslag
Om den kontaktpunkt som utses i enlighet med andra stycket inte är en domare ska den berörda medlemsstaten utse en domare som ska bistå kontaktpunkten i dess förbindelser med lokala rättsliga myndigheter.
Domaren ska vara fullvärdig medlem av nätverket.
Om en kontaktpunkt som utses i enlighet med andra stycket inte är en domare kan kontaktpunkten i fråga begära att en eller flera domare utses att bistå kontaktpunkten i dess förbindelser med lokala rättsliga myndigheter.
Domaren eller domarna i fråga kan utses till fullvärdiga eller tillfälliga medlemmar av nätverket.
Ändringsförslag
14
Förslag till beslut – ändringsakt
Kommissionens förslag
Ändringsförslag
ba) Följande punkt ska införas som punkt 2a:
” 2a.
Ändringsförslag
15
Förslag till beslut – ändringsakt
Beslut 2001/470/EG
Kommissionens förslag
Ändringsförslag
ca) Följande punkt 4a ska införas:
” 4a.
De ska i detta syfte utverka de berörda organisationernas samtycke till att ingå i nätverket. ”
Ändringsförslag
16
Förslag till beslut – ändringsakt
Beslut 2001/470/EG
Kommissionens förslag
Ändringsförslag
a) I punkt 1 ska led b ersättas med följande:
utgår
Ändringsförslag
17
Förslag till beslut – ändringsakt
Beslut 2001/470/EG
Kommissionens förslag
Ändringsförslag
ba) Följande led ba ska läggas till:
Ändringsförslag
18
Förslag till beslut – ändringsakt
Beslut 2001/470/EG
Kommissionens förslag
Ändringsförslag
ca) informera allmänheten om det rättsliga samarbetet på privaträttens område inom Europeiska unionen, om de relevanta gemenskapsrättsliga och internationella instrumenten och om medlemsstaternas nationella lagstiftning, särskilt när det gäller tillgång till domstolsprövning ,
ca) ge allmänheten möjlighet att få tillgång till information om det rättsliga samarbetet på privaträttens område inom Europeiska unionen, om de relevanta gemenskapsrättsliga och internationella instrumenten och om medlemsstaternas nationella lagstiftning, särskilt genom att förse de nationella justitieministeriernas webbplatser med en länk till det europeiska rättsliga nätverkets webbplats ,
Ändringsförslag
19
Förslag till beslut – ändringsakt
Beslut 2001/470/EG
Kommissionens förslag
Ändringsförslag
ba) Följande punkt 2a ska införas:
” 2a.
– främja det mellanstatliga samarbetet på privaträttens område,
– göra det lättare för jurister att på ett ändamålsenligt och konkret sätt tillämpa gemenskapsrättsliga instrument och gällande konventioner mellan två eller fler medlemsstater,
– underlätta möjligheterna till rättslig prövning, särskilt genom att medverka, när detta är nödvändigt, i utarbetandet och uppdateringen av de faktablad som avses i artikel 15.
För att fullgöra dessa uppgifter och se till att deras respektive erfarenheter får så stor spridning som möjligt ska kontaktpunkterna stå i regelbunden kontakt med de berörda yrkesorganisationerna.
Kontaktpunkterna ska därför tillhandahålla allmänna upplysningar om genomförandet av gemenskapens lagstiftning eller internationella instrument om samarbete på privaträttens område, varvid inga uppgifter ska överlämnas som rör specifika fall.
Ändringsförslag
20
Förslag till beslut – ändringsakt
Beslut 2001/470/EG
Kommissionens förslag
Ändringsförslag
f) vartannat år utarbeta en rapport om sin verksamhet och lägga fram den vid ett möte med nätverkets medlemmar.
f) vartannat år utarbeta en rapport om sin verksamhet och lägga fram den vid ett möte med nätverkets medlemmar.
Denna rapport ska innehålla förslag om bästa praxis och särskilt påpeka brister i nätverket.
Ändringsförslag
21
Förslag till beslut – ändringsakt
Kommissionens förslag
Ändringsförslag
1.
Nätverket ska ha förbindelser med andra europeiska nätverk som har samma mål, särskilt det europeiska rättsliga nätverket på straffrättens område och det europeiska nätverket för utbildning av domare.
1.
Nätverket ska ha förbindelser med andra europeiska nätverk som har samma mål, särskilt det europeiska rättsliga nätverket på straffrättens område , det europeiska notariatnätverket och det europeiska nätverket för utbildning av domare.
Motivering
Det europeiska notariatnätverket (”European Notarial Network”) är det första och hittills enda nätverk som skapats av en juridisk yrkeskår.
Man bör uttryckligen hänvisa till det i texten till beslutet såsom ett exempel på god praxis och i syfte att påskynda de juridiska yrkeskårernas integrering i det europeiska rättsliga nätverket.
Ändringsförslag
22
Förslag till beslut – ändringsakt
Beslut 2001/470/EG
Artikel 13a
Kommissionens förslag
Ändringsförslag
Genom den bäst lämpade tekniska utrustningen ska allmänheten stegvis få tillgång till kontaktpunkterna i nätverket , som ska informera om innehållet i och tillämpningen av gemenskapsrättsliga eller internationella instrument rörande rättsligt samarbete på privaträttens område samt vid behov hänvisa till de myndigheter som ansvarar för den konkreta tillämpningen av instrumenten, särskilt de myndigheter som avses i artikel 6 .
Genom den bäst lämpade tekniska utrustningen för att informera om innehållet i och tillämpningen av gemenskapsrättsliga eller internationella instrument rörande rättsligt samarbete på privaträttens område ska allmänheten stegvis få tillgång till den information som finns att hämta på det europeiska rättsliga nätverket .
Ändringsförslag
23
Förslag till beslut – ändringsakt
Beslut 2001/470/EG
Artikel 19
Kommissionens förslag
Ändringsförslag
Senast den […] [tre år efter det att detta beslut har blivit tillämpligt], och därefter vart tredje år, ska kommissionen lägga fram en rapport om nätverkets verksamhet för Europaparlamentet, rådet och Europeiska ekonomiska och sociala kommittén.
Rapporten ska vid behov åtföljas av förslag till anpassningar .
Senast den […] [tre år efter det att detta beslut har blivit tillämpligt], och därefter vart tredje år, ska kommissionen lägga fram en rapport om nätverkets verksamhet för Europaparlamentet, rådet och Europeiska ekonomiska och sociala kommittén.
Rapporten ska vid behov åtföljas av förslag till anpassning och ska särskilt uppmärksamma det arbete som bedrivs inom nätverket för att föra utformningen, utvecklingen och införandet av europeisk e-juridik vidare, i första hand i syfte att förbättra medborgarnas tillgång till domstolsprövning .
ÄRENDETS GÅNG
Titel
Inrättande av ett europeiskt rättsligt nätverk på privaträttens område
Referensnummer
KOM(2008)0380 – C6-0248/2008 – 2008/0122(COD)
Ansvarigt utskott
LIBE
Yttrande
Tillkännagivande i kammaren
JURI
10.7.2008
Föredragande av yttrande
Utnämning
Diana Wallis
9.9.2008
Antagande
4.11.2008
Slutomröstning: resultat
+:
–:
0:
25
Slutomröstning: närvarande ledamöter
Carlo Casini, Titus Corlăţean, Bert Doorn, Monica Frassoni, Giuseppe Gargani, Lidia Joanna Geringer de Oedenberg, Neena Gill, Othmar Karas, Klaus-Heiner Lehne, Katalin Lévai, Antonio López-Istúriz White, Antonio Masip Hidalgo, Hans-Peter Mayer, Manuel Medina Ortega, Aloyzas Sakalas, Francesco Enrico Speroni, Diana Wallis, Jaroslav Zvěřina, Tadeusz Zwiefka
Slutomröstning: närvarande suppleanter
Sharon Bowles, Eva Lichtenberger, Rareş-Lucian Niculescu, Georgios Papastamkos, József Szájer, Jacques Toubon, Renate Weber
ÄRENDETS GÅNG
Titel
Inrättande av ett europeiskt rättsligt nätverk på privaträttens område
Referensnummer
KOM(2008)0380 – C6-0248/2008 – 2008/0122(COD)
Framläggande för parlamentet
23.6.2008
Ansvarigt utskott
Tillkännagivande i kammaren
LIBE
10.7.2008
Rådgivande utskott
Tillkännagivande i kammaren
JURI
10.7.2008
Föredragande
Utnämning
Ona Juknevičienė
15.9.2008
Bestridande av den rättsliga grunden
JURI:s yttrande
JURI
17.11.2008
Behandling i utskott
9.9.2008
7.10.2008
5.11.2008
17.11.2008
Antagande
17.11.2008
Slutomröstning: resultat
+:
–:
0:
43
Slutomröstning: närvarande ledamöter
Alexander Alvaro, Catherine Boursier, Emine Bozkurt, Kathalijne Maria Buitenweg, Maddalena Calia, Giusto Catania, Jean-Marie Cavada, Fabio Ciani, Carlos Coelho, Elly de Groen-Kouwenhoven, Panayiotis Demetriou, Gérard Deprez, Agustín Díaz de Mera García Consuegra, Claudio Fava, Armando França, Kinga Gál, Patrick Gaubert, Jeanine Hennis-Plasschaert, Wolfgang Kreissl-Dörfler, Stavros Lambrinidis, Roselyne Lefrançois, Baroness Sarah Ludford, Maria Grazia Pagano, Martine Roure, Sebastiano Sanzarello, Vladimir Urutchev, Ioannis Varvitsiotis, Manfred Weber, Tatjana Ždanoka
Slutomröstning: närvarande suppleanter
Marco Cappato, Carlo Casini, Elisabetta Gardini, Monica Giuntini, Genowefa Grabowska, Luis Herrero-Tejedor, Sophia in ‘t Veld, Ona Juknevičienė, Sylvia-Yvonne Kaufmann, Jörg Leichtfried, Nicolae Vlad Popa, Luca Romagnoli, Stefano Zappalà
Slutomröstning: närvarande suppleanter (art.
178.2)
Inés Ayala Sender
A6-0485/2008
Fiskeriutskottet
Föredragande:
Pedro Guerreiro
PE 414.313v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING..........................................................................................................................10
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................13
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om den gemensamma fiskeripolitiken och fiskeriförvaltningens ekosystemansats
( 2008/2178(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av Förenta Nationernas havsrättskonvention av den 10 december 1982,
– med beaktande av rådets förordning (EG) nr 2371/2002 av den 20 december 2002 om bevarande och hållbart utnyttjande av fiskeresurserna inom ramen för den gemensamma fiskeripolitiken
EGT L 358, 31.12.2002, s.
59.
(GFP),
– med beaktande av kommissionens meddelande om den gemensamma fiskeripolitikens roll för att genomföra en ekosystemansats i havsförvaltningen ( KOM(2008)0187 ),
– med beaktande av resultaten vid rådets möte (jordbruk och fiske) den 29 och 30 september 2008 om ovannämnda meddelande från kommissionen,
– med beaktande av artikel 45 i arbetsordningen,
– med beaktande av betänkandet från fiskeriutskottet ( A6‑0485/2008 ), och av följande skäl:
A. I ett geografiskt område är alla levande organismer (människor, växter, djur och mikroorganismer), deras fysiska miljö (såsom jord, vatten och luft) och de naturliga cykler som håller dem vid liv, sammanlänkade med varandra.
C. En ekosystemansats för fisket är för närvarande den bästa grunden för ett helhetsomfattande system för förvaltning och beslutsfattande som beaktar samtliga berörda aktörer och element, deras krav och behov, samt framtida konsekvenser för systemet och samverkan mellan systemet och övriga faktorer.
D. Fisket i vattnen i varje medlemsstats exklusiva ekonomiska zon (EEZ) är viktigt för deras självförsörjning och oberoende, särskilt när det gäller livsmedel.
F. Den vetenskapliga forskningen om fiskeresursernas hållbarhet förutsätter att alla antaganden som grundar sig på förutfattade meningar förkastas, vilket innebär att ekosystemanalysen av fiskeresurserna är verkligt ekosystemisk endast om den grundar sig på vetenskapliga fakta.
G. En sådan ekosystemansats måste vara dynamisk och flexibel då information ges och beslut fattas, eftersom nya vetenskapliga rön och samspel ständigt kan leda till att denna ansats måste anpassas.
H. Allvarliga och oroväckande överträdelser av reglerna för den gemensamma fiskeripolitiken förekommer ofta, vilket även fastställdes i kommissionens meddelande KOM(2008)0670 , trots försök att minska gemenskapens flotta.
I. Bedömningen av fiskeresurserna är inriktad på vattnens hållbarhet, vilken är fundamental för fiskerinäringen och något som medlemsstaterna måste bevara.
J. Fiskeripolitikens huvudsyfte, som alla stater som deltog i världstoppmötet för en hållbar utveckling i Johannesburg 2002 var överens om, är maximal hållbar fångst.
K. Fiskerinäringens kraftigt minskade avkastning beror på att många fiskbestånd med kommersiellt värde fiskats ut, något som gjort det nödvändigt att belägga fiskeriaktiviteterna med restriktioner, att priserna i första ledet har stagnerat/minskat, samt att produktionsfaktorerna (diesel och bensin) har ökat lavinartat, något som slår hårdare mot länder där dessa kostnader är högre, särskilt på grund av bristen på stödåtgärder i denna näring, jämfört med dem som vidtagits i andra länder.
L. Kommissionen har lagt fram ett förslag om att börja diskutera en eventuell reform av den gemensamma fiskeripolitiken.
Europaparlamentet fäster uppmärksamheten på fiskesektorns stora ekonomiska, sociala och kulturella betydelse i vissa kustsamhällen i EU.
Europaparlamentet insisterar på behovet av att tillämpa stöd- eller ersättningsmekanismer för de fiskare som drabbas av fleråriga återhämtnings- och förvaltningsplaners ekonomiska och sociala återverkningar, liksom på behovet av skyddsåtgärder för ekosystemen.
Europaparlamentets och rådets direktiv 2008/56/EG av den 17 juni 2008 om upprättande av en ram för gemenskapens åtgärder på havsmiljöpolitikens område (Ramdirektiv om en marin strategi) (EUT L 164, 25.6.2008, s.
Europaparlamentet uppmanar kommissionen att studera och föreslå öppnare system för övervakning och kontroll av lossning av fiske, illegala fångster och kassering av oönskade fiskar.
Europaparlamentet anser att det är olämpligt att mäta alla fiskeansträngningar på ett och samma sätt, utan att hänsyn tas till olika slags fiskeflottor och fiskeredskap, och anser att hänsyn måste tas till olika fiskarter, fiskeredskap och den påverkan fångsterna av varje fiskart har på vattnen vid kontrollen av fiskeansträngningarna.
Europaparlamentet anser att de rumsliga begränsningarna (avgränsade eller skyddade områden, till exempel skyddade marina områden) kräver ett tvärvetenskapligt underlag som stöder dem, särskilt i fråga om de olika aktiviteternas och faktorernas faktiska effekt på ekosystemen och begränsningarnas faktiska fördelar, vilket omfattar djupgående specifika studier av deras miljöpåverkan och socioekonomiska effekt för fiskesamhällena.
Europaparlamentet anser därför att en av de främsta uppgifterna på fiskeriförvaltningens område är att vetenskapligt utvärdera om det finns överdimensionerade fiskeflottor och överexploaterade fiskeresurser, och vilka de i så fall är, för att kunna vidta lämpliga och specifika åtgärder.
44.
Europaparlamentet menar att införandet av industriella trålningsredskap har gett upphov till ökad fiskerelaterad dödlighet, vilket har gjort det nödvändigt att kontrollera denna fångstmetod separat, till exempel genom att behålla de gränser som gäller för fiskeområde (närhet eller avstånd till kusten).
Europaparlamentet uppmanar kommissionen att så mycket som möjligt påskynda den ekologiska certifieringen av fisket i syfte att främja ett renare fiske som i större utsträckning beaktar miljön.
53.
MOTIVERING
Kommissionens meddelande om den gemensamma fiskeripolitikens roll för att genomföra en ekosystemansats i havsförvaltningen ingår i de initiativ som kommissionen lägger fram för att inleda en debatt om en eventuell reform av den gemensamma fiskeripolitiken före 2012.
När det gäller de många varierande och komplexa frågor som kommissionen ställer anser föredraganden att det är viktigt att understryka några väsentliga aspekter.
Fiskerinäringen är en verksamhet av yttersta vikt för att förse människan med föda och garantera hennes överlevnad vilket är all fiskeripolitiks huvudsakliga syfte.
Därför måste betydelsen av fisket i medlemsstaternas exklusiva ekonomiska zoner för deras självförsörjning och oberoende understrykas, särskilt i fråga om livsmedel.
En fiskeripolitik måste sätta fångsten av fiskeresurserna i första rummet, utan att glömma föregående och efterföljande näringsled och den mycket viktiga vetenskapliga forskningen, särskilt utvärderingen och planeringen av fångsterna och fiskeresursernas biomassa.
Med andra ord är en fiskeripolitik inte, och får inte vara, en politik avsedd för haven eller den marina miljön.
Havspolitiken bör ge företräde åt haven på samma sätt som fiskeripolitiken gör det åt fiskeriet.
Förutom detta måste man alltid beakta de vetenskapliga resultaten i stället för att förlita sig på gissningar grundade på förutfattade meningar om att fisket är orsaken till systemens ohållbarhet.
Förslaget om en ekosystemanalys av utvärderingen av fiskeresurserna kan godtas om det grundar sig på vetenskapliga fakta om vattnens hållbarhet och tar hänsyn till de många olika faktorer vid sidan av fiskeriet som påverkar ekosystemet.
Det är viktigt att understryka att den gemensamma fiskeripolitiken måste främja en modernisering och en hållbar utveckling av fiskerinäringen som dels gör den socioekonomiskt möjlig och ger hållbara fiskeresurser, och dels garanterar livsmedelssäkerhet, allmänhetens självförsörjning av fisk och livsmedel, bibehållna arbetstillfällen och förbättrade livsvillkor för fiskare.
Hänsyn måste vidare tas till att den kraftigt minskade avkastningen beror på fiskeaktiviteternas inskränkningar och att priserna i första ledet har stagnerat/minskat, samt att produktionskostnaderna (diesel och bensin) har ökat lavinartat.
Fiskeripolitiken förutsätter att hänsyn tas till många olika dimensioner – sociala, ekologiska och ekonomiska – vilket kräver ett integrerat och balanserat synsätt, oförenligt med den rådande uppfattningen om en i förväg fastställd prioriteringsordning.
Detta innebär att fiskeripolitiken inte får vara underordnad någon annan gemenskapspolitik – det som snarare krävs är att den senare bevarar och integrerar fiskeripolitikens mål.
En fiskeripolitik måste utgå från antagandet om det ömsesidiga beroendet mellan fiskesamhällenas välbefinnande och hållbarheten hos de ekosystem i vilka de ingår, bland annat genom att erkänna det småskaliga kustfiskets och det icke-kommersiella fiskets särskilda egenskaper och betydelse.
Ett införande av en ekosystemansats i havsförvaltningen kräver med nödvändighet tvärvetenskapliga och sektorsövergripande åtgärder bland de olika åtgärder och politiska riktlinjer som påverkar de marina ekosystemen – åtgärder som är mer långtgående och kommer före dem som fastställts för fiskerinäringen, annars går det inte att uppnå de uppställda målen.
Det är för övrigt nödvändigt att erkänna att det finns stora skillnader mellan de olika marina områdena och de resurser som finns i dem, de olika fiskeflottorna och fiskeredskapen och deras effekt på ekosystemen, vilket kräver varierande fiskeriförvaltningsåtgärder, specifika och anpassade till varje fall, som vid behov ersätter fiskarna för uppkomna socioekonomiska följder.
Fiskeriförvaltningens första och främsta uppgift, som ju är en näring som exploaterar en självförnyande resurs, består i att (direkt eller indirekt) kontrollera de totala fiskeansträngningarna så att de begränsas till maximal hållbar fångst.
Fiskeriförvaltningens befintliga instrument, som grundar sig på totala tillåtna fångstmängder (TAC), anses hittills vara den bästa metoden för att kontrollera de totala fiskeansträngningarna, i så måtto att den direkt kontrollerar fångsten och indirekt fiskeansträngningarna.
Fördelningen av TAC per flotta och fiskeredskap, när det gäller principen om relativ stabilitet, är varje medlemsstats exklusiva behörighet.
Det är mycket viktigt att medlemsstaterna utövar sitt självbestämmande över sitt territorium, inklusive de tolv sjömilen territorialvatten – som, i förhållande till dess geografiska beskaffenhet, kan utökas – och ger sina inhemska flottor rätten till självbestämmande, med förbehåll för befintliga mellanstatliga överenskommelser.
På samma sätt är det viktigt att de exklusiva ekonomiska zoner som avser de yttre randområdena permanent betraktas som ”område för exklusiv tillgång”, för att de marina ekosystemen, fiskeaktiviteterna och de lokala fiskesamhällena ska bli hållbara.
I den meningen kan man med oro se på de förslag som gäller tillträdet till resurserna och som syftar till att införa ett system med överföringsbara individuella kvoter, vilket medför en koncentration av fiskeaktiviteterna och enskildas tillägnande av fiskerättigheter.
När det gäller fiskeansträngningarna bör det påpekas att alla inte bör mätas efter samma mått – hänsyn måste tas till de olika fiskemetoderna och fiskeredskapen och till den biologiska mångfalden.
När det gäller de rumsliga begränsningarna (avgränsade eller skyddade områden, till exempel skyddade marina områden) är det viktigt att påpeka att det krävs ett tvärvetenskapligt underlag som stöder dem.
Vidare är det viktigt att understryka att det är olämpligt och oberättigat att driva en politik som uppmuntrar en urskillningslös fartygsskrotning utan hänsyn till flottornas beskaffenhet, fiskeresurser, varje medlemsstats konsumtionsbehov och dess socioekonomiska betydelse.
Därför är det nödvändigt att vetenskapligt utvärdera om det finns överdimensionerade fiskeflottor och i så fall vilka de är och vilka fiskeresurser som är överexploaterade.
Slutligen måste det understrykas att det är mycket viktigt att låta fiskerinäringen medverka vid definitionen, införandet och utvärderingen av den gemensamma fiskeripolitikens olika åtgärder.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
2.12.2008
Slutomröstning: resultat
+:
–:
0:
17
3
Slutomröstning: närvarande ledamöter
Stavros Arnaoutakis, Elspeth Attwooll, Niels Busk, Luis Manuel Capoulas Santos, David Casa, Emanuel Jardim Fernandes, Carmen Fraga Estévez, Ioannis Gklavakis, Pedro Guerreiro, Ian Hudghton, Heinz Kindermann, Willy Meyer Pleite, Rosa Miguélez Ramos, Philippe Morillon, Seán Ó Neachtain, Struan Stevenson, Catherine Stihler, Margie Sudre
Slutomröstning: närvarande suppleanter
Raül Romeva i Rueda, Thomas Wise
A6-0488/2008
Budgetkontrollutskottet
Föredragande:
Véronique Mathieu
Rådgivande utskotts föredragande (*):
Nickolay Mladenov , utskottet för utrikesfrågor
Csaba Őry , utskottet för utveckling
(*) Förfarande med associerade utskott – artikel 47 i arbetsordningen
PE 412.305v02-00
INNEHÅLL
(*) Förfarande med associerade utskott – artikel 47 i arbetsordningen
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om budgetkontrollen av EU-medlen i Afghanistan
( 2008/2152(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av sina tidigare resolutioner om Afghanistan och, särskilt, sin resolution av den 8 juli 2008
Antagna texter, P6_TA(2008)0337 . ,
– med beaktande av konferenserna i Bonn 2001, Tokyo 2002 och Berlin 2004 under vilka Förenta nationerna, Europeiska unionen och det internationella samfundet lovade att lämna ett internationellt bistånd på totalt över 8 000 000 000 EUR till Afghanistan och med beaktande av konferensen i London 2006, under vilken Afghanistanöverenskommelsen undertecknades,
– med beaktande av den nationella utvecklingsstrategin, som den afghanska regeringen antog i början av 2008 och som också är strategin för att minska fattigdomen i landet,
– med beaktande av konferensen i Paris den 12 juni 2008 under vilken givarländerna lovade mer än 21 000 000 000 USD i bistånd till Afghanistan,
– med beaktande av de åtaganden som unionen ingått i samband med den tidigare nämnda Pariskonferensen om effektiviteten i biståndet till Afghanistan samt den uppförandekod som Europeiska unionen antog 2007,
– med beaktande av sin resolution av den 22 april 2008 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2006, avsnitt III – kommissionen
Antagna texter, P6_TA(2008)0133 . , och särskilt punkterna 181‑200 (externa åtgärder, humanitärt bistånd och utveckling),
– med beaktande av landsstrategidokumentet 2003–2006 som antagits av kommissionen i samförstånd med parlamentets där stabiliteten och minskningen av fattigdomen betonades,
– med beaktande av landsstrategidokumentet 2007–2013 samt det fleråriga vägledande programmet 2007–2010 som antogs av kommissionen i samförstånd med Europaparlamentet och som föreskriver ett belopp på 610 000 000 EUR för Islamiska republiken Afghanistan under budgetåren 2007–2010.
– med beaktande av parlamentets delegation som besökte Afghanistan mellan den 26 april och den 1 maj 2008 för att undersöka förutsättningarna för att genomföra EU-biståndet och det internationella biståndet samt rapporten från detta besök,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1. , och särskilt artikel 53 och dess genomförandebestämmelser,
– med beaktande av artiklarna 285–287 i fördraget om Europeiska unionens funktionssätt
EUT C 115, 9.5.2008, s.
47. om revisionsrätten och artiklarna 310–325 i nämnda fördrag om finansiella bestämmelser, som kommer att träda i kraft efter att ratificeringsprocessen slutförts för Lissabonfördraget om ändring av fördraget om Europeiska unionen och fördraget om upprättandet av Europeiska gemenskapen
EUT C 306, 17.12.2007, s.
1. .
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1073/1999 av den 25 maj 1999 om utredningar som utförs av Europeiska byrån för bedrägeribekämpning (OLAF)
EGT L 136, 31.5.1999, s.
1. ,
– med beaktande av millennieutvecklingsmålen och målen i millenniedeklarationen som antogs av FN den 8 september 2000 och undertecknades av 189 länder,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1905/2006 av den 18 december 2006 om upprättande av ett finansieringsinstrument för utvecklingssamarbete
EUT L 378, 27.12.2006, s.
41. ,
– med beaktande av artikel 45 i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet och yttrandena från utskottet för utrikesfrågor, utskottet för utveckling och budgetutskottet ( A6‑0488/2008 ), och av följande skäl:
A. Afghanistan är i en nästan kontinuerlig konflikt- eller krigssituation sedan flera årtionden och vid sidan av narkotikahandel och en latent korruption, som återfinns på alla förvaltningsnivåer, plågas centralregeringen sedan länge av svaga strukturer och bristfällig kapacitet och sakkunskap samt kroniskt otillräckliga medel där statens budgetinkomster täcker knappt 30 procent av de totala utgifterna.
B. Den allvarliga situation som Afghanistan står inför kräver en skyndsam förbättring av styrelseformerna så att det uppstår en starkare stat som kan garantera befolkningen säkerhet och respekt för lagarna samt kan skapa nödvändiga förutsättningar för en hållbar utveckling av landet.
C. I det nuvarande läget med global ekonomisk nedgång är det mycket viktigt att man ser till att kontrollen av EU:s finansiering av utvecklingssamarbete är effektiv.
D. I artikel 25.1 b i instrumentet för utvecklingssamarbete fastställs villkoren för budgetstöd till partnerländerna.
2.
Europaparlamentet konstaterar att unionens bistånd består av direktstöd och indirekt stöd.
Mellan 2002 och 2007 genomfördes gemenskapens direktstöd, som utgör 70 procent (970 000 000 EUR) av gemenskapens totala stöd, genom kommissionen i form av finansieringsavtal med den afghanska staten, kontrakt med leverantörer av tjänster, varor och anläggningsarbeten och avtal om bidrag med internationella organisationer och europeiska eller lokala icke-statliga organisationer medan det indirekta stödet främst förvaltades av Förenta nationerna (13 procent av medlen) och Världsbanken (17 procent av medlen).
Prioriterade sektorer för biståndet
Europaparlamentet konstaterar att för att förverkliga de två långsiktiga prioriterade mål som ställts upp för perioden 2007–2013 är följande sektorer prioriterade för biståndstilldelningen: styrelseformer, landsbygdsutveckling och hälsovård medan andra åtgärdsområden som inte prioriterats är socialt skydd, regionalt samarbete och minröjning.
Sammanfattning av utnyttjandet av Europeiska unionens medel
Europaparlamentet anser att den afghanska regeringen måste göra inrättandet av en rättsstat och kampen mot korruption och narkotikahandel till en av sina politiska prioriteringar och anser att utan adekvata styrelseformer kommer inga hållbara framsteg att göras i Afghanistan.
Europaparlamentet noterar kommissionens ansträngningar att ge ökat värde åt sina insatser i sina afghanska samarbetsparters ögon, men beklagar att medlemsstaterna nästan inte alls stöder kommissionen när den försöker ta fram projekt.
Europaparlamentet understryker att bidragsgivarnas verksamhet i Afghanistan måste samordnas bättre under ledning av FN:s biståndsuppdrag i Afghanistan, och anser att kommissionen bör stärka samordningen av bidrag bland medlemsstaterna och på så sätt göra EU:s stöd både mer verkningsfullt och mer synligt.
Rekommendationer
När det gäller det internationella biståndets samordning och synlighet
31.
32.
När det gäller biståndets prioriterade sektorer
När det gäller kontrollen av unionens medel
Europaparlamentet begär tillräcklig finansiering av säkerhetskostnaderna i projekt som leds av kommissionen, så att hjälparbetarna skyddas och medel inte avleds av den legitima säkerhetshanteringen från projektens målsättningar och resultat.
När det gäller bistånd till utveckling av den afghanska förvaltningens kapacitet
Europaparlamentet begär att utbildningar liknande dem som anordnades av OLAF och EuropeAid för afrikanska statstjänstemän under temat ”skydd och optimering av allmänna medel - samarbete mellan nationella och internationella institutioner” ska organiseras i Afghanistan.
Europaparlamentet uppmanar kommissionen och medlemsstaterna samt den afghanska regeringen att se till att deras program och verksamheter, särskilt på provinsnivå, till fullo samordnas med Afghanistans nationella utvecklingsstrategi och ligger i linje med de åtaganden som samtliga parter gjorde vid Pariskonferensen.
Europaparlamentet uppmuntrar varje initiativ som syftar till att öka kontakterna mellan Europaparlamentets interparlamentariska delegationer och Wolesi Jirga och Meshrano Jirga, de två kammarna i det afghanska parlamentet, för att främja goda parlamentariska styrelseformer.
Europaparlamentet påminner om sin rekommendation till rådet av den 25 oktober 2007 om opiumproduktion för medicinska ändamål i Afghanistan
Antagna texter, P6_TA(2007)0485 . , där rådet uppmanades att motsätta sig användningen av desinfektion som ett sätt att utrota vallmoodlingar i Afghanistan inom ramen för integrerade utvecklingsprogram och att ge sitt stöd till en diskussion om möjligheterna för och genomförbarheten av ett vetenskapligt pilotprojekt för ”Vallmo för medicin”.
o
o o
MOTIVERING
Europeiska unionens stöd och dess användning
Europeiska unionen ger direkt och indirekt stöd.
Mellan 2002 och 2007 uppgick det direkta gemenskapsstödet till 70 procent (970 miljoner euro) av det totala gemenskapsstödet medan det indirekta gemenskapsstödet, som förvaltas av internationella organisationer, uppgick till 30 procent av gemenskapsstödet (422 miljoner euro).
Stödet har avsatts till förvaltningsfonder med flera givare (trust funds) som förvaltas av FN (13 procent av fonderna) eller Världsbanken (17 procent av fonderna).
- Lofta (Fonden för lag och ordning i Afghanistan), med ett stöd på 180,5 miljoner som förvaltas av UNDP, där Europeiska unionen är den största givaren med 38 procent.
Det aktuella gemenskapsstödet regleras i ett strategidokument för perioden 2007–2013 och i ett flerårigt vägledande program i vilket de stora dragen och de prioriterade områdena för gemenskapens åtgärder fastställts för perioden 2007–2010.
Preliminär utvärdering av gemenskapsstödet
Sedan Afghanistanöverenskommelsen undertecknades i början av 2006 har stora framsteg gjorts i fråga om givarländernas utbetalning av stöd, vilket har gjort det möjligt att minska överlappande kostnader och korruption.
Den nya strategi för direkt utbetalning av medel till den afghanska regeringen som tillämpats av de internationella organisationerna, däribland Världsbanken, tycks vara en lovande metod som gör ministerierna direkt ansvariga.
Störst framsteg har bland annat gjorts inom hälso- och sjukvård, utbildning och infrastruktur (framför allt väginfrastruktur), där resultaten varit lovande efter talibanernas fall.
Följaktligen kan det konstateras att barnadödligheten minskat avsevärt (från 22 procent år 2001 till 12,9 procent år 2006), att en större procentandel afghaner har fått direkt tillgång till primärvård (65 procent år 2006 jämfört med 9 procent år 2001) och att utbildningssektorn börjar uppvisa positiva tecken på utveckling, eftersom allt fler barn, framför allt flickor, elever och lärare återvänt till skolan (andelen barn som deltar i skolundervisning har således ökat från 5 procent år 2001 till över 60 procent år 2007).
Den pågående återuppbyggnaden av grundskolan och utbildningen av lärare kan också nämnas.
Även de afghanska myndigheternas insatser för att utarbeta initiativ för jämställdhet mellan könen bör betonas.
Det finns dock en brist på samordning mellan givarländerna på internationell nivå, och även mellan de olika EU‑medlemsstaterna och Europeiska kommissionen, trots att den skulle kunna ha en enande funktion.
Därav följer att kostnadseffektiviteten är mycket lägre än vad den borde vara och det är tydligt att den afghanska befolkningen skulle ha kunnat dra mycket större direkt nytta av de internationella medel och gemenskapsmedel som tilldelats landet.
Kontrollsystemet för det direkta och indirekta gemenskapsstödet
Med tanke på den afghanska förvaltningens strukturella brister ska alla viktiga faser i fråga om urval, ingående av avtal, godkännande av avtal och betalningar för projekt som finansieras med gemenskapsmedel i allmänhet godkännas och undertecknas på förhand av kommissionens avdelningar (delegationerna och/eller huvudkontoret i förekommande fall) och alla projekt och program ska genomgå åtminstone en granskning före slutbetalning.
Enligt information från kommissionens behöriga avdelningar ska avtal ingås och betalningar överenskommas, godkännas, undertecknas och kontrolleras direkt av kommissionens avdelningar vid direkt central projektförvaltning genom leverantörer, tjänsteleverantörer och andra tjänstetillhandahållare (artikel 53a i budgetförordningen och artikel 36 i genomförandebestämmelserna).
Vid icke-styrkta eller icke-godkända utgifter ska kommissionen enligt samma källor omedelbart återkräva motsvarande belopp genom indrivning, genom att utnyttja bankgarantierna för avtalen eller genom avräkning från andra utbetalningar som ska göras till de berörda avtalsslutande parterna inom andra avtal.
Vid direkt central förvaltning av bidragsavtal med icke-statliga organisationer (NGO) gäller samma förfaranden och system (artikel 53a i budgetförordningen och artikel 36 i genomförandebestämmelserna).
Vid anlitande av internationella organisationer för gemensamt utarbetande och genomförande av gemensamma projekt som endast finansieras med gemenskapsstöd ingår kommissionens avdelningar ett direkt avtal i vilket de berörda internationella organisationernas uppgifter och skyldigheter fastställs.
Gemenskapsstöd kan utbetalas via förvaltningsfonder med flera givare.
När kommissionen betalar ut gemenskapsstöd via en förvaltningsfond med flera givare som förvaltas av en internationell organisation sköts genomförandeförfarandet för gemenskapsstödet gemensamt.
Gemenskapsmedlen läggs ihop med medlen från andra givare för att finansiera de program och projekt som den berörda förvaltningsfondens styrelse har beslutat om.
Det är därför svårt att koppla ett särskilt projekt till gemenskapsstödet, eftersom de olika givarnas medel är utbytbara och alla finansierar samma verksamhet.
Dessutom deltar kommissionen systematiskt i givarkommittéerna som kontrollerar varje förvaltningsfond, och i de olika arbetsgrupper som fastställer de sektorsvisa prioriteringar som styr projektens utformning.
Enligt bestämmelserna i ramavtalen och de upplysningar som erhållits genomför kommissionen dessutom som grund för gemenskapens utbetalningar och motsvarande utgifter finansiella stickprovskontroller av räkenskaperna och verifikationerna vid förvaltnings- och finansavdelningarna hos de internationella organisationer som sammanställer motsvarande dokument.
Inom ramen för tillämpningen av artikel 53d i budgetförordningen ska kommissionen innan den betalar ut ett finansiellt bidrag till en internationell organisation kontrollera att denna vederbörligt uppfyller internationella standarder för bokföring, revision, internkontroll och offentlig upphandling.
Kampen mot korruption och narkotikahandel
Föredraganden påminner om att Afghanistan är en av de största producenterna av vallmo och anser att det är absolut nödvändigt att aktivt bekämpa all narkotikahandel och utarbeta program som syftar till att införa alternativa grödor, vilket visat sig effektivt i den gyllene triangeln i Thailand.
6.11.2008
Föredragande (*):
Nickolay Mladenov
(*) Förfarande med associerade utskott – artikel 47 i arbetsordningen
FÖRSLAG
Utskottet för utrikesfrågor uppmanar budgetkontrollutskottet att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet erinrar om att Afghanistanöverenskommelsen, som ingicks mellan Islamiska republiken Afghanistan och världssamfundet vid Londonkonferensen 2006, är den ömsesidigt bindande ramen för återuppbyggnad och statsbyggande i Afghanistan.
Europaparlamentet uppmanar kommissionen och medlemsstaterna samt den afghanska regeringen att se till att deras program och verksamheter, särskilt på provinsnivå, till fullo samordnas med Afghanistans nationella utvecklingsstrategi och ligger i linje med de åtaganden som samtliga parter gjort vid Pariskonferensen.
Europaparlamentet erinrar om att det i 2008 års budget tog initiativ till att stödja demokratisk uppbyggnad av parlament i tredjeländer och åtar sig att använda de avsedda resurserna för att stärka det afghanska parlamentets förmåga att stifta lagar, övervaka den verkställande makten och vara fullt representativt för det afghanska folket.
EUT C 263 E, 16.10.2008, s.
651. , där rådet uppmanades att motsätta sig användningen av desinfektion som ett sätt att utrota vallmoodlingar i Afghanistan inom ramen för integrerade utvecklingsprogram och att ge sitt stöd till en diskussion om möjligheterna för och genomförbarheten av ett vetenskapligt pilotprojekt för ”Vallmo för medicin”.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
6.11.2008
Slutomröstning: resultat
+:
–:
0:
45
5
Slutomröstning: närvarande ledamöter
Vittorio Agnoletto, Roberta Alma Anastase, André Brie, Philip Claeys, Véronique De Keyser, Giorgos Dimitrakopoulos, Michael Gahler, Georgios Georgiou, Ana Maria Gomes, Jana Hybášková, Jelko Kacin, Metin Kazak, Maria Eleni Koppa, Joost Lagendijk, Vytautas Landsbergis, Johannes Lebech, Francisco José Millán Mon, Philippe Morillon, Pasqualina Napoletano, Annemie Neyts-Uyttebroeck, Baroness Nicholson of Winterbourne, Janusz Onyszkiewicz, Ria Oomen-Ruijten, Ioan Mircea Paşcu, João de Deus Pinheiro, Hubert Pirker, Samuli Pohjamo, Bernd Posselt, Libor Rouček, Christian Rovsing, Flaviu Călin Rus, Jacek Saryusz-Wolski, Inese Vaidere, Geoffrey Van Orden, Marcello Vernola, Kristian Vigenin, Andrzej Wielowieyski, Jan Marinus Wiersma, Zbigniew Zaleski, Josef Zieleniec
Slutomröstning: närvarande suppleanter
Árpád Duka-Zólyomi, Kinga Gál, Milan Horáček, Marie Anne Isler Béguin, Tunne Kelam, Miloš Koterec, Nickolay Mladenov, Inger Segelström
Slutomröstning: närvarande suppleanter (art.
178.2)
Wolfgang Bulfon, Rosa Miguélez Ramos
10.11.2008
över budgetkontrollen av EU-medlen i Afghanistan
Föredragande (*):
Csaba Őry
(*) Förfarande med associerade utskott – artikel 47 i arbetsordningen
FÖRSLAG
Utskottet för utveckling uppmanar budgetkontrollutskottet att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
- med beaktande av Europaparlamentets och rådets förordning (EG) nr 1905/2006 av den 18 december 2006 om upprättande av ett finansieringsinstrument för utvecklingssamarbete (instrument för utvecklingssamarbete – DCI)
41. ,
- med beaktande av Förenta nationernas millenniemål och målen i millenniedeklarationen, som undertecknats av 189 länder i september 2000.
A. I det nuvarande läget med global ekonomisk nedgång är det mycket viktigt att man ser till att kontrollen av EU:s finansiering av utvecklingssamarbete är effektiv.
B. I artikel 25.1 b i instrumentet för utvecklingssamarbete fastställs villkoren för budgetstöd till partnerländerna.
2.
Europaparlamentet betonar behovet av bättre övervakning av genomförandet av EU:s utvecklingssamarbete.
4.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
5.11.2008
Slutomröstning: resultat
+:
–:
0:
29
Slutomröstning: närvarande ledamöter
Josep Borrell Fontelles, Danutė Budreikaitė, Marie-Arlette Carlotti, Corina Creţu, Nirj Deva, Alexandra Dobolyi, Beniamino Donnici, Fernando Fernández Martín, Juan Fraile Cantón, Alain Hutchinson, Romana Jordan Cizelj, Filip Kaczmarek, Glenys Kinnock, Maria Martens, Gay Mitchell, Toomas Savi, Pierre Schapira, Frithjof Schmidt, Jürgen Schröder, Feleknas Uca, Johan Van Hecke, Anna Záborská, Jan Zahradil, Mauro Zani
Slutomröstning: närvarande suppleanter
Miguel Angel Martínez Martínez, Manolis Mavrommatis, Csaba Őry, Renate Weber, Gabriele Zimmer
Föredragande:
Laima Liucija Andrikienė
FÖRSLAG
Parlamentet understryker i detta sammanhang betydelsen av kommissionens program för ett effektivt bistånd och noterar Europeiska rådets slutsatser från mötet den 26 maj 2008 när det gäller EU-biståndets effektivitet i Afghanistan.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
10.11.2008
Slutomröstning: resultat
+:
–:
0:
17
Slutomröstning: närvarande ledamöter
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
2.12.2008
Slutomröstning: resultat
+:
–:
0:
13
Slutomröstning: närvarande ledamöter
Jean-Pierre Audy, Herbert Bösch, Paulo Casaca, Antonio De Blasio, Szabolcs Fazakas, Aurelio Juri, Dan Jørgensen, Rodi Kratsa-Tsagaropoulou, Bogusław Liberadzki, Jan Mulder, Bart Staes
Slutomröstning: närvarande suppleanter
Véronique Mathieu, Gabriele Stauner
A6-0085/2009
om millennieutvecklingsmålavtalen
(2008/2128(INI))
Utskottet för utveckling
Föredragande:
Alain Hutchinson
PE 418.116v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING..........................................................................................................................14
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................16
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om millennieutvecklingsmålavtalen
( 2008/2128(INI) )
Europaparlamentet utfärdar denna resolution
- med beaktande av FN:s millenniedeklaration av den 18 september 2000 genom vilken det internationella samfundet åtagit sig att uppfylla millennieutvecklingsmålen för att fram till 2015 halvera fattigdomen i världen; denna deklaration har också bekräftats under flera av FN:s konferenser, bland annat konferensen i Monterrey om utvecklingsfinansiering,
- med beaktande av de åtaganden som medlemsstaterna gjorde under Europeiska rådets möte i Barcelona den 14 mars 2002,
- med beaktande av sin resolution av den 20 juni 2007 om millennieutvecklingsmålen i halvtid
Antagna texter från detta sammanträde, P6_TA(2007)0274 . ,
- med beaktande av den gemensamma förklaringen från rådet och företrädarna för medlemsstaternas regeringar, församlade i rådet, Europaparlamentet och kommissionen om Europeiska unionens utvecklingspolitik: ”Europeiskt samförstånd”
EUT C 46, 24.2.2006, s.
1. som undertecknades den 20 december 2005,
- med beaktande av kommissionens ”millennieutvecklingsmålspaket” från 2005,
- med beaktande av kommissionens meddelande om snabbare framsteg i strävan att nå millennieutvecklingsmålen – utvecklingsfinansiering och effektivitet i biståndet ( KOM(2005)0133 ),
- med beaktande av meddelandet om att hålla Europas löften om utvecklingsfinansiering ( KOM(2007)0164 ),
- med beaktande av kommissionens meddelande om EU:s bistånd: Mer, bättre och snabbare ( KOM(2006)0087 ),
- med beaktande av sin resolution av den 23 september 2008 om uppföljningen av Monterreykonferensen 2002 om finansieringen av utvecklingsinsatser
Antagna texter från detta sammanträde, P6_TA(2008)0420 . ,
- med beaktande av resultatet av och slutdokumentet om den internationella konferensen om utvecklingsfinansiering för att se över genomförandet av Monterreykonferensen (Doha, Qatar, den 29 november–2 december 2008)
A/Conf.212/L.1/Rev1 av den 9 december 2008. ,
- med beaktande av sin resolution av den 22 maj 2008 om uppföljningen av Parisförklaringen från 2005 om biståndseffektivitet
Antagna texter från detta sammanträde, P6_TA(2008)0237 . ,
- med beaktande av kommissionens dokument av den 19 juni 2007 om millennieutvecklingsmålsavtal – en strategi för ett långsiktigare och förutsägbarare budgetstöd,
- med beaktande av det nya strategiska partnerskapet Afrika–EU,
- med beaktande av sin resolution av den 25 oktober 2007 om läget i förbindelserna mellan EU och Afrika
Antagna texter från detta sammanträde, P6_TA(2007)0483 . ,
- med beaktande av Parisförklaringen om biståndseffektivitet av den 2 mars 2005 och slutsatserna från högnivåforumet i Accra som ägde rum den 2–4 september 2008 om uppföljningen av denna förklaring,
- med beaktande av sin resolution av den 6 april 2006 om biståndets effektivitet och korruptionen i utvecklingsländerna
EUT C 293 E, 2.12.2006, s.
316. ,
- med beaktande av sin resolution av den 4 september 2008 om mödradödlighet inför FN:s högnivåmöte den 25 september 2008 om översyn av millennieutvecklingsmålen
Antagna texter från detta sammanträde, P6_TA(2008)0406 . ,
- med beaktande av ”The Aid Delivery Methods.
Guidelines of the Programming, Design & Management of General Budget Support”
Offentliggjord på engelska i januari 2007 av kommissionen, byrån för samarbete EuropeAid – generaldirektoratet för bistånd – generaldirektoratet för yttre förbindelser. ,
- med beaktande av bestämmelserna i Cotonouavtalet av den 23 juni 2000, särskilt artikel 58 i 2005 års version som räknar upp de institutioner som är berättigade till stöd,
- med beaktande av OECD:s rekommendationer beträffande god sed för budgetstöd i dokumentet om att harmonisera biståndet för att förbättra dess effektivitet
DAC Reference Document, Volume 2, 2006. ,
- med beaktande av revisionsrättens särskilda rapport nr 2/2005 om EUF:s budgetstöd till AVS-länderna: kommissionens förvaltning av området ”reformen av de offentliga finanserna”
EUT C 249, 7.10.2005, s.
1. ,
- med beaktande av revisionsrättens särskilda rapport nr 10/2008 om EG:s utvecklingsbistånd till hälso- och sjukvård i Afrika söder om Sahara, samt kommissionens svar,
- med beaktande av granskningsrapporten utarbetad av IDD and Associates, med en utvärdering av det allmänna budgetstödet
IDD and Associates, maj 2006. , maj 2006,
- med beaktande av sin resolution av den 13 februari 2006 om en ny finansieringsmekanism för millenniemålen
EUT C 290 E, 29.11.2006, s.
396. ,
- med beaktande av Europeiska gemenskapens och EU ländernas undertecknande av FN:s konvention om rättigheter för personer med funktionshinder av den 13 december 2006,
- med beaktande av artikel 45 i arbetsordningen,
- med beaktande av betänkandet från utskottet för utveckling och yttrandet från budgetutskottet ( A6–0085/2009 ), och av följande skäl:
A. Genom att ansluta sig till 2000 års millenniedeklaration åtog sig Europeiska unionen att tillsammans med hela det internationella samfundet halvera den extrema fattigdomen i världen fram till 2015, och att därvid särskilt inrikta sig på att uppnå de åtta millennieutvecklingsmålen,
B. Det uppskattas att omkring 1,4 miljarder personer fortfarande lever under fattigdomsgränsen (det vill säga 1,25 US‑dollar per dag), vilket motsvarar en fjärdedel av utvecklingsvärldens befolkning.
C. Kommissionen och EU:s medlemsstater har under 2007 gjort nya åtaganden för att i hög grad bidra till att inhämta förseningar när det gäller att uppfylla dessa mål.
D. Bristen på tillgång till hälsovård och bastjänster orsakar flera miljoner dödsfall och befäster fattigdomen, medan tillgången till dessa tjänster och till en utbildning utgör en mänsklig rättighet, regeringarna är skyldiga att garantera att den respekteras och tillämpas.
E. Möjligheten finns att millennieutvecklingsmålavtalen ska utgöra ett instrument bland andra som svar på de utmaningar som uppstår i utvecklingsländerna till följd av den globala livsmedelkrisen, särskilt inom jordbrukssektorn.
F. Trots de stora ansträngningar som utvecklingsländerna samtyckt till hittills, har de flesta av utvecklingsländerna inte de resurser som krävs för att ta itu med utmaningarna vad gäller hälsa och utbildning, och därför krävs det stöd utifrån.
G. Europaparlamentet bör bevilja Europeiska utvecklingsfonden (EUF) ansvarsfrihet.
H. Kommissionen har för avsikt att avsevärt öka användningen av budgetstödet under den tionde EUF för att göra stödet effektivare och uppnå de fastställda målen.
I. Lärare inom hälso- och sjukvården och sjukvårdsanställda i utvecklingsländerna arbetar för närvarande under beklagliga förhållanden, och det behövs närmare två miljoner lärare och mer än fyra miljoner sjukvårdsanställda för att nå millennieutvecklingsmålen.
Ett tillräckligt budgetstöd, i form av budgetstöd knutet till ett millennieutvecklingsmålavtal, skulle kunna göra det möjligt att anställa och utbilda dem.
K. EU har för avsikt att fortsätta att höja sina utgifter för budgetstöd, bland annat genom att avsevärt höja det sektorsinriktade budgetstödet för hälsa och utbildning, särskilt i de afrikanska länderna.
L. I millennieutvecklingsmålavtalen fastställs konkreta resultat som ska uppnås i fråga om millennieutvecklingsmålen rörande hälsa och grundutbildning, men millennieutvecklingsmålavtal kan också komma att ingås för andra prioriterade sektorer.
M. Enligt den officiella hållning om utvecklingsstöd som parlamentet gav uttryck för i sin resolution av den 13 februari 2006 om en ny finansieringsmekanism för millenniemålen
EUT C 290 E, 29.11.2006, s.
396, punkt 6. måste ökad kvantitet ”gå hand i hand med ökad kvalitet.
N. Ett förutsägbart och långsiktigt biståndsflöde kan på ett direkt och effektivt sätt bidra till det konkreta genomförandet av de strategier för avskaffandet av fattigdom, som fastställs i millennieutvecklingsmålen.
O. Trots de åtaganden som gjorts vid konferenserna i Monterrey (2002), Gleneagles (2005), Paris (2005) och Accra (2008) för att öka kvantiteten och höja kvaliteten hos utvecklingsbidraget, beviljar fortfarande ett fåtal av unionens medlemsstater allt det stöd som de har åtagit sig att tillhandahålla, och när det tillhandahålls visar sig en del av detta stöd vara olämpligt.
P. Det verkar som om utbetalningar av budgetstöd som tillhandahålls av kommissionen försenas i 30 procent av fallen på grund av dess orimliga administrativa bördor.
Q. Budgetstödets oförutsägbarhet framgår bland annat av det faktum att de flesta villkor för tillhandahållande av detta stöd är årliga, och denna oförutsägbarhet tvingar ibland mottagarländerna att använda stödet innan det faktiskt har tillhandahållits och utan att med bestämdhet veta om stödet kommer fram.
R. EU:s oförutsägbara utvecklingsstöd berör också mottagarländer med en viss rättssäkerhet och en stabil lagstiftning.
S. Kommissionen är den främsta multilaterala givaren av utvecklingsstöd, och en av de största givarna av budgetstöd, och den använder sig i allt större utsträckning av denna stödform som har styrt en femtedel av det stöd som kommissionen har gett under de senaste åren.
T. Om budgetstödet redan är ett av de instrument som möjliggör ett förbättrat stöd från unionen, bör det vara mer synligt och beviljas på längre sikt.
U. Det budgetstöd som kommissionen för närvarande tillhandahåller planeras vanligen för en treårsperiod i taget, eller för ett år i taget för vissa byråer.
V. Förslaget till millennieutvecklingsmålavtal påverkar inte budgeten och millennieutvecklingsmålavtalet är inte ett nytt instrument, utan ett sätt att genomföra de befintliga instrumenten.
W. För närvarande är det inte klart vilken status kommissionens dokument om millennieutvecklingsmålavtal ska ha.
X. Kommissionen anser att det har blivit dags att genomföra idén om ett avtal som knyts till märkbara resultat i fråga om millennieutvecklingsmålen, i stället för att varje år kontrollera att varje enskild givares villkor uppfylls.
Y. Avtalets löptid innebär ett finansiellt åtagande som ger givarlandet större förutsägbarhet i utbyte mot ett djupare engagemang från mottagarlandets sida i fråga om de konkreta resultat som måste uppnås.
Z. Kommissionen planerar att ingå de första millennieutvecklingsmålavtalen för en sexårsperiod, det vill säga fram till slutet av den tionde EUF.
Ett av kriterierna för att kunna ingå ett millennieutvecklingsmålavtal är att landet respekterar Cotonouavtalets artikel 9 om de mänskliga rättigheterna, de demokratiska principerna och rättsstaten.
Som millennieutvecklingsmålavtalen är utformade idag avser de endast AVS-länderna.
Den grundläggande principen för utvecklingsstöd är att det ska tillhandahålla stöd för dem som behöver det mest och till de platser där det kan användas på det mest effektiva sättet.
När det gäller budgetstöd har avtal redan ingåtts mellan kommissionen och Burkina Faso (2005–2008), Etiopien (2003–2006), Ghana (2007–2009), Kenya (2004–2006), Madagaskar (2005–2007), Malawi (2006–2008), Mali (2003–2007), Moçambique (2006–2008), Tanzania (2006–2008), Uganda (2005–2007) samt Zambia (2007–2008).
Enligt de ”allmänna skyldigheterna”, och särskilt artikel 32 i FN:s konvention om rättigheter för personer med funktionshinder, är de parter som har undertecknat skyldiga att beakta funktionshinder i sitt utvecklingssamarbete.
Millenniemål – Utvecklingssamarbete
Europaparlamentet bekräftar att för att uppnå millennieutvecklingsmålen måste givarländerna respektera alla sina åtaganden och förbättra kvaliteten på det stöd de tillhandahåller.
Europaparlamentet påminner om målet i Abujaförklaringen, där det fastställs att 15 procent av statsbudgeten ska anslås till hälso- och sjukvård, och målet i den världsomfattande kampanjen för utbildning, där det fastställs att 20 procent av statsbudgeten ska anslås till utbildningssektorn.
Prioriterade sektorer
Effektivt stöd – Stabilitet och förutsägbarhet
Millennieutvecklingsmålavtal
Europaparlamentet konstaterar att det huvudsakliga syftet med millennieutvecklingsmålavtalen är att bidra till ett effektivt stöd och skynda på framstegen vad gäller att uppfylla millennieutvecklingsmålen i de länder som behöver det mest.
Europaparlamentet ber kommissionen och mottagarländerna att se till att deras parlament och civila samhällen, inbegripet handikappsorganisationer, engageras i samtliga steg i dialogen om budgetstöd, inbegripet utarbetandet, genomförandet och utvärderingen av planeringen som fastställs i millennieutvecklingsmålavtalen.
För att förbättra insynen anser Europaparlamentet att villkoren för utbetalning av den del som kan variera bör grundas på uppnådda resultat, om detta uppmuntrar givarländerna och mottagarländerna att analysera den verkliga effekten som de använda medlen har medfört, och om det förbättrar insynen vad gäller användningen av allmänna medel.
Urvalskriterier – Kreativitet och flexibilitet
26.
Utvärdering – Resultatindikatorer
0 0
MOTIVERING
2005 konstaterade kommissionen officiellt att EU:s samarbete med sina partner i utvecklingsländerna var ineffektivt.
Tillgång till hälsovård och grundutbildning utgör till exempel en dröm för miljontals människor i världen och i synnerhet för kvinnorna.
Varje dag är det 72 miljoner barn, i huvudsak flickor, som inte går till skolan.
Varje minut dör en kvinna till följd av komplikationer i samband med graviditet eller förlossning, och ett barn dör var tredje sekund på grund av en sjukdom som en läkare hade kunnat förebygga.
Samtidigt utgör tillgång till hälsovård och grundutbildning en mänsklig rättighet som regeringarna är skyldiga att respektera.
Under de tio senaste åren har ett många av utvecklingsländernas regeringar gjort enorma ansträngningar i detta hänseende, men de har helt enkelt inte tillräckliga resurser för att klara det själva.
Under tiden är Afrika söder om Sahara den region i världen där situationen utan tvekan är allra värst, och med tanke på hur utvecklingen ser ut riskerar den katastrofala situationen i regionen att vara under många år framöver.
Nästan hälften av alla afrikaner lever på mindre än 0,78 euro (1 dollar) per dag, 75 procent av alla aidsoffer är afrikaner och cirka 42 procent av den afrikanska befolkningen har inte alltid tillgång till dricksvatten.
Utöver länderna i Afrika söder om Sahara är samtliga utvecklingsländer som samarbetar med Europeiska unionen i desperat behov av statligt samarbete för en effektivare utveckling.
Budgetstöd är ett av de samarbetsinstrument som under vissa omständigheter gör det möjligt att tillhandahålla ett mer förutsägbart och långsiktigare stöd genom mottagarländernas statliga finanser, för att bland annat finansiera deras behov i fråga om hälsovård, utbildning och andra prioriterade områden.
Kommissionen är en av de viktigaste givarna när det gäller denna typ av stöd.
Föredraganden påminner om att Europaparlamentet sedan länge har begärt att man (via gemenskapsbudgeten) ska lägga större vikt vid EU:s utvecklingssamarbete när det gäller hälsovård och grundutbildning.
Enligt parlamentets beräkningar i samband med ansvarsfrihetsförfarandet för budgeten 2007 användes var det mindre än 7 procent av gemenskapens budgetmedel för utvecklingssamarbete som användes inom dessa områden.
Europaparlamentet välkomnar kommissionens förklaring i samband med förhandlingarna om finansieringsinstrumentet för utvecklingssamarbete, om att kommissionen åtar sig att ”avsätta ett riktmärke på 20 procent av det beviljade stödet till de nationella program som omfattas av instrumentet för utvecklingssamarbete senast 2009 till grundskole- och gymnasieutbildning och grundläggande hälsovård genom projekt-, program- och budgetstöd med anknytning till dessa sektorer”.
Parlamentet anser att tillämpningsområdet för millennieutvecklingsmålavtalen skulle kunna utökas till de länder som omfattas av finansieringsinstrumentet för utvecklingssamarbete, och att detta vore ett utmärkt sätt för kommissionen att nå det uppsatta målet.
För utvecklingsländerna vore detta ett intressant och önskvärt initiativ, men för kommissionen kvarstår en serie frågor att klargöra.
Det rör till exempel de kriterier som tillämpas för att fastställa vilka utvecklingsländer som kan ingå denna typ av avtal.
Detta rör fortfarande frågan om hur lång tid initiativet är tänkt att vara och hur det är tänkt att genomföras rent generellt.
Även om kommissionens budgetstöd är positivt på många sätt, bland genom att det är knutet till uppvisade resultat i fråga om hälsovård och utbildning och genom att det generellt ska planeras för tre år i taget, är det således långt ifrån perfekt.
För det första kan budgetstödet påverka utvecklingen i mottagarländerna negativt.
För det andra, även om kommissionen väljer att tillhandahålla ett långsiktigt budgetstöd finns det ingen garanti för att stödet blir mer förutsägbart på kort sikt, eftersom de administrativa förfarandena ofta är så omfattande att de leder till stora förseningar i utbetalningarna.
För det tredje är insynen mycket bristfällig när det gäller kommissionens budgetstöd, och de berörda länderna och deras befolkningar har mycket svårt att anpassa sig efter villkoren.
Finansieringsavtalen offentliggörs sällan och kommissionen låter inte alltid de civila samhällsorganisationerna och parlamenten delta i dialogen med utvecklingsländernas regeringar.
Idag råder det emellertid bred enighet om att man uppnår bättre effektivitet genom att göra utvecklingen till en fråga för inte bara utvecklingsländernas regeringar, utan även för deras medborgare.
En förutsättning för att förslaget om millennieutvecklingsmålavtal ska kunna utgöra en lämplig lösning för att effektivisera gemenskapssamarbetet är att man klart och tydligt fastställer en definition och villkor för att få ingå avtal samt villkor för genomförandet och utvärderingen av avtalet.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
17.2.2009
Slutomröstning: resultat
+:
–:
0:
23
Slutomröstning: närvarande ledamöter
Alessandro Battilocchio, Thijs Berman, Thierry Cornillet, Alexandra Dobolyi, Fernando Fernández Martín, Alain Hutchinson, Romana Jordan Cizelj, Filip Kaczmarek, Glenys Kinnock, Maria Martens, Gay Mitchell, Luisa Morgantini, José Javier Pomés Ruiz, José Ribeiro e Castro, Toomas Savi, Frithjof Schmidt, Jürgen Schröder, Feleknas Uca
Slutomröstning: närvarande suppleanter
Miguel Angel Martínez Martínez, Manolis Mavrommatis, Renate Weber, Gabriele Zimmer
Slutomröstning: närvarande suppleanter (art.
178.2)
Emilio Menéndez del Valle
A6-0248/2009
*
BETÄNKANDE
om förslaget till rådets direktiv om djurhälsovillkor vid förflyttning och import av hästdjur från tredjeland (kodifierad version)
(KOM(2008)0715 – C6‑0479/2008 – 2008/0219(CNS))
Utskottet för rättsliga frågor
Föredragande:
Lidia Joanna Geringer de Oedenberg
(Kodifiering – artikel 80 i arbetsordningen)
PE 423.758v01-00
Teckenförklaring
* Samrådsförfarandet
majoritet av de avgivna rösterna
**I Samarbetsförfarandet (första behandlingen)
majoritet av de avgivna rösterna
**II Samarbetsförfarandet (andra behandlingen)
*** Samtyckesförfarandet
majoritet av parlamentets samtliga ledamöter utom i de fall som avses i artiklarna 105, 107, 161 och 300 i EG-fördraget och artikel 7 i EU-fördraget
***I Medbeslutandeförfarandet (första behandlingen)
majoritet av de avgivna rösterna
***II Medbeslutandeförfarandet (andra behandlingen)
majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten
majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
***III Medbeslutandeförfarandet (tredje behandlingen)
majoritet av de avgivna rösterna för att godkänna det gemensamma utkastet
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
BILAGA: YTTRANDE FRÅN DEN RÅDGIVANDE GRUPPEN, SAMMANSATT AV DE JURIDISKA AVDELNINGARNA VID EUROPAPARLAMENTET, RÅDET OCH KOMMISSIONEN 6
ÄRENDETS GÅNG....................................................................................................................8
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till rådets direktiv om djurhälsovillkor vid förflyttning och import av hästdjur från tredjeland (kodifierad version)
( KOM(2008)0715 – C6‑0479/2008 – 2008/0219(CNS) )
(Samrådsförfarandet – kodifiering)
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till rådet ( KOM(2008)0715 ),
– med beaktande av artikel 37 i EG-fördraget, i enlighet med vilken rådet har hört parlamentet ( C6‑0479/2008 ),
– med beaktande av det interinstitutionella avtalet av den 20 december 1994 om en påskyndad arbetsmetod för officiell kodifiering av texter till rättsakter
EGT C 102, 4.4.1996, s.
2. ,
– med beaktande av artiklarna 80 och 51 i arbetsordningen,
– med beaktande av betänkandet från utskottet för rättsliga frågor ( A6‑0248/2009 ).
Europaparlamentet godkänner kommissionens förslag såsom det anpassats till rekommendationerna från den rådgivande gruppen, sammansatt av de juridiska avdelningarna vid Europaparlamentet, rådet och kommissionen.
BILAGA: YTTRANDE FRÅN DEN RÅDGIVANDE GRUPPEN, SAMMANSATT AV DE JURIDISKA AVDELNINGARNA VID EUROPAPARLAMENTET, RÅDET OCH KOMMISSIONEN
DE JURIDISKA AVDELNINGARNAS
RÅDGIVANDE GRUPP
Bryssel den 23 februari 2009
YTTRANDE
TILL EUROPAPARLAMENTET
RÅDET
KOMMISSIONEN
I enlighet med det interinstitutionella avtalet av den 20 december 1994 om en påskyndad arbetsmetod för officiell kodifiering av texter till rättsakter, särskilt punkt 4, sammanträdde den rådgivande gruppen, sammansatt av de juridiska avdelningarna vid Europaparlamentet, rådet och kommissionen, den 3 december 2008 för att bland annat granska ovannämnda förslag från kommissionen.
Vid sammanträdet
Den rådgivande gruppen hade 22 språkversioner av förslaget till sitt förfogande och arbetade utifrån den engelska versionen, som utgör den ursprungliga språkversionen för texten under diskussion. behandlade gruppen förslaget till rådets direktiv som syftar till att kodifiera rådets direktiv 90/426/EEG av den 26 juni 1990 om djurhälsovillkor vid förflyttning och import av hästdjur från tredjeland, och konstaterade enhälligt följande:
1) I skäl 3 bör ordalydelsen ” förflyttning av hästdjur mellan medlemsstaterna ” ändras till ” förflyttning av hästdjur inom och mellan medlemsstaterna ”.
Gruppen anser att denna skillnad synbarligen behöver rättas till.
6) I artikel 15 a bör orden ” och typen av import ” strykas.
8) I artikel 19 a bör orden ” eller typer av import ” strykas.
C. Pennera J.-C. Piris C.-F. Durand
Juridisk rådgivare Juridisk rådgivare Generaldirektör
ÄRENDETS GÅNG
Titel
Djurhälsovillkor vid förflyttning och import av hästdjur från tredjeland (kodifierad version)
Referensnummer
KOM(2008)0715 – C6-0479/2008 – 2008/0219(CNS)
Begäran om samråd med parlamentet
8.12.2008
Ansvarigt utskott
Tillkännagivande i kammaren
JURI
15.12.2008
Föredragande
Utnämning
Lidia Joanna Geringer de Oedenberg
3.11.2008
Antagande
31.3.2009
A7-0072/2009
*
BETÄNKANDE
om Konungariket Belgiens, Republiken Tjeckiens, Förbundsrepubliken Tysklands, Konungariket Spaniens, Republiken Frankrikes, Republiken Ungerns, Konungariket Nederländernas, Republiken Slovakiens, Republiken Finlands, Konungariket Sveriges och Förenade konungariket Storbritannien och Nordirlands initiativ inför antagandet av rådets beslut om inrättande av ett europeiskt nätverk för förebyggande av brottslighet (EUCPN) och om upphävande av beslut 2001/427/RIF
(11421/2009 – C7‑0109/2009 – 2009/0812(CNS))
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
Föredragande: Sonia Alfano
PE 430.474v03-00
Teckenförklaring
* Samrådsförfarandet
majoritet av de avgivna rösterna
**I Samarbetsförfarandet (första behandlingen)
majoritet av de avgivna rösterna
**II Samarbetsförfarandet (andra behandlingen)
*** Samtyckesförfarandet
majoritet av parlamentets samtliga ledamöter utom i de fall som avses i artiklarna 105, 107, 161 och 300 i EG-fördraget och artikel 7 i EU-fördraget
***I Medbeslutandeförfarandet (första behandlingen)
majoritet av de avgivna rösterna
***II Medbeslutandeförfarandet (andra behandlingen)
majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten
majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
***III Medbeslutandeförfarandet (tredje behandlingen)
majoritet av de avgivna rösterna för att godkänna det gemensamma utkastet
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Parlamentets ändringar markeras med fetkursiv stil .
I samband med ändringsakter ska de delar av en återgiven befintlig rättsakt som inte ändrats av kommissionen, men som parlamentet önskar ändra, markeras med fet stil .
Eventuella strykningar ska i sådana fall markeras enligt följande: [...].
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING............................................................................................................................7
ÄRENDETS GÅNG..................................................................................................................10
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om Konungariket Belgiens, Republiken Tjeckiens, Förbundsrepubliken Tysklands, Konungariket Spaniens, Republiken Frankrikes, Republiken Ungerns, Konungariket Nederländernas, Republiken Slovakiens, Republiken Finlands, Konungariket Sveriges och Förenade konungariket Storbritannien och Nordirlands initiativ inför antagandet av rådets beslut om inrättande av ett europeiskt nätverk för förebyggande av brottslighet (EUCPN) och om upphävande av beslut 2001/427/RIF
(11421/2009 – C7‑0109/2009 – 2009/0812(CNS) )
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
– med beaktande av Konungariket Belgiens, Republiken Tjeckiens, Förbundsrepubliken Tysklands, Konungariket Spaniens, Republiken Frankrikes, Republiken Ungerns, Konungariket Nederländernas, Republiken Slovakiens, Republiken Finlands, Konungariket Sveriges och Förenade konungariket Storbritannien och Nordirlands initiativ (11421/2009),
1.
2.
Europaparlamentet uppmanar rådet att inte anta initiativet formellt före Lissabonfördragets ikraftträdande, så att slutakten hinner slutföras och EG-domstolen, kommissionen och parlamentet garanteras en fullständig roll och kan utöva full kontroll (protokoll till Lissabonfördraget om övergångsbestämmelser).
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen och Konungariket Belgiens, Republiken Tjeckiens, Förbundsrepubliken Tysklands, Konungariket Spaniens, Republiken Frankrikes, Republiken Ungerns, Konungariket Nederländernas, Republiken Slovakiens, Republiken Finlands, Konungariket Sveriges och Förenade konungariket Storbritannien och Nordirlands regeringar parlamentets ståndpunkt.
MOTIVERING
Det europeiska nätverket för förebyggande av brottslighet
Det europeiska nätverket för förebyggande av brottslighet (EUCPN, nedan: nätverket) inrättades 2001 på grundval av rådets beslut (2001/427/RIF)
2001/427/RIF: Rådets beslut av den 28 maj 2001 om inrättande av ett europeiskt nätverk för förebyggande av brottslighet.
http://eur-lex.europa.eu/LexUriServ/LexUriServ.do?uri=CELEX:32001D0427:SV:HTML .
I beslutet bekräftas det att nätverket ska
– samla in och analysera information om detta område i syfte att utbyta bästa praxis,
– anordna konferenser, seminarier, sammanträden, initiativ och verksamhet som främjar utbyte av erfarenheter och bästa praxis,
– ställa sin sakkunskap om brottsförebyggande till rådets och kommissionens förfogande.
I detta syfte anges det i beslutet att nätverket ska ha en struktur, grundad på kontaktpunkter som utses av kommissionen (en kontaktpunkt) och de enskilda medlemsstaterna (högst tre nationella kontaktpunkter per medlemsstat).
Kontaktpunkterna ska omfatta åtminstone en företrädare för de nationella myndigheter som är behöriga för förebyggande av brottslighet i alla dess aspekter, medan de övriga kontaktpunkterna får utses av specialiserade forskare och universitetslärare eller andra aktörer inom området för brottsförebyggande verksamhet.
Medlemsstaterna ska dock se till att man involverar forskare, universitetslärare och andra aktörer på det brottsförebyggande området, t.ex. icke-statliga organisationer, lokala myndigheter och den privata sektorn.
Europol och Europeiska centrumet för kontroll av narkotika och narkotikamissbruk bör medverka i arbetet, liksom övriga behöriga organ.
2005 genomfördes en intern översyn av nätverkets struktur, som ledde till att det inrättades två ständiga utskott, en för arbetsprogrammet och en för forskning, medan kommissionen överlät förvaltningen av webbplatsen åt Storbritannien, som därefter haft som uppgift att se till att den hålls uppdaterad
Nätverkets webbplats: http://www.eucpn.org/ .
I mars 2009 offentliggjordes en extern utvärdering av hur nätverket fungerar, där man å ena sidan betonade betydelsen av de mål och uppgifter som nätet fått och genomfört, och å andra sidan avslöjade att organisationen hade misslyckats och därför inte klarat av att utveckla nätverkets potential och inverkan fullt ut.
Till de problem som den externa utvärderingen avslöjade hör bristen på lämpliga resurser, ett ineffektivt sekretariat, avsaknaden av engagemang bland de nationella företrädarna, ett bristfälligt arbetsprogram samt utläggning av kriminologisk forskning på entreprenad (till universitetet i Wien, där man har en forskare som arbetar på halvtid, två av fem arbetsdagar).
Utvärderingen omfattade även möjligheten att lägga ned nätverket.
Därför tillsatte nätverket en arbetsgrupp för att undersöka rekommendationerna från den externa utvärderingen i mars 2009 och fastställde att ändringar var nödvändiga när det gäller inrättandet av nätverket.
Även om vissa medlemsstater också övervägde möjligheten att lägga ned nätverket med tanke på det allmänna missnöjet över att målen inte uppnåtts, lade en grupp medlemsstater fram ett förslag om översyn av nätverket, och EU:s ordförandeland Sverige tog med förslaget bland de prioriteringar som ska antas under det halvår som Sverige innehar ordförandeskapet, och i vilket fall som helst innan Lissabonfördraget träder i kraft.
Förslaget till rådets beslut om inrättande av ett europeiskt nätverk
för förebyggande av brottslighet (EUCPN) och om upphävande av beslut 2001/427/RIF
Det berörda förslaget omfattar upphävande av beslut 2001/427/RIF.
Bland de få ändringar som föreslås i dokumentet finns en begränsad omstrukturering av nätverket genom inrättandet av ett externt sekretariat samt ett försök att förtydliga uppgifterna, rollerna och ansvarsområdena för nätverket samt de organ som är verksamma inom det.
Den nya och komplicerade struktur som föreslås innebär att nätverket ska bestå av ett sekretariat, kontaktpunkter som ska utses av varje medlemsstat och en styrelse.
Styrelsen ska bestå av nationella företrädare som medlemsstaterna utser och ha en ordförande (som utses bland de nationella företrädarna).
Ordföranden ska leda en verkställande kommitté (bestående av högst sex ytterligare styrelsemedlemmar och en företrädare för kommissionen).
Man bör notera att det nya förslaget leder till sammanblandning av kontaktpunkter och nationella företrädare.
Dessutom avskaffas delvis hänvisningarna till att sakkunniga, vetenskapsmän, icke-statliga organisationer och det civila samhället ska göras delaktiga både på EU-nivå och nationell nivå.
Vissa av de strukturella förbindelserna mellan nätverket och de övriga gemenskapsinstitutioner och -organ som arbetar med brott och brottsförebyggande avskaffas också.
Beslutet omfattar i synnerhet inte någon form av samarbete med Europaparlamentet, och dessutom bortser man från det tidigare kravet på språkkunskaper.
I de diskussioner som kommissionen och medlemsstaterna, församlade i rådet, har fört om förslaget rörde den mest omdiskuterade och kontroversiella frågan sekretariatet, dess finansiering, möjligheten att lägga ut det på entreprenad, sekretariatets oberoende och styrande roll gentemot kommissionen och rådet samt personalrelaterade problem.
Föredragandens ståndpunkt
Föredraganden är extremt besviken över att nätverket inte kunnat fungera i enlighet med beslutet om dess inrättande eller leva upp till förväntningarna, och inte heller kunnat bidra till uppnåendet av det synnerligen viktiga målet att förebygga brottslighet i Europeiska unionen.
Bristen på samarbete mellan kommissionen, rådet och medlemsstaterna har bidragit till att skapa en situation där nätverket faktiskt saboteras, liksom EU:s mer generella mål att bekämpa brottslighet, medräknat organiserad brottslighet, genom förebyggande verksamhet.
Bristande involvering av det civila samhället, universitetsvärlden och icke-statliga organisationer, avsaknaden av översättningar och information på nätverkets webbplats samt bristfälligt utarbetande av material om brottsförebyggande (t.ex. dokument för skolor, lärare och elever) har bland annat medverkat till att nätverket överskuggas av andra institutioner och relevanta aktörer inom denna sektor.
Föredraganden fördömer vissa medlemsstaters motvillighet i detta sammanhang, och befarar att en sådan attityd i själva verket döljer en oro som man inte vill medge för att man då måste ta itu med det problem som det innebär att brottsliga organisationer vinner mark på ett allt mer oroväckande sätt i fler och fler medlemsstater.
Ur interinstitutionell synpunkt vill man alltså att Europaparlamentet ska avstå från de institutionella befogenheter som det nya fördraget medger parlamentet inom området för brottsförebyggande, nämligen medbeslutande.
Föredraganden skulle endast ha kunnat acceptera detta tillvägagångssätt om kommissionen och rådet högtidligen hade försäkrat att de ska lägga fram ett ambitiöst förslag genast efter Lissabonfördragets ikraftträdande med utgångspunkt i diskussionerna om inrättande av ett observationsorgan om brottslighet, särskilt organiserad brottslighet, vilket skulle ha fullständiga befogenheter och en exakt avgränsad behörighet när det gäller att samla in, jämföra och utvärdera data och information samt avge rekommendationer.
ÄRENDETS GÅNG
Titel
Inrättande av ett europeiskt nätverk för förebyggande av brottslighet
Referensnummer
11421/2009 – C7-0109/2009 – 2009/0812(CNS)
Begäran om samråd med parlamentet
28.7.2009
Ansvarigt utskott
Tillkännagivande i kammaren
LIBE
14.9.2009
Föredragande
Utnämning
Sonia Alfano
29.9.2009
Behandling i utskott
5.11.2009
12.11.2009
Antagande
12.11.2009
Slutomröstning: resultat
+:
–:
0:
41
2
Slutomröstning: närvarande ledamöter
Jan Philipp Albrecht, Sonia Alfano, Vilija Blinkevičiūtė, Louis Bontes, Emine Bozkurt, Simon Busuttil, Carlos Coelho, Cornelis de Jong, Agustín Díaz de Mera García Consuegra, Cornelia Ernst, Kinga Gál, Kinga Göncz, Sylvie Guillaume, Jeanine Hennis-Plasschaert, Salvatore Iacolino, Lívia Járóka, Teresa Jiménez-Becerril Barrio, Timothy Kirkhope, Juan Fernando López Aguilar, Monica Luisa Macovei, Claude Moraes, Antigoni Papadopoulou, Georgios Papanikolaou, Jacek Protasiewicz, Carmen Romero López, Judith Sargentini, Csaba Sógor, Renate Sommer, Rui Tavares, Axel Voss, Manfred Weber, Tatjana Ždanoka
Slutomröstning: närvarande suppleanter
Alexander Alvaro, Andrew Henry William Brons, Ioan Enciu, Ana Gomes, Nadja Hirsch, Monika Hohlmeier, Ramón Jáuregui Atondo, Franziska Keller, Petru Constantin Luhan, Cecilia Wikström
Slutomröstning: närvarande suppleanter (art.
187.2)
Algirdas Saudargas
A7-0076/2009
***II
ANDRABEHANDLINGS-REKOMMENDATION
om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets förordning om märkning av däck vad gäller drivmedelseffektivitet och andra väsentliga parametrar
(14639/6/2009 – C7‑0287/2009 – 2008/0221(COD))
Utskottet för industrifrågor, forskning och energi
Föredragande:
Ivo Belet
PE 430.733v01-00
Teckenförklaring
* Samrådsförfarandet
majoritet av de avgivna rösterna
**I Samarbetsförfarandet (första behandlingen)
majoritet av de avgivna rösterna
**II Samarbetsförfarandet (andra behandlingen)
*** Samtyckesförfarandet
majoritet av parlamentets samtliga ledamöter utom i de fall som avses i artiklarna 105, 107, 161 och 300 i EG-fördraget och artikel 7 i EU-fördraget
***I Medbeslutandeförfarandet (första behandlingen)
majoritet av de avgivna rösterna
***II Medbeslutandeförfarandet (andra behandlingen)
majoritet av de avgivna rösterna för att godkänna den gemensamma ståndpunkten
majoritet av parlamentets samtliga ledamöter för att avvisa eller ändra den gemensamma ståndpunkten
***III Medbeslutandeförfarandet (tredje behandlingen)
majoritet av de avgivna rösterna för att godkänna det gemensamma utkastet
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Parlamentets ändringar markeras med fetkursiv stil .
I samband med ändringsakter ska de delar av en återgiven befintlig rättsakt som inte ändrats av kommissionen, men som parlamentet önskar ändra, markeras med fet stil .
Eventuella strykningar ska i sådana fall markeras enligt följande: [...].
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
ÄRENDETS GÅNG....................................................................................................................6
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets förordning om märkning av däck vad gäller drivmedelseffektivitet och andra väsentliga parametrar
(14639/6/2009 – C7‑0287/2009 – 2008/0221(COD) )
(Medbeslutandeförfarandet: andra behandlingen)
Europaparlamentet utfärdar denna resolution
– med beaktande av rådets gemensamma ståndpunkt (14639/6/2009 – C7‑0287/2009 ),
– med beaktande av parlamentets ståndpunkt vid första behandlingen av ärendet
Antagna texter från sammanträdet 22.4.2009, P7_TA(2009)0248 . , en behandling som avsåg kommissionens förslag till Europaparlamentet och rådet ( KOM(2008)0779 ),
– med beaktande av kommissionens ändrade förslag ( KOM(2009)0348 ),
– med beaktande av artikel 72 i arbetsordningen,
– med beaktande av andrabehandlingsrekommendationen från utskottet för industrifrågor, forskning och energi ( A7‑0076/2009 ).
1.
4.
ÄRENDETS GÅNG
Titel
Märkning av däck avseende bränsleeffektivitet*
Referensnummer
14639/6/2009 – C7-0287/2009 – 2008/0221(COD)
Parlamentets första behandling – P ‑ nummer
22.4.2009 T6-0248/2009
Kommissionens förslag
KOM(2008)0779 – C6-0411/2008
Kommissionens ändrade förslag
KOM(2009)0348
Ansvarigt utskott
Tillkännagivande i kammaren
ITRE
Föredragande
Utnämning
Ivo Belet
17.12.2008
Antagande
23.11.2009
Slutomröstning: resultat
+:
–:
0:
37
Slutomröstning: närvarande ledamöter
Slutomröstning: närvarande suppleanter
Ilda Figueiredo, Françoise Grossetête, Yannick Jadot, Werner Langen, Hermann Winkler
Slutomröstning: närvarande suppleanter (art.
187.2)
Anna Záborská
A7-0107/2010
BETÄNKANDE
om begäran om upphävande av Miloslav Ransdorfs immunitet
(2009/2208(IMM))
Utskottet för rättsliga frågor
Föredragande:
Francesco Enrico Speroni
PE 439.329v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT...........................................................3
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.......................................................9
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
om begäran om upphävande av Miloslav Ransdorfs immunitet
( 2009/2208(IMM) )
Europaparlamentet fattar detta beslut
– med beaktande av den begäran om upphävande av Miloslav Ransdorfs immunitet som översändes av den behöriga tjeckiska myndigheten den 16 september 2009 och som tillkännagavs i kammaren den 23 november 2009,
– med beaktande av Europeiska unionens domstols domar av den 12 maj 1964 och den 10 juli 1986
Dom av den 12 maj 1964 i mål 101/63, Wagner mot Fohrmann och Krier, REG 1964, s.
383; svensk specialutgåva, volym 1, s.
203, och dom av den 10 juli 1986 i mål 149/85, Wybot mot Faure m.fl., REG 1986, s.
703. ,
– med beaktande av betänkandet från utskottet för rättsliga frågor ( A7‑0107/2010 ), och av följande skäl:
A. Miloslav Ransdorf är ledamot i Europaparlamentet.
Europaparlamentet beslutar att upphäva Miloslav Ransdorfs immunitet.
2.
1.
2.
3.
Genom sin handling bröt Ransdorf mot bestämmelserna i artikel 5/1h i vägtrafiklagen (lag nr 361/2000).
Det föreligger ett fall av grundad misstanke om att en straffbar handling – förorsakande av kroppsskada – begicks, i enlighet med artikel 223 i lag nr 140/1961 (brottsbalken), där följande anges: ” En person som skadar en annans hälsa genom oaktsamhet, genom att bryta mot en viktig skyldighet till följd av anställning, yrke, ställning eller tjänst, eller en skyldighet enligt lagen, ska straffas med frihetsberövande i högst ett år eller förbud att utöva en (särskild) verksamhet. ”
Enligt artikel 9 i brottsbalken ska den som bryter mot lagen ställas till svars för detta.
Artikel 65 i brottsbalken om upphörande av samhällsfara på grund av straffbar handling – enligt vilken ” den straffbara handling som utgjorde en fara för samhället när den begicks upphör att vara straffbar när den fara för samhället som handlingen medförde undanröjs, till följd av händelsernas utveckling eller genom gärningsmannens egen försorg ” – är inte tillämplig i detta fall.
II.
LAGSTIFTNINGEN OCH ALLMÄNNA ÖVERVÄGANDEN SOM RÖR IMMUNITETEN FÖR LEDAMÖTERNA AV EUROPAPARLAMENTET
1.
Artiklarna 8 och 9 i protokollet om Europeiska gemenskapernas immunitet och privilegier av den 8 april 1965 lyder som följer:
Artikel 8:
Europaparlamentets ledamöter får inte förhöras, kvarhållas eller lagföras på grund av yttranden de gjort eller röster de avlagt under utövandet av sitt ämbete.
Artikel 9:
Under Europaparlamentets sessioner ska dess ledamöter åtnjuta,
a) vad avser deras egen stats territorium, den immunitet som beviljas parlamentsledamöter i deras land,
b) vad avser alla andra medlemsstaters territorium, immunitet vad gäller alla former av kvarhållande och lagföring.
Immuniteten skall även vara tillämplig på ledamöterna under resan till och från Europaparlamentets mötesplats.
Immuniteten kan inte åberopas av en ledamot som tas på bar gärning och kan inte hindra Europaparlamentet att utöva sin rätt att upphäva en av dess ledamöters immunitet.
2.
Förfarandet i Europaparlamentet styrs av artiklarna 6 och 7 i arbetsordningen.
De relevanta bestämmelserna lyder som följer:
Artikel 6 – Upphävande av immunitet
1.
Parlamentet ska vid utövandet av sina befogenheter i frågor som rör immunitet och privilegier i första hand försöka upprätthålla parlamentets integritet som en demokratisk lagstiftande församling och befästa ledamöternas oberoende när dessa fullgör sina åligganden.
(...)
3.
Varje begäran om fastställelse av immunitet och privilegier som en ledamot eller före detta ledamot lämnar in till talmannen ska tillkännages i kammaren och hänvisas till behörigt utskott.
(...)
Artikel 7 – Immunitetsförfaranden:
1.
Behörigt utskott ska utan dröjsmål, och i den ordning de inkommit, pröva varje begäran om upphävande av immunitet och varje begäran om fastställelse av immunitet eller privilegier.
2.
Utskottet ska lägga fram ett förslag till beslut, i vilket utskottet endast ska rekommendera huruvida en begäran om upphävande av immuniteten eller en begäran om fastställelse av immunitet och privilegier ska bifallas eller avslås.
3.
Utskottet kan uppmana den berörda myndigheten att förse utskottet med alla upplysningar och preciseringar som det anser sig behöva för att kunna ta ställning till om immuniteten bör upphävas eller fastställas.
De har rätt att låta sig företrädas av en annan ledamot.
4.
Om en begäran om upphävande av immunitet hänför sig till flera gärningar kan upphävande av immuniteten beträffande var och en av dessa gärningar bli föremål för ett enskilt beslut.
I utskottets betänkande kan det i undantagsfall föreslås att upphävandet av immuniteten endast ska beröra åtalet och att ledamoten, så länge som det inte finns någon lagakraftvunnen dom varken kan gripas, anhållas, häktas eller utsättas för någon annan åtgärd som skulle förhindra ledamoten att utföra sina åligganden i enlighet med uppdraget som ledamot av Europaparlamentet.
(...)
6.
7.
Utskottet får emellertid under inga omständigheter uttala sig i skuldfrågan, eller på annat sätt yttra sig över ledamoten eller om det riktiga i att väcka åtal för de uttalanden eller handlingar som tillskrivs ledamoten, inte ens vid tillfällen där utskottet genom prövning av en begäran erhåller detaljerad kunskap i fallet.
(...)
III.
MOTIVERING TILL DET FÖRESLAGNA BESLUTET
1.
Först och främst är tillämpligheten av artikel 8 i protokollet självfallet inte aktuell, av det uppenbara skälet att personskada som orsakats av en bilist på intet sätt kan jämställas med yttranden som gjorts eller röster som avlagts under utövandet av ämbetet som ledamot av Europaparlamentet.
2.
När det gäller artikel 9 är det, med tanke på att klagomålet mot Ransdorf avser handlingar som begicks i Tjeckien och att han var tjeckisk medborgare då de begicks, endast följande del som är tillämplig: ” Under Europaparlamentets sessioner ska dess ledamöter åtnjuta, a) vad avser deras egen stats territorium, den immunitet som beviljas parlamentsledamöter i deras land ” .
3.
Räckvidden för den parlamentariska immuniteten i Tjeckien är mycket lik den som säkrar Europaparlamentets sätt att fungera, som grundar sig på protokollet om immunitet och privilegier.
I lag nr 141/1961 (dvs. brottsbalken), artikel 10 om uteslutande från domsrätten för de organ som är behöriga för straffrättsliga förfaranden, anges följande: ” Personer som har privilegier eller immunitet enligt nationell eller internationell lagstiftning ska uteslutas från domsrätten för de organ som är behöriga för straffrättsliga förfaranden enligt denna lag ”.
Om respektive kammare inte ger sitt samtycke är straffrättsliga åtgärder uteslutna för all framtid. ”
Med andra ord kan ett straffrättsligt förfarande mot Ransdorf enligt gällande tjeckisk lagstiftning inledas endast om hans immunitet upphävs.
IV.
SLUTSATS
Med ovanstående överväganden som underlag och efter att ha övervägt skälen för och emot upphävande av ledamotens immunitet rekommenderar utskottet för rättsliga frågor att Europaparlamentet ska upphäva Miloslav Ransdorfs parlamentariska immunitet.
Om respektive kammare inte ger sitt samtycke är straffrättsliga åtgärder uteslutna för all framtid.”
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
22.3.2010
Slutomröstning: resultat
+:
–:
0:
19
Slutomröstning: närvarande ledamöter
Raffaele Baldassarre, Luigi Berlinguer, Marielle Gallo, Gerald Häfner, Klaus-Heiner Lehne, Jiří Maštálka, Bernhard Rapkay, Evelyn Regner, Francesco Enrico Speroni, Dimitar Stoyanov, Alexandra Thein, Diana Wallis, Cecilia Wikström, Zbigniew Ziobro, Tadeusz Zwiefka
Slutomröstning: närvarande suppleanter
Sajjad Karim, Vytautas Landsbergis, Kurt Lechner, Eva Lichtenberger
A7-0142/2010
*
BETÄNKANDE
om förslaget till rådets förordning om gemenskapens ekonomiska stöd till avvecklingen av enheterna 1–4 i kärnkraftverket Kozloduj i Bulgarien - ”Kozloduj-programmet”
(KOM(2009)0581 – C7‑0289/2009 – 2009/0172(NLE))
Utskottet för industrifrågor, forskning och energi
Föredragande:
Rebecca Harms
PE 438.485v02-00
Teckenförklaring
* Samrådsförfarandet
*** Samtyckesförfarandet
***I Medbeslutandeförfarandet (första behandlingen)
***II Medbeslutandeförfarandet (andra behandlingen)
***III Medbeslutandeförfarandet (tredje behandlingen)
(Angivet förfarande baseras på den rättsliga grund som kommissionen föreslagit.)
Ändringsförslag till lagtexter
Eventuella strykningar ska i sådana fall markeras enligt följande: [...].
Kursiv stil används för att uppmärksamma berörda avdelningar på eventuella problem i texten.
Kursiveringen används för att markera ord eller textavsnitt som det finns skäl att korrigera innan den slutliga texten produceras (exempelvis om en språkversion innehåller uppenbara fel eller saknar textavsnitt).
Dessa förslag underställs berörda avdelningar för godkännande.
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING..........................................................................................................................22
YTTRANDE från budgetutskottet ............................................................................27
YTTRANDE från utskottet för miljö, folkhälsa och livsmedelssäkerhet 32
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................46
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till rådets förordning gemenskapens ekonomiska stöd till avvecklingen av enheterna 1–4 i kärnkraftverket Kozloduj i Bulgarien - ”Kozloduj-programmet”
( KOM(2009)0581 – C7‑0289/2009 – 2009/0172(NLE) )
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till rådet ( KOM(2009)0581 ),
– med beaktande av artikel 30 i akten om villkoren för Republiken Bulgariens och Rumäniens anslutning till de fördrag som ligger till grund för Europeiska Unionen och om anpassning av fördragen, med avseende på reaktorerna 1–4 i kärnkraftverket Kozloduj i Bulgarien,
– med beaktande av meddelandet från kommissionen till rådet och Europaparlamentet ”Kärnteknisk säkerhet i Europeiska unionen” ( KOM(2002)0605 ),
– med beaktande av artikel 203 i Euratomfördraget, i enlighet med vilken rådet har hört parlamentet ( C7‑0289/2009 ),
– med beaktande av artikel 55 i arbetsordningen,
– med beaktande av betänkandet från utskottet för industrifrågor, forskning och energi och yttrandena från budgetutskottet och utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A7‑0142/2010 ).
Europaparlamentet påpekar att det årliga beloppet för programmet för avveckling av kärnkraftverket Kozloduj kommer att fastställas under det årliga budgetförfarandet i enlighet med bestämmelserna i punkt 38 i det interinstitutionella avtalet av den 17 maj 2006.
5.
Ändringsförslag
1
Förslag till förordning
Skäl 1
Kommissionens förslag
Ändringsförslag
(1) Bulgarien lovade att stänga enheterna 1 och 2 samt 3 och 4 i kärnkraftverket Kozloduj till den 31 december 2002 respektive den 31 december 2006, och att därefter avveckla dessa enheter.
Europeiska unionen har förklarat sig vara villig att fram till 2009 ge fortsatt ekonomiskt stöd till Bulgariens avvecklingsverksamhet som en förlängning av föranslutningsstödet inom ramen för Phareprogrammet.
(1) Under anslutningsförhandlingarna 2005 gick Bulgarien med på att stänga enheterna 1 och 2 samt 3 och 4 i kärnkraftverket Kozloduj till den 31 december 2002 respektive den 31 december 2006, och att därefter avveckla dessa enheter.
Europeiska unionen har förklarat sig vara villig att fram till 2009 ge fortsatt ekonomiskt stöd till Bulgariens avvecklingsverksamhet som en förlängning av föranslutningsstödet inom ramen för Phareprogrammet.
Vid tiden för anslutningsförhandlingarna försäkrade EU också att det ekonomiska stödet skulle övervägas i en övergripande översyn av gemenskapsstödet för perioden 2007–2013.
Ändringsförslag
2
Förslag till förordning
Skäl 2
Kommissionens förslag
Ändringsförslag
(2) I 2005 års fördrag om Republiken Bulgariens och Rumäniens anslutning till Europeiska unionen, och särskilt i artikel 30 i akten om villkoren för Republiken Bulgariens och Rumäniens anslutning till de fördrag som ligger till grund för Europeiska Unionen och om anpassning av fördragen föreskrivs med anledning av Bulgariens åtagande att stänga enheterna 3 och 4 i kärnkraftverket Kozloduj ett stödprogram (nedan kallat Kozloduj-programmet) med en budget på 210 miljoner euro för perioden 2007–2009.
(2) I 2005 års fördrag om Republiken Bulgariens och Rumäniens anslutning till Europeiska unionen, och särskilt i artikel 30 i akten om villkoren för Republiken Bulgariens och Rumäniens anslutning till de fördrag som ligger till grund för Europeiska Unionen och om anpassning av fördragen föreskrivs med anledning av Bulgariens åtagande att stänga enheterna 3 och 4 i kärnkraftverket Kozloduj ett stödprogram (nedan kallat Kozloduj‑programmet) med en budget på 210 miljoner euro för perioden 2007–2009 .
I programmet ingår stöd för att täcka kapacitetsförlusten till följd av stängningen av kärnkraftverket Kozloduj .
Motivering
Syftet med det ekonomiska stödet är att som ett led i Bulgariens integration i Europeiska unionen lösa den svåra frågan om stängningen av kärnkraftverket Kozloduj med den ekonomiska belastning som detta innebär för Bulgarien.
Ändringsförslag
3
Förslag till förordning
Skäl 2a (nytt)
Kommissionens förslag
Ändringsförslag
(2a) Gemenskapens principer om solidaritet och likabehandling kräver ett rättvist tillvägagångssätt, nu som förr, gentemot medlemsstater i behov av ekonomiskt stöd för att avveckla kärnkraftverk, enligt åtaganden i deras anslutningsfördrag eller tilläggsprotokoll om a tt stänga enheter vid kärnkraft verk.
Ändringsförslag
4
Förslag till förordning
Skäl 4
Kommissionens förslag
Ändringsförslag
(4) EU har noterat de insatser och stora framsteg som Bulgarien har gjort med förberedelsefasen för avvecklingen inom ramen för Kozloduj-programmet, där de gemenskapsmedel som anslagits fram till 2009 har använts; likaså har EU noterat behovet av ytterligare ekonomiskt stöd efter 2009 för att fortsätta med den konkreta nedmonteringen.
(4) EU har noterat de insatser och stora framsteg som Bulgarien har gjort med förberedelsefasen för avvecklingen inom ramen för Kozloduj-programmet, där de gemenskapsmedel som anslagits fram till 2009 har använts; likaså har EU noterat behovet av ytterligare ekonomiskt stöd efter 2009 för att fortsätta med den konkreta nedmonteringen i enlighet med anslutningsfördraget från 2005, samtidigt som man tillämpar högsta möjliga säkerhetsstandarder .
Ändringsförslag
5
Förslag till förordning
Skäl 5
Kommissionens förslag
Ändringsförslag
(5) Det är också viktigt att använda kärnkraftverket Kozlodujs egna resurser, eftersom man därigenom bibehåller den nödvändiga expertisen och samtidigt lindrar de sociala och ekonomiska följderna av den tidigarelagda stängningen genom att sysselsätta personal från det stängda kärnkraftverket.
Fortsatt ekonomiskt stöd är därför en förutsättning för att den nödvändiga s äkerhetsstandarden ska kunna upprätthållas.
(5) Det är också viktigt att använda kärnkraftverket Kozlodujs egna resurser, eftersom man därigenom bibehåller den nödvändiga expertisen , förbättrar kunskapen och kompetensen och samtidigt lindrar de sociala och ekonomiska följderna av den tidigarelagda stängningen genom att sysselsätta personal från det stängda kärnkraftverket.
Fortsatt ekonomiskt stöd är därför en förutsättning för att nödvändiga säkerhets-, folkhälso- och miljökrav ska kunna upprätthållas.
Ändringsförslag
6
Förslag till förordning
Skäl 6
Kommissionens förslag
Ändringsförslag
(6) Europeiska unionen noterar också behovet av ekonomiskt stöd för att fortsätta lindringsåtgärderna inom energisektorn med tanke på den omfattande kapacitetsförlusten till följd av kärnkraftsenheternas stängning, och de följder för regionens försörjningstrygghet som detta medför .
(6) Europeiska unionen noterar också behovet och nödvändigheten av ekonomiskt stöd till fortsatta framsteg på väg mot en energieffektivare ekonomi, något som kommer att positivt påverka försörjningstryggheten, elpriserna och mängden utsläppta växthusgaser i Bulgarien.
Eftersom Bulgarien måste komma längre med slutförvaringen av bestrålade bränsleelement och högaktivt avfall och eftersom slutförvaringen av alla de radioaktiva ämnen som uppstått i samband med stängningen av kärnkraftverket Kozloduj är mycket viktig och kräver noggrann planering bör unionen hjälpa Bulgarien med att hitta lösningar på slutförvaringsfrågan, vilket vid behov kan ske utgående från en utredning som bulgariska staten gjort om slutförvaringen av alla de radioaktiva ämnen som uppstått i samband med avvecklingen .
Ändringsförslag
7
Förslag till förordning
Skäl 6a (nytt)
Kommissionens förslag
Ändringsförslag
(6a) Förlusten av produktionskapacitet till följd av den tidigarelagda stängningen av kärnkraftverket Kozlodujs enheter 1–4 har lett till en betydande ökning av utsläppsvolymen för växthusgaser, beräknad till 15 TWh för perioden 2011 ‑2013 med koldioxidekvivalenter på cirka 1,2 Gg/GWh, vilket för Bulgariens del har betytt ytterligare påverkan av omkring 18 000 Gg eller 18 000 kt koldioxidekvivalenter.
Koldioxidutsläppen måste därför minskas ännu mer .
Ändringsförslag
8
Förslag till förordning
Skäl 6b (nytt)
Kommissionens förslag
Ändringsförslag
(6b) Unionen erkänner behovet av att dämpa skadeverkningarna på miljön och minska utsläpp en som har ökat eftersom den ersättande kapaciteten mestadels kommit från brunkolskraftverk.
Ändringsförslag
9
Förslag till förordning
Skäl 6c (nytt)
Kommissionens förslag
Ändringsförslag
(6c) Ekonomiskt stöd från EU kan behövas till åtgärder som lindrar de sociala och ekonomiska följderna av stängningen av kärnkraftverket Kozlodujs enheter 1–4, såsom omskolningsprogram för att berörd personal ska kunna använda sin kompetens i andra sektorer, till exempel inom industriell forskning eller förnybar energi.
Ändringsförslag
10
Förslag till förordning
Skäl 7
Kommissionens förslag
Ändringsförslag
(7) Under perioden 2010–2013 bör därför ett belopp på 300 miljoner euro avsättas i Europeiska unionens allmänna budget för finansieringen av nedläggningen av kärnkraftverket Kozloduj.
Av detta belopp bör 180 miljoner euro användas till stöd för avvecklingsprogrammet och återstoden, 120 miljoner euro, till stöd för både energieffektivitets- och energisparåtgärder.
Ändringsförslag
11
Förslag till förordning
Skäl 7a (nytt)
Kommissionens förslag
Ändringsförslag
Uppgraderingen av anläggnings infrastrukturen enligt projekt 4 får innefatta endast åtgärder som hänför sig till avvecklingen av enheterna 1–4.
__________
1 SE K(2009) 1431.
Ändringsförslag
12
Förslag till förordning
Skäl 8
Kommissionens förslag
Ändringsförslag
(8) Gemenskapens budgetanslag för avveckling bör inte leda till snedvridning av konkurrensen för energiförsörjningsföretag på energimarknaden i unionen.
Dessa anslag bör även användas för att finansiera åtgärder för att kompensera den minskade produktionskapaciteten i linje med det relevanta regelverket.
(8) Gemenskapens budgetanslag för avveckling bör inte leda till snedvridning av konkurrensen för energiförsörjningsföretag på energimarknaden i unionen.
Dessa anslag bör även användas för att finansiera åtgärder för energieffektivitet och energisparande i linje med det relevanta regelverket samt bestämmelserna för den gemensamma europeiska energimarknadens funktion .
Ändringsförslag
13
Förslag till förordning
Skäl 10
Kommissionens förslag
Ändringsförslag
(10) EBRD har bland annat till uppgift att förvalta de offentliga medel som har anslagits till programmen för avveckling av kärnkraftverk och att följa upp programmens ekonomiska förvaltning för att se till att de offentliga medlen används på bästa möjliga sätt.
(10) EBRD har bland annat till uppgift att förvalta de offentliga medel som har anslagits till programmen för avveckling av de enheter vid kärnkraftverk som omfattades av avtal om stängning i samband med anslutningen.
EBRD följer upp programmens ekonomiska förvaltning för att se till att de offentliga medlen används på bästa möjliga sätt.
Ändringsförslag
14
Förslag till förordning
Skäl 11
Kommissionens förslag
Ändringsförslag
(11) För att största möjliga effektivitet ska garanteras bör bästa tillgängliga tekniska expertis användas vid avvecklingen av kärnkraftverket Kozloduj, med hänsyn tagen till vilken typ av reaktorer som ska stängas och de tekniska specifikationer som gäller för dem.
(11) För att största möjliga effektivitet ska garanteras och de eventuella konsekvenserna för miljön minimeras bör bästa tillgängliga tekniska expertis användas vid avvecklingen av enheterna 1–4 i kärnkraftverket Kozloduj, med hänsyn tagen till vilken typ av reaktorer som ska stängas och de tekniska specifikationer som gäller för dem.
Ändringsförslag
15
Förslag till förordning
Skäl 11a (nytt)
Kommissionens förslag
Ändringsförslag
__________
1 EUT L 124, 17.5.2005, s.
1.
Ändringsförslag
16
Förslag till förordning
Skäl 12
Kommissionens förslag
Ändringsförslag
(12) Avvecklingen av kärnkraftverket Kozloduj bör ske i enlighet med relevant miljölagstiftning, bland annat rådets direktiv 85/337/EEG av den 27 juni 1985 om bedömning av inverkan på miljön av vissa offentliga och privata projekt.
(12) Avvecklingen av enheterna 1–4 i kärnkraftverket Kozloduj bör ske i enlighet med Bulgariens nationella lagstiftning, dess licensavtal och relevant miljölagstiftning, bland annat rådets direktiv 85/337/EEG av den 27 juni 1985 om bedömning av inverkan på miljön av vissa offentliga och privata projekt.
Ändringsförslag
17
Förslag till förordning
Skäl 12a (nytt)
Kommissionens förslag
Ändringsförslag
De lindrande åtgärderna inom energisektorn i form av energieffektivitet och förnybar energi bör stödjas genom en särskild bulgarisk nationell strategi.
__________
1 EGT L 159, 29.6.1996, s.
1.
Ändringsförslag
18
Förslag till förordning
Skäl 12b (nytt)
Kommissionens förslag
Ändringsförslag
(12b) Principerna om ekonomi, effektivitet och ändamålsenlighet för de anslagna medlen kan säkras genom utvärdering och effektivitetsrevisioner av de program som tidigare finansierats.
Motivering
Det behövs garantier för att man vid tilldelningen av medel genom projekten under 2007‑2009 har tagit hänsyn till sund ekonomisk förvaltning såsom denna definieras i budgetförordningen.
Ändringsförslag
19
Förslag till förordning
Skäl 13a (nytt)
Kommissionens förslag
Ändringsförslag
(13a) De villkor som gäller metoden för gemensam förvaltning vid genomförandet av budgeten fastställs i artiklarna 53d, 108a och 165 i rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget 1 , och i artiklarna 35 och 43 i kommissionens förordning (EG, Euratom) nr 2342/2002 av den 23 december 2002 om genomförandebestämmelser för rådets förordning (EG, Euratom) nr 1605/2002 med budgetförordning för Europeiska gemenskapernas allmänna budget 2 .
__________
1 EGT L 248, 16.9.2002, s.
1.
2 EGT L 357, 31.12.2002, s.
1.
Motivering
Enligt budgetförordningen och genomförandebestämmelserna har kommissionen rätt att genomföra sin budget genom gemensam förvaltning med internationella organisationer om dessa organisationer tillämpar standarder som ger garantier som motsvarar internationellt godkända standarder för, som ett minimum, reglerna för räkenskaper, revision, intern kontroll och upphandling.
Ändringsförslag
20
Förslag till förordning
Skäl 13b (nytt)
Kommissionens förslag
Ändringsförslag
(13b) Fallet med Kozloduj bör tjäna som exempel och kommissionen bör utarbeta en fullständig och exakt avvecklingsbudget för att en analys och beräkning av kostnaderna för framtida avveckling av kärnkraftverk ska kunna göras.
Ändringsförslag
21
Förslag till förordning
Artikel 1
Kommissionens förslag
Ändringsförslag
I denna förordning fastställs ett program med detaljerade genomförandebestämmelser för gemenskapens ekonomiska bidrag till avvecklingen av enheterna 1–4 i kärnkraftverket Kozloduj, och följderna för Bulgarien av stängningen av dessa enheter (nedan kallat Kozloduj-programmet).
I denna förordning fastställs ett program med detaljerade genomförandebestämmelser för gemenskapens ekonomiska bidrag till det fortsatta arbetet med avvecklingen av enheterna 1–4 i kärnkraftverket Kozloduj, och följderna för miljön, ekonomin och försörjningstryggheten i Bulgarien av den tidiga stängningen av dessa enheter (nedan kallat Kozloduj-programmet).
Motivering
Någon kompensation skulle inte behövas om alla kraftverk fortsatte vara i drift under hela den livslängd de konstruerats för.
Ändringsförslag
22
Förslag till förordning
Artikel 2
Kommissionens förslag
Ändringsförslag
Syftet med gemenskapens stöd till Kozloduj-programmet i enlighet med denna förordning är att ekonomiskt stödja åtgärder inom ramen för avvecklingen av kärnkraftverket Kozloduj , åtgärder för miljöuppgradering i linje med regelverket och för modernisering av den konventionella produktionskapaciteten för att ersätta produktionskapaciteten för de fyra reaktorerna vid kärnkraftverket Kozloduj samt andra åtgärder som följer av beslutet att stänga och avveckla detta kärnkraftverk och som bidrar till den nödvändiga omstruktureringen, miljöuppgraderingen och moderniseringen av energiproduktionen och överförings- och distributionssektorerna i Bulgarien samt till att förbättra energiförsörjningstryggheten och energieffektiviteten i Bulgarien.
Syftet med gemenskapens stöd till Kozloduj-programmet i enlighet med denna förordning är i första hand att ekonomiskt stödja åtgärder inom ramen för avvecklingen av enheterna 1–4 i kärnkraftverket Kozloduj .
Stödet ska också inriktas på åtgärder för miljöuppgradering i linje med regelverket och för modernisering av produktionskapaciteten för att ersätta produktionskapaciteten för de fyra reaktorerna vid kärnkraftverket Kozloduj samt andra åtgärder som följer av beslutet att stänga och avveckla dessa enheter och som bidrar till den nödvändiga omstruktureringen, miljöuppgraderingen och moderniseringen och förstärkningen av energiproduktionen och överförings- och distributionssektorerna i Bulgarien samt till att förbättra energiförsörjningstryggheten , försörjningsnormerna, energieffektiviteten och användningen av förnybar energi i Bulgarien och samtidigt uppmuntra till energisparande och främja förnybar energi .
Ekonomiskt stöd kan också ges för att lindra de sociala och ekonomiska följder som övergången för med sig för de berörda samhällena, exempelvis genom att skapa nya hållbara arbetstillfällen och industrier.
Ändringsförslag
23
Kommissionens förslag
Ändringsförslag
1.
Det finansiella referensbelopp som krävs för genomförandet av Kozloduj‑programmet för perioden 1 januari 2010–31 december 2013 fastställs härmed till 300 miljoner euro.
1.
Det finansiella referensbelopp enligt punkt 38 i IIA av den 17 maj 2006 som krävs för genomförandet av Kozloduj‑programmet för perioden 1 januari 2010–31 december 2013 fastställs härmed till 300 miljoner euro.
Ändringsförslag
24
Kommissionens förslag
Ändringsförslag
2.
De årliga anslagen ska beviljas av budgetmyndigheten inom ramen för budgetplanen.
2.
De årliga anslagen ska beviljas av budgetmyndigheten inom ramen för budgetplanen och enligt kraven i avvecklingsprocessen .
Motivering
Genomförandet av avtalet om Kozloduj-programmet bör vara en smidig och framgångsrik process, där Republiken Bulgarien är ekonomiskt och socialt delaktig i EU.
Ändringsförslag
25
Kommissionens förslag
Ändringsförslag
3.
3.
Anslagen för Kozloduj-programmet ska ses över under perioden 1 januari 2010–31 december 2013 för att man ska kunna ta hänsyn till gjorda framsteg under programmets genomförande och till de långsiktiga effekterna på och konsekvenserna för miljön, ekonomin och försörjningstryggheten av den tidiga stängningen av enheterna 1–4 i kärnkraftverket Kozloduj , och för att man ska kunna se till att programplaneringen och fördelningen av resurserna grundas på faktiska betalningsbehov och faktisk absorberingskapacitet.
Ändringsförslag
26
Kommissionens förslag
Ändringsförslag
2.
2.
De ska följa EU:s regler för offentlig upphandling.
Ändringsförslag
27
Kommissionens förslag
Ändringsförslag
1.
Kommissionen får, direkt genom sina anställda eller genom någon annan behörig organisation den valt, utföra en granskning av hur bidraget har använts.
Granskningen får utföras under hela löptiden för avtalet mellan gemenskapen och EBRD om att tillhandahålla gemenskapsmedel till internationella fonden för avvecklingsstöd till Kozloduj samt under fem år efter dagen för utbetalning av den sista bidragsdelen.
I förekommande fall kan revisionens resultat leda till att kommissionen beslutar om återkrav.
1.
Kommissionen ska övervaka och får, direkt genom sina anställda eller genom någon annan behörig organisation den valt, utföra en granskning av hur bidraget har använts.
Granskningen får utföras under hela löptiden för avtalet mellan gemenskapen och EBRD om att tillhandahålla gemenskapsmedel till internationella fonden för avvecklingsstöd till Kozloduj samt under fem år efter dagen för utbetalning av den sista bidragsdelen.
I förekommande fall kan granskningens resultat leda till att kommissionen beslutar om återkrav.
Finansieringen av sådana granskningar och eventuella andra bedömningar omfattas inte av budgeten för avvecklingsstöd .
Ändringsförslag
28
Kommissionens förslag
Ändringsförslag
2.
Kommissionens personal och extern personal med fullmakt från kommissionen ska ges lämplig tillgång till mottagarens kontorslokaler och till alla upplysningar, även i elektronisk form, som behövs för att utföra granskningen.
2.
Kommissionens personal och extern personal med fullmakt från kommissionen ska ges lämplig tillgång till mottagarens kontorslokaler och till alla upplysningar, även i elektronisk form, som behövs för att utföra granskningen.
I granskningen ska också ingå en undersökning av rådande tillståndsläge för avvecklingen.
Motivering
För att garantera att resurserna sätts in i rätt tid och att det bättre övervakas att de används till det de är avsedda för.
Ändringsförslag
29
Kommissionens förslag
Ändringsförslag
Revisionsrätten ska ha samma rättigheter som kommissionen, särskilt när det gäller tillträde.
Revisionsrätten och Europaparlamentet ska ha samma rättigheter som kommissionen, särskilt när det gäller tillträde.
Ändringsförslag
30
Förslag till förordning
Artikel 7
Kommissionens förslag
Ändringsförslag
Kommissionen ska se till att denna förordning tillämpas och regelbundet rapportera till Europaparlamentet och rådet.
Efterhandsutvärderingen ska innehålla en fullständig och exakt kostnadsbudget för avvecklingen av ett kärnkraftverk så att man kan planera för framtida avvecklingsprojekt.
Den ska också analysera ekonomiska, sociala och miljömässiga kostnader, med fokus på frigjord reststrålning och konsekvenser för försörjningstryggheten.
Ändringsförslag
31
Förslag till förordning
Artikel 7a (ny)
Kommissionens förslag
Ändringsförslag
Artikel 7a
Kommissionen ska utgående från internationellt godkända standarder göra en överensstämmelsebedömning av åtminstone reglerna för räkenskaper, revision, intern kontroll och upphandling vid Europeiska banken för återuppbyggnad och utveckling, innan de sammanlagda överenskomna bidragen undertecknas.
Motivering
Enligt budgetförordningen och genomförandebestämmelserna har kommissionen rätt att genomföra sin budget genom gemensam förvaltning med internationella organisationer om dessa organisationer tillämpar standarder som ger garantier som motsvarar internationellt godkända standarder åtminstone för reglerna för räkenskaper, revision, intern kontroll och upphandling.
MOTIVERING
I samband med de central- och östeuropeiska staternas anslutning blev frågan om hur kärnkraften användes där samt om hur det radioaktiva avfallet hanterades aktuell inom Europeiska unionen.
Anslutningsländerna hade objektivt sett mindre rigorösa normer för säkerhet och detta gav anledning till påverkan och ekonomiskt stöd för att förbättra skyddet för människor och miljö.
Det var mestadels först efter anslutningen som man började införa olika juridiska och tekniska bestämmelser för kärnkraftsavveckling.
Och nu liksom förr finns det endast en begränsad kapacitet att tillgå för omhändertagande av det avfall som uppkommer i samband med avvecklingen.
Somliga av de stater som anslutit sig har inte ens i dag, lika litet som förr, fastställt om de bestrålade bränsleelementen ska upparbetas eller gå till direkt geologisk slutförvaring.
KOM(2008)0542 .
Detta kommer utan tvivel att påverka hur energiskt man i dessa stater driver på framstegen i frågan om slutförvaring, framför allt av högaktivt avfall och bestrålade bränsleelement.
Detta gäller framför allt också för Bulgarien.
Inte heller har dessa stater någon obligatorisk planering av hur mer långlivat låg- och medelaktivt avfall ska hanteras.
Den nuvarande strategin går ut på att bestrålade bränsleelement från Bulgarien i huvudsak upparbetas i Ryssland.
Republiken Bulgarien: Third National Report on Fulfilment of the Obligations on the Joint Convention on the safety of Spent Fuel Management and on the Safety of Radioactive Waste Management, Sofia, september 2008.
Detta innebär att belastningen av människor och miljö vid hanteringen av den farligaste produkten från användningen av kärnkraft väsentligen förläggs till en stat som inte är medlem av EU.
Upparbetningen innefattar dels stora säkerhetstekniska risker (mycket höga utsläpp vid normal drift och risk för svåra olyckor) och dels en stor risk för kärnvapenspridning, alltså för att kärnkraften används för militära ändamål.
Upparbetning kan inte accepteras som metod för bortskaffning av bestrålade bränsleelement.
De bristfälligheter som beskrivits i det föregående tangerar också Europeiska unionens säkerhetsintressen.
Därför är det viktigt att de central- och östeuropeiska staterna snabbt gör framsteg med slutförvaringen av bestrålade bränsleelement och högaktivt avfall.
Det förslag till förordning som kommissionen lagt fram i dokument KOM(2009)0581 syftar till att trygga ekonomiskt stöd till nedläggningen av reaktorerna 1–4 i kärnkraftverket i Kozloduj i Bulgarien samt till hanteringen av de radioaktiva ämnen som blir aktuella i samband med denna.
Kommissionen motiverar sitt förslag med att republiken Bulgarien av historiska skäl inte avsatt tillräckliga resurser för nedmonteringen av reaktorerna samt med de skyldigheter i fråga om förtida stängning av Kozloduj 1–4, vilka ingår i anslutningsakten.
Föredraganden instämmer med denna motivering och betonar att vardera parten måste rätta sig efter anslutningsaktens bestämmelser om nedläggning av reaktorerna Kozloduj 1–4.
Om det inte ges något ekonomiskt stöd från gemenskapen kan följden enligt kommissionen bli att säkerheten på ort och ställe ytterligare försämras och att enheterna 3 och 4 åter tas i bruk och detta är något vi måste undvika.
Kommissionen hade fastställt att det i fråga om enheterna Kozloduj 1–4 ”inte är sannolikt att man kommer att kunna uppnå en hög kärnteknisk säkerhetsnivå” och under 2002 bekräftat att de måste avvecklas
KOM(2002)0605 . , vilket än en gång bekräftats 2009
SEK(2009)1431 . .
Föredraganden stöder denna uppfattning, men konstaterar dessutom att just denna reaktortyp visserligen utmärks av särskilt otillräcklig säkerhet, men att säkerheten också för alla andra reaktortyper är begränsad och att svåra olyckor inte går att utesluta för någon enda reaktortyp eller i något enda land.
Enheterna 1–2 i Kozloduj stängdes som ett led i förberedelserna inför avveckling vid utgången av 2002 och samma skedde med enheterna 3–4 vid utgången av 2006.
I de båda enheterna som stängdes 2002 kunde avvecklingsåtgärderna inför en omedelbar nedmontering genomföras utan avbrott.
I enheterna 3–4 kan avvecklingsåtgärder vidtas endast i begränsad skala, eftersom det fortfarande finns bestrålade bränsleelement i lagringsbassängerna.
För att öka säkerheten vid anläggningen och förhindra att dessa bägge enheter eventuellt åter tas i bruk måste man så fort som möjligt överföra bränsleelementen till extern mellanlagring och nedmonteringen sättas i gång med detsamma.
Detta uppskattade värde kan jämföras exempelvis med kostnaderna för två anläggningar i Greifswald i Tyskland, som vardera hade två reaktorer av samma reaktortyp.
Utgående från de kostnader som angetts för Greifswald kan man härleda sig till en kostnad på 1 780 miljoner EUR för fyra reaktorer, med hänsyn tagen till att villkoren delvis är annorlunda
Förbundsrepubliken Tysklands strålskyddsverk: Undersökning av sparpotentialen i samband med avveckling och nedmontering av tyska kärnanläggningar, projekt O2 S 7778, på uppdrag från förbundsrepublikens ministerium för utbildning och forskning. .
Republiken Bulgariens regering hade ursprungligen yrkat på 202 miljoner EUR för nästa fas inom avvecklingen av de fyra reaktorerna.
Kommissionen har för perioden 2010–2013 föreslagit 180 miljoner EUR i stöd till avvecklingen.
Det internationella samfundet (i allt väsentligt EU) ställde fram till 2006 340 miljoner EUR till förfogande (Phare), under 2007 och 2008 253 miljoner EUR (EBRD) och för 2009 89,5 miljoner EUR.
Fram till 2013 kommer sammanlagt ca 860 miljoner EUR att ha getts som stöd till avvecklingen.
Också fast man i dagens läge inte exakt känner till hur stort stödet var fram till 2006 samt under 2009 måste man utgå från att kostnaderna fram till 2013 för avvecklingen samt för hanteringen av det radioaktiva avfallet och den hittills planerade mellanlagringen av bestrålade bränsleelement i stort sett är täckta.
Med beaktande av att Bulgarien självt ska stå för en del av kostnaderna får det bidrag på 180 miljoner EUR som kommissionen föreslagit för den fortsatta avvecklingen anses som lämpligt.
Det ovannämnda finansieringsbehovet på 1 800 miljoner EUR innefattar inga kostnader för och det av kommissionen föreslagna ekonomiska stödet på 300 miljoner EUR inget projekt för slutförvaring av bränsleelementen.
Bulgariens aktuella strategi för upparbetning utanför Europeiska unionen kan, såsom det påtalats i det föregående, inte accepteras, vare sig av omsorg om kärnsäkerheten eller säkerhetsskyddet.
I den tredje rapporten i anslutning till den gemensamma konventionen angavs som grunder till beslutet om upparbetning i stället för direkt slutförvaring dels att det inte fanns tillräckliga ekonomiska resurser att tillgå och dels att man ville undvika att utsätta kommande generationer för en oskälig belastning.
Argumentet om en belastning av kommande generationer håller inte streck.
Vid upparbetningen förintas ju inga av de ämnen som uppkommer vid användningen av kärnkraft: alltså finns de också kvar för kommande generationer.
För att upparbetningen ska kunna frångås så fort som möjligt bör de ekonomiska resurser som saknas ställas till förfogande av EU.
Enligt uppgifter från kommissionen
Den budget på 120 miljoner EUR som ställts till förfogande för hanteringen av bestrålade bränsleelement fram till 2013 bör användas till åtgärder för att den sammanlagda mellanlagringskapaciteten snabbare ska kunna ställas till förfogande samt för att arbetet med att välja slutförvaringsplats snabbt slutföras, liksom också till åtgärder för undersökning av geologisk lämplighet.
I kommissionens förslag till förordning om ekonomiskt stöd inom ramen för Kozloduj‑projektet ingår också stöd till energiprojekt.
Detta tillbakavisas av föredraganden.
Republiken Bulgarien har fram till 2009 redan fått över 259 miljoner EUR från Europeiska banken för återuppbyggnad och utveckling som stöd till energiprojekt.
Enligt kommissionen har det i huvudsak varit frågan om förbättring av energieffektiviteten och användning av förnybar energi.
KOM(2009)0581 .
På det sättet kunde Bulgarien producera el med mindre utsläpp av koldioxid och överlag på ett miljövänligare sätt.
Bulgarien har dock för sin del beslutat att öka elproduktionskapaciteten genom att använda kärnkraft.
Om man samtidigt frångår kol som bränsle skulle detta i begränsad omfattning kunna minska koldioxidutsläppen, men det innebär dock en ökad belastning på människor och miljö till följd av radioaktiviteten och ökade risker för säkerheten till följd av eventuella incidenter.
Nu är det dock så, att varje euro som investeras i energieffektivitet avsevärt snabbare minskar koldioxidutsläppen avsevärt mera än varje euro som investeras i kärnkraft och därför blir följden i själva verket större utsläpp om man har kvar kärnkraften än om man följer andra strategier.
Nu har det redan gått åtta år sedan enheterna 1–2 stängdes och enheterna 3–4 stängdes för mer än tre år sedan, alltså bara fem år före den tidpunkt som ursprungligen inplanerats.
Man hade alltså tillräckligt med tid på sig för att hinna planera och förverkliga en ersättande kapacitet och tack vare stödet från Europeiska banken för återuppbyggnad och utveckling fanns det också möjligheter till detta.
Ytterligare stöd skulle snedvrida konkurrensen till skada för andra stater eller producenter.
Sådant är inte tillåtet enligt gemenskapslagstiftningen.
Efter 2007 (det år då enheterna 1–4 i kärnkraftverket Kozloduj stängdes) hade Bulgarien inga problem med sin elförsörjning.
ENTSOE 2009.
Alltså behövs det ingen ersättande produktionskapacitet för att landet i fortsättningen ska klara elförsörjningen.
Om begreppet ”region” i kommissionens förslag också avser områden utanför Bulgarien, då skulle det först och främst behövas undersökningar av elförsörjningen i dessa stater.
Eftersom grannländerna, med undantag för Rumänien och Grekland, inte är medlemmar av EU, skulle man dessutom få lov att se efter i vad mån det vore tillåtet att stödja deras elförsörjning med medel från EU.
De driftsansvariga för kraftverken i Bulgarien får dessutom intäkter genom exporten.
Denna export får inte finansieras med EU-medel.
Med hänsyn tagen till att 120 miljoner EUR ställts till förfogande för den fortsatta hanteringen av bestrålade bränsleelement förefaller kommissionens förslag i fråga om avvecklingen att vara ändamålsenligt.
Fortsatt stöd ur EU:s budget motsvarar EU:s intresse av säkerhet vid användningen av kärnkraft.
Det är på sin plats att stödmedlen tilldelas via Europeiska banken för återuppbyggnad och utveckling.
Om det inte gavs något stöd skulle man inte kunna utesluta att enheterna Kozloduj 3–4 togs i bruk på nytt, vilket skulle innebära avsevärda risker för incidenter.
Svåra incidenter skulle få konsekvenser inte bara för Bulgarien.
Bulgarien har hittills inte avsatt tillräckligt med resurser för avvecklingen.
Utan EU-medel finns det troligen inga garantier för att avvecklingsåtgärderna till skydd för människor och miljö fortsätts i den utsträckning som behövs.
Eftersom anslagen i dagens läge är så pass små bidrar EU-medlen till att det i samband med avvecklingsåtgärderna uppnås en hög nivå av säkerhet till skydd för människor och miljö.
EU-medlen får inte användas till något annat än till avvecklingen av enheterna Kozloduj 1–4 och då till de projekt som fastställts och till att bränsleelementen snabbt ska kunna föras över till torr mellanlagring och till slutförvaring.
De ändringar och kompletteringar som föreslagits i skälen och artiklarna preciserar hur medlen bör användas och anknyter användningen till EU:s prioriterade mål, nämligen till att rigorösa normer för säkerhet ska iakttas vid avvecklingen samt att den liberaliserade energimarknaden ska förverkligas genom att konkurrenssnedvridningar på längre sikt undviks.
Artikel 6 i förordningen bör möjliggöra en effektiv kontroll av vad EU-medlen används till och likaså att de tas i bruk vid lämpliga tidpunkter.
Med tanke på detta är det till nytta om man hela tiden känner till den aktuella situationen inom tillståndsförfarandet.
YTTRANDE från budgetutskottet
till utskottet för industrifrågor, forskning och energi
över förslaget till rådets förordning om gemenskapens ekonomiska stöd till avvecklingen av enheterna 1–4 i kärnkraftverket Kozloduj i Bulgarien - ”Kozloduj-programmet”
( KOM(2009)0581 – C7‑0289/2009 – 2009/0172(NLE) )
Föredragande:
Helga Trüpel
KORTFATTAD MOTIVERING
Litauen, Slovakien och Bulgarien får ekonomiskt stöd från gemenskapen för sina insatser för att uppfylla åtagandet att stänga första generationens kärnreaktorer.
Stödet till Bulgarien har reglerats genom anslutningsfördraget och skulle vara avslutat i slutet av 2009, medan stödet till Litauen och Slovakien kommer att fortsätta till 2013.
I slutet av förhandlingarna om den fleråriga budgetramen var Bulgarien ännu inte medlemsstat och landet fattade dessutom beslutet om avveckling rätt sent.
Därför infördes inga anslag i den fleråriga budgetramen 2007–2013 för finansiering efter 2009.
Det ekonomiska stöd som tillhandahölls före 2009 för avvecklingen var främst avsett för förberedelser.
Förslaget om förlängning syftar till att förlänga stödet till Bulgarien för att följa upp och garantera säkert underhåll och avveckling av kärnkraftverket Kozloduj enligt den plan som fastställts.
Förslaget innehåller även lindrande åtgärder för energisektorn.
Det anslag som begärs av gemenskapen kommer att vara sammanlagt 300 miljoner euro för perioden 2010–2013.
Stödet kommer att göras tillgängligt som ett gemenskapsbidrag till den internationella stödfond för avvecklingen av Kozloduj som förvaltas av EBRD.
Kommissionen lade fram sitt förslag för fortsatt stöd till avvecklingen av Kozloduj i oktober 2009, mitt i budgetförfarandet för 2010.
Budgetförslaget för 2010 ingick i ändringsskrivelse 2.
Förslaget kom mycket sent och innebar en stor utmaning för budgetmyndigheten eftersom budgetbehoven för avvecklingen av Kozloduj skulle omfattas av rubrik 1a, precis som återhämtningsplanen för Europa som krävde en finansiering på nästan 2 miljarder euro 2010.
Med hänsyn till de politiska åtaganden som ingicks i samband med anslutningsförhandlingarna, samt det odiskutabla behovet av att garantera en säker avveckling av föråldrad kärnteknik, måste finansieringen av Kozloduj tryggas.
I slutändan tillhandahölls de budgetmedel som behövdes 2010, 75 miljoner euro, genom utnyttjande av flexibilitetsmekanismen.
Finansieringen på 225 miljoner euro för perioden 2011–2013 bör i princip hämtas från rubrik 1a.
Kommissionen har tagit med de nödvändiga beloppen i budgetplaneringen för denna period.
Tillsammans med de övriga förändringar som väntas minskar marginalen i rubrik 1a hastigt och närmar sig 34 miljoner euro 2012.
Marginalen skulle bli något större 2011 och 2013.
I den finansieringsöversikt som bifogas förslaget erkänner kommissionen att förslaget kan komma att kräva att bestämmelserna i det interinstitutionella avtalet tillämpas.
Enligt punkt 38 i det interinstitutionella avtalet kommer det finansiella referensbelopp som rådet eventuellt vill införa inte att påverka budgetmyndighetens befogenheter eftersom detta program inte omfattas av medbeslutandeförfarandet.
Beloppen kommer därför att fastställas i det årliga budgetförfarandet.
Med tanke på den begränsade marginalen och de eventuella kommande behoven kommer det att vara viktigt att på förhand eller, om ingen flerårig lösning nås, i samband med varje budgetförfarande, avgöra vilken som skulle vara den bästa finansieringskällan för Kozloduj.
När detta förslag till yttrande presenteras har föredraganden inte bestämt sig för vilken hon anser vara den lämpligaste lösningen när det gäller kommissionens förslag och dess förenlighet med budgeten.
Därför lägger hon fram två olika alternativ:
– I alternativ A (som representeras av ändringsförslag 1) anges att förslaget är förenligt med budgeten.
– I alternativ B (som representeras av ändringsförslag 2) anges att förslaget är oförenligt med budgeten.
ÄNDRINGSFÖRSLAG
Budgetutskottet uppmanar utskottet för industrifrågor, forskning och energi att som ansvarigt utskott infoga följande ändringsförslag i sitt betänkande:
Ändringsförslag
1
Förslag till lagstiftningsresolution
Punkt 1a (ny)
Förslag till lagstiftningsresolution
Ändringsförslag
Ändringsförslag
2
Förslag till lagstiftningsresolution
Punkt 1b (ny)
Förslag till lagstiftningsresolution
Ändringsförslag
Ändringsförslag
3
Förslag till lagstiftningsresolution
Punkt 1c (ny)
Förslag till lagstiftningsresolution
Ändringsförslag
Ändringsförslag
4
Kommissionens förslag
Ändringsförslag
1.
Det finansiella referensbelopp som krävs för genomförandet av Kozloduj‑programmet för perioden 1 januari 2010–31 december 2013 fastställs härmed till 300 miljoner euro.
1.
Det finansiella referensbelopp enligt punkt 38 i IIA av den 17 maj 2006 som krävs för genomförandet av Kozloduj‑programmet för perioden 1 januari 2010–31 december 2013 fastställs härmed till 300 miljoner euro.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
8.4.2010
Slutomröstning: resultat
+:
–:
0:
30
1
1
Slutomröstning: närvarande ledamöter
Slutomröstning: närvarande suppleanter
YTTRANDE från utskottet för miljö, folkhälsa och livsmedelssäkerhet
till utskottet för industrifrågor, forskning och energi
över förslaget till rådets förordning om gemenskapens ekonomiska stöd till avvecklingen av enheterna 1–4 i kärnkraftverket Kozloduj i Bulgarien - ”Kozloduj-programmet”
( KOM(2009)0581 – C7‑0289/2009 – 2009/0172(NLE) )
Föredragande:
Antonyia Parvanova
KORTFATTAD MOTIVERING
Bulgarien har fullgjort sina åtaganden och stängt enheterna 1–4 i kärnkraftverket Kozloduj i enlighet med artikel 30 i protokollet till anslutningsfördraget för Bulgarien och Rumänien.
Bulgarien ska nu avveckla dessa fyra enheter.
Den ändrade strategin för nedmontering och avveckling och den nödvändiga finansiering som detta medför samt efterlevnaden och fullgörandet av åtaganden kopplade till kärnkraftverket Kozloduj utgör skäl för en förlängning av gemenskapens ekonomiska stöd, så att högsta möjliga nivå garanteras när det gäller säkerhet och miljö i samband med nedmonteringen och avvecklingen av enheterna 1–4.
Dessutom har andra medlemsstater, t.ex.
Slovakien och Litauen, kunnat dra nytta av ett liknande stödprogram för avveckling av kärnkraftverk som pågår ända fram till 2013, medan stödet till Bulgarien upphör 2009.
Tillämpningen av gemenskapens principer om solidaritet och likabehandling utgör ytterligare ett skäl för att förlänga gemenskapens ekonomiska stöd.
Gemenskapsstödet för avvecklingen av enheterna 1–4 i kärnkraftverket Kozloduj bör riktas mot ett enda mål: att se till att nedmonteringen sker på ett säkert sätt och inom utsatt tid samtidigt som högsta möjliga standard garanteras i fråga om insyn och miljöskydd.
Därför bör man under varje fas i avvecklingen lägga särskild tonvikt vid säkerhets- och miljöskyddsnormer i enlighet med gällande lagstiftning, såsom rådets direktiv 96/29/Euratom om fastställande av grundläggande säkerhetsnormer för skydd av arbetstagarnas och allmänhetens hälsa mot de faror som uppstår till följd av joniserande strålning.
Man bör även rikta särskild uppmärksamhet mot hälsoskyddet för de arbetstagare som deltar i avvecklingen, och uppföljande hälsokontroller bör göras under en längre period.
Insyn är också ytterst viktigt för att se till att allmänheten känner till och kan engagera sig i de beslut som tas om avvecklingen samt i framtida frågeställningar som hör samman med avvecklingen, t.ex. slutförvaringen av radioaktivt avfall.
Det är därför oerhört viktigt med efterlevnad av internationella konventioner där nödvändiga krav redan fastställs på nationell, internationell och gränsöverskridande nivå, såsom Århuskonventionen av den 25 juni 1998, så att tillgång till information, allmänhetens deltagande och insyn garanteras.
När man betraktar bestämmelserna i förslaget till förordning till stöd för åtgärderna inom energisektorn för att dämpa effekterna av den tidigarelagda stängningen av enheterna 1–4 i kärnkraftverket Kozloduj måste man givetvis beakta att energi- och kärnkraftssektorn samt miljön påverkas betydligt mer än väntat.
Till exempel beräknas förlusten av produktionskapacitet till följd av den tidigarelagda stängningen av de fyra enheterna leda till en ännu större ökning av utsläppsvolymen för växthusgaser, 15 TWh för perioden 2011–2013 med koldioxidekvivalenter på cirka 1,2 Gg/GWh, vilket för Bulgariens del kommer att betyda ytterligare påverkan av omkring 18 000 Gg eller 18 000 kt koldioxidekvivalenter.
Koldioxidutsläppen måste därför minskas ännu mer.
De övergripande och långsiktiga konsekvenserna av den tidigarelagda stängningen av de fyra reaktorerna innebar ett åsidosättande av de huvudsakliga principer som ligger till grund för unionens nuvarande energistrategi: hållbarhet och minskning av koldioxidutsläpp, trygg energiförsörjning och en konkurrenskraftig energisektor.
Förlusten av produktionskapaciteten från kärnkraftverket Kozlodujs fyra enheter måste till stor del kompenseras med import av primära energikällor och med importerade och inhemska fossila energikällor.
Av hänsyn till miljön, ekonomin och energiförsörjningstryggheten i regionen är det viktigt att förlänga gemenskapsstödet till den bulgariska energisektorn så att de långsiktiga konsekvenserna av den tidigarelagda stängningen av de fyra reaktorerna kan hanteras.
Konsekvens och enhetlighet med EU:s miljö- och energistrategier måste säkerställas så att genomförandet av gemenskapens ekonomiska stöd leder till en effektiv och optimal avveckling av enheterna 1–4 i kärnkraftverket Kozloduj.
ÄNDRINGSFÖRSLAG
Utskottet för miljö, folkhälsa och livsmedelssäkerhet uppmanar utskottet för industrifrågor, forskning och energi att som ansvarigt utskott infoga följande ändringsförslag i sitt betänkande:
Ändringsförslag
1
Förslag till förordning
Skäl 1
Kommissionens förslag
Ändringsförslag
(1) Bulgarien lovade att stänga enheterna 1 och 2 samt 3 och 4 i kärnkraftverket Kozloduj till den 31 december 2002 respektive den 31 december 2006, och att därefter avveckla dessa enheter.
Europeiska unionen har förklarat sig vara villig att fram till 2009 ge fortsatt ekonomiskt stöd till Bulgariens avvecklingsverksamhet som en förlängning av föranslutningsstödet inom ramen för Phareprogrammet.
(1) Bulgarien lovade att stänga enheterna 1 och 2 samt 3 och 4 i kärnkraftverket Kozloduj till den 31 december 2002 respektive den 31 december 2006, och att därefter avveckla dessa enheter.
Europeiska unionen har förklarat sig vara villig att fram till 2009 ge fortsatt ekonomiskt stöd till Bulgariens avvecklingsverksamhet som en förlängning av föranslutningsstödet inom ramen för Phareprogrammet.
EU har dessutom gett politiska garantier för att ett fortsatt gemenskapsstöd ska övervägas vid den allmänna översynen av budgetplanen 2007–2013.
Ändringsförslag
2
Förslag till förordning
Skäl 2a (nytt)
Kommissionens förslag
Ändringsförslag
(2a) Gemenskapens principer om solidaritet och likabehandling kräver ett rättvist tillvägagångssätt, nu som förr, gentemot medlemsstater i behov av ekonomiskt stöd för att avveckla kärnkraftverk, enligt åtaganden i deras anslutningsfördrag eller tilläggsprotokoll om att stänga enheter vid kärnkraftsverk.
Ändringsförslag
3
Förslag till förordning
Skäl 5
Kommissionens förslag
Ändringsförslag
(5) Det är också viktigt att använda kärnkraftverket Kozlodujs egna resurser, eftersom man därigenom bibehåller den nödvändiga expertisen och samtidigt lindrar de sociala och ekonomiska följderna av den tidigarelagda stängningen genom att sysselsätta personal från det stängda kärnkraftverket.
Fortsatt ekonomiskt stöd är därför en förutsättning för att den nödvändiga s äkerhetsstandarden ska kunna upprätthållas.
(5) Det är också viktigt att använda kärnkraftverket Kozlodujs egna resurser, eftersom man därigenom bibehåller den nödvändiga expertisen , förbättrar kunskapen och kompetensen och samtidigt lindrar de sociala och ekonomiska följderna av den tidigarelagda stängningen genom att sysselsätta personal från det stängda kärnkraftverket.
Fortsatt ekonomiskt stöd är därför en förutsättning för att nödvändiga säkerhets-, folkhälso- och miljökrav ska kunna upprätthållas.
Ändringsförslag
4
Förslag till förordning
Skäl 6
Kommissionens förslag
Ändringsförslag
(6) Europeiska unionen noterar också behovet av ekonomiskt stöd för att fortsätta lindringsåtgärderna inom energisektorn med tanke på den omfattande kapacitetsförlusten till följd av kärnkraftsenheternas stängning, och de följder för regionens försörjningstrygghet som detta medför.
(6) Europeiska unionen noterar också behovet av ekonomiskt stöd för att fortsätta lindringsåtgärderna inom energisektorn med tanke på den omfattande kapacitetsförlusten till följd av kärnkraftsenheternas stängning, och de följder för miljön, konsumentpriserna på energi samt regionens försörjningstrygghet som detta medför , och för utsläppsvolymen av växthusgaser, eftersom bortfallet av produktionskapaciteten hos enheterna 1–4 i kärnkraftverket Kozloduj till stor del måste kompenseras med import av primära energikällor och med importerade och inhemska fossila energikällor, varvid behovet att öka energieffektiviteten och utveckla sektorn för förnybar energ i särskilt ska uppmärksammas .
Ändringsförslag
5
Förslag till förordning
Skäl 6a (nytt)
Kommissionens förslag
Ändringsförslag
Ändringsförslag
6
Förslag till förordning
Skäl 6b (nytt)
Kommissionens förslag
Ändringsförslag
(6b) Ekonomiskt stöd från EU kan behövas till åtgärder som lindrar de sociala och ekonomiska följderna av stängningen av kärnkraftverket Kozlodujs enheter 1–4, såsom omskolningsprogram för att berörd personal ska kunna använda sin kompetens i andra sektorer, till exempel inom industriell forskning eller förnybar energi.
Ändringsförslag
7
Förslag till förordning
Skäl 7
Kommissionens förslag
Ändringsförslag
(7) Under perioden 2010–2013 bör därför ett belopp på 300 miljoner euro avsättas i Europeiska unionens allmänna budget för finansieringen av nedläggningen av kärnkraftverket Kozloduj.
(7) Under perioden 2010–2013 bör därför ett belopp på 300 miljoner euro avsättas i Europeiska unionens allmänna budget för finansieringen av nedläggningen av kärnkraftverket Kozloduj och för lindringsåtgärderna inom energisektorn .
Ändringsförslag
8
Förslag till förordning
Skäl 8
Kommissionens förslag
Ändringsförslag
(8) Gemenskapens budgetanslag för avveckling bör inte leda till snedvridning av konkurrensen för energiförsörjningsföretag på energimarknaden i unionen.
Dessa anslag bör även användas för att finansiera åtgärder för att kompensera den minskade produktionskapaciteten i linje med det relevanta regelverket.
(8) Gemenskapens budgetanslag för avveckling bör inte leda till snedvridning av konkurrensen för energiförsörjningsföretag på energimarknaden i unionen.
Dessa anslag bör även användas för att finansiera åtgärder för att kompensera den minskade produktionskapaciteten i linje med det relevanta regelverket , uppmuntra til l energisparande och främja förnybar energi .
Ändringsförslag
9
Förslag till förordning
Skäl 11
Kommissionens förslag
Ändringsförslag
(11) För att största möjliga effektivitet ska garanteras bör bästa tillgängliga tekniska expertis användas vid avvecklingen av kärnkraftverket Kozloduj, med hänsyn tagen till vilken typ av reaktorer som ska stängas och de tekniska specifikationer som gäller för dem.
(11) För att största möjliga effektivitet ska garanteras och för att minska eventuella miljökonsekvenser bör bästa tillgängliga tekniska expertis användas vid avvecklingen av kärnkraftverket Kozloduj, med hänsyn tagen till vilken typ av reaktorer som ska stängas och de tekniska specifikationer som gäller för dem.
Ändringsförslag
10
Förslag till förordning
Skäl 11a (nytt)
Kommissionens förslag
Ändringsförslag
Ändringsförslag
11
Förslag till förordning
Skäl 12a (nytt)
Kommissionens förslag
Ändringsförslag
__________
1 EGT L 159, 29.6.1996, s.
1.
Ändringsförslag
12
Förslag till förordning
Skäl 13a (nytt)
Kommissionens förslag
Ändringsförslag
(13a) De villkor som gäller metoden för gemensam förvaltning vid genomförandet av budgeten fastställs i artiklarna 53d, 108a och 165 i rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget 1 , och i artiklarna 35 och 43 i kommissionens förordning (EG, Euratom) nr 2342/2002 av den 23 december 2002 om genomförandebestämmelser för rådets förordning (EG, Euratom) nr 1605/2002 med budgetförordning för Europeiska gemenskapernas allmänna budget 2 .
__________
1 EGT L 248, 16.9.2002, s.
1.
2 EGT L 357, 31.12.2002, s.
1.
Motivering
Enligt budgetförordningen och genomförandebestämmelserna har kommissionen rätt att genomföra sin budget genom gemensam förvaltning med internationella organisationer om dessa organisationer tillämpar standarder som ger garantier som motsvarar internationellt godkända standarder för, som ett minimum, reglerna för räkenskaper, revision, intern kontroll och upphandling.
Ändringsförslag
13
Förslag till förordning
Skäl 13b (nytt)
Kommissionens förslag
Ändringsförslag
(13b) Fallet med Kozloduj bör tjäna som exempel och kommissionen bör utarbeta en fullständig och exakt avvecklingsbudget för att en analys och beräkning av kostnaderna för framtida avveckling av kärnkraftverk ska kunna göras.
Ändringsförslag
14
Förslag till förordning
Artikel 1
Kommissionens förslag
Ändringsförslag
I denna förordning fastställs ett program med detaljerade genomförandebestämmelser för gemenskapens ekonomiska bidrag till avvecklingen av enheterna 1–4 i kärnkraftverket Kozloduj, och följderna för Bulgarien av stängningen av dessa enheter (nedan kallat Kozloduj‑programmet).
I denna förordning fastställs ett program med detaljerade genomförandebestämmelser för gemenskapens ekonomiska bidrag till avvecklingen av enheterna 1–4 i kärnkraftverket Kozloduj, och följderna för miljön, ekonomin och energiförsörjningstryggheten i regionen av att dessa enheter i Bulgarien stängs (nedan kallat Kozloduj-programmet).
Ändringsförslag
15
Förslag till förordning
Artikel 2
Kommissionens förslag
Ändringsförslag
Syftet med gemenskapens stöd till Kozloduj-programmet i enlighet med denna förordning är att ekonomiskt stödja åtgärder inom ramen för avvecklingen av kärnkraftverket Kozloduj, åtgärder för miljöuppgradering i linje med regelverket och för modernisering av den konventionella produktionskapaciteten för att ersätta produktionskapaciteten för de fyra reaktorerna vid kärnkraftverket Kozloduj samt andra åtgärder som följer av beslutet att stänga och avveckla detta kärnkraftverk och som bidrar till den nödvändiga omstruktureringen, miljöuppgraderingen och moderniseringen av energiproduktionen och överförings- och distributionssektorerna i Bulgarien samt till att förbättra energiförsörjningstryggheten och energieffektiviteten i Bulgarien.
Syftet med gemenskapens stöd till Kozloduj-programmet i enlighet med denna förordning är att ekonomiskt stödja åtgärder inom ramen för avvecklingen av kärnkraftverket Kozloduj, åtgärder för miljöuppgradering i linje med regelverket och för modernisering av den konventionella produktionskapaciteten för att ersätta produktionskapaciteten för de fyra reaktorerna vid kärnkraftverket Kozloduj samt andra åtgärder som följer av beslutet att stänga och avveckla detta kärnkraftverk och som bidrar till den nödvändiga omstruktureringen, miljöuppgraderingen och moderniseringen av energiproduktionen och överförings- och distributionssektorerna i Bulgarien samt till att förbättra energiförsörjningstryggheten och energieffektiviteten i Bulgarien , samtidigt som energibesparande åtgärder måste uppmuntras och förnybar energi främjas .
Ekonomiskt stöd kan också ges för att lindra den socioekonomiska övergången i de berörda kommunerna, till exempel genom utvecklande av nya hållbara arbetstillfällen och industrier.
Ändringsförslag
16
Kommissionens förslag
Ändringsförslag
3.
Anslagen för Kozloduj-programmet kan ses över under perioden 1 januari 2010– 31 december 2013 för att man ska kunna ta hänsyn till gjorda framsteg under programmets genomförande och för att man ska kunna se till att programplaneringen och fördelningen av resurserna grundas på faktiska betalningsbehov och faktisk absorberingskapacitet.
3.
Anslagen för Kozloduj-programmet ska ses över årligen under perioden 1 januari 2010–31 december 2013 för att man ska kunna ta hänsyn till gjorda framsteg under programmets genomförande och till de långsiktiga effekterna på och konsekvenserna för miljön, ekonomin och försörjningstryggheten till följd av den tidigarelagda stängningen av kärnkraftverket Kozlodujs enheter 1–4, och för att man ska kunna se till att programplaneringen och fördelningen av resurserna grundas på faktiska betalningsbehov och faktisk absorberingskapacitet.
Ändringsförslag
17
Kommissionens förslag
Ändringsförslag
1.
Kommissionen får, direkt genom sina anställda eller genom någon annan behörig organisation den valt, utföra en granskning av hur bidraget har använts.
Granskningen får utföras under hela löptiden för avtalet mellan gemenskapen och EBRD om att tillhandahålla gemenskapsmedel till internationella fonden för avvecklingsstöd till Kozloduj samt under fem år efter dagen för utbetalning av den sista bidragsdelen.
I förekommande fall kan revisionens resultat leda till att kommissionen beslutar om återkrav.
1.
Kommissionen ska övervaka och får, direkt genom sina anställda eller genom någon annan behörig organisation den valt, utföra en granskning av hur bidraget har använts.
Granskningen får utföras under hela löptiden för avtalet mellan gemenskapen och EBRD om att tillhandahålla gemenskapsmedel till internationella fonden för avvecklingsstöd till Kozloduj samt under fem år efter dagen för utbetalning av den sista bidragsdelen.
I förekommande fall kan granskningens resultat leda till att kommissionen beslutar om återkrav.
Ändringsförslag
18
Kommissionens förslag
Ändringsförslag
2.
Kommissionens personal och extern personal med fullmakt från kommissionen ska ges lämplig tillgång till mottagarens kontorslokaler och till alla upplysningar, även i elektronisk form, som behövs för att utföra granskningen.
2.
Kommissionens personal och extern personal med fullmakt från kommissionen ska ges lämplig tillgång till mottagarens kontorslokaler och till alla upplysningar, även i elektronisk form, som behövs för att utföra granskningen.
I granskningen ska också ingå en undersökning om hur långt man kommit i tillståndsgivningen för avveckling.
Motivering
Syftet är att garantera att resurserna används när de ska och att mer noggrant se till att de används för det de är avsedda.
Ändringsförslag
19
Förslag till förordning
Artikel 7
Kommissionens förslag
Ändringsförslag
Kommissionen ska se till att denna förordning tillämpas och årligen rapportera till Europaparlamentet och rådet.
Efterhandsutvärderingen ska innehålla en fullständig och exakt kostnadsbudget för avvecklingen av ett kärnkraftverk så att man kan planera för framtida avvecklingsprojekt.
Den ska också analysera ekonomiska, sociala och miljömässiga kostnader, med fokus på frigjord reststrålning och konsekvenser för försörjningstryggheten.
Ändringsförslag
20
Förslag till förordning
Artikel 7a (ny)
Kommissionens förslag
Ändringsförslag
Artikel 7a
Kommissionen ska göra en bedömning av överensstämmelsen med internationellt godkända standarder , åtminstone i fråga om reglerna för räkenskaper, revision, intern kontroll och upphandling vid Europeiska banken för återuppbyggnad och utveckling, innan de sammanlagda överenskomna bidragen undertecknas.
Motivering
Enligt budgetförordningen och genomförandebestämmelserna har kommissionen rätt att genomföra sin budget genom gemensam förvaltning med internationella organisationer om dessa organisationer tillämpar standarder som ger garantier som motsvarar internationellt godkända standarder för, som ett minimum, reglerna för räkenskaper, revision, intern kontroll och upphandling.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
7.4.2010
Slutomröstning: resultat
+:
–:
0:
47
7
1
Slutomröstning: närvarande ledamöter
János Áder, Elena Oana Antonescu, Kriton Arsenis, Pilar Ayuso, Paolo Bartolozzi, Sergio Berlato, Milan Cabrnoch, Martin Callanan, Nessa Childers, Chris Davies, Esther de Lange, Anne Delvaux, Bas Eickhout, Edite Estrela, Jill Evans, Elisabetta Gardini, Julie Girling, Françoise Grossetête, Cristina Gutiérrez-Cortines, Satu Hassi, Jolanta Emilia Hibner, Dan Jørgensen, Christa Klaß, Holger Krahmer, Jo Leinen, Peter Liese, Kartika Tamara Liotard, Linda McAvan, Radvilė Morkūnaitė-Mikulėnienė, Miroslav Ouzký, Vladko Todorov Panayotov, Gilles Pargneaux, Antonyia Parvanova, Andres Perello Rodriguez, Mario Pirillo, Pavel Poc, Frédérique Ries, Anna Rosbach, Oreste Rossi, Horst Schnellhardt, Richard Seeber, Theodoros Skylakakis, Bogusław Sonik, Catherine Soullie, Salvatore Tatarella, Anja Weisgerber, Glenis Willmott, Sabine Wils
Slutomröstning: närvarande suppleanter
Bill Newton Dunn, Justas Vincas Paleckis, Alojz Peterle, Bart Staes, Michail Tremopoulos, Thomas Ulmer, Marita Ulvskog
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
28.4.2010
Slutomröstning: resultat
+:
–:
0:
47
4
1
Slutomröstning: närvarande ledamöter
Jean-Pierre Audy, Zigmantas Balčytis, Bendt Bendtsen, Jan Březina, Reinhard Bütikofer, Maria Da Graça Carvalho, Giles Chichester, Christian Ehler, Lena Ek, Ioan Enciu, Gaston Franco, Adam Gierek, Norbert Glante, Fiona Hall, Jacky Hénin, Sajjad Karim, Arturs Krišjānis Kariņš, Philippe Lamberts, Bogdan Kazimierz Marcinkiewicz, Angelika Niebler, Jaroslav Paška, Aldo Patriciello, Anni Podimata, Miloslav Ransdorf, Herbert Reul, Teresa Riera Madurell, Jens Rohde, Paul Rübig, Amalia Sartori, Francisco Sosa Wagner, Konrad Szymański, Britta Thomsen, Patrizia Toia, Niki Tzavela, Marita Ulvskog, Vladimir Urutchev, Adina-Ioana Vălean, Alejo Vidal-Quadras
Slutomröstning: närvarande suppleanter
Matthias Groote, Cristina Gutiérrez-Cortines, Rebecca Harms, Oriol Junqueras Vies, Ivailo Kalfin, Ivari Padar, Vladko Todorov Panayotov, Markus Pieper, Mario Pirillo, Vladimír Remek, Frédérique Ries, Theodoros Skylakakis, Silvia-Adriana Ţicău, Hermann Winkler
A7-0154/2010
om sakernas Internet
(2009/2224(INI))
Utskottet för industrifrågor, forskning och energi
Föredragande:
Maria Badia i Cutchet
PE 438.414v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING..........................................................................................................................14
YTTRANDE från utskottet för internationell handel ...............................16
YTTRANDE från utskottet för den inre marknaden och konsumentskydd 20
YTTRANDE från utskottet för rättsliga frågor ...........................................24
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................28
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om sakernas Internet
( 2009/2224(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens meddelande till Europaparlamentet, rådet, Europeiska ekonomiska och sociala kommittén och Regionkommittén av den 18 juni 2009 ”Sakernas Internet – En handlingsplan för Europa” ( KOM(2009)0278 ),
– med beaktande av det arbetsprogram som det spanska EU-ordförandeskapet lade fram den 27 november 2009, särskilt målsättningen att utveckla framtidens Internet,
– med beaktande av kommissionens meddelande av den 28 januari 2009 ”Investera nu i morgondagens Europa” ( KOM(2009)0036 ),
– med beaktande av kommissionens rekommendation om genomförandet av principerna om integritets- och dataskydd i tillämpningar som stöds av radiofrekvensidentifiering (RFID) (K(2009)3200),
– med beaktande av Europaparlamentets och rådets direktiv 95/46/EG av den 24 oktober 1995 om skydd för enskilda personer med avseende på behandling av personuppgifter och om det fria flödet av sådana uppgifter,
– med beaktande av Europaparlamentets och rådets direktiv 2002/58/EG av den 12 juli 2002 om behandling av personuppgifter och integritetsskydd inom sektorn för elektronisk kommunikation,
– med beaktande av den ekonomiska återhämtningsplanen för Europa ( KOM(2008)0800 ),
– med beaktande av betänkandet från utskottet för industrifrågor, forskning och energi om fastställandet av en ny digital agenda för Europa: 2015.eu
2009/2225(INI) , betänkande av Del Castillo, A7-0066/2010 . ,
– med beaktande av artikel 48 i arbetsordningen,
– med beaktande av betänkandet från utskottet för industrifrågor, forskning och energi och yttrandena från utskottet för internationell handel, utskottet för den inre marknaden och konsumentskydd och utskottet för rättsliga frågor ( A7‑0154/2010 ), och av följande skäl:
A. Internet har utvecklats snabbt under de senaste 25 åren, och denna utveckling väntas fortsätta, vilket kommer att medföra att Internet sprids ytterligare – genom utbyggnaden av bredbandsnätet – och att nya tillämpningar skapas.
B. Sakernas Internet kan leva upp till samhällets och medborgarnas förväntningar, men det krävs forskning för att klargöra hur dessa förväntningar ser ut och för att ringa in de områden där hänsynen till och oron över skyddet av den personliga integriteten och personuppgifterna kan leda till att tillämpningar blockeras.
C. Informations- och kommunikationstekniken (IKT) är viktig för att främja social utveckling och ekonomisk tillväxt och stimulera forskning, innovation och kreativitet inom offentliga och privata organ i EU.
D. Unionen bör ta fram en gemensam referensram för att kunna utforma och skärpa reglerna när det gäller förvaltningen av systemet, sekretessen, informationssäkerheten, hanteringen av etikfrågor, skyddet av privatlivet, insamlingen och lagringen av personuppgifter samt konsumentupplysningen.
E. Med begreppet sakernas Internet avses den övergripande tanken om föremål (både elektroniska föremål och vardagsföremål) som kan läsas, uppfattas, sändas, nås och/eller styras på distans via Internet.
G. Framtidens Internet kommer att överskrida de nuvarande traditionella gränserna för den virtuella världen genom att vara kopplat till de fysiska föremålens värld.
I. RFID-tekniken kan betraktas som en katalysator och en accelerator för den ekonomiska utvecklingen inom informations- och kommunikationssektorn.
K. Som i alla e-hälsovårdssystem krävs det att hälso- och sjukvårdspersonal, patienter och relevanta nämnder (t.ex. uppgiftsskydds- och etiknämnder) deltar aktivt i arbetet med att utforma, utveckla och genomföra system med RFID-teknik.
L. RFID kan bidra till att öka energieffektiviteten, minska utsläppen av växthusgaser och möjliggöra koldioxidredovisning på produktnivå.
M. RFID-tekniken och annan teknik i samband med sakernas Internet kan ge medborgarna fördelar i form av ökad livskvalitet, trygghet, säkerhet och välfärd, förutsatt att man på rätt sätt hanterar frågorna om skyddet av privatlivet och personuppgifterna.
N. Det behövs hållbara, energieffektiva kommunikationsstandarder som är inriktade på säkerhet och integritet och använder kompatibla eller identiska protokoll på olika frekvenser.
Q. Arbetet med att skapa miniatyrprodukter för sakernas Internet innebär tekniska utmaningar, t.ex. när det gäller att integrera elektronik, sensorer och system för inmatning och överföring av RFID-uppgifter i ett chip som inte är större än några millimeter.
T. Det är viktigt att göra EU-medborgarna mer medvetna om ny teknik och därtill hörande tillämpningar, bl.a. om konsekvenserna för samhället och miljön, och att främja konsumenternas digitala kompetens och e-kompetens.
U. Utvecklingen av sakernas Internet bör vara öppen och tillgänglig för alla EU-medborgare samt stödjas genom effektiv politik som syftar till att överbrygga den digitala klyftan i EU och att ge fler medborgare e-kompetens och kunskap om sin digitala omgivning.
Det kan hända att den nuvarande digitala klyftan vidgas, eller så kan en ny digital klyfta skapas.
Europaparlamentet anser att de kommande årens utveckling av sakernas Internet och därtill hörande tillämpningar kommer att få avgörande konsekvenser för EU‑medborgarnas vardag och vanor, vilket kommer att medföra en lång rad ekonomiska och sociala förändringar.
Kommissionen bör därför genomföra fler och mer utförliga undersökningar av denna teknik.
· miljökonsekvenserna och återvinningen av chippen,
· användarnas personliga integritet och förtroende,
· de ökade it-säkerhetsriskerna,
· förekomsten av smarta chip i vissa produkter,
· rätten till ”chippens tystnad”, som innebär delaktighet och kontrollmöjligheter för användarna,
· medborgarnas garantier när det gäller skydd vid insamling och bearbetning av personuppgifter,
· behovet av att utveckla ytterligare en nätstruktur och infrastruktur för tillämpningar av och maskinvara för sakernas Internet,
· garantierna för bästa möjliga skydd mot alla slags it-angrepp för medborgarna och företagen i EU,
· de elektromagnetiska fältens inverkan på djur, särskilt på fåglar i städerna,
· harmoniseringen av regionala standarder,
· utvecklingen av öppna tekniska standarder och driftskompabilitet mellan olika system.
Parlamentet noterar i detta sammanhang yttrandet från Europeiska datatillsynsmannen.
Europaparlamentet uppmanar operatörerna av RFID-tillämpningar att vidta alla rimliga åtgärder för att se till att uppgifterna i fråga inte kan knytas till en identifierad eller identifierbar fysisk person genom något medel som sannolikt kan användas av antingen operatören av RFID-tillämpningar eller någon annan person, såvida dessa uppgifter inte behandlas i enlighet med de tillämpliga principerna och rättsliga dataskyddsbestämmelserna.
• De sätt som finns att möjliggöra identifiering och spårbarhet ska nämnas uttryckligen.
• Säkerhetsåtgärder ska vidtas som garanti för att endast behöriga användare får tillgång till data.
• Konsumenterna och de myndigheter som ansvarar för tilldelningen ska få möjlighet att kontrollera uppgifternas läsbarhet och systemets funktioner.
Parlamentet påminner i detta sammanhang om att Europeiska byrån för nät- och informationssäkerhet (ENISA) spelar en avgörande roll för nätsäkerheten och informationssäkerheten och följaktligen för säkerheten i samband med sakernas Internet, vilket kommer att bidra till att skapa en högre grad av acceptans och förtroende från konsumenternas sida.
Europaparlamentet understryker att forskningen kommer att spela en central roll för att skapa konkurrens mellan leverantörerna om att kunna erbjuda den datorkraft som krävs för att tillämpningar av sakernas Internet ska fungera i realtid.
Det är dessutom mycket viktigt att analysera aspekter som gäller säkerhetssystem för trådlösa nätverk.
MOTIVERING
Det har gått mer än 40 år sedan de första Internetapplikationerna, vilket uppfinnaren av World Wide Web, Tim Berners-Lee, påminde om vid sitt besök nyligen i Europaparlamentet
Den åttonde årliga STOA-föreläsningen, 1 december 2009. .
Under årens lopp har Internet genomgått en ständig och oavbruten utveckling, särskilt under de senaste 25 åren.
I dag förbinder nätet ca 1,5 miljard människor, och dess öppna struktur, som bygger på en standardiserad teknik, har lett till en världsvid spridning och driftskompatibilitet.
Sakernas Internet, ett projekt som inleddes 1999 i USA, blir allt populärare och kommer under de följande tio-femton åren att revolutionera interagerandet mellan människor och föremål och mellan själva föremålen tack vare den ökande användningen av RFID-tekniken (radiofrekvensidentifikation).
Den beståndsdel som karaktäriserar RFID-tekniken är transpondern (eller etiketten), det vill säga en elektronisk komponent som utgörs av ett chip och en antenn.
Chippet, som är några millimeter stort per sida, kan trådlöst innehålla, ta emot och överföra information om karaktären och sammansättningen av den produkt som den är placerad på.
Experter på området menar att chippet i framtiden kommer att ersätta de streckkoder som är i bruk i dag.
Fördelen med RFID-tekniken jämfört med dagens teknik är att chippet inte behöver vara i kontakt med avläsaren för att bli avläst, såsom fallet är med magnetband, och det behöver inte vara synligt, vilket gäller för streckkoder.
Dessutom ska man beakta de särskilda uppgifter och den mängd uppgifter som chippen kan innehålla om de föremål som de är förbundna med, och som denna teknik ger möjlighet till.
Nuvarande tillämpningar av sakernas Internet och framtida utveckling
Det finns redan konkreta exempel inom en rad sektorer:
· Inom bilbranschen kan chip skicka information i realtid till föraren om däcktryck.
· Inom livsmedelsbranschen gör RFID-tekniken det möjligt att garantera en hög standard när det gäller varornas hygiensäkerhet samt deras kemiska, fysiska och organoleptiska egenskaper.
Med hjälp av chippen kan varan dessutom oftare och snabbare spåras.
Många andra tillämpningar har redan utvecklats och tagits i bruk inom logistik- och transportsektorn med mycket positiva resultat.
Några länder (Storbritannien och USA) har infört ett chip i sina nationella pass.
I framtiden kommer RFID-tekniken tillsammans med en IP-adress att göra det möjligt att skapa ett enormt trådlöst sakernas Internet.
Det exempel som oftast anges är kylskåp som, om det programmeras på lämpligt sätt, kommer att kunna känna igen varor som har passerat eller närmar sig bästföredatum, och sänder uppgifterna vidare till konsumenten.
Ytterligare utveckling planeras när systemet förbinds med Galileo.
I kommissionens meddelande av den 18 juni 2009
KOM(2009)0278 . , som detta initiativbetänkande utgår från, föreslås en handlingsplan med 14 initiativ, som bl.a. syftar till att utveckla sakernas Internet och främja dess spridning.
Föredragandens ståndpunkt
– radiovågornas inverkan på hälsan,
– chippens elektromagnetiska inverkan,
– återvinning av chippen,
– konsumenternas rätt till skydd av sitt privatliv,
– förekomsten av smarta chip i en viss produkt,
– rätten till ”chippens tystnad”,
– medborgarnas garantier när det gäller skydd av personuppgifter.
Som föredraganden ser det kommer utvecklingen av nya tillämpningar och funktionssättet för sakernas Internet och dess starka påverkan på EU-medborgarnas vardag och deras vanor att gå hand i hand med det förtroende som konsumenterna i EU har för systemet.
Det är därför viktigt att det finns ett regelverk och en rättslig ram som dels skyddar konsumenterna, dels stimulerar till offentliga och privata investeringar i sakernas Internet.
Sakernas Internet innebär stora ekonomiska möjligheter, eftersom det gör det möjligt att optimera produktionsmetoderna och energiförbrukningen, skapa nya arbetstillfällen och nya tjänster för allt fler medborgare och företag i EU.
YTTRANDE från utskottet för internationell handel
till utskottet för industrifrågor, forskning och energi
över sakernas Internet
( 2009/2224(INI) )
Föredragande: William (The Earl of) Dartmouth
FÖRSLAG
Utskottet för internationell handel uppmanar utskottet för industrifrågor, forskning och energi att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet uppmanar kommissionen att utvärdera de eventuella effekterna av dess föreslagna strategi för de europeiska företagens produktivitet och konkurrenskraft på den internationella marknaden.
Europaparlamentet menar att sakernas Internet kan bidra till att främja handelsflödena mellan EU och tredjeländer genom att marknaderna utvidgas och kvalitetsgarantier för handelsvarorna säkerställs.
Europaparlamentet uppmanar kommissionen att aktivt bidra till att bestämma och fastställa principer och regler för förvaltningen av sakernas Internet med sina handelsparter i internationella forum, såsom Världshandelsorganisationen.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
28.4.2010
Slutomröstning: resultat
+:
–:
0:
17
1
Slutomröstning: närvarande ledamöter
Kader Arif, Daniel Caspary, Joe Higgins, Yannick Jadot, Metin Kazak, Bernd Lange, Emilio Menéndez del Valle, Vital Moreira, Niccolò Rinaldi, Helmut Scholz, Peter Šťastný, Gianluca Susta, Jan Zahradil, Pablo Zalba Bidegain, Paweł Zalewski
Slutomröstning: närvarande suppleanter
YTTRANDE från utskottet för den inre marknaden och konsumentskydd
till utskottet för industrifrågor, forskning och energi
över sakernas Internet
( 2009/2224(INI) )
Föredragande: Christian Engström
FÖRSLAG
Utskottet för den inre marknaden och konsumentskydd uppmanar utskottet för industrifrågor, forskning och energi att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet välkomnar kommissionens planer på att under 2010 offentliggöra ett meddelande om personlig integritet och förtroende i informationssamhället och att fortsätta övervaka aspekterna beträffande skydd av personuppgifter för att trygga konsumenternas rättigheter och intressen.
Europaparlamentet betonar att konsumenterna behöver öppenhet beträffande följdkostnader, till exempel när det gäller strömförbrukning vid inkoppling och användning av saker.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
28.4.2010
Slutomröstning: resultat
+:
–:
0:
27
1
Slutomröstning: närvarande ledamöter
Cristian Silviu Buşoi, Lara Comi, Anna Maria Corazza Bildt, António Fernando Correia De Campos, Jürgen Creutzmann, Christian Engström, Evelyne Gebhardt, Louis Grech, Małgorzata Handzlik, Malcolm Harbour, Sandra Kalniete, Alan Kelly, Eija-Riitta Korhola, Edvard Kožušník, Giovanni La Via, Kurt Lechner, Toine Manders, Hans-Peter Mayer, Mitro Repo, Dominique Riquet, Robert Rochefort, Zuzana Roithová, Heide Rühle, Andreas Schwab, Róża Gräfin Von Thun Und Hohenstein, Kyriacos Triantaphyllides, Bernadette Vergnaud
Slutomröstning: närvarande suppleanter
YTTRANDE från utskottet för rättsliga frågor
till utskottet för industrifrågor, forskning och energi
över sakernas Internet
( 2009/2224(INI) )
Föredragande:
Eva Lichtenberger
FÖRSLAG
Utskottet för rättsliga frågor uppmanar utskottet för industrifrågor, forskning och energi att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
A. Framtidens Internet kommer att överskrida dagens traditionella gränser för den virtuella världen genom att kopplas till de fysiska föremålens värld.
Europaparlamentet uppskattar det faktum att kommissionen reagerar i god tid på den nya utvecklingen inom denna sektor så att det politiska systemet kan fastställa regler tillräckligt tidigt.
Europaparlamentet framhåller att det är viktigt att främja säkerhetsnormer genom att se till att alla eventuella personuppgifter som lagras i chippet inte kan avläsas av tredje part utan att de berörda personerna är medvetna om detta.
10.
Europaparlamentet begär att största möjliga vaksamhet iakttas när det gäller respekten för de grundläggande rättigheterna vid användningen av RFID-chip, eftersom varje person som har tillgång till en lämplig läsare kan avläsa innehållet i dessa chip, vilka kan innehålla personuppgifter som gör det möjligt att identifiera den berörda personen på avstånd.
Europaparlamentet betonar att uppgiftsskyddet – som har blivit nödvändigt i vårt moderna och demokratiska europeiska samhälle, där allt större volymer av personuppgifter samlas in, tas fram och analyseras – bör betraktas som en princip av författningsmässigt värde.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
28.4.2010
Slutomröstning: resultat
+:
–:
0:
22
1
Slutomröstning: närvarande ledamöter
Raffaele Baldassarre, Luigi Berlinguer, Sebastian Valentin Bodu, Françoise Castex, Christian Engström, Lidia Joanna Geringer de Oedenberg, Daniel Hannan, Klaus-Heiner Lehne, Antonio López-Istúriz White, Antonio Masip Hidalgo, Alajos Mészáros, Bernhard Rapkay, Evelyn Regner, Francesco Enrico Speroni, Kay Swinburne, Alexandra Thein, Diana Wallis, Rainer Wieland, Cecilia Wikström, Tadeusz Zwiefka
Slutomröstning: närvarande suppleanter
Piotr Borys, Sergio Gaetano Cofferati, Kurt Lechner, Eva Lichtenberger, József Szájer
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
4.5.2010
Slutomröstning: resultat
+:
–:
0:
47
Slutomröstning: närvarande ledamöter
Slutomröstning: närvarande suppleanter
António Fernando Correia De Campos, Andrzej Grzyb, Rebecca Harms, Ivailo Kalfin, Silvana Koch-Mehrin, Bernd Lange, Werner Langen, Marian-Jean Marinescu, Vladimír Remek, Silvia-Adriana Ţicău, Catherine Trautmann, Lambert van Nistelrooij, Hermann Winkler
A7-0181/2010
BETÄNKANDE
om förslaget till Europaparlamentets och rådets beslut om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
(KOM(2010)0196 – C7‑0116/2010 – 2010/2067(BUD))
Budgetutskottet
Föredragande: Barbara Matera
PE 441.290v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
BILAGA: EUROPAPARLAMENTETS OCH RÅDETS BESLUT..............................................6
MOTIVERING............................................................................................................................8
BILAGA: SKRIVELSE FRÅN UTSKOTTET FÖR SYSSELSÄTTNING OCH SOCIALA FRÅGOR 11
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................14
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om förslaget till Europaparlamentets och rådets beslut om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
( KOM(2010)0196 – C7‑0116/2010 – 2010/2067(BUD) )
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2010)0196 – C7‑0116/2010 ),
– med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
EUT C 139, 14.6.2006, s.
1. , särskilt punkt 28,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1927/2006 av den 20 december 2006 om upprättande av Europeiska fonden för justering för globaliseringseffekter
EUT L 406, 30.12.2006, s.
1. ,
– med beaktande av betänkandet från budgetutskottet ( A7‑0181/2010 ), och av följande skäl:
A. Europeiska unionen har inrättat lagstiftningsinstrument och budgetinstrument för att kunna ge kompletterande stöd till arbetstagare som blivit arbetslösa till följd av genomgripande strukturförändringar inom världshandeln och för att underlätta deras återinträde på arbetsmarknaden.
B. Tillämpningsområdet för fonden har utvidgats för ansökningar om stöd från fonden som inges från och med den 1 maj 2009 och omfattar nu stöd till arbetstagare som har blivit uppsagda som en direkt följd av den globala finansiella och ekonomiska krisen.
C. Unionens ekonomiska stöd till arbetstagare som har blivit uppsagda bör vara dynamiskt och ges så snabbt och effektivt som möjligt, i enlighet med Europaparlamentets, rådets och kommissionens gemensamma uttalande, som antogs vid förlikningsmötet den 17 juli 2008, och med vederbörlig hänsyn till bestämmelserna i det interinstitutionella avtalet av den 17 maj 2006 om antagandet av beslut rörande fondens utnyttjande.
D. Irland har ansökt om ekonomiskt bidrag ur fonden till följd av uppsägningar vid Waterford Crystal och tre av dess underleverantörer (Thomas Fennell Engineering Ltd, RPS Engineering Services och Abbey Electric) som är verksamma inom kristallglasbranschen
EGF/2009/012 IE/Waterford Crystal. .
E. Ansökan uppfyller kriterierna för berättigande till stöd enligt förordningen om upprättande av Europeiska fonden för justering för globaliseringseffekter.
Europaparlamentet påminner kommissionen om att den i samband med utnyttjandet av Europeiska fonden för justering för globaliseringseffekter inte systematiskt ska överföra betalningsbemyndiganden från ESF, eftersom Europeiska fonden för justering för globaliseringseffekter inrättades som ett enskilt och särskilt instrument med sina egna mål och tidsfrister.
Europaparlamentet välkomnar det nya formatet för kommissionens förslag, där det i motiveringsdelen läggs fram tydliga och detaljerade uppgifter om ansökan med en analys av kriterier för stödberättigande och en förklaring av orsakerna till att ansökan godkänts, vilket ligger i linje med parlamentets krav.
BILAGA: EUROPAPARLAMENTETS OCH RÅDETS BESLUT
av den ... maj 2010
om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av fördraget om Europeiska unionens funktionssätt,
med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
EUT C 139, 14.6.2006, s.
1. , särskilt punkt 28,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1927/2006 av den 20 december 2006 om upprättande av Europeiska fonden för justering av globaliseringseffekter
EUT L 406, 30.12.2006, s.
1. , särskilt artikel 12.3,
EUT C (…), (…), s. (…). ,
och av följande skäl:
(2) Fondens tillämpningsområde utvidgades, när det gäller ansökningar som lämnades från och med den 1 maj 2009, till att omfatta stöd för arbetstagare som sagts upp som en direkt följd av den globala ekonomiska krisen.
(3) Det interinstitutionella avtalet av den 17 maj 2006 gör det möjligt att utnyttja medel från fonden inom den årliga övre gränsen på 500 miljoner euro.
Denna ansökan uppfyller kraven för ekonomiska bidrag i artikel 10 i förordning (EG) nr 1927/2006.
Kommissionen föreslår därför att ett belopp på 2 570 853 euro ska anslås.
(5) Fonden bör därför utnyttjas för att tillhandahålla ett ekonomiskt bidrag för den ansökan som Irland lämnat in.
HÄRIGENOM FÖRESKRIVS FÖLJANDE:
Artikel 1
Europeiska fonden för justering av globaliseringseffekter ska tas i anspråk för att tillhandahålla beloppet 2 570 853 euro för åtagande- och betalningsbemyndiganden i Europeiska unionens allmänna budget för budgetåret 2010.
Artikel 2
Ordförande Ordförande
MOTIVERING
Europeiska fonden för justering för globaliseringseffekter har inrättats för att ge kompletterande stöd till arbetstagare som drabbats av konsekvenserna av större strukturella förändringar i världshandelsmönstren.
Enligt bestämmelserna i punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 om budgetdisciplin och sund ekonomisk förvaltning
EUT C 139, 14.6.2006, s.
1. och artikel 12 i förordning (EG) nr 1927/2006
EUT L 406, 30.12.2006, s.
1. får det årliga belopp som avdelas för fonden inte överstiga 500 miljoner euro som tas från eventuella marginaler under det samlade utgiftstaket för det föregående året och/eller från outnyttjade åtagandebemyndiganden som frigjorts under de två senaste åren, med undantag för sådana som ingår under budgetrubrik 1b.
Anslagen förs in i budgeten i form av en avsättning så snart kommissionen har funnit tillräckliga marginaler och/eller frigjort åtaganden.
Förfarandet går till så att kommissionen efter en positiv bedömning av en ansökan lägger fram ett förslag till budgetmyndigheten om att utnyttja fonden och samtidigt gör en begäran om överföring av medel.
Parallellt kan ett trepartsförfarande anordnas för att nå en överenskommelse om utnyttjandet av fonden och de belopp som krävs.
Trepartsförfarandet kan genomföras i förenklad form.
II.
Nuläget: Kommissionens förslag
Den 6 maj 2010 antog kommissionen tre nya förslag till beslut om utnyttjande av Europeiska fonden för globaliseringseffekter till förmån för Irland och Spanien för att stödja återintegrering på arbetsmarknaden av arbetstagare som har blivit uppsagda som en följd av den globala finansiella och ekonomiska krisen.
Detta förslag gäller Irlands ansökan till följd av uppsägningar i Waterford Crystal och tre av dess underleverantörer.
Detta är den sjunde ansökan som ska behandlas inom ramen för budgeten för 2010.
Denna ansökan, ärende EGF/2009/012 IE/Waterford Crystal, lämnades in till kommissionen den 7 augusti 2009.
Kommissionens bedömning baserades på en analys av sambandet mellan uppsägningarna och genomgripande strukturförändringar inom världshandeln eller finanskrisen, den oförutsägbara karaktären på de aktuella uppsägningarna, belägg för antalet uppsagda och uppfyllande av kriterierna i artikel 2, förklaring till uppsägningarnas oförutsägbara karaktär, uppgift om vilka företag som tvingas avskeda personal och vilka arbetstagare som stödet ska riktas till, en beskrivning av det berörda territoriet och dess myndigheter och övriga aktörer, de förväntade konsekvenserna av uppsägningarna för den lokala, regionala eller nationella sysselsättningen, det samordnade paketet med individanpassade tjänster som ska finansieras tillsammans med uppgifter om hur det kompletterar åtgärder som finansieras genom strukturfonderna, det eller de datum då man började eller planerar att börja tillhandahålla individanpassade tjänster till de berörda arbetstagarna, förfaranden för samråd med arbetsmarknadens parter samt system för ledning och kontroll.
Enligt kommissionens bedömning har kriterierna för berättigande till stöd enligt förordningen om upprättande av Europeiska fonden för justering för globaliseringseffekter uppfyllts i ansökan.
För att utnyttja fonden har kommissionen överlämnat en begäran om överföring (DEC 09/2010) till budgetmyndigheten om ett sammanlagt belopp på 2 570 853 euro från reserven för Europeiska fonden för justering för globaliseringseffekter (40 02 43) för åtagandebemyndiganden och från ESF:s budgetpost (04 02 17 – ESF konvergens) för betalningsbemyndiganden till budgetposten för Europeiska fonden för justering för globaliseringseffekter (04 05 01).
När det gäller alternativa källor till betalningsanslagen har kommissionen förklarat att man hittills har tagit de nödvändiga betalningsanslagen från Europeiska socialfondens budget eftersom det rör sig om närliggande politikområden och med tanke på att det årliga kravet för betalningsanslag från Europeiska fonden för justering av globaliseringseffekter än så länge har legat på omkring 1 procent av Europeiska socialfondens betalningskapital.
Såhär i början av budgetåret är det svårt att hitta alternativa källor.
För att kunna tillgodose denna begäran i samband med framtida ärenden som rör fonden är kommissionen dock villig att söka efter alternativa källor till betalningsanslagen, när så är möjligt och lämpligt, och när det inte finns någon risk för att behandlingen av begäran om överföring försenas.
Enligt det interinstitutionella avtalet får fonden utnyttjas upp till det årliga taket på 500 miljoner EUR.
Under 2010 har budgetmyndigheten redan godkänt fem förslag till utnyttjande av fonden, för ett totalbelopp på 16 338 363 euro för Tyskland (Karmann) och Litauen (Snaige, byggande av hus, möbel- och klädestillverkning), vilket innebär att det kvarstår 483 661 637 euro.
III.
Förfarande
Kommissionen har inkommit med en begäran om överföring
DEC 09/2010 av den 6 maj 2010. för att föra in specifika åtagande- och betalningsbemyndiganden i 2010 års budget i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006.
Enligt en intern överenskommelse ska utskottet för sysselsättning och sociala frågor delta i processen för att konstruktivt stödja och bidra till bedömningen av ansökningarna från fonden.
Efter sin bedömning lade Europaparlamentets utskott för sysselsättning och sociala frågor fram sina synpunkter på utnyttjandet av fonden, vilka beskrivs i det yttrande som bifogas detta betänkande.
I Europaparlamentets, rådets och kommissionens gemensamma uttalande, som antogs under förlikningsmötet den 17 juli 2008, bekräftades vikten av att säkerställa ett snabbt förfarande, med vederbörlig respekt för det interinstitutionella avtalet, för att anta beslut om utnyttjande av fonden.
BILAGA: SKRIVELSE FRÅN UTSKOTTET FÖR SYSSELSÄTTNING OCH SOCIALA FRÅGOR
ES/sg
D(2010)27788
Alain Lamassoure
Ordförande för budgetutskottet
ASP 13E158
Ärende: Yttrande över utnyttjandet av Europeiska fonden för justering för globaliseringseffekter för ärende EGF/2009/012 IE/Waterford Crystal, Irland ( KOM(2010)0196 )
EMPL-utskottet och arbetsgruppen för Europeiska fonden för justering för globaliseringseffekter är positiva till att utnyttja fonden för denna ansökan.
I detta sammanhang vill EMPL-utskottet framföra vissa synpunkter, utan att därför ifrågasätta överföringen av betalningsbemyndiganden.
EMPL-utskottets synpunkter grundar sig på följande överväganden:
b) De irländska myndigheterna påpekar i ansökan att företaget drabbades hårt av finanskrisen i oktober 2008 då det höll på att omstrukturera sina skulder och att de anser att om Waterford Crystal hade fått denna ytterligare finansiering skulle företaget ha lyckats omstrukturera sina skulder och kunnat fortsätta sin verksamhet genom att fokusera på sina huvudprodukter och fortsätta sina investeringar i nya produkter och processen att förlägga produktionen till lågkostnadsländer.
c) Mer än 72 procent av de arbetstagare som avskedats är äldre än 45 år och har aldrig arbetat vid något annat företag än Waterford Crystal.
d) Utbildningsministeriet inom den irländska regeringen ansvarar nu för ansökan om bidrag från Europeiska fonden för justering av globaliseringseffekter.
f) Det fanns företag i andra EU-medlemsstater som var direkt beroende av Waterford Wedgewood-gruppen.
g) Åtgärder till stöd för företagandet är mycket viktiga eftersom de innebär verkliga möjligheter för en ny yrkesmässig framtid för arbetstagare som blivit uppsagda och de utgör generellt grunden för inrättandet av nya arbetstillfällen.
Utskottet för sysselsättning och sociala frågor uppmanar därför budgetutskottet att som ansvarigt utskott infoga följande i sitt resolutionsförslag när det gäller Irlands ansökan:
Europaparlamentet beklagar emellertid att det gått så lång tid mellan den sista kompletterande informationen till ansökan mottogs den 3 november 2009 och kommissionens slutliga beslut den 6 maj 2010.
Europaparlamentet upprepar därför sin uppmaning till kommissionen att i sin årsrapport ta med uttömmande information om komplementariteten mellan Europeiska fonden för justering för globaliseringseffekter och åtgärder som stöds av andra strukturfonder i överensstämmelse med artikel 6 i förordningen om Europeiska fonden för justering för globaliseringseffekter.
Med vänlig hälsning
Pervenche Berès
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
2.6.2010
Slutomröstning: resultat
+:
–:
0:
26
Slutomröstning: närvarande ledamöter
Marta Andreasen, Francesca Balzani, Lajos Bokros, Jean-Luc Dehaene, José Manuel Fernandes, Eider Gardiazábal Rubial, Salvador Garriga Polledo, Jens Geier, Ivars Godmanis, Estelle Grelier, Carl Haglund, Jutta Haug, Sidonia Elżbieta Jędrzejewska, Jan Kozłowski, Alain Lamassoure, Vladimír Maňka, Miguel Portas, Dominique Riquet, László Surján, Derek Vaughan, Angelika Werthmann, Jacek Włosowicz
Slutomröstning: närvarande suppleanter
Paul Rübig
Slutomröstning: närvarande suppleanter (art.
187.2)
Peter Jahr, Andres Perello Rodriguez, Britta Reimers
A7-0318/2010
om förslaget till Europaparlamentets och rådets beslut om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
(KOM(2010)0529 – C7‑0309/2010 – 2010/2225(BUD))
Budgetutskottet
Föredragande: Barbara Matera
PE 450.599v02-00
INNEHÅLL
BILAGA: SKRIVELSE FRÅN UTSKOTTET FÖR SYSSELSÄTTNING OCH SOCIALA FRÅGOR 11
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om förslaget till Europaparlamentets och rådets om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
( KOM(2010)0529 – C7‑0309/2010 – 2010/2225(BUD) )
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2010)0529 – C7‑0309/2010 ),
– med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
EUT C 139, 14.6.2006, s.
1. , särskilt punkt 28,
EUT L 406, 30.12.2006, s.
1. ,
– med beaktande av skrivelsen från utskottet för sysselsättning och sociala frågor,
– med beaktande av betänkandet från budgetutskottet ( A7‑0318/2010 ), och av följande skäl:
A. Europeiska unionen har inrättat lagstiftningsinstrument och budgetinstrument för att kunna ge kompletterande stöd till arbetstagare som blivit arbetslösa till följd av genomgripande strukturförändringar inom världshandeln och för att underlätta deras återinträde på arbetsmarknaden.
B. Tillämpningsområdet för fonden har utvidgats för ansökningar om stöd från fonden som inges från och med den 1 maj 2009 och omfattar nu stöd till arbetstagare som har blivit uppsagda som en direkt följd av den globala finansiella och ekonomiska krisen.
C. Unionens ekonomiska stöd till arbetstagare som har blivit uppsagda bör vara dynamiskt och ges så snabbt och effektivt som möjligt, i enlighet med Europaparlamentets, rådets och kommissionens gemensamma uttalande, som antogs vid förlikningsmötet den 17 juli 2008, och med vederbörlig hänsyn till bestämmelserna i det interinstitutionella avtalet av den 17 maj 2006 om antagandet av beslut rörande fondens utnyttjande.
D. Nederländerna har ansökt om ekonomiskt bidrag från fonden till följd av 821 uppsägningar vid 70 företag som är verksamma inom sektorn Nace rev 2 huvudgrupp 18 (Grafisk produktion och reproduktion av inspelningar) i de två till varandra gränsande Nuts II-regionerna Noord Brabant och Zuid Holland.
E. Ansökan uppfyller kriterierna för berättigande till stöd enligt förordningen om upprättande av Europeiska fonden för justering för globaliseringseffekter.
Europaparlamentet välkomnar det nya formatet för kommissionens förslag, där det i motiveringsdelen läggs fram tydliga och detaljerade uppgifter om ansökan med en analys av kriterier för stödberättigande och en förklaring av orsakerna till att ansökan godkänts, vilket ligger i linje med parlamentets krav.
9.
BILAGA: EUROPAPARLAMENTETS OCH RÅDETS BESLUT
av den ...
om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning (ansökan EGF/2009/027 NL/ Noord Brabant och Zuid Holland huvudgrupp 18 från Nederländerna)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av fördraget om Europeiska unionens funktionssätt,
med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
EUT C 139, 14.6.2006, s.
1. , särskilt punkt 28,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1927/2006 av den 20 december 2006 om upprättande av Europeiska fonden för justering för globaliseringseffekter
EUT L 406, 30.12.2006, s.
med beaktande av Europeiska kommissionens förslag
EUT C […], […], s. […]. , och
av följande skäl:
(2) Tillämpningsområdet för fonden har utvidgats, och från och med den 1 maj 2009 är det möjligt att söka stöd för åtgärder som riktas till arbetstagare som har blivit uppsagda som en direkt följd av den globala finansiella och ekonomiska krisen.
(3) Det interinstitutionella avtalet av den 17 maj 2006 gör det möjligt att använda medel från fonden upp till ett belopp på högst 500 miljoner euro per år.
(4) Nederländerna lämnade den 30 december 2009 in en ansökan om medel från fonden med anledning av uppsägningar vid 70 företag som är verksamma inom huvudgrupp 18 (Grafisk produktion och reproduktion av inspelningar) enligt Nace rev 2, i de angränsande Nuts II-regionerna Noord Brabant (NL41) och Zuid Holland (NL33), och kompletterade ansökan med ytterligare uppgifter fram till den 11 maj 2010.
Ansökan uppfyller villkoren för fastställande av det ekonomiska stödet enligt artikel 10 i förordning (EG) nr 1927/2006.
Kommissionen föreslår därför att ett belopp på 2 890 027 euro ska anslås.
(5) Fonden bör därför utnyttjas för att bevilja det ekonomiska stöd som Nederländerna ansökt om.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Europeiska fonden för justering för globaliseringseffekter ska belastas med 2 890 027 euro i åtagande- och betalningsbemyndiganden ur Europeiska unionens allmänna budget för 2010.
Artikel 2
Detta beslut ska offentliggöras i Europeiska unionens officiella tidning .
Utfärdat i
På Europaparlamentets vägnar På rådets vägnar
Ordförande Ordförande
MOTIVERING
Europeiska fonden för justering för globaliseringseffekter har inrättats för att ge kompletterande stöd till arbetstagare som drabbats av konsekvenserna av större strukturella förändringar i världshandelsmönstren.
Enligt bestämmelserna i punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 om budgetdisciplin och sund ekonomisk förvaltning
EUT C 139, 14.6.2006, s.
1. och artikel 12 i förordning (EG) nr 1927/2006
EUT L 406, 30.12.2006, s.
1. får det årliga belopp som avdelas för fonden inte överstiga 500 miljoner euro som tas från eventuella marginaler under det samlade utgiftstaket för det föregående året och/eller från outnyttjade åtagandebemyndiganden som frigjorts under de två senaste åren, med undantag för sådana som ingår under budgetrubrik 1b.
Anslagen förs in i budgeten i form av en avsättning så snart kommissionen har funnit tillräckliga marginaler och/eller frigjort åtaganden.
Förfarandet går till så att kommissionen efter en positiv bedömning av en ansökan lägger fram ett förslag till budgetmyndigheten om att utnyttja fonden och samtidigt gör en begäran om överföring av medel.
Parallellt kan ett trepartsförfarande anordnas för att nå en överenskommelse om utnyttjandet av fonden och de belopp som krävs.
Trepartsförfarandet kan ske i förenklad form.
II.
Aktuellt läge: Kommissionens förslag
Den 1 oktober 2010 antog kommissionen ett nytt förslag till beslut om utnyttjande av Europeiska fonden för globaliseringseffekter till förmån för Nederländerna för att stödja återintegrering på arbetsmarknaden av arbetstagare som har blivit uppsagda som en följd av den globala finansiella och ekonomiska krisen.
Detta är den artonde ansökan som ska behandlas inom ramen för budgeten för 2010 och avser utnyttjande av ett totalbelopp på 2 890 027 euro från fonden till förmån för Nederländerna.
Ansökan avser 821 uppsägningar i 70 företag som är verksamma i sektorn Nace rev 2 huvudgrupp 18 (Grafisk produktion och reproduktion av inspelningar) inom de två till varandra gränsande Nuts II-regionerna Noord Brabant och Zuid Holland under referensperioden på nio månader från den 1 april 2009 till den 29 december 2009.
Denna ansökan, ärende EGF/2009/027 NL/Noord Brabant och Zuid Holland, lämnades in till kommissionen den 30 december 2009 och kompletterades med ytterligare uppgifter fram till den 11 maj 2010.
Enligt kommissionens bedömning har kriterierna för berättigande till stöd enligt förordningen om upprättande av Europeiska fonden för justering för globaliseringseffekter uppfyllts i ansökan.
Föredraganden är glad att kunna konstatera att kommissionen har pekat ut en alternativ källa till betalningsbemyndiganden, utöver oanvända medel från Europeiska socialfonden, i enlighet med upprepade krav från Europaparlamentet.
Hon anser dock att valet i detta fall (budgetpost avsedd för stöd till företagande och innovation) inte är tillfredsställande med tanke på de allvarliga brister som kommissionen stöter på vid genomförande av programmen för konkurrenskraft och innovation.
Under en period av ekonomisk kris bör dessa anslag faktiskt snarast höjas.
Föredraganden uppmanar därför kommissionen att fortsätta ansträngningarna för att hitta mera lämpliga budgetposter för betalningar i framtiden.
Enligt det interinstitutionella avtalet får fonden utnyttjas upp till det årliga taket på 500 miljoner EUR.
III.
Förfarande
Kommissionen har inkommit med en begäran om överföring
DEC 31/2010 av den 1 september 2010. för att föra in specifika åtagande- och betalningsbemyndiganden i 2010 års budget i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006.
Enligt en intern överenskommelse ska utskottet för sysselsättning och sociala frågor delta i processen för att konstruktivt stödja och bidra till bedömningen av ansökningarna ur fonden.
Efter sin bedömning lade Europaparlamentets utskott för sysselsättning och sociala frågor fram sina synpunkter på utnyttjandet av fonden, vilka beskrivs i det yttrande som bifogas detta betänkande.
I Europaparlamentets, rådets och kommissionens gemensamma uttalande, som antogs under förlikningsmötet den 17 juli 2008, bekräftades vikten av att säkerställa ett snabbt förfarande, med vederbörlig respekt för det interinstitutionella avtalet, för att anta beslut om utnyttjande av fonden.
BILAGA: SKRIVELSE FRÅN UTSKOTTET FÖR SYSSELSÄTTNING OCH SOCIALA FRÅGOR
ES/jm
D(2010)52566
Alain Lamassoure
Ordförande för budgetutskottet
ASP 13E158
Ärende: Yttrande om ianspråktagandet av Europeiska fonden för justering för globaliseringseffekter i ärendet EGF/2009/027 NL/Noord Brabant och Zuid Holland huvudgrupp 18 ( KOM(2010)0529 )
Utskottet för sysselsättning och sociala frågor och arbetsgruppen för Europeiska fonden för justering för globaliseringseffekter är positiva till att utnyttja fonden för denna ansökan.
I detta sammanhang vill utskottet för sysselsättning och sociala frågor framföra vissa synpunkter, utan att därför ifrågasätta överföringen av betalningsbemyndigandena.
EMPL-utskottets synpunkter grundar sig på följande överväganden:
A) Denna ansökan är baserad på artikel 2c i förordningen om Europeiska fonden för justering för globaliseringseffekter och omfattar 821 uppsägningar som inträffade under referensperioden på nio månader mellan den 1 april och den 29 december 2009 i 70 företag som arbetar med inom grafisk produktion och reproduktion av inspelningar, i enlighet med huvudgrupp 18 i förordning (EG) nr 1893/2006.
C) Denna sektor drabbades hårt av finanskrisen vilket ledde till ett fall i efterfrågan på tjänster och produkter från förlags- och tryckeribranschen med cirka 32 procent för tryckt reklammaterial och mellan 7,5 och 18,2 procent för tidskrifter och tidningar.
D) Den nederländska förlags- och tryckeribranschen genomgick en kostsam omstrukturering för att förbli tekniskt konkurrenskraftig i förhållande till företag från länder utanför EU, särskilt Turkiet, Kina och Indien och risken är att den på grund av krisen inte kan dra nytta av de stora investeringar och satsningar som gjorts.
H) Flera utbildningsprojekt som finansieras av Europeiska socialfonden och som är avsedda för arbetstagare i den grafiska sektorn har inrättats och utbildningen sammanfaller tidsmässigt med de åtgärder som ska finansieras genom fonden.
I) Nederländerna ansöker om stöd för alla arbetstagare som blivit uppsagda, inklusive de som är över 65 år gamla.
Utskottet för sysselsättning och sociala frågor uppmanar därför budgetutskottet att som ansvarigt utskott infoga följande förslag i sitt resolutionsförslag avseende Nederländernas ansökan:
Parlamentet beklagar dock att denna ansökan inte särskilt anger vilket mervärde som åtgärder från globaliseringsfonden skulle ge.
Med vänlig hälsning
Pervenche Berès
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
9.11.2010
Slutomröstning: resultat
+:
–:
0:
19
1
1
Slutomröstning: närvarande ledamöter
Alexander Alvaro, Reimer Böge, Lajos Bokros, Giovanni Collino, Göran Färm, José Manuel Fernandes, Eider Gardiazábal Rubial, Salvador Garriga Polledo, Jutta Haug, Jiří Havel, Ivailo Kalfin, Sergej Kozlík, Jan Kozłowski, Barbara Matera, Claudio Morganti, Miguel Portas, Dominique Riquet, László Surján, Helga Trüpel, Derek Vaughan, Angelika Werthmann
A7-0014/2011
***II
ANDRABEHANDLINGS-REKOMMENDATION
om rådets ståndpunkt vid första behandlingen inför antagandet av Europaparlamentets och rådets förordning om ändring av förordning (EG) nr 1889/2006 om inrättandet av ett finansieringsinstrument för främjande av demokrati och mänskliga rättigheter i hela världen
(16446/1/2010 – C7‑0427/2010 – 2009/0060B(COD))
Utskottet för utrikesfrågor
Föredragande:
Kinga Gál och Barbara Lochbihler
PE 456.703v02-00
Teckenförklaring
* Samrådsförfarande
*** Godkännandeförfarande
***I Ordinarie lagstiftningsförfarande (första behandlingen)
***II Ordinarie lagstiftningsförfarande (andra behandlingen)
***III Ordinarie lagstiftningsförfarande (tredje behandlingen)
(Det angivna förfarandet baseras på den rättsliga grund som angetts i förslaget till akt.)
Ändringsförslag till ett förslag till akt
Parlamentets ändringsförslag till ett förslag till akt ska markeras med fetkursiv stil .
De berörda avdelningarna tar sedan ställning till dessa korrigeringsförslag.
Om parlamentet önskar ändra delar av en bestämmelse i en befintlig akt som inte ändrats i förslaget till akt, ska dessa markeras med fet stil .
Eventuella strykningar ska i sådana fall markeras enligt följande: [...] .
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
ÄRENDETS GÅNG..................................................................................................................10
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om rådets ståndpunkt vid första behandlingen inför antagandet av Europaparlamentets och rådets förordning om ändring av förordning (EG) nr 1889/2006 om inrättandet av ett finansieringsinstrument för främjande av demokrati och mänskliga rättigheter i hela världen
(16446/1/2010 – C7‑0427/2010 – 2009/0060B(COD) )
(Ordinarie lagstiftningsförfarande: andra behandlingen)
Europaparlamentet utfärdar denna resolution
– med beaktande av rådets ståndpunkt vid första behandlingen (16446/1/2010 – C7‑0427/2010 ),
– med beaktande av sin ståndpunkt vid första behandlingen av ärendet
Antagna texter från sammanträdet 21.10.2010, P7_TA(2010)0380 . en behandling som avsåg kommissionens förslag till Europaparlamentet och rådet ( KOM(2009)0194 ),
– med beaktande av artikel 66 i arbetsordningen,
– med beaktande av andrabehandlingsrekommendationen från utskottet för utrikesfrågor ( A7‑0014/2011 ).
1.
EUROPAPARLAMENTETS STÅNDPUNKT
VID ANDRA BEHANDLINGEN
* Ändringar: ny text eller text som ersätter tidigare text markeras med fetkursiv stil och strykningar med symbolen ▌. *
---------------------------------------------------------
EUROPAPARLAMENTETS OCH RÅDETS FÖRORDNING
om ändring av förordning (EG) nr 1889/2006 om inrättandet av ett finansieringsinstrument för främjande av demokrati och mänskliga rättigheter i hela världen.
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europeiska kommissionens förslag,
i enlighet med det ordinarie lagstiftningsförfarandet
Europaparlamentets ståndpunkt av den 21 oktober 2010 (ännu ej offentliggjord i EUT) och rådets ståndpunkt vid första behandlingen av den 10 december 2010 (ännu ej offentliggjord i EUT).
Europaparlamentets ståndpunkt av den ... (ännu ej offentliggjord i EUT). ,
av följande skäl:
1) En ny ram för planeringen och tillhandahållandet av gemenskapens externa bistånd fastställdes 2006 i syfte att göra biståndet effektivare och öppnare.
Ramen omfattar rådets förordning (EG) nr 1085/2006 av den 17 juli 2006 om upprättande av ett instrument för stöd inför anslutningen
EUT L 210, 31.7.2006, s.
82. , Europaparlamentets och rådets förordning (EG) nr 1638/2006 av den 24 oktober 2006 om fastställande av allmänna bestämmelser för upprättandet av ett europeiskt grannskaps- och partnerskapsinstrument
EUT L 310, 9.11.2006, s.
1. , rådets förordning (EG) nr 1934/2006 av den 21 december 2006 om inrättande av ett finansieringsinstrument för samarbete med industriländer och andra höginkomstländer och territorier
EUT L 405, 30.12.2006, s.
41. , Europaparlamentets och rådets förordning (EG) nr 1717/2006 av den 15 november 2006 om upprättande av ett stabilitetsinstrument
EUT L 327, 24.11.2006, s.
1. , rådets förordning (Euratom) nr 300/2007 av den 19 februari 2007 om upprättande av ett instrument för kärnsäkerhetssamarbete
EUT L 81, 22.3.2007, s.
1. , Europaparlamentets och rådets förordning (EG) nr 1889/2006
EUT L 386, 29.12.2006, s.
1. och Europaparlamentets och rådets förordning (EG) nr 1905/2006 av den 18 december 2006 om upprättande av ett finansieringsinstrument för utvecklingssamarbete
EUT L 378, 27.12.2006, s.
41. .
2) Vid genomförandet av dessa förordningar har det framkommit inkonsekvenser när det gäller undantag till principen om att utgifter i samband med skatter, tullar och andra avgifter inte berättigar till unionsfinansiering.
Det föreslås därför att de relevanta bestämmelserna i förordning (EG) nr 1889/2006 ändras i syfte att anpassa den till de övriga instrumenten.
3a) Kommissionen bör ha befogenhet att anta delegerade akter i enlighet med artikel 290 i fördraget om Europeiska unionens funktionssätt när det gäller strategidokument, eftersom dessa kompletterar förordning (EG) nr 1889/2006 och gäller generellt.
Det är särskilt viktigt att kommissionen genomför lämpliga samråd under sitt förberedande arbete, inklusive på expertnivå.
4) Förordning (EG) nr 1889/2006 bör därför ändras i enlighet med detta.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 1889/2006 ska ändras på följande sätt:
1) Artikel 5.3 ska ersättas med följande:
”3.
Strategidokumenten och eventuella ändringar eller förlängningar av dessa ska antas av kommissionen genom delegerade akter i enlighet med artikel 17 och enligt villkoren i artiklarna 17a och 17b.”
2) Artikel 6.3 ska ersättas med följande:
”3.
De årliga handlingsprogrammen och eventuella ändringar eller förlängningar av dessa ska antas av kommissionen under beaktande av Europaparlamentets och rådets yttranden.”
3) Artikel 7.3 och 7.4 ska ersättas med följande:
”3.
Om utgifterna för de särskilda åtgärderna är lika med eller överstiger 3 000 000 EUR ska de antas av kommissionen under beaktande av Europaparlamentets och rådets yttranden.
4.
Om utgifterna för de särskilda åtgärderna understiger 3 000 000 EUR ska kommissionen underrätta Europaparlamentet och rådet om åtgärderna inom tio arbetsdagar efter antagandet av dess beslut.”
4) Artikel 9.2 ska ersättas med följande:
”2.
Kommissionen ska regelbundet underrätta Europaparlamentet och rådet om de ad hoc-åtgärder som vidtas.”
5) Artikel 13.6 ska ersättas med följande:
”6.
Stöd från unionen får i princip inte användas för att betala skatter, tullar eller andra avgifter i de stödmottagande länderna.”
6) Artikel 16.2 ska ersättas med följande:
”2.
Kommissionen ska för kännedom överlämna utvärderingsrapporterna till Europaparlamentet och rådet.
Resultaten ska användas för att förbättra utformningen av programmen och tilldelningen av resurser.”
7) Artikel 17 ska ersättas med följande:
”Artikel 17
Utövande av delegering
1.
2.
När kommissionen antar en delegerad akt, ska den samtidigt underrätta Europaparlamentet och rådet.
3.
Befogenheten att anta delegerade akter ges till kommissionen med förbehåll för de villkor som anges i artiklarna 17a och 17b.”
Artikel 17a
Återkallande av delegering
1.
Den delegering av befogenhet som avses i artikel 5 får när som helst återkallas av Europaparlamentet eller rådet.
2.
Den institution som har inlett ett internt förfarande för att besluta huruvida en delegering av befogenhet ska återkallas, ska sträva efter att underrätta den andra institutionen och kommissionen i rimlig tid innan det slutliga beslutet fattas, och ange vilken delegerad befogenhet som kan komma att återkallas samt skälen för återkallandet.
3.
Beslutet om återkallande innebär att delegeringen av de befogenheter som anges i beslutet upphör att gälla.
Det får verkan omedelbart, eller vid ett senare, i beslutet angivet datum.
Det påverkar inte giltigheten av delegerade akter som redan trätt i kraft.
Detta beslut ska offentliggöras i Europeiska unionens officiella tidning.
Artikel 17b
Invändning mot delegerade akter
1.
Europaparlamentet eller rådet får invända mot en delegerad akt inom en frist på två månader från delgivningsdagen.
På Europaparlamentets eller rådets initiativ ska fristen förlängas med två månader.
2.
Om varken Europaparlamentet eller rådet vid utgången av den frist som avses i punkt 1 har invänt mot den delegerade akten, ska den offentliggöras i Europeiska unionens officiella tidning och träda i kraft den dag som anges i den.
Den delegerade akten får offentliggöras i Europeiska unionens officiella tidning och träda i kraft före utgången av denna frist om både Europaparlamentet och rådet har underrättat kommissionen om att de har beslutat att inte göra invändningar.
3.
Om antingen Europaparlamentet eller rådet inkommer med invändningar mot en delegerad akt inom den frist som anges i punkt 1 ska akten inte träda i kraft.
Den institution som gör invändningar ska ange skälen till sina invändningar mot den delegerade akten.”
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Utfärdad i
På Europaparlamentets vägnar På rådets vägnar
Ordförande Ordförande
ÄRENDETS GÅNG
Titel
Finansieringsinstrument för främjande av demokrati och mänskliga rättigheter i hela världen (ändring av förordning (EG) nr 1889/2006)
Referensnummer
16446/1/2010 – C7-0427/2010 – 2009/0060B(COD)
Par lamentets första behandling – P ‑ nummer
21.10.2010 T7-0380/2010
Kommissionens förslag
KOM(2009)0194 - C7-0158/2009
Mottagande av rådets ståndpunkt vid första behandlingen: tillkännagivande i kammaren
16.12.2010
Ansvarigt utskott
Tillkännagivande i kammaren
AFET
16.12.2010
Föredragande
Utnämning
Barbara Lochbihler
13.1.2011
Kinga Gál
13.1.2011
Antagande
26.1.2011
Slutomröstning: resultat
+:
–:
0:
56
1
1
Slutomröstning: närvarande ledamöter
Gabriele Albertini, Pino Arlacchi, Sir Robert Atkins, Dominique Baudis, Franziska Katharina Brantner, Frieda Brepoels, Elmar Brok, Arnaud Danjean, Mário David, Michael Gahler, Andrzej Grzyb, Takis Hadjigeorgiou, Heidi Hautala, Anna Ibrisagic, Anneli Jäätteenmäki, Jelko Kacin, Tunne Kelam, Nicole Kiil-Nielsen, Maria Eleni Koppa, Andrey Kovatchev, Wolfgang Kreissl-Dörfler, Alexander Graf Lambsdorff, Vytautas Landsbergis, Ryszard Antoni Legutko, Sabine Lösing, Barry Madlener, Mario Mauro, Kyriakos Mavronikolas, Francisco José Millán Mon, Alexander Mirsky, María Muñiz De Urquiza, Annemie Neyts-Uyttebroeck, Norica Nicolai, Raimon Obiols, Ria Oomen-Ruijten, Pier Antonio Panzeri, Ioan Mircea Paşcu, Vincent Peillon, Alojz Peterle, Bernd Posselt, Hans-Gert Pöttering, Cristian Dan Preda, Libor Rouček, José Ignacio Salafranca Sánchez-Neyra, Nikolaos Salavrakos, Jacek Saryusz-Wolski, Werner Schulz, Adrian Severin, Marek Siwiec, Ernst Strasser, Hannes Swoboda, Charles Tannock, Inese Vaidere, Geoffrey Van Orden, Kristian Vigenin, Graham Watson, Boris Zala
Slutomröstning: närvarande suppleanter
Laima Liucija Andrikienė, Elena Băsescu, Emine Bozkurt, Nikolaos Chountis, Véronique De Keyser, Kinga Gál, Liisa Jaakonsaari, Evgeni Kirilov, Georgios Koumoutsakos, Barbara Lochbihler, Norbert Neuser, Doris Pack, Marietje Schaake, György Schöpflin, Alf Svensson, Ivo Vajgl, Renate Weber
Ingivande
28.1.2011
A7-0020/2011
***III
BETÄNKANDE
om förlikningskommitténs gemensamma utkast till Europaparlamentets och rådets förordning om passagerares rättigheter vid busstransport och om ändring av förordning (EG) nr 2006/2004
(PE-CONS 00063/2010 – C7‑0015/2011 – 2008/0237(COD))
Europaparlamentets delegation till förlikningskommittén
Delegationsordförande:
Rodi Kratsa-Tsagaropoulou
Föredragande: Antonio Cancian
PE 454.601v03-00
Teckenförklaring
* Samrådsförfarande
*** Godkännandeförfarande
***I Ordinarie lagstiftningsförfarande (första behandlingen)
***II Ordinarie lagstiftningsförfarande (andra behandlingen)
***III Ordinarie lagstiftningsförfarande (tredje behandlingen)
(Det angivna förfarandet baseras på den rättsliga grund som angetts i förslaget till akt.)
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING............................................................................................................................7
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förlikningskommitténs gemensamma utkast till Europaparlamentets och rådets förordning om passagerares rättigheter vid busstransport och om ändring av förordning (EG) nr 2006/2004
(PE-CONS 00063/2010 – C7‑0015/2011 – 2008/0237(COD) )
(Ordinarie lagstiftningsförfarande: tredje behandlingen)
Europaparlamentet utfärdar denna resolution
– med beaktande av förlikningskommitténs gemensamma utkast (PE-CONS 00063/2010 – C7‑0015/2011 ),
– med beaktande av yttrandet från Europeiska ekonomiska och sociala kommittén av den 16 juli 2009
EUT C 317, 23.12.2009, s.
99. ,
– med beaktande av sin ståndpunkt vid första behandlingen av ärendet
EUT C 184, 8.7.2010, s.
312. , en behandling som avsåg kommissionens förslag till Europaparlamentet och rådet ( KOM(2008)0817 ),
– med beaktande av parlamentets ståndpunkt vid andra behandlingen av ärendet
Antagna texter från sammanträdet 6.7.2010, P7_TA(2010)0256 . , en behandling som avsåg rådets ståndpunkt vid första behandlingen
EUT C 122 E, 11.5.2010, s.
1. ,
– med beaktande av kommissionens yttrande över parlamentets ändringar i rådets ståndpunkt vid första behandlingen ( KOM(2010)0469 ),
– med beaktande av artikel 69 i arbetsordningen,
– med beaktande av betänkandet från parlamentets delegation till förlikningskommittén ( A7‑0020/2011 ).
1.
Europaparlamentet godkänner det gemensamma utkastet.
2.
Europaparlamentet uppdrar åt talmannen att tillsammans med rådets ordförande underteckna akten i enlighet med artikel 297.1 i fördraget om Europeiska unionens funktionssätt.
MOTIVERING
Bakgrund
Den 4 december 2008 lade kommissionen fram ett förslag till förordning om passagerares rättigheter vid busstransport.
Med tanke på den stadiga tillväxten inom denna transportbransch var syftet med förslaget att upprätta EU-övergripande rättigheter för skydd av passagerare som är jämförbara med de som gäller för andra transportslag och att säkerställa en rättvis konkurrens mellan dels transportörer från olika medlemsstater, dels olika transportslag.
Det ordinarie lagstiftningsförfarandet och förlikningsförfarandet
Efter parlamentets ståndpunkt vid första behandlingen från den 23 april 2009 antog rådet sin ståndpunkt vid första behandlingen den 11 mars 2010.
I denna ändrade rådet centrala delar av förslaget till förordning genom att urvattna eller helt ta bort flera viktiga bestämmelser som fanns i både kommissionens förslag och parlamentets ståndpunkt vid första behandlingen.
Vid sin andra behandling den 6 juli 2010 antog parlamentet 50 ändringsförslag till rådets ståndpunkt.
De frågor som det rådde mest oenighet om var: förordningens tillämpningsområde och tidsplanen för att införa den, regler om ansvar, skadestånd och assistans, rättigheter för personer med funktionshinder eller nedsatt rörlighet, passagerares rättigheter vid inställda resor eller förseningar samt hantering av klagomål och nationella tillsynsorgan.
Eftersom rådet inte kunde godta alla parlamentets ändringar krävdes det ett förlikningsförfarande.
Parlamentets delegation höll sitt konstituerande sammanträde den 8 september 2010 i Strasbourg.
Delegationen gav Kratsa-Tsagaropoulou, vice talman och ordförande för delegationen, Simpson, ordförande för utskottet för transport och turism och Cancian, föredragande, mandat att förhandla med rådet.
Det hölls trepartsmöten den 13 september, 13 oktober och 16 november, som följdes upp av möten med parlamentets delegation den 19 oktober och 23 november.
Trepartsmötena ledde till vissa framsteg i ett antal frågor men frågan om förordningens tillämpningsområde visade sig vara den stora stötestenen.
Förlikningskommittén hade ett möte i Europaparlamentet kvällen den 30 november 2010 i syfte att formellt öppna förlikningsförfarandet och eventuellt nå en överenskommelse i alla återstående frågor.
Efter flera timmars förhandlingar nådde man en övergripande överkommelse under natten.
Denna överenskommelse godkändes av parlamentets delegation med arton röster för, en röst emot och tre nedlagda röster.
Huvudpunkterna i överenskommelsen
Överenskommelsens huvudpunkter kan sammanfattas på följande sätt:
Tillämpningsområde
Förordningen ska gälla för all nationell och gränsöverskridande linjetrafik på en sträcka om minst 250 kilometer (fjärrtrafik).
Passagerare som endast reser en del av en sådan fjärrtrafiksträcka omfattas också.
Dessutom kommer tolv grundläggande rättigheter som förordningen ger även att gälla för passagerare som reser reguljärt på kortare sträckor.
Dessa gäller framför behoven hos personer med funktionshinder eller nedsatt rörlighet, såsom icke-diskriminerande tillgång till transporter, rätt att kompenseras för förlust av eller skada på rullstolar och annan rörlighetsutrustning, inlämnande och hantering av klagomål, utbildning om funktionshinder för busspersonal, information som ska ges under resan osv.
Avviskelser från tidsplanen
Förutom dessa grundläggande rättigheter får medlemsstaterna undanta inhemsk reguljärtrafik från tillämpningen av förordningen under en period om högst fyra år, vilket kan förlängas en gång.
Medlemsstaterna får också under fyra år med möjlighet till förlängning en gång, undanta vissa sträckor om en betydande del av sträckan går utanför unionen.
Ersättning och assistans i händelse av olyckor
Passagerare har rätt till ersättning vid dödsfall, inklusive för rimliga begravningskostnader, eller personskada och för bagage som förlorats eller skadats på grund av olyckor.
Taken för sådana ersättningar får i den nationella lagstiftningen inte understiga de minimibelopp som fastställs i förordningen, dvs. 220 000 euro per passagerare och 1 200 euro per bagagekolli.
Skada på hjälpmedel såsom rullstolar ska ersättas i sin helhet.
Vid en olycka har passagerarna dessutom rätt till assistans för att täcka sina omedelbara praktiska behov, däribland mat och kläder, transporter, hjälp med inledande assistans och logi för upp till 80 euro per natt och passagerare för högst två nätter.
Passagerares rättigheter vid inställda resor eller förseningar
Om en reguljär bussavgång är inställd, försenad med mer än 120 minuter eller överbokad ska passagerarna omedelbart ges rätt att välja mellan att fortsätta resan, att utan extra kostnad ombokas till sin slutstation eller att få biljettpriset återbetalat.
Om transportören inte erbjuder denna möjlighet ska passageraren ha rätt till kompensation motsvarande 50 procent av biljettpriset, utöver att biljettpriset återbetalas.
I de fall då bussen blir köroduglig under en resa, ska transportören tillhandahålla antingen vidareresa med annat fordon eller transport till en lämplig väntplats eller terminal, varifrån resan kan fortsätta.
Rättigheter för personer med funktionshinder eller nedsatt rörlighet
Bussföretag måste ge assistans till personer med funktionshinder eller nedsatt rörlighet förutsatt att passageraren informerar företaget om sina behov senast 36 timmar före avgång.
Om transportören inte kan ge lämplig assistans har den passagerare som har nedsatt rörlighet rätt att utan extra kostnad ledsagas av en person som han eller hon själv utser.
Alla förluster av och skador på rullstolar och annan hjälputrusning måste kompenseras av företaget eller ledningsorganet vid den ansvariga stationen.
Slutsats
Den slutliga texten är en mycket tillfredsställande och välbalanserad kompromiss eftersom den säkerställer passagerarnas rättigheter utan att utgöra en stor belastning för transportörerna, som ofta är små och medelstora företag.
Framför allt kan resultatet av förlikningsförfarandet ses som en framgång för parlamentet med tanke på följande:
a) För tillämpningsområdet var rådets ursprungliga förhandlingsståndpunkt 500 kilometer medan kompromissen blev 250 kilometer.
b) I sin ursprungliga ståndpunkt angav rådet tre grundläggande passagerarrättigheter som ska gälla oavsett avstånd medan den slutliga kompromissen innehåller tolv sådana rättigheter, där man särskilt fokuserar på behoven hos personer med funktionshinder eller nedsatt rörlighet.
c) För undantagen ville rådet ursprungligen se 15 år för inhemsk trafik och en obegränsad tid för internationell trafik, medan den slutliga kompromissen innebär högst åtta år i båda fall (en period om fyra år som kan förnyas en gång).
d) Vid en olycka eller om en avgång ställs in eller försenas med mer än 90 minuter ska varje passagerare vid behov ha rätt till hotellogi till en total kostnad av 80 euro per natt under högst två nätter, medan rådets ursprungliga ståndpunkt var 50 euro.
e) Vid en olycka ska passagerarna ha rätt till omedelbar assistans, däribland logi (se ovan), mat, kläder, transporter och hjälp med inledande assistans.
f) Om en avgång är inställd, försenad med mer än 120 minuter eller överbokad, ska passagerarna ha rätt till ersättning motsvarande 50 procent av biljettpriset, utöver rätten att välja mellan att fortsätta resan eller att ombokas till sin slutstation eller att återbetalas biljettpriset.
g) Avtalet ger möjlighet för passagerare att på elektronisk väg få uppdaterad information i realtid.
Parlamentets delegation till förlikningskommittén rekommenderar därför att det gemensamma utkastet antas vid tredje behandlingen.
ÄRENDETS GÅNG
Titel
Förslag till Europaparlamentets och rådets förordning om passagerares rättigheter vid busstransport och om ändring av förordning (EG) nr 2006/2004
Referensnummer
PE-CONS 63/2010 – C7‑0015/2011 – 2008/0237(COD)
Delegationsordförande: vice talman
Rodi Kratsa-Tsagaropoulou
Ansvarigt utskott
Ordförande
TRAN
Brian Simpson
Föredragande
Antonio Cancian
Förslag till akt – första behandlingen
KOM(2008)0817 – C6‑0469/2008
Parlamentets första behandling – P ‑nummer
23.04.2009
P6_TA(2009)0281
Kommissionens ändrade förslag
Rådets ståndpunkt vid första behandlingen
Tillkännagivande i kammaren
05218/3/2010 – C7‑0077/2010
Kommissionens ståndpunkt (artikel 294.6 i fördraget om Europeiska unionens funktionssätt,
KOM(2010)0121
Parlamentets andra behandling – P ‑nummer
06.07.2010
P7_TA(2010)0256
KOM(2010)0469
Datum för rådets mottagande av parlamentets ståndpunkt vid andra behandlingen
09.08.2010
Datum för rådets skrivelse om icke godkännande av parlamentets ändringar
25.11.2010
Förlikningskommitténs sammanträden
30.11.2010
Omröstning i parlamentets delegation
30.11.2010
Slutomröstning: resultat
+:
–:
0:
18
1
3
Närvarande ledamöter
Rodi Kratsa-Tsagaropoulou, Antonio Cancian, Brian Simpson, Georges Bach, Mathieu Grosch, Dieter-Lebrecht Koch, Ádám Kósa, Marian-Jean Marinescu, Inés Ayala Sender, Saïd El Khadraoui, Debora Serracchiani, Izaskun Bilbao Barandica, Michael Cramer, Eva Lichtenberger
Närvarande suppleanter
Carlo Fidanza, Werner Kuhn, Bogdan Kazimierz Marcinkiewicz, Hella Ranner, Spyros Danellis, Ismail Ertug, Nathalie Griesbeck, Vilja Savisaar-Toomast; Guido Milana
Närvarande suppleanter (art.
Datum för enighet i förlikningskommittén
30.11.2010
Enighet efter skriftväxling
0.0.0000
0.0.0000
Datum då ordförandena förklarade det gemensamma utkastet för godkänt och översände det till parlamentet och rådet
24.1.2011
Ingivande
2.2.2011
...
A7-0029/2011
om jämställdhet mellan kvinnor och män i Europeiska unionen – 2010
(2010/2138(INI))
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
Föredragande: Mariya Nedelcheva
PE 450.870v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING..........................................................................................................................18
YTTRANDE från utskottet för sysselsättning och sociala frågor ...20
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................26
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om jämställdhet mellan kvinnor och män i Europeiska unionen – 2010
( 2010/2138(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av artikel 23 i Europeiska unionens stadga om de grundläggande rättigheterna,
– med beaktande av Europeiska konventionen om skydd för de mänskliga rättigheterna och de grundläggande friheterna,
– med beaktande av Stockholmsprogrammet
Europeiska unionens råds dokument nr 5731/10 av den 3 mars 2010. ,
– med beaktande av rådets direktiv 2000/43/EG av den 29 juni 2000 om genomförandet av principen om likabehandling av personer oavsett deras ras eller etniska ursprung
EGT L 180, 19.7.2000, s.
22. , rådets direktiv 2000/78/EG av den 27 november 2000 om inrättande av en allmän ram för likabehandling
EGT L 303, 2.12.2000, s.
16. och rådets direktiv 2004/113/EG av den 13 december 2004 om genomförande av principen om likabehandling av kvinnor och män när det gäller tillgång till och tillhandahållande av varor och tjänster
EUT L 373, 21.12.2004, s.
37. ,
– med beaktande av kommissionens årliga rapporter om jämställdhet mellan kvinnor och män i Europeiska unionen 2000, 2001, 2002, 2004, 2005, 2006, 2007 och 2008 ( KOM(2001)0179 , KOM(2002)0258 , KOM(2003)0098 , KOM(2004)0115 , KOM(2005)0044 , KOM(2006)0071 , KOM(2007)0049 respektive KOM(2008)0010 ),
– med beaktande av kommissionens rapport av den 18 december 2009 om jämställdhet mellan kvinnor och män – 2010 ( KOM(2009)0694 ),
– med beaktande av Europaparlamentets och rådets direktiv 2006/54/EG av den 5 juli 2006 om genomförandet av principen om lika möjligheter och likabehandling av kvinnor och män i arbetslivet (omarbetning)
EUT L 204, 26.7.2006, s.
23. ,
EUT L 180, 15.7.2010, s.
EUT L 68, 18.3.2010, s.
– med beaktande av direktiv 89/552/EEG, ”Television utan gränser”,
– med beaktande av kommissionens rapport av den 3 oktober 2008 ”Förverkligande av Barcelonamålen avseende barnomsorg före den obligatoriska skolåldern” ( KOM(2008)0638 ),
– med beaktande av kommissionens meddelande av den 21 september 2010 ”Strategi för jämställdhet 2010–2015” ( KOM(2010)0491 ),
– med beaktande av FN:s konvention om avskaffande av all slags diskriminering av kvinnor från 1979 och FN:s handlingsplattform från Peking,
– med beaktande av den europeiska jämställdhetspakt som Europeiska rådet antog den 23−24 mars 2006,
– med beaktande av Europeiska kommissionens rådgivande kommitté för lika möjligheter för kvinnor och män och av dess yttrande av den 22 mars 2007 om löneskillnader mellan könen,
– med beaktande av Europarådets människorättskommissaries dokument om mänskliga rättigheter och könsidentitet (2009),
– med beaktande av rapporten från byrån för grundläggande rättigheter om homofobi, transfobi och diskriminering på grund av sexuell läggning och könsidentitet (2010),
– med beaktande av sin resolution av den 6 maj 2009 om aktiv inkludering av människor som är utestängda från arbetsmarknaden
P6_TA(2009)0371 . ,
– med beaktande av sin resolution av den 10 februari 2010 om jämställdhet mellan kvinnor och män – 2009
P7_TA(2010)0021 . ,
– med beaktande av sin resolution av den 17 juni 2010 om jämställdhetsaspekterna av den ekonomiska och finansiella krisen
P7_TA(2010)0231 . ,
– med beaktande av sin resolution av den 17 juni 2010 om utvärderingen av resultaten från färdplanen för jämställdhet 2006–2010 och rekommendationer för framtiden
P7_TA(2010)0232 . ,
– med beaktande av sin resolution av den 19 oktober 2010 om kvinnor med otrygga anställningsförhållanden,
– med beaktande av sin resolution av den 13 mars 2007 om en färdplan för jämställdhet 2006–2010
EUT C 301 E, 13.12.2007, s.
56. ,
– med beaktande av sin resolution av den 3 september 2008 om jämställdhet mellan kvinnor och män – 2008
EUT C 259 E, 4.12.2009, s.
35. ,
– med beaktande av sin resolution av den 18 november 2008 med rekommendationer till kommissionen om tillämpningen av principen om likalön för kvinnor och män
EUT C 16 E, 22.1.2010, s.
21. ,
– med beaktande av sin resolution av den 15 december 2010 om reklamens inverkan på konsumenternas beteende
P7_TA(2010)0484 . ,
– med beaktande av artikel 48 i arbetsordningen,
– med beaktande av betänkandet från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män och yttrandet från utskottet för sysselsättning och sociala frågor ( A7‑0029/2011 ), och av följande skäl:
A. Enligt fördraget om Europeiska unionen och Europeiska unionens stadga om de grundläggande rättigheterna är jämställdhet en av EU:s grundläggande principer, men det råder fortfarande stor brist jämställdhet.
B. EU har inte förskonats från den ekonomiska och finansiella krisen, som har visat sig vara förödande för både kvinnors och mäns sysselsättning, i synnerhet för kvinnors ekonomiska ställning, men som på lång sikt riskerar att påverka kvinnornas sysselsättning mer.
C. Jämställdhet har en positiv inverkan på produktiviteten och den ekonomiska tillväxten och ökar kvinnornas deltagande på arbetsmarknaden, vilket i sin tur ger många sociala och ekonomiska fördelar.
E. Arbetslöshetsnivån bland kvinnor underskattas ofta på grund av den stora andel kvinnor som inte förvärvsarbetar (två tredjedelar av 63 miljoner kvinnor mellan 25 och 64 år) eller är deltidsarbetslösa.
I. Moderskap borde inte utgöra ett hinder för kvinnors karriärmöjligheter, men statistiken visar tydligt att kvinnor som har barn ägnar färre timmar åt förvärvsarbete än kvinnor utan barn, i motsats till män som har barn, som förvärvsarbetar mer än män utan barn.
J. Vid Europeiska rådets möte i Barcelona i mars 2002 uppmanades medlemsstaterna att se till att det senast 2010 fanns barnomsorg för minst 90 procent av alla barn mellan tre år och den obligatoriska skolåldern och för minst 33 procent av alla barn under tre år, men i många länder saknas det fortfarande tillräcklig offentligfinansierad barnomsorg, vilket drabbar familjer som har det dåligt ställt extra hårt.
L. Tillgången till barnomsorg, äldreomsorg och omsorgstjänster för andra behövande personer är av grundläggande vikt för att lika många kvinnor som män ska arbeta och studera.
M. Ansvaret för hushållsarbetet vilar i betydligt högre grad på kvinnor än på män och värderas inte i ekonomiska termer eller i form av ett erkännande av dess värde, trots att omsorg i hemmet om barn, sjuka och äldre är ett svårt och obetalt arbete.
O. Antalet kvinnor och flickor som slår in på den naturvetenskapliga banan – särskilt matematik och IT – är fortfarande mycket lågt, vilket leder till en kraftig snedfördelning mellan kvinnor och män på detta område.
P. Krisen kan förvärra den sneda könsfördelningen ytterligare inom olika branscher och yrken, ett problem som ökar i stället för att minska i vissa länder.
R. Fler kvinnor än män tar universitetsexamen (58,9 procent av examina), men kvinnor har fortfarande i genomsnitt 18 procent lägre lön än männen och är underrepresenterade på de ledande befattningarna inom näringslivet, förvaltningen och politiken.
S. Det europeiska nätverk för kvinnor i beslutsfattande ställning inom politik och näringsliv som skapades i juni 2008 kan bidra till en mer jämnare könsfördelning på beslutsfattande nivå.
U. Positiva åtgärder till förmån för kvinnor har visat sig vara av grundläggande vikt för deras fullständiga deltagande på arbetsmarknaden och i samhället i stort.
W. Europaåret 2011 avser frivilligarbete och det är viktigt att betona den positiva inverkan som jämställdhetsprincipen kan ha på program för frivilligarbete.
X. Kvinnor som tillhör minoriteter, i synnerhet romska kvinnor, utsätts regelbundet för flerfaldig diskriminering på flera olika områden och missgynnas inte bara jämfört med kvinnor som tillhör majoritetsbefolkningen, utan även jämfört med män som tillhör etniska minoriteter, samt löper särskilt stor risk för att drabbas av utestängning.
Kvinnor utsätts för flera olika typer av diskriminering och löper större risk att drabbas av social utestängning, fattigdom och extrema människorättskränkningar, t.ex. människohandel, i synnerhet om de inte tillhör majoritetsbefolkningen.
Europaparlamentet uppmanar medlemsstaterna att med kommissionens stöd uppmuntra kvinnors deltagande i yrkesutbildning inom ramen för livslångt lärande genom att intensifiera redan befintliga åtgärder, mot bakgrund av omställningen till en hållbar ekonomi med fokus på små och medelstora företag, och därigenom öka kvinnliga arbetstagares anställbarhet.
Europaparlamentet uppmanar kommissionen att främja en dialog med arbetsmarknadens parter om frågor som insyn i lönesättningen och deltids- och visstidsavtal för kvinnor samt hur man ska uppmuntra kvinnor att arbeta inom gröna och innovativa branscher.
Europaparlamentet insisterar på att undanröjandet av löneklyftan är en prioriterad fråga och beklagar därför att kommissionen inte gjort tillräckligt för att återuppliva den europeiska debatten om detta, i synnerhet genom en översyn av den befintliga lagstiftningen om tillämpning av principen om lika lön för kvinnor och män, något som Europaparlamentet efterfrågade i sin resolution av den 18 november 2009.
Europaparlamentet uppmanar kommissionen att försäkra sig om att medlemsstaterna på ett korrekt sätt tillämpar de olika EU-bestämmelserna om möjligheterna att förena arbete och privatliv genom att anpassa arbetsförhållandena för kvinnor och män.
Europaparlamentet uppmanar offentliga och privata organ att införa jämställdhetsplaner i sina interna bestämmelser, att förse dem med strikta målsättningar på kort, medellång och lång sikt och att göra årliga utvärderingar av hur målsättningarna har förverkligats.
Europaparlamentet understryker att ungdomar måste få välja yrkesbana fritt och påpekar därför vikten av att lärarna inte automatiskt leder in sina elever på yrkesbanor utifrån könsstereotyper och att alla möjliga yrkesbanor framhålls.
Europaparlamentet påpekar att medlemsstaterna måste vidta åtgärder, särskilt genom lagstiftning, för att fastställa bindande mål om en jämn könsfördelning på högre befattningar inom näringslivet, den offentliga förvaltningen och politiken.
Europaparlamentet välkomnar den allmänna debatten om att öka andelen kvinnor med ledande befattningar i näringslivet och uppmanar företagen att på frivillig basis införa en kvot för detta, på grundval av könsfördelningen bland personalen.
Europaparlamentet betonar vikten av att medlemsstaterna och de regionala och lokala myndigheterna vidtar åtgärder för att med hjälp av instrument som Europeiska socialfonden (ESF) eller programmet Progress göra det lättare för kvinnor som utsatts för könsrelaterat våld att komma tillbaka in på arbetsmarknaden.
MOTIVERING
Den rådande finansiella, ekonomiska och sociala krisen har en katastrofal inverkan på arbetslösheten, medborgarnas levnadsvillkor och samhället i allmänhet.
I sin årliga rapport från 2010 anger kommissionen med rätta de utmaningar som väntar i krisens kölvatten när det gäller jämställdhet.
Föredraganden understryker att man måste ringa in de verkliga följderna av krisen för kvinnor.
Detta gäller framför allt kvinnors sysselsättning.
Kvinnorna har i detta sammanhang generellt sett drabbats senare än män på grund av att de främst är sysselsatta inom sektorer som har stått emot effekterna av krisen längre (vård, skola, omsorg osv.).
Det finns dock risk för att dessa sektorer drabbas mer varaktigt, vilket skulle göra kvinnornas sysselsättning mer långvarigt osäker än männens.
Vare sig det gäller arbets- och anställningsvillkor eller tillträde till arbetsmarknaden har kvinnorna således drabbats hårt, och om konkreta åtgärder inte vidtas omgående riskerar deras situation att förvärras ytterligare.
Kvinnor missgynnas i hög grad på arbetsmarknaden eftersom de är förpassade till deltidsanställningar och tidsbegränsade anställningar, ofta med otillräckliga löner.
Jämställdhet i arbetslivet borde inte längre vara bara något som eftersträvas, utan måste bli verklighet.
Därför är det viktigt att medlemsstaternas regeringar och kommissionen upprätthåller jämställdhetspolitiken och sörjer för att de avsatta medlen inte minskar.
Krisen får dock inte enbart uppfattas som något negativt.
Den måste ses som ett tillfälle för makthavarna att ställa de rätta frågorna och betrakta sin egen politik ur en ny synvinkel.
Mot bakgrund av krisen måste vi ompröva mäns och kvinnors respektive roller i samhället, bland annat via en fullständig jämställdhetsintegrering på alla politikområden.
Detta jämställdhetsideal bör uppnås genom konkreta och varaktiga åtgärder, i synnerhet inom utbildningen.
För att förhindra att könsstereotyper består måste barn tidigt lära sig om principen om jämställdhet.
Utbildning av unga utgör nyckeln till jämställdhet, oavsett om det sker via kontinuerlig information, informationskampanjer eller vägledning för att orientera pojkar och flickor mot andra yrken än traditionella mans- eller kvinnoyrken.
Föredraganden framhåller vikten av kvinnor i beslutsfattande ställning – en traditionellt manlig miljö.
Kvinnor måste få tillgång till befattningar som motsvarar deras kompetens, oavsett om det rör sig om de börsnoterade bolagens styrelser eller deras representation i politiken.
Trots att de ofta har högre kvalifikationer nekas kvinnor ibland tillträde till ledande ansvarstunga poster, vilket skapar en förskjutning mellan deras utbildningsnivå och deras ställning.
Det är också viktigt att stärka jämställdhetsperspektivet inom fattigdomsbekämpningen.
De mest utsatta grupperna av kvinnor borde ägnas särskild uppmärksamhet under Europaåret för bekämpning av fattigdom 2010.
Det bör vidtas åtgärder för att förhindra att kvinnor som är utsatta på grund av de är funktionshindrade, invandrare eller tillhör en minoritet hamnar i en osäker situation samt för att underlätta deras integration i samhället.
Föredraganden rekommenderar därför kommissionen att inom ramen för EU:s strategi för integration av romerna ägna betydande insatser åt integration av romska kvinnor.
Jämställdhet främjas även genom bekämpning av våld mot kvinnor.
Alla typer av fysiskt, psykologiskt och sexuellt våld, oavsett hur grovt det är, måste bekämpas och fördömas.
I bekämpningen av könsrelaterat våld ingår att man genomför informationskampanjer och undervisar barn och ungdomar om hur avskyvärt detta våld är.
Att fördöma könsrelaterat våld innebär att man måste definiera det ur juridisk synvinkel och föreskriva straff som står i proportion till brottet.
Till exempel syraattacker en typ av våld som dessvärre fortfarande förekommer i vissa medlemsstater.
Det finns fortfarande tabun i våra samhällen när det gäller vissa typer av våld mot kvinnor.
YTTRANDE från utskottet för sysselsättning och sociala frågor
till utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
över jämställdhet mellan kvinnor och män i Europeiska unionen – 2010
( 2010/2138(INI) )
Föredragande: Nadja Hirsch
FÖRSLAG
Utskottet för sysselsättning och sociala frågor uppmanar utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet uppmanar kommissionen att uppdatera jämställdhetsindikatorerna, utöka dem med kriteriet civilstånd och tillämpa indikatorerna för att regelbundet bedöma ojämlikheter mellan kvinnor och män.
Europaparlamentet välkomnar meddelandet ”Strategi för jämställdhet 2010–2015” som antogs av kommissionen den 21 september 2010.
Europaparlamentet betonar att tillvaratagandet av den kvinnliga arbetskraftens potential även är i linje med Europa 2020-strategins mål om minskad fattigdom samt att tillgång till sysselsättning utgör en hörnsten i ansträngningarna för att bekämpa fattigdom.
Europaparlamentet uppmanar medlemsstaterna att med kommissionens stöd och genom att intensifiera redan befintliga åtgärder uppmuntra kvinnors deltagande i yrkesutbildning inom ramen för livslångt lärande, mot bakgrund av omställningen till en hållbar ekonomi med fokus på små och medelstora företag, och därigenom öka kvinnliga arbetstagares anställbarhet.
Europaparlamentet uppmanar medlemsstaterna att stödja sysselsättningen för ”gravida kvinnor och mödrar med ensamt ansvar för familjen”, som är en missgynnad grupp, och underlätta dessa kvinnors tillgång till ett värdigt och fast arbete så att de ska kunna förena familj och arbete.
Europaparlamentet uppmanar kommissionen att främja en dialog med arbetsmarknadens parter för att granska frågor som insyn i lönesättningen och deltids- och visstidsavtal för kvinnor samt hur man ska uppmuntra kvinnor att delta i gröna och innovativa branscher.
Europaparlamentet understryker vikten av förhandlingar och kollektivavtal för att bekämpa diskriminering av kvinnor, särskilt i fråga om sysselsättning, lön, arbetsvillkor, karriärmöjligheter och utbildning.
Europaparlamentet välkomnar den allmänna debatten om att öka andelen kvinnor med ledande befattningar i näringslivet och uppmanar företagen att på frivillig basis införa en kvot på grundval av könsfördelningen bland personalen.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
25.1.2011
Slutomröstning: resultat
+:
–:
0:
40
1
2
Slutomröstning: närvarande ledamöter
Regina Bastos, Edit Bauer, Jean-Luc Bennahmias, Pervenche Berès, Philippe Boulland, Alejandro Cercas, Ole Christensen, Marije Cornelissen, Tadeusz Cymański, Frédéric Daerden, Karima Delli, Proinsias De Rossa, Frank Engel, Sari Essayah, Richard Falbr, Ilda Figueiredo, Nadja Hirsch, Stephen Hughes, Danuta Jazłowiecka, Martin Kastler, Ádám Kósa, Jean Lambert, Veronica Lope Fontagné, Olle Ludvigsson, Elizabeth Lynne, Thomas Mann, Elisabeth Morin-Chartier, Csaba Őry, Siiri Oviir, Rovana Plumb, Konstantinos Poupakis, Licia Ronzulli, Elisabeth Schroedter, Joanna Katarzyna Skrzydlewska, Jutta Steinruck, Traian Ungureanu
Slutomröstning: närvarande suppleanter
Raffaele Baldassarre, Kinga Göncz, Richard Howitt, Jan Kozłowski, Gesine Meissner, Cecilia Wikström
Slutomröstning: närvarande suppleanter (art.
187.2)
Claudio Morganti
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
27.1.2011
Slutomröstning: resultat
+:
–:
0:
22
2
Slutomröstning: närvarande ledamöter
Regina Bastos, Edit Bauer, Emine Bozkurt, Andrea Češková, Marije Cornelissen, Edite Estrela, Ilda Figueiredo, Teresa Jiménez-Becerril Barrio, Nicole Kiil-Nielsen, Rodi Kratsa-Tsagaropoulou, Siiri Oviir, Raül Romeva i Rueda, Joanna Katarzyna Skrzydlewska, Marc Tarabella, Britta Thomsen, Marina Yannakoudakis
Slutomröstning: närvarande suppleanter
Anne Delvaux, Christa Klaß, Mariya Nedelcheva, Norica Nicolai, Antigoni Papadopoulou, Rovana Plumb, Joanna Senyszyn
Slutomröstning: närvarande suppleanter (art.
187.2)
Stanimir Ilchev
A7-0074/2011
BETÄNKANDE
om grönboken om bolagsstyrning i finansinstitut
(2010/2303(INI))
Utskottet för ekonomi och valutafrågor
Föredragande: Ashley Fox
Rådgivande utskotts föredragande (*): Alexandra Thein, utskottet för rättsliga frågor
(*) Förfarande med associerat utskott – artikel 50 i arbetsordningen
PE 454.525v05-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
YTTRANDE från utskottet för rättsliga frågor ...........................................11
YTTRANDE från utskottet för den inre marknaden och konsumentskydd 17
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................21
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om grönboken om bolagsstyrning i finansinstitut
( 2010/2303(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av artikel 48 i arbetsordningen,
– med beaktande av Europaparlamentets och rådets direktiv 2010/76/EU av den 24 november 2010 om ändring av direktiv 2006/48/EG och 2006/49/EG i fråga om kapitalkrav för handelslager och omvärdepapperisering samt samlad tillsynsbedömning av ersättningspolitik
EUT L 329, 14.12.2010, s.
3. ,
– med beaktande av betänkandet från utskottet för ekonomi och valutafrågor och yttrandena från utskottet för rättsliga frågor och utskottet för den inre marknaden och konsumentskydd ( A7‑0074/2011 ).
Tillvägagångssätt
1.
Risk
Europaparlamentet betonar att det yttersta ansvaret för riskstyrning ligger hos styrelsen, som också måste ta ansvaret för att uppvisa regelefterlevnad och för att upprätta återhämtningsplaner.
Europaparlamentet påpekar att systemet för kommunikation mellan riskhanteringsfunktioner och styrelsen bör förbättras genom att inrätta ett förfarande för att hänföra konflikter och problem till rätt nivå i hierarkin så att de kan lösas.
Europaparlamentet föreslår också att det bör upprättas förfaranden för att protokollföra situationer då riskkommitténs synpunkter inte beaktas och att dessa protokoll överlämnas till revisorer och tillsynsmyndigheter.
Europaparlamentet anser att mer uppmärksamhet bör fästas vid genomförande av åtgärder som höjer riskmedvetandet i finansinstitut, eftersom ett stärkt riskmedvetande på alla nivåer i företaget – också bland de anställda – är avgörande för en bättre riskhantering.
Styrelser
34.
Europaparlamentet betonar att företagsledningen och ersättningspolicyn måste respektera och främja den princip om lika löner och lika behandling av kvinnor och män som är fastslagen genom fördragen och EU:s direktiv.
Ersättning
Europaparlamentet noterar att frågan om ersättning i finansinstitut har behandlats inom ramen för den tredje översynen av kapitalkravsdirektivet (CRD III).
Europaparlamentet anser att aktieägarna bör bidra till att bestämma en hållbar ersättningspolicy och bör ges möjlighet att uttrycka sina synpunkter om ersättningspolicyn, med rätt att avvisa den ersättningspolicy som ersättningskommittén har föreslagit vid bolagsstämman.
Tillsynsmyndigheter, revisorer och institut
Europaparlamentet betonar att offentliga myndigheter, inbegripet de europeiska tillsynsmyndigheterna och nationella tillsynsmyndigheter, måste uppfylla höga standarder för oberoende och för bolagsstyrning.
Europaparlamentet uppmanar institutionella aktieägare att inta en aktivare roll när det gäller att ställa styrelsen till svars och få den att på ett lämpligt sätt förklara sin strategi i syfte att återspegla förmånstagarnas långsiktiga intressen.
65.
till utskottet för ekonomi och valutafrågor
över bolagsstyrning i finansinstitut och ersättningspolicy
( 2010/2303(INI) )
Rådgivande utskotts föredragande (*): Alexandra Thein
(*) Förfarande med associerat utskott – artikel 50 i arbetsordningen
KORTFATTAD MOTIVERING
Bakgrund
Denna grönbok syftar till att dra lärdomar av den globala finanskrisen som utlöstes genom banken Lehman Brothers konkurs hösten 2008 efter en orimlig värdepapperisering av amerikanska subprime-bolån.
Inte minst med tanke på de nya finansiella instrumenten i en globaliserad värld görs nu en kritisk granskning av soliditeten i finansinstituten och hela finanssystemet liksom av regleringen av och tillsynen över dessa så att en upprepning av en sådan situation ska kunna undvikas i framtiden.
En förstärkning av bolagsstyrningen ses av kommissionen som kärnpunkten i dess program för finansmarknadsreform och krisförebyggande.
Kommissionen konstaterar i synnerhet att bolagsstyrningen i finanstjänstesektorn, på grund av många aktörers systemvikt, måste ta hänsyn till andra intressenter (insättare, sparare, livförsäkringsinnehavare, osv.) och finanssystemets stabilitet.
De förslag som tas upp i grönboken bör stödja och komplettera de rättsliga arrangemang som införts eller planterats för att konsolidera finanssystemet, särskilt inom ramen för den europeiska tillsynsstrukturen, kapitalkravsdirektivet (CRD III), Solvens II-direktivet för försäkringsbolag, översynen av företag för kollektiva investeringar i överlåtbara värdepapper (UCITS) och bestämmelserna för förvaltare av alternativa investeringsfonder (AIF‑förvaltare).
Grönboken fokuserar på en snäv definition av bolagsstyrning där också externa revisorers roll ingår.
Andra viktiga aspekter av bolagsstyrningen – t.ex. separation av olika funktioner inom finansföretag, de interna kontrollernas funktion och redovisningens oberoende – behandlas inte i grönboken.
Föredragandens ståndpunkter
Att ta finansiella risker är en central uppgift för finansbranschen och nödvändig för att den ska lyckas i sina affärer och för att den ska fylla sina funktioner för ekonomin som helhet.
Det ligger i allmänhetens intresse att man inte inkräktar på dessa funktioner mer än vad som krävs för att förhindra systemkriser.
Det bör också i detta sammanhang förtydligas att finansinstitut måste kunna försättas i konkurs på ett kontrollerat sätt så länge detta inte skulle innebära någon systemrisk och det genom de finansiella sammankopplingarna inte skulle kunna leda till dominoeffekter på marknaden.
Föredraganden ser det som en grundläggande och avgörande fråga att mer än tidigare utveckla en ordning och en kultur av hållbar och fullt ut ansvarstagande riskhantering i finansinstituten liksom en övervakning av detta.
Denna lika viktiga som komplexa utmaning bör mötas med en uppsättning direkta eller indirekta åtgärder.
Många sådana åtgärder vidtogs redan förra året på EU- eller medlemsstatsnivå, särskilt när det gäller ersättning till ledande personer.
Vetenskapliga studier visar att inte minst åtgärder som syftar till att professionalisera styrelser och öka mångfalden i dessa utifrån ett antal kriterier verkar vara välmotiverat och lovande.
Hur styrelseledamöternas ansvar och förpliktelser utformas måste visserligen definieras klart, men rent konkret också hanteras med stor urskillning så att man inte äventyrar finansinstitutens vilja att ta affärschanser, vilket är en positiv aspekt av deras verksamhet, eller kvaliteten på de personer som står till förfogande.
En annan central uppgift är enligt föredraganden är att eliminera eller åtminstone minska den roll som intressekonflikter spelar för finansiella kriser.
När det gäller konflikterna mellan traditionell bankverksamhet i form av kreditgivning och investmentbanktjänster inom finansinstitut förefaller en tvingande lag som föreskriver att ett visst finansinstitut endast får fylla en av dessa båda funktioner vara en tänkvärd möjlighet, men med tanke på möjliga effektivitetsförluster och den europeiska finansbranschens globala konkurrenskraft är den knappast värd att genomföra.
Kompromisslösa åtgärder är däremot påkallade för att utesluta intressekonflikter hos personer som spelar en avgörande roll vid övervakningen av risker, framför allt styrelseledamöter.
Den brittiska ”Stewardship Code” skulle kunna fungera som förebild för en enhetlig EU-kod för institutionella investerare.
FÖRSLAG
Utskottet för rättsliga frågor uppmanar utskottet för ekonomi och valutafrågor att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet betonar hur viktigt det är med arbetstagarföreträdare i styrelserna, särskilt på grund av deras långsiktiga intresse av en hållbar företagsledning liksom deras erfarenhet och kunskaper om företagets interna struktur.
Europaparlamentet anser att om det skulle vara obligatoriskt för en eller flera ledamöter av revisionskommittén att vara ledamöter av riskkommittén och vice versa, skulle detta kunna leda till att kompetensen splittras och förmågan att fokusera på ett enda uppdrag går förlorad.
Europaparlamentet noterar att ordföranden för riskkommittén bör rapportera till bolagsstämman, eller att han eller hon under inga omständigheter ska kunna avsättas av den verkställande ledningen eller styrelsen.
Europaparlamentet anser att mer uppmärksamhet bör fästas vid genomförande av åtgärder som höjer riskmedvetandet i finansinstitut, eftersom ett stärkt riskmedvetande på alla nivåer i företaget – också bland de anställda – är avgörande för en bättre riskhantering.
Europaparlamentet påpekar att systemet för kommunikation mellan riskhanteringsfunktioner och styrelsen bör förbättras genom att inrätta ett förfarande för att hänföra konflikter och problem till rätt nivå i hierarkin så att de kan lösas.
Europaparlamentet anser att det är nödvändigt med en klart definierad europeisk minimistandard för det ansvar som ledamöter i finansinstituts styrelser bär.
23.
Europaparlamentet betonar att det är nödvändigt med fullständig transparens för att aktieägare ska kunna få en fullständig uppsikt över ersättningspolicyn, vilket bland annat innebär att antalet anställda som erhåller mer än 500 000 EUR, i intervaller på 500 000 EUR, bör offentliggöras.
Europaparlamentet anser att det är nödvändigt, med beaktande av dagens olika rättsliga och ekonomiska modeller, att harmonisera det övergripande innehållet och de närmare uppgifterna i gemenskapens regler för intressekonflikter så att olika finansinstitut blir föremål för liknande regler, i enlighet med vilka de måste tillämpa reglerna i MiFID, kapitalkravsdirektivet (CRD), UCITS-direktivet eller Solvens II-direktivet.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
28.2.2011
Slutomröstning: resultat
+:
–:
0:
19
Slutomröstning: närvarande ledamöter
Raffaele Baldassarre, Sebastian Valentin Bodu, Françoise Castex, Christian Engström, Klaus-Heiner Lehne, Antonio Masip Hidalgo, Alajos Mészáros, Bernhard Rapkay, Evelyn Regner, Francesco Enrico Speroni, Alexandra Thein, Cecilia Wikström, Zbigniew Ziobro, Tadeusz Zwiefka
Slutomröstning: närvarande suppleanter
Piotr Borys, Sergio Gaetano Cofferati, Sajjad Karim, Eva Lichtenberger, Toine Manders
till utskottet för ekonomi och valutafrågor
över bolagsstyrning i finansiella institut
( 2010/2303(INI) )
Föredragande:
Othmar Karas
FÖRSLAG
Utskottet för den inre marknaden och konsumentskydd uppmanar utskottet för ekonomi och valutafrågor att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet är medvetet om att det efter finanskrisen står klart att det behövs påtagliga och betydande förbättringar av konsumentskyddets kvalitet och av garantierna på området för finansiella tjänster, särskilt i fråga om kontroll och tillsyn.
Europaparlamentet anser att finanssektorn måste rätta sig efter realekonomins behov, bidra till en hållbar utveckling och ta största möjliga samhällsansvar.
Parlamentet betonar att företagsledningen och ersättningspolicyn måste respektera och främja den princip om lika löner och lika behandling av kvinnor och män som är fastslagen genom fördragen och EU:s direktiv.
Europaparlamentet anser att både företagsledning och styrelse bör hållas rättsligt ansvariga, de facto och personligen, för att bolagsstyrningsprinciperna upprättas och genomförs korrekt på alla nivåer inom företaget och koncernen.
Direktiv 2010/76/EU (EUT L 329, 14.12.2010, s.
3). och Solvens II, och förväntar sig att denna liksom andra lagstiftningsåtgärder som redan vidtagits snabbt ska genomföras från och med januari 2011.
EUT L 294, 10.11.2001, s.
22. om komplettering av stadgan för europabolag ska genomföras effektivt.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
28.2.2011
Slutomröstning: resultat
+:
–:
0:
30
Slutomröstning: närvarande ledamöter
Pablo Arias Echeverría, Cristian Silviu Buşoi, Anna Maria Corazza Bildt, António Fernando Correia De Campos, Jürgen Creutzmann, Christian Engström, Louis Grech, Małgorzata Handzlik, Philippe Juvin, Eija-Riitta Korhola, Mitro Repo, Robert Rochefort, Zuzana Roithová, Heide Rühle, Christel Schaldemose, Andreas Schwab, Catherine Stihler, Kyriacos Triantaphyllides, Bernadette Vergnaud, Barbara Weiler
Slutomröstning: närvarande suppleanter
Damien Abad, Cornelis de Jong, María Irigoyen Pérez, Constance Le Grip, Emma McClarkin, Antonyia Parvanova, Konstantinos Poupakis, Sylvana Rapti, Olga Sehnalová, Wim van de Camp
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
16.3.2011
Slutomröstning: resultat
+:
–:
0:
37
3
2
Slutomröstning: närvarande ledamöter
Burkhard Balz, Sharon Bowles, Udo Bullmann, Pascal Canfin, Nikolaos Chountis, George Sabin Cutaş, Rachida Dati, Leonardo Domenici, Derk Jan Eppink, Diogo Feio, Vicky Ford, Ildikó Gáll-Pelcz, José Manuel García-Margallo y Marfil, Jean-Paul Gauzès, Sven Giegold, Sylvie Goulard, Liem Hoang Ngoc, Wolf Klinz, Philippe Lamberts, Astrid Lulling, Hans-Peter Martin, Íñigo Méndez de Vigo, Ivari Padar, Antolín Sánchez Presedo, Olle Schmidt, Edward Scicluna, Peter Simon, Peter Skinner, Theodor Dumitru Stolojan, Ivo Strejček, Marianne Thyssen, Corien Wortmann-Kool
Slutomröstning: närvarande suppleanter
Sophie Auconie, Elena Băsescu, Saïd El Khadraoui, Ashley Fox, Danuta Jazłowiecka, Olle Ludvigsson, Thomas Mann, Miguel Portas, Catherine Stihler
Slutomröstning: närvarande suppleanter (art.
187.2)
David Campbell Bannerman
A7-0116/2011
BETÄNKANDE
om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2009, avsnitt VIII – Europeiska ombudsmannen
(C7‑0218/2010 – 2010/2149(DEC))
Budgetkontrollutskottet
Föredragande: Crescenzio Rivellini
PE 450.686v02-00
INNEHÅLL
1.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT.......................................................3
2.
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.............................................4
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.......................................................6
1.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2009, avsnitt VIII – Europeiska ombudsmannen
( C7‑0218/2010 – 2010/2149(DEC) )
Europaparlamentet fattar detta beslut
EUT L 69, 13.3.2009. ,
– med beaktande av Europeiska unionens slutliga årsredovisning för budgetåret 2009 ( SEK(2010)0963 – C7-0218/2010 )
EUT C 308, 12.11.2010, s.
1. ,
– med beaktande av Europeiska ombudsmannens årsrapport om de internrevisioner som genomförts under 2009,
– med beaktande av revisionsrättens årsrapport om genomförandet av budgeten för budgetåret 2009, samt de granskade institutionernas svar
EUT C 303, 9.11.2010, s.
1. ,
– med beaktande av förklaringen om räkenskapernas tillförlitlighet och de underliggande transaktionernas laglighet och korrekthet som avges av revisionsrätten i enlighet med artikel 287 i fördraget om Europeiska unionens funktionssätt
129. ,
– med beaktande av artiklarna 272.10, 274, 275 och 276 i EG-fördraget och artiklarna 314.10, 317, 318 och 319 i fördraget om Europeiska unionens funktionssätt,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1. , särskilt artiklarna 50, 86, 145, 146 och 147,
– med beaktande av artikel 77 och bilaga VI i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet ( A7‑0116/2011 ) och av följande skäl:
2.
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2009, avsnitt VIII – Europeiska ombudsmannen
( C7‑0218/2010 – 2010/2149(DEC) )
Europaparlamentet utfärdar denna resolution
EUT L 69, 13.3.2009. ,
– med beaktande av Europeiska unionen slutliga årsredovisning för budgetåret 2009 ( SEK(2010)0963 – C7-0218/2010 )
EUT C 308, 12.11.2010, s.
1. ,
– med beaktande av Europeiska ombudsmannens årsrapport om de internrevisioner som genomförts under 2009,
– med beaktande av revisionsrättens årsrapport om genomförandet av budgeten för budgetåret 2009, samt de granskade institutionernas svar
EUT C 303, 9.11.2010, s.
1. ,
– med beaktande av förklaringen om räkenskapernas tillförlitlighet och de underliggande transaktionernas laglighet och korrekthet som avges av revisionsrätten i enlighet med artikel 287 i fördraget om Europeiska unionens funktionssätt
129. ,
– med beaktande av artiklarna 272.10, 274, 275 och 276 i EG-fördraget och artiklarna 314.10, 317, 318 och 319 i fördraget om Europeiska unionens funktionssätt,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1. , särskilt artiklarna 50, 86, 145, 146 och 147,
– med beaktande av artikel 77 och bilaga VI i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet ( A7‑0116/2011 ), och av följande skäl:
4.
Europaparlamentet noterar att revisionsrätten i sin årsrapport angav att granskningen inte föranledde några ytterligare stora anmärkningar när det gäller ombudsmannen.
Europaparlamentet konstaterar att ombudsmannens kansli omorganiserades den 1 januari 2010, och uppmanar ombudsmannen att rapportera om effekten av dessa förändringar i den årliga verksamhetsrapporten.
Europaparlamentet välkomnar genomförandet av centrala resultatindikatorer i den årliga förvaltningsplanen, och att målen för 2009 uppnåtts.
10.
11.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
22.3.2011
Slutomröstning: resultat
+:
–:
0:
19
1
Slutomröstning: närvarande ledamöter
Marta Andreasen, Jean-Pierre Audy, Inés Ayala Sender, Zigmantas Balčytis, Andrea Češková, Andrea Cozzolino, Luigi de Magistris, Tamás Deutsch, Martin Ehrenhauser, Jens Geier, Gerben-Jan Gerbrandy, Ingeborg Gräßle, Ville Itälä, Iliana Ivanova, Bogusław Liberadzki, Monica Luisa Macovei, Jan Olbrycht, Aldo Patriciello, Crescenzio Rivellini, Christel Schaldemose, Bart Staes, Georgios Stavrakakis, Søren Bo Søndergaard
Slutomröstning: närvarande suppleanter
Chris Davies, Derk Jan Eppink, Christofer Fjellner, Véronique Mathieu
A7-0127/2011
BETÄNKANDE
om ansvarsfrihet för genomförandet av budgeten för Europeiska kemikaliemyndigheten för budgetåret 2009
(C7‑0245/2009 – 2010/2185(DEC))
Budgetkontrollutskottet
Föredragande: Georgios Stavrakakis
PE 450.710v02-00
INNEHÅLL
1.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT.......................................................3
2.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT.......................................................5
3.
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.............................................6
YTTRANDE från utskottet för miljö, folkhälsa och livsmedelssäkerhet 10
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................13
1.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
om ansvarsfrihet för genomförandet av budgeten för Europeiska kemikaliemyndigheten för budgetåret 2009
( C7‑0245/2009 – 2010/2185(DEC) )
Europaparlamentet fattar detta beslut
– med beaktande av den slutliga årsredovisningen för Europeiska kemikaliemyndigheten för budgetåret 2009,
– med beaktande av revisionsrättens rapport om årsredovisningen för Europeiska kemikaliemyndigheten för budgetåret 2009, samt myndighetens svar
EUT C 338, 14.12.2010, s.
34. ,
– med beaktande av rådets rekommendation av den 15 februari 2011 (5892/2011 – C7‑0052/2011 ),
– med beaktande av artikel 276 i EG-fördraget och artikel 319 i fördraget om Europeiska unionens funktionssätt,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1. , särskilt artikel 185,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 om inrättande av en europeisk kemikaliemyndighet
EUT L 396, 30.12.2006, s.
1. , särskilt artikel 97,
– med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002
EGT L 357, 31.12.2002, s.
72. av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002, särskilt artikel 94,
– med beaktande av artikel 77 och bilaga VI i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A7‑0127/2011 ).
2.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
om avslutande av räkenskaperna för Europeiska kemikaliemyndigheten för budgetåret 2009
( C7‑0245/2009 – 2010/2185(DEC) )
Europaparlamentet fattar detta beslut
– med beaktande av den slutliga årsredovisningen för Europeiska kemikaliemyndigheten för budgetåret 2009,
– med beaktande av revisionsrättens rapport om årsredovisningen för Europeiska kemikaliemyndigheten för budgetåret 2009, samt myndighetens svar
EUT C 338, 14.12.2010, s.
34. ,
– med beaktande av rådets rekommendation av den 15 februari 2011 (5892/2011 – C7‑0052/2011 ),
– med beaktande av artikel 276 i EG-fördraget och artikel 319 i fördraget om Europeiska unionens funktionssätt,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1. , särskilt artikel 185,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 om inrättande av en europeisk kemikaliemyndighet
EUT L 396, 30.12.2006, s.
1. , särskilt artikel 97,
– med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002
EGT L 357, 31.12.2002, s.
72. , särskilt artikel 94,
– med beaktande av artikel 77 och bilaga VI i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A7‑0127/2011 ).
3.
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska kemikaliemyndigheten för budgetåret 2009
( C7‑0245/2009 – 2010/2185(DEC) )
Europaparlamentet utfärdar denna resolution
– med beaktande av den slutliga årsredovisningen för Europeiska kemikaliemyndigheten för budgetåret 2009,
– med beaktande av revisionsrättens rapport om årsredovisningen för Europeiska kemikaliemyndigheten för budgetåret 2009, samt myndighetens svar
EUT C 338, 14.12.2010, s.
34. ,
– med beaktande av rådets rekommendation av den 15 februari 2011 (5892/2011 – C7‑0052/2011 ),
– med beaktande av artikel 276 i EG-fördraget och artikel 319 i fördraget om Europeiska unionens funktionssätt,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1. , särskilt artikel 185,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 om inrättande av en europeisk kemikaliemyndighet
EUT L 396, 30.12.2006, s.
1. , särskilt artikel 97,
– med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002
EGT L 357, 31.12.2002, s.
72. av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002, särskilt artikel 94,
– med beaktande av artikel 77 och bilaga VI i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A7‑0127/2011 ).
A. Revisionsrätten har förklarat att den har uppnått en rimlig säkerhet om att räkenskaperna för budgetåret 2009 är tillförlitliga och att de underliggande transaktionerna är lagliga och korrekta.
B. År 2009 var myndighetens andra verksamhetsår.
C. Den 5 maj 2010 beviljade Europaparlamentet den verkställande direktören för Europeiska kemikaliemyndigheten ansvarsfrihet för genomförandet av myndighetens budget för budgetåret 2008
EUT L 252, 25.9.2010, s.
146. , och i sin resolution som åtföljde beslutet om ansvarsfrihet framförde parlamentet bland annat följande synpunkter:
– Europaparlamentet påpekar att revisionsrätten har konstaterat förseningar i driften på grund av problem med införandet av IT-systemet och bristen på kvalificerad personal.
– Europaparlamentet uttrycker sin tillfredsställelse över myndighetens första framgångsrika självständiga verksamhetsår, eftersom kommissionen (GD Näringsliv) ansvarade för myndighetens budgetförvaltning 2007.
Europaparlamentet noterar att myndigheten 2008 finansierades genom ett bidrag från gemenskapen på 62 200 000 EUR i enlighet med artikel 185 i den allmänna budgetförordningen och i mindre utsträckning av avgifter som industrin erlägger vid registrering av kemikalier i enlighet med Reach-förordningen (Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 om registrering, utvärdering, godkännande och begränsning av kemikalier (Reach), och om inrättande av en europeisk kemikaliemyndighet
EUT L 396, 30.12.2006, s.
1. ).
Europaparlamentet konstaterar att ökningen under avdelning III (driftsutgifter) främst är ett resultat av ökade kostnader för programvaruutveckling, eftersom stora investeringar har krävts för att förbättra IT-systemet för Reach och för ytterligare utveckling av ett omfattande verktyg för kemikaliesäkerhetsbedömning/kemikaliesäkerhetsrapport.
Verksamhetsresultat
Överföring av anslag mellan budgetår
Internrevision
Europaparlamentet uppmanar myndigheten att informera den ansvarsfrihetsbeviljande myndigheten om de steg som vidtagits för att förbättra dess kontrollsystem genom att stärka dess finansiella rutiner, arbetsflöde, granskningar, handlingsplaner och riskbedömningar.
– alla delar i finansieringsbesluten finns på plats (t.ex. standardformat för myndighetens program och finansiella beslut),
– den information som krävs på varje nivå inom organisationen är tillbörligt fastställd och hanterad,
– programmet visar samtliga resurser som görs tillgängliga genom budgeten, samt att
– dokumentationen över de finansiella förfarandena och checklistorna slutförs och uppdateras.
o
o o
16.
När det gäller övriga övergripande iakttagelser som utgör en del av beslutet om ansvarsfrihet hänvisar Europaparlamentet till sin resolution av den … maj 2011
Antagna texter, P7_TA-PROV(2011). om byråernas verksamhetsresultat, ekonomiska förvaltning och kontroll.
till budgetkontrollutskottet
över ansvarsfrihet för genomförandet av Europeiska kemikaliemyndighetens budget för budgetåret 2009
( C7-0245/2010 – 2010/2185(DEC) )
Föredragande: Jutta Haug
FÖRSLAG
EUT L 396, 30.12.2006, s.
Europaparlamentet konstaterar att ökningen under avdelning III (driftsutgifter) främst beror på ökade kostnader för programvaruutveckling, eftersom stora investeringar har krävts för att förbättra IT-systemet för Reach och för ytterligare utveckling av ett omfattande verktyg för kemikaliesäkerhetsbedömning/kemikaliesäkerhetsrapport.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
16.3.2011
Slutomröstning: resultat
+:
–:
0:
49
7
Slutomröstning: närvarande ledamöter
János Áder, Kriton Arsenis, Pilar Ayuso, Paolo Bartolozzi, Sandrine Bélier, Sergio Berlato, Martin Callanan, Nessa Childers, Chris Davies, Bairbre de Brún, Bas Eickhout, Edite Estrela, Karl-Heinz Florenz, Elisabetta Gardini, Julie Girling, Cristina Gutiérrez-Cortines, Satu Hassi, Jolanta Emilia Hibner, Dan Jørgensen, Karin Kadenbach, Christa Klaß, Holger Krahmer, Jo Leinen, Corinne Lepage, Linda McAvan, Radvilė Morkūnaitė-Mikulėnienė, Miroslav Ouzký, Vladko Todorov Panayotov, Gilles Pargneaux, Antonyia Parvanova, Andres Perello Rodriguez, Sirpa Pietikäinen, Mario Pirillo, Pavel Poc, Vittorio Prodi, Frédérique Ries, Anna Rosbach, Oreste Rossi, Dagmar Roth-Behrendt, Daciana Octavia Sârbu, Horst Schnellhardt, Richard Seeber, Theodoros Skylakakis, Bogusław Sonik, Salvatore Tatarella, Åsa Westlund, Glenis Willmott, Sabine Wils, Marina Yannakoudakis
Slutomröstning: närvarande suppleanter
Jutta Haug, Marisa Matias, Bill Newton Dunn, Bart Staes, Eleni Theocharous, Thomas Ulmer, Anna Záborská
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
21.3.2011
Slutomröstning: resultat
+:
–:
0:
16
2
Slutomröstning: närvarande ledamöter
Marta Andreasen, Jean-Pierre Audy, Inés Ayala Sender, Jorgo Chatzimarkakis, Tamás Deutsch, Martin Ehrenhauser, Jens Geier, Ingeborg Gräßle, Iliana Ivanova, Elisabeth Köstinger, Monica Luisa Macovei, Aldo Patriciello, Crescenzio Rivellini, Bart Staes, Georgios Stavrakakis, Søren Bo Søndergaard
Slutomröstning: närvarande suppleanter
A7-0131/2011
BETÄNKANDE
om ansvarsfrihet för genomförandet av budgeten för det europeiska gemensamma företaget för ITER och utveckling av fusionsenergi för budgetåret 2009
(C7‑0247/2010 – 2010/2187(DEC))
Budgetkontrollutskottet
Föredragande: Georgios Stavrakakis
PE 450.716v02-00
INNEHÅLL
1.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT.......................................................3
2.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT.......................................................5
3.
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.............................................6
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.......................................................9
1.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
om ansvarsfrihet för genomförandet av budgeten för det europeiska gemensamma företaget för ITER och utveckling av fusionsenergi för budgetåret 2009
( C7‑0247/2010 – 2010/2187(DEC) )
– med beaktande av den slutliga årsredovisningen för det europeiska gemensamma företaget för ITER och utveckling av fusionsenergi för budgetåret 2009,
– med beaktande av revisionsrättens rapport om den slutliga årsredovisningen för det europeiska gemensamma företaget för ITER och utveckling av fusionsenergi för budgetåret 2009, samt det europeiska gemensamma företagets svar
EUT C 342, 16.12.2010, s.
22. ,
– med beaktande av rådets rekommendation av den 15 februari 2011 (5894/2011 – C7‑0051/2011 ),
– med beaktande av artikel 276 i EG-fördraget och artikel 319 i fördraget om Europeiska unionens funktionssätt,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1. , särskilt artikel 185,
– med beaktande av rådets beslut 2007/198/Euratom av den 27 mars 2007 om inrättande av ett europeiskt gemensamt företag för ITER och utveckling av fusionsenergi samt om beviljande av förmåner till detta företag
EUT L 90, 30.3.2007, s.
58. , särskilt artikel 5,
– med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002
EGT L 357, 31.12.2002, s.
72. av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002, särskilt artikel 94,
– med beaktande av artikel 77 och bilaga VI i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet ( A7‑0131/2011 ).
2.
FÖRSLAG TILL EUROPAPARLAMENTETS BESLUT
om avslutande av räkenskaperna för det europeiska gemensamma företaget för ITER och utveckling av fusionsenergi för budgetåret 2009
( C7‑0247/2010 – 2010/2187(DEC) )
Europaparlamentet fattar detta beslut
– med beaktande av den slutliga årsredovisningen för det europeiska gemensamma företaget för ITER och utveckling av fusionsenergi för budgetåret 2009,
– med beaktande av revisionsrättens rapport om den slutliga årsredovisningen för det europeiska gemensamma företaget för ITER och utveckling av fusionsenergi för budgetåret 2009, samt det europeiska gemensamma företagets svar
EUT C 342, 16.12.2010, s.
22. ,
– med beaktande av rådets rekommendation av den 15 februari 2011 (5894/2011 – C7‑0051/2011 ),
– med beaktande av artikel 276 i EG-fördraget och artikel 319 i fördraget om Europeiska unionens funktionssätt,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1. , särskilt artikel 185,
EUT L 90, 30.3.2007, s.
58. , särskilt artikel 5,
– med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002
EGT L 357, 31.12.2002, s.
72. av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002, särskilt artikel 94,
– med beaktande av artikel 77 och bilaga VI i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet ( A7‑0131/2011 ).
3.
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för det europeiska gemensamma företaget för ITER och utveckling av fusionsenergi för budgetåret 2009
( C7‑0247/2010 – 2010/2187(DEC) )
Europaparlamentet utfärdar denna resolution
– med beaktande av den slutliga årsredovisningen för det europeiska gemensamma företaget för ITER och utveckling av fusionsenergi för budgetåret 2009,
– med beaktande av revisionsrättens rapport om den slutliga årsredovisningen för det europeiska gemensamma företaget för ITER och utveckling av fusionsenergi för budgetåret 2009, samt det europeiska gemensamma företagets svar
EUT C 342, 16.12.2010, s.
22. ,
– med beaktande av rådets rekommendation av den 15 februari 2011 (5894/2011 – C7‑0051/2011 ),
– med beaktande av artikel 276 i EG-fördraget och artikel 319 i fördraget om Europeiska unionens funktionssätt,
– med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget
EGT L 248, 16.9.2002, s.
1. , särskilt artikel 185,
EUT L 90, 30.3.2007, s.
58. , särskilt artikel 5,
– med beaktande av budgetförordningen för det europeiska gemensamma företaget för ITER och utveckling av fusionsenergi, som antogs genom ett beslut i ITERS styrelse den 22 oktober 2007 (nedan kallad det gemensamma företagets budgetförordning),
– med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002
EGT L 357, 31.12.2002, s.
72. av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002, särskilt artikel 94,
– med beaktande av artikel 77 och bilaga VI i arbetsordningen,
– med beaktande av betänkandet från budgetkontrollutskottet ( A7‑0131/2011 ).
A. Revisionsrätten har förklarat att den har uppnått en rimlig säkerhet om att räkenskaperna för budgetåret 2009 är tillförlitliga och att de underliggande transaktionerna är lagliga och korrekta.
B. Det gemensamma företaget är i ett inledningsskede och hade inte till fullo inrättat sina system för interna kontroller och ekonomisk information vid utgången av 2009.
C. Det gemensamma företagets budgetförordning är baserad på rambudgetförordningen, som nyligen ändrats för att överensstämma med de ändringar som gjorts i den allmänna budgetförordningen.
D. Den 9 oktober 2008 avgav revisionsrätten sitt yttrande nr 4/2008 om det gemensamma företagets budgetförordning.
Genomförande av budgeten
Europaparlamentet noterar att det gemensamma företagets banktillgodohavanden i slutet av året uppgick till 42 000 000 EUR, vilket strider mot principen om balans i budgeten.
Årsredovisningar
5.
Internkontrollsystem
7.
Budgetförordningen
– undantag från budgetprinciperna,
– rollen för kommissionens internrevisionstjänst,
– inrättandet av en revisionskommitté,
– sen inbetalning av medlemmarnas årsavgifter,
– villkoren för beviljande av bidrag,
– de övergångsregler som föreskrivs i artikel 133 i det gemensamma företagets budgetförordning.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
21.3.2011
Slutomröstning: resultat
+:
–:
0:
20
3
Slutomröstning: närvarande ledamöter
Marta Andreasen, Jean-Pierre Audy, Inés Ayala Sender, Andrea Češková, Jorgo Chatzimarkakis, Tamás Deutsch, Martin Ehrenhauser, Jens Geier, Ingeborg Gräßle, Iliana Ivanova, Elisabeth Köstinger, Monica Luisa Macovei, Aldo Patriciello, Crescenzio Rivellini, Bart Staes, Georgios Stavrakakis, Søren Bo Søndergaard
Slutomröstning: närvarande suppleanter
A7-0179/2011
*
BETÄNKANDE
om förslaget till rådets förordning om ändring av förordning (EG) nr 1467/97 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott
(KOM(2010)0522 – C7‑0396/2010 – 2010/0276(CNS))
Utskottet för ekonomi och valutafrågor
Föredragande: Diogo Feio
PE 454.690v03-00
Teckenförklaring
* Samrådsförfarande
*** Godkännandeförfarande
***I Ordinarie lagstiftningsförfarande (första behandlingen)
***II Ordinarie lagstiftningsförfarande (andra behandlingen)
***III Ordinarie lagstiftningsförfarande (tredje behandlingen)
(Det angivna förfarandet baseras på den rättsliga grund som angetts i förslaget till akt.)
Ändringsförslag till ett förslag till akt
Parlamentets ändringsförslag till ett förslag till akt ska markeras med fetkursiv stil .
De berörda avdelningarna tar sedan ställning till dessa korrigeringsförslag.
Om parlamentet önskar ändra delar av en bestämmelse i en befintlig akt som inte ändrats i förslaget till akt, ska dessa markeras med fet stil .
Eventuella strykningar ska i sådana fall markeras enligt följande: [...] .
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
YTTRANDE FRÅN utskottet för rättsliga frågor ...........................................26
YTTRANDE från utskottet för sysselsättning och sociala frågor ...35
ÄRENDETS GÅNG..................................................................................................................51
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till rådets förordning om ändring av förordning (EG) nr 1467/97 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott
( KOM(2010)0522 – C7‑0396/2010 – 2010/0276(CNS) )
(Särskilt lagstiftningsförfarande – samråd)
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till rådet ( KOM(2010)0522 ),
– med beaktande av yttrandet från utskottet för rättsliga frågor över den föreslagna rättsliga grunden,
– med beaktande av yttrandet av Europeiska centralbanken av den 16 februari 2011
Ännu ej offentliggjort i EUT. .
– med beaktande av artiklarna 55 och 37 i arbetsordningen,
– med beaktande av betänkandet från utskottet för ekonomi och valutafrågor och yttrandet från utskottet för sysselsättning och sociala frågor ( A7‑0179/2011 ).
1.
PARLAMENTETS ÄNDRINGAR
* Ändringar: ny text eller text som ersätter tidigare text markeras med fetkursiv stil och strykningar med symbolen ▌. *
till kommissionens förslag till
---------------------------------------------------------
RÅDETS FÖRORDNING (EU) nr …/…
om ändring av förordning (EG) nr 1467/97 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Europeiska kommissionens förslag,
efter översändande av utkastet till lagstiftningsakt till de nationella parlamenten,
med beaktande av Europaparlamentets yttrande
EUT C , , s.. ,
i enlighet med det ordinarie lagstiftningsförfarandet, och
av följande skäl:
(1) Samordningen av medlemsstaternas ekonomiska politik inom unionen bör enligt fördraget om Europeiska unionens funktionssätt (EUF-fördraget) innebära att man följer riktlinjerna om stabila priser, sunda och balanserade offentliga finanser och monetära förhållanden samt en stabil betalningsbalans , i syfte att uppnå en hållbar tillväxt och social sammanhållning, samt måle n som fastställts i EU- och EUF ‑ fördragen, samtidigt som fördragens övergripande klausuler respekteras .
(2) Inledningsvis utgick stabilitets- och tillväxtpakten från rådets förordning (EG) nr 1466/97 av den 7 juli 1997 om förstärkning av övervakningen av de offentliga finanserna samt övervakningen och samordningen av den ekonomiska politiken, rådets förordning (EG) nr 1467/97 av den 7 juli 1997 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott samt Europeiska rådets resolution av den 17 juni 1997 om stabilitets- och tillväxtpakten.
Förordningarna (EG) nr 1466/97 och (EG) nr 1467/97 ändrades år 2005 genom förordningarna (EG) nr 1055/2005 respektive (EG) nr 1056/2005.
Dessutom antogs rådets rapport av den 20 mars 2005 om ”Att förbättra genomförandet av stabilitets- och tillväxtpakten”.
(2b) En heltäckande och integrerad lösning på euroområdets skuldkris är nödvändig eftersom en punktinsatsmetod hittills inte har fungerat.
(2c) Medlemsstaternas politiska svar på bedömningar, beslut, rekommendationer och varningar från kommissionen eller rådet inom ramen för den europeiska planeringsterminen bör beaktas i) i förfarandena för kontroll av efterlevnaden av stabilitets- och tillväxtpaktens förebyggande och korrigerande delar, ii) i verkställighetsåtgärderna för att korrigera alltför stora makroekonomiska obalanser i euroområdet, iii) för att säkerställa att villkor relaterade till anslag från Europeiska valutafonden är korrekt anpassade till medlemsstaternas särdrag och att den ekonomiska politiken är på rätt spår, och iv) för att säkerställa att det finansiella stödet från Europeiska valutafonden till medlemsstaterna kommer att lindra de ekonomiska anpassningschockerna, hjälpa medlemsstaterna att undvika statsbankrutt, förhindra kostnader för andra länder genom spridning och garantera finansiell stabilitet i euroområdet som helhet.
(2d) Kommissionen bör få en starkare och mer oberoende roll i förfarandet för förstärkt övervakning.
Detta gäller medlemsstatsspecifika bedömningar, övervakningsinsatser, övervakningsbesök, rekommendationer och varningar.
Dessutom måste rådets roll minskas i de etapper som leder till potentiella sanktioner, och omröstningen med omvänd kvalificerad majoritet i rådet måste användas där så är möjligt i enlighet med EUF-fördraget.
Den rådsmedlem som företräder den berörda medlemsstaten och företrädarna för de medlemsstater som inte följer rådets rekommendationer att vidta korrigerande åtgärder i enlighet med stabilitets- och tillväxtpakten eller åtgärder vid alltför stora makroekonomiska obalanser bör inte delta i omröstningen.
(3) Stabilitets- och tillväxtpakten grundas på målet om sunda och hållbara offentliga finanser, som ett sätt att stärka förutsättningarna för prisstabilitet och stark varaktig tillväxt som kan bidra till ökad sysselsättning.
Genomförandet bör därför mätas i jämförelse med förmågan att uppnå dessa mål.
(4a) Den ekonomiska utvecklingen i unionen har skapat nya problem för den nationella finanspolitiken och har särskilt belyst behovet av enhetliga minimikrav för reglerna och förfarandena i medlemsstaternas budgetstruktur.
(4b) Ramen för förbättrad ekonomisk styrning bör bygga på flera sammanlänkade politiska åtgärder för hållbar tillväxt och sysselsättning, vilka måste vara inbördes samstämda, i synnerhet en unionsstrategi för tillväxt och sysselsättning som särskilt är inriktad på att utveckla och förstärka den inre marknaden, främja internationella handelsförbindelser och konkurrenskraft, en effektiv ram för att förebygga och korrigera alltför stora underskott i de offentliga finanserna (stabilitets- och tillväxtpakten), en stabil ram för att förebygga och korrigera makroekonomiska obalanser, minimikrav för nationella budgetramar, förstärkt reglering och tillsyn av finansmarknaderna (inbegripet Europeiska systemrisknämndens makrotillsyn) och en trovärdig permanent krislösningsmekanism.
(4c) Att uppnå och upprätthålla en dynamisk inre marknad bör betraktas som en central aspekt av en ekonomisk och monetär union som fungerar väl och friktionsfritt.
(4d) Stabilitets- och tillväxtpakten och unionens ram för ekonomisk styrning som helhet bör komplettera och vara förenliga med en unionsstrategi för tillväxt och skapande av sysselsättning som syftar till att stärka unionens konkurrenskraft.
Miljöansvar, sociala framsteg och stabilitet, samt utveckling och stärkande av den inre marknaden bör också omfattas av denna ram.
Dessa samband bör i princip inte medge undantag från stabilitets- och tillväxtpaktens bestämmelser.
(4e) En förstärkt ekonomisk styrning bör åtföljas av en större demokratisk legitimitet för ekonomisk styrning i unionen, vilket bör uppnås genom att Europaparlamentet och de nationella parlamenten i högre grad och i ett tidigare skede involveras i all samordning av den ekonomiska politiken.
(4f) Medlemsstaterna bör föreskriva budgetåtgärder, såsom nationella budgetbestämmelser, som respekterar principerna i rådets direktiv 2011/…/EU [om krav på medlemsstaternas budgetramar], och att offentliga institutioner, som är helt oberoende, deltar i budgetprocessen och i den medelfristiga budgetramen.
Nationella budgetbestämmelser bör komplettera medlemsstaternas åtaganden inom stabilitets- och tillväxtpakten.
Nationella institutioner bör spela en mer framträdande roll i budgetövervakningen för att stärka det nationella ansvaret, stärka kontrollen av efterlevnaden genom den nationella allmänheten och komplettera den ekonomiska och politiska analys som görs på EU-nivå.
Transparens, ansvars- och redovisningsskyldighet och oberoende tillsyn är centrala delar av en förstärkt ekonomisk styrning.
Rådet och kommissionen bör offentliggöra och förklara skälen för sina ståndpunkter och beslut vid lämpliga tidpunkter under samordningen av den ekonomiska politiken.
De nationella budgetramarna bör inbegripa upprättandet och stärkandet av rollen för oberoende budgetorgan och säkerställa att transparent budgetstatistik publiceras.
(4h) Utan att det påverkar rättigheterna och skyldigheterna enligt EUF-fördraget, bör de medlemsstater som inte har euron som valuta ha rätt att tillämpa lagstiftningen om ekonomisk styrning.
(4i) Erfarenheterna och misstagen från det första årtiondet med den ekonomiska och monetära unionen visar att det behövs en förbättrad ekonomisk styrning inom unionen, som bör bygga på ett större nationellt ansvar för gemensamt överenskomna regler och åtgärder och på solid are ramar för övervakning på EU ‑ nivå av den nationella ekonomiska politiken.
(4j) Kommissionen och rådet bör vid tillämpningen av denna förordning beakta alla relevanta faktorer och den ekonomiska och budgetmässiga situationen i de berörda medlemsstaterna, särskilt huruvida de är föremål för ett EU/IMF ‑ anpassningsprogram.
Dessutom bör en övergångsperiod införas så att medlemsstaterna kan anpassa sin politik till vissa bestämmelser i denna förordning.
(4k) I artikel 3 i protokollet (nr 12) om förfarandet vid alltför stora underskott som är fogat till fördragen föreskrivs att medlemsstaterna ska säkerställa att nationella förfaranden på budgetområdet gör det möjligt för dem att uppfylla de förpliktelser inom detta område som följer av fördragen.
De medlemsstater som har euron som valuta bör därför förankra målen för unionens budgetpolitik i nationell lagstiftning, och bör tillse att adekvata budgetförfaranden finns på plats för att uppfylla dessa mål.
(4l) Den permanenta krismekanismen bör antas i enlighet med det ordinarie lagstiftningsförfarandet och bygga på unionsmetoden i syfte att, å ena sidan, stärka parlamentets deltagande och förbättra den demokratiska ansvars- och redovisningsskyldigheten och, å andra sidan, stödja sig på kommissionens sakkunskaper, oberoende och opartiskhet.
(4m) Med tanke på marknadsvolatiliteten och nivåerna på räntedifferenserna mellan statsobligationer från vissa medlemsstater som har euron som valuta bör resoluta åtgärder vidtas för att försvara eurons stabilitet.
(4n) Europeiska valutafonden bör ha tre syften: den bör täcka en andel av medlemsstaternas statsskuld som kan betalas utan hot mot den finansiella stabiliteten i någon annan medlemsstat eller i euroområdet som helhet (eurovärdepapper), den bör hjälpa en medlemsstat som möter finansiella svårigheter med att lösa den kris som medlemsstaten har hamnat i (permanent krislösningsmekanism) och slutligen bör den uppbåda resurser för att finansiera investeringar som kan främja ekonomisk tillväxt (projektobligationer).
(4o) Medlemsstater som har euron som valuta bör sammanföra upp till [...] procent av statsskulden på basis av solidariskt ansvar (eurovärdepapper).
Medan gemensamma emissioner skulle öka likviditeten för obligationerna på kapitalmarknaden, skulle det gemensamma ansvaret hjälpa de stater som möter allt större svårigheter att anskaffa kapital.
Eurovärdepapper bör vara prioriterade i förhållande till nationella statspapper.
De skulle kunna bidra till att främja euron som reservvaluta.
(4p) För att förbättra budgetdisciplinen bör länder med en trovärdig ekonomisk politik och budgetpolitik tillåtas låna upp till [...] procent av sin BNP, medan länder med en svagare ekonomisk eller budgetmässig situation skulle tvingas betala en premie/extra räntesats eller endast kunna låna en mindre andel av BNP i eurovärdepapper.
I extrema fall, dvs. om ett medverkande land konsekvent för en ohållbar ekonomisk politik eller budgetpolitik bör dess deltagande i emissionen av eurovärdepapper avbrytas.
(4q) En europeisk valutafond, som förvaltas enligt unionsregler och finansieras i synnerhet med bötesintäkter, bör inrättas i syfte att säkra hela euroområdets finansiella stabilitet.
Denna fond bör grundas på rådets beslut av den 9–10 maj 2010 och uttalandet från Eurogruppen av den 28 november 2010.
(5) Reglerna om budgetdisciplin och om hur den ska respekteras och efterlevnaden kontrolleras bör stärkas, särskilt genom att ge skuldernas och den övergripande hållbarhetens nivå och utveckling en mer framträdande roll.
(5a) Skuldkriterierna, inbegripet privata skulder om de implicit utgör eventualförpliktelser för den offentliga sektorn, bör integreras bättre i varje steg av förfarandet vid alltför stora underskott så att de offentliga finansernas hållbarhet kan garanteras samtidigt som en lämplig nivå för offentliga investeringar bibehålls.
(5b) Konsolideringen av den inre marknaden är en grundläggande förutsättning för att den ekonomiska och monetära unionen ska kunna fungera korrekt och förstärkas .
I detta hänseende måste man avlägsna de befintliga rättsliga och fysiska hindren för att skapa ett gemensamt europeiskt järnvägsområde, särskilt för godstrafiken.
(5c) Större balans bör säkerställas mellan ekonomiska hänsyn och det politiska handlingsutrymmet men reglerna bör även i fortsättningen vara enkla, transparenta och genomförbara.
(5d) En bedömning av de offentliga finansernas hållbarhet, bland annat skuldnivån, skuldprofilen (inbegripet löptid) och skuldutvecklingen ska mer eftertryckligt beaktas när det gäller konvergenstakten mot medlemsstatsspecifika budgetmål på medellång sikt som ska inkluderas i stabilitets- och konvergensprogrammen.
(5e) Som ett komplement till förfarandet vid alltför stora underskott bör det fastställas en tydlig, harmoniserad ram för att bedöma och övervaka skuldutvecklingen, inbegripet implicita skyldigheter och ansvarsförbindelser, t.ex. pensionsåtaganden och offentliga garantier (t.ex. avseende kapital, räntor eller inkomstflöden) för investeringar i finanssektorn och i offentlig-privata partnerskap samt sådana investeringars kostnader för den nationella budgeten under åren.
(5f) Strukturen för att kontrollera offentliga och privata skulder bör främja långsiktig tillväxt, ta vederbörlig hänsyn till budgetpolitikens konjunkturdämpande roll och förbättra investeringsvillkor och utveckla den inre marknaden, samtidigt som medlemsstatsspecifika prioriteringar och behov respekteras.
(6) För att det nuvarande förfarandet vid alltför stora underskott ska kunna genomföras utifrån både underskotts- och skuldkriteriet, krävs ▌ett numeriskt riktmärke som tar hänsyn till konjunkturcykeln för bedömningen av om den offentliga skuldens andel av bruttonationalprodukten minskar i tillräcklig utsträckning och närmar sig referensvärdet i tillfredsställande takt , eller anses befinna sig i en situation av övergående avvikelse från den tillräckliga minskningstakten .
Alla faktorer av betydelse bör beaktas vid bedömningen.
(6a) En försiktig och hållbar finanspolitik bör leda till att det medelfristiga målet för de offentliga finanserna uppnås och att det även i fortsättningen respekteras.
De medlemsstater som håller fast vid det medelfristiga budgetmålet bör därigenom få en säkerhetsmarginal gentemot referensvärdet för det offentliga underskottet på 3 % av BNP, vilket innebär snabba framsteg mot hållbara offentliga finanser, och samtidigt få budgetmässigt manöverutrymme, särskilt med tanke på behovet av offentliga investeringar.
(7a) Inom ramen för stabilitets- och tillväxtpaktens förebyggande del bör incitamentet för en försiktig och hållbar finanspolitik bestå i att en medlemsstat i euroområdet som inte genomför en tillräcklig budgetkonsolidering måste lämna en tillfällig räntebärande deposition.
(8a) Även när förekomsten av ett alltför stort underskott har fastställts bör alla relevanta faktorer beaktas under de följande skedena i förfarandet.
Genomförandet av åtgärder för att öka den potentiella tillväxttakten på medellång sikt inom ramen för unionens gemensamma tillväxtstrategi bör i synnerhet beaktas på ett lämpligt sätt när man fastställer, och eventuellt förlänger, tidsfristen för att korrigera det alltför stora överskottet.
(8b) När man beaktar reformer av pensionssystemen bland de relevanta faktorerna bör huvudkriteriet vara huruvida de förbättrar hållbarheten på lång sikt i pensionssystemet generellt, utan att öka riskerna för budgetsituationen på medellång sikt.
Man bör därvid även ta hänsyn till de minimikrav som fastställs i rådets direktiv [om krav på medlemsstaternas budgetramar] liksom andra överenskomna önskvärda krav på budgetdisciplin.
(10) Övervakningen av om rådets rekommendationer om korrigering av alltför stora överskott följs bör underlättas genom att dessa specificerar årliga finanspolitiska mål, som överensstämmer med den begärda förbättringen av de offentliga finanserna i konjunkturrensade termer, exklusive finanspolitiska engångsåtgärder och andra tillfälliga åtgärder.
I detta sammanhang bör det årliga riktmärket motsvarande 0,5 % av BNP uppfattas som årsmedelvärde.
(11) Vid bedömningen av effektiva åtgärder vore det en fördel att använda följandet av offentliga utgiftsmål som utgångspunkt tillsammans med genomförandet av andra planerade särskilda åtgärder på intäktssidan.
(12) Vid bedömningen av om tidsfristen exceptionellt bör förlängas för att korrigera ett alltför stort underskott, bör ▌hänsyn tas till omfattande och allvarliga konjunkturnedgångar eller exceptionella omständigheter i en medlemsstat .
(14) För att säkerställa att deltagande medlemsstater följer unionens ramverk för den finanspolitiska tillsynen, bör regelbaserade incitament och sanktioner utformas utifrån artikel 136 i EUF-fördraget för att åstadkomma rättvisa, punktliga och effektiva mekanismer för följande av stabilitets- och tillväxtpaktens regler.
(14a) Ekonomiskt och politiskt känsligare incitament och sanktioner bör ta vederbörlig hänsyn till det nationella underskottets och den nationella skuldens struktur (inbegripet implicita skyldigheter), ”konjunkturcykeln”, i syfte att undvika en konjunkturförstärkande finanspolitik, samt den strukturella sammansättningen av de offentliga inkomster och utgifter som behövs för tillväxtfrämjande strukturreformer.
Om medlemsstaterna uppfyller kriterierna för att använda sådana mekanismer kan kommissionen och rådet uppmana dem att lämna in den ansökan som behövs.
(14c) Incitament för och sanktioner mot medlemsstater i euroområdet bör genomdrivas och tillämpas med hänsyn till de mycket nära kopplingarna till medlemsstater utanför euroområdet, särskilt de medlemsstater som förväntas bli en del av detta område, som en del av det nya multilaterala tillsynssystemet och stabilitets- och tillväxtpaktens förstärkta instrument, särskilt tydligare fokus på budgetmål på medellång sikt.
(14d) Rådet och kommissionen bör offentliggöra sina ståndpunkter och beslut vid lämpliga tidpunkter under samordningen av den ekonomiska politiken – alltid med vederbörligt iakttagande av bestämmelserna i fördraget – så att ett effektivt kollegialt tryck kan åstadkommas, och Europaparlamentet bör kunna uppmana den berörda medlemsstaten att förklara sina beslut och politiska åtgärder inför parlamentets ansvariga utskott.
(14e) Kommissionens årliga politiska rekommendationer bör diskuteras i Europaparlamentet innan diskussionerna i rådet inleds.
(14f) De böter som indrivits i enlighet med artikel 12 i denna förordning bör utgöra sådana andra inkomster som avses i artikel 311 i EUF-fördraget, och bör föras till en permanent krismekanism för de medlemsstater som har euron som valuta.
Tills denna mekanism har inrättats bör böterna avsättas till finansieringsinstrument med riskdelning för EU-relevanta projekt som finansieras av Europeiska investeringsbanken i enlighet med bestämmelserna i det till fördragen fogade protokollet (nr 5) om Europeiska investeringsbankens stadga.
(15) Vid hänvisningarna i förordning (EG) nr 1467/97 bör det beaktas att artikelnumreringen i fördraget om Europeiska unionens funktionssätt är ny och att rådets förordning (EG) nr 3605/93 ersatts med rådets förordning (EG) nr 479/2009 av den 25 maj 2009 om tillämpningen av protokollet om förfarandet vid alltför stora underskott som är fogat till fördraget om upprättandet av Europeiska gemenskapen.
(16) Förordning (EG) nr 1467/97 bör därför ändras i enlighet med detta.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 1467/97 ska ändras på följande sätt.
1.
Artikel 1 ska ersättas med följande:
”Artikel 1
1.
Bestämmelserna i denna förordning ska påskynda och förtydliga tillämpningen av förfarandet vid alltför stora underskott .
Syftet med förfarandet vid alltför stora underskott är att förhindra alltför stora underskott i den offentliga sektorns finanser och att i de fall underskott uppstår bidra till att de omgående korrigeras, varvid iakttagandet av budgetdisciplin granskas med utgångspunkt från kriterierna offentliga underskott och offentliga skulder.
Rådet ska använda omröstning med omvänd kvalificerad majoritet när det fattar beslut om antagande av rekommendationer och förelägganden utifrån kommissionens formella ståndpunkter enligt artikel 126 i EUF-fördraget.
▐
2.
En medlemsstat med undantag får tillämpa de bestämmelser som gäller för deltagande medlemsstater i enlighet med denna förordning, och ska i sådant fall meddela kommissionen detta.
Ett sådant meddelande ska offentliggöras i Europeiska unionens officiella tidning.
Den berörda medlemsstaten ska vid tillämpningen av denna förordning anses som deltagande medlemsstat från och med dagen efter ett sådant offentliggörande.”
2.
Artikel 2 ska ändras på följande sätt:
a) I punkt 1 ska första stycket ersättas med följande:
”1.
b) Följande punkt ▌ska läggas till:
”1a.
Kravet enligt skuldkriteriet ska också anses vara uppfyllt om budgetprognoserna från kommissionen anger att den föreskrivna minskningen i differensen kommer att inträffa under en treårsperiod som omfattar två år efter det sista året för vilket uppgifterna finns tillgängliga.
För en medlemsstat som är föremål för förfarandet vid alltför stora underskott [datum för antagande av denna förordning - ska införas] och under en treårsperiod från korrigeringen av det alltför stora underskottet ska kravet enligt skuldkriteriet anses vara uppfyllt om den berörda medlemsstaten gör tillräckliga framsteg när det gäller att uppfylla det enligt bedömningen i rådets yttranden om dess stabilitets- eller konvergensprogram.
Vid tillämpningen av riktmärket för skuldanpassning ska de relevanta faktorerna för varje land i enlighet med punkt 3 beaktas.
I denna bedömning ska särskild uppmärksamhet fästas vid den fas av konjunkturcykeln som en medlemsstat befinner sig i.”
c) Punkt 3 ska ersättas med följande:
”3.
Rapporten ska på lämpligt sätt ta upp
– Det ekonomiska lägets utveckling på medellång sikt , särskilt tillväxtpotential och konjunkturutveckling , inflation, politiskt genomförande av unionens gemensamma tillväxtstrategi, och andra mål i enlighet med EUF-fördraget, förhindrande och korrigering av alltför stora makroekonomiska obalanser och den privata sektorns nettosparande.
– Utvecklingen avseende anpassningsbanan för att uppnå budgetmålen på medellång sikt (särskilt primära utgifter, offentliga investeringar ▌och de offentliga finansernas allmänna kvalitet, särskilt då de nationella budgetramarnas ändamålsenlighet), enligt artikel 5 i förordning (EG) nr 1466/97 .
– Utvecklingen av de offentliga löpande utgifterna på medellång sikt ska också beaktas, särskilt deras stabilitet i reala termer.
– Rapporten ska ▌också innehålla en analys av den offentliga skuldställningen på medellång sikt , dess dynamik och hållbarhet (särskilt ▌riskfaktorer ▌ inklusive skuldernas löptids- och valutastruktur, stock-/flödesjusteringar och deras sammansättning , ackumulerade reserver och andra finansiella tillgångar; garantier särskilt till finanssektorn; och alla implicit relaterade skulder såsom privata skulder om de implicit utgör eventualförpliktelser för den offentliga sektorn).
– Dessutom ska kommissionen vederbörligen och uttryckligen beakta eventuella andra faktorer som enligt den berörda medlemsstaten har betydelse för en samlad bedömning av om underskotts- och skuldkriterierna uppfylls och som medlemsstaten har förelagt rådet och kommissionen ▌.
I detta sammanhang ska särskild hänsyn tas till budgetmässiga ansträngningar för att främja internationell solidaritet och uppnå unionens politiska mål, och framför allt skuld som uppstått i form av bilateralt och multilateralt stöd mellan medlemsstaterna i samband med åtgärder för att trygga den finansiella stabiliteten .
Särskild och uttrycklig hänsyn ska också tas till den finansiella bördan från rekapitaliseringsåtgärder och andra tillfälliga statliga stödåtgärder för den finansiella sektorn vid allvarliga finansiella störningar samt lån och garantier som beviljats andra medlemsstater och den europeiska finansiella stabiliseringsfaciliteten och den europeiska stabiliseringsmekanismen.
När kommissionen utarbetar en rapport får den begära ytterligare information från den berörda medlemsstaten.
d) Punkt 4 ska ersättas med följande:
”4.
da) Punkt 5 ska ersättas med följande:
”5.
db) Följande punkt ska införas:
”5a.
Dessa faktorer ska dock beaktas under de steg som föregår beslutet om förekomsten av ett alltför stort underskott vid bedömningen av om skuldkriteriet uppfylls.”
dc) Punkt 6 ska ersättas med följande:
”6.
e) Punkt 7 ska ersättas med följande:
”7.
2a.
Följande avsnitt ska införas:
”AVSNITT 1a
EKONOMISK DIALOG
Artikel 2a
3.
Artikel 3 ska ändras på följande sätt:
(-a) Punkt 1 ska ersättas med följande:
1.
a) Punkt 2 ska ersättas med följande:
”2.
b) ▌Punkt 3 ska ersättas med följande:
” 3.
c) Punkt 4 ska ersättas med följande:
”4.
Om omständigheterna är allvarliga får tidsfristen för effektiva åtgärder förkortas till tre månader.
I rådets rekommendation ska det även fastställas en tidsfrist för korrigeringen av det alltför stora underskottet, vilken ska slutföras under det år som följer på året då underskottet fastställdes, om inte särskilda omständigheter föreligger.
I sin rekommendation ska rådet begära att medlemsstaten uppnår årliga budgetmål som enligt rekommendationens underliggande prognos som ett riktmärke motsvarar en minskning av underskottet med minst 0,5 % av BNP av sitt konjunkturrensade saldo, utan engångsåtgärder och tillfälliga åtgärder som direkt eller indirekt påverkar budgeten , för att korrigera det alltför stora underskottet inom tidsfristen i rekommendationen.”
d) Följande punkt ▌ska läggas till:
”4a.
Kommissionen får begära ytterligare rapportering från den berörda medlemsstaten.
Rapporten ska offentliggöras.”
da) Följande punkt ska införas:
”4b.
Europaparlamentets behöriga utskott kan bjuda in en företrädare för den berörda medlemsstaten för att inför utskottet förklara den ekonomiska politiken och budgetpolitiken och ange vilka åtgärder man avser att vidta för att komma tillrätta med det alltför stora underskottet.
Medlemsstaten får också av samma skäl begära att bli inbjuden till Europaparlamentet.”
e) Punkt 5 ska ersättas med följande:
”5.
Rådet ska bedöma om det, jämfört med de ekonomiska prognoserna i sin rekommendation, föreligger oväntade negativa ekonomiska händelser med stora negativa effekter för de offentliga finanserna.
4.
Artikel 4 ska ändras på följande sätt:
a) Punkt 1 ska ersättas med följande:
” 1.
b) Punkt 2 ska ersättas med följande:
”2.
Kommissionen kan genomföra övervakningsbesök på plats i enlighet med artikel 10a.
För deltagande medlemsstater, och medlemsstater som deltar i ERM2, ska sådana besök genomföras i samarbete med Europeiska centralbanken.
Kommissionen ska rapportera till Europaparlamentet och rådet om resultatet av besöket, och ska offentliggöra resultatet.
2a.
Europaparlamentet ska underrättas om de förhållanden som beskrivs i punkterna 1 och 2.”
5.
Artikel 5 ska ändras på följande sätt:
a) Punkt 1 ska ersättas med följande:
”1.
I föreläggandet ska rådet begära att medlemsstaten uppnår årliga budgetmål som enligt rekommendationens underliggande prognos som ett riktmärke motsvarar en årlig minskning av underskottet med minst 0,5 % av BNP av sitt konjunkturrensade saldo, utan engångsåtgärder och tillfälliga åtgärder som direkt eller indirekt påverkar budgeten , för att korrigera det alltför stora underskottet inom tidsfristen i rekommendationen.
Rådet ska också ange åtgärder som främjar att dessa mål uppnås.”
b) Följande punkt 1a ska läggas till:
”1a.
Kommissionen ska genom övervakningsbesök i enlighet med artikel 10a följa och utvärdera de anpassningsåtgärder som vidtagits för att tackla det alltför stora underskottet, och utarbeta en rapport till rådet.
Rapporten ska offentliggöras.”
ba) Följande punkt ska införas:
”1b.
Europaparlamentets behöriga utskott kan bjuda in den berörda medlemsstaten för att inför utskottet förklara den ekonomiska politiken och budgetpolitiken och ange vilka åtgärder man avser att vidta för att komma till rätta med det alltför stora underskottet.
Medlemsstaten får också av samma skäl begära att bli inbjuden till Europaparlamentet.”
c) Punkt 2 ska ersättas med följande:
”2.
Rådet ska bedöma om det, jämfört med de ekonomiska prognoserna i sin rekommendation, föreligger oväntade negativa ekonomiska händelser med stora negativa effekter för de offentliga finanserna.
6.
Artikel 6 ska ersättas med följande:
”Artikel 6
1.
2.
”Artikel 7
Ett påskyndat förfarande ska användas om det rör sig om ett avsiktligt planerat underskott som enligt rådets beslut är alltför stort.
Europaparlamentets behöriga utskott får uppmana medlemsstaten att rapportera inför parlamentets behöriga utskott.”
7a.
Följande artikel ska införas:
”Artikel 7a
Möten mellan parlament
Alltid när det anordnas ett möte mellan Europaparlamentets behöriga utskott och en medlemsstat för att förklara en ståndpunkt, en begärd åtgärd eller avvikelser från kraven i denna, ska mötet hållas under överinseende av antingen
a) Europaparlamentet,
b) medlemsstatens parlament, eller
c) parlamentet i den medlemsstat som för tillfället innehar ordförandeskapet för unionen.”
8.
Artikel 8 ska ersättas med följande:
”Artikel 8
9.
10.
Artikel 10 ska ändras på följande sätt:
a) Inledningsfrasen till punkt 1 ska ersättas med följande:
”1.
Kommissionen och rådet ska regelbundet övervaka genomförandet av de åtgärder som har vidtagits.”
aa) Följande punkt ska införas:
”1a.
Kommissionen och rådet ska rapportera sina resultat i enlighet med punkt 1 till Europaparlamentet.
b) I punkt 3 ska hänvisningen till ”förordning (EG) nr 3605/93” ersättas med en hänvisning till ”förordning (EG) nr 479/2009”.
10a.
Följande artikel ska införas:
”Artikel 10a
1.
Kommissionen ska se till att det förs en ständig dialog med medlemsstaternas myndigheter i enlighet med målen i denna förordning.
I detta syfte ska kommissionen genomföra besök i alla medlemsstater för en regelbunden dialog och, vid behov, övervakning.
Kommissionen får, om den anser det lämpligt, inbjuda företrädare för Europeiska centralbanken eller andra relevanta institutioner att delta i dialog- och övervakningsbesöken.
2.
När kommissionen organiserar dialog- och övervakningsbesök, ska den när så är lämpligt översända sina preliminära resultat till den berörda medlemsstaten för synpunkter.
3.
Kommissionen ska i samband med dialogbesök granska den aktuella ekonomiska situationen i medlemsstaten och fastställa eventuella risker och svårigheter när det gäller att uppfylla målen i denna förordning.
4.
Kommissionen ska i samband med övervakningsbesök följa upp processerna och kontrollera att åtgärder vidtagits i överensstämmelse med rådets och kommissionens beslut i enlighet med målen i denna förordning.
Övervakningsbesök ska enbart genomföras i undantagsfall och bara då det föreligger betydande risker eller svårigheter när det gäller att uppnå dessa mål.
5.
Kommissionen ska informera Ekonomiska och finansiella kommittén om orsakerna till övervakningsbesöken.
6.
Medlemsstaterna ska vidta alla åtgärder som krävs för att underlätta dialog- och övervakningsbesöken.
Medlemsstaterna ska på begäran av kommissionen och på frivillig basis se till att alla relevanta nationella myndigheter bistår vid förberedelsen och genomförandet av dialog- och övervakningsbesök.”
11.
”Artikel 11
När rådet beslutar att tillämpa sanktioner mot en deltagande medlemsstat i enlighet med artikel 126.11 i EUF-fördraget, ska som regel böter åläggas.
Europaparlamentets behöriga utskott får, inom tre månader från det datum då de sanktioner som avses i punkt 1 tillkännagavs, uppmana den berörda medlemsstaten att inför utskottet förklara varför den trots utfärdade varningar inte har åtgärdat det alltför stora underskottet.
Medlemsstaten får också av samma skäl begära att bli inbjuden till Europaparlamentet.”
12.
Artikel 12 ska ersättas med följande:
”Artikel 12
Fastställandet av den rörliga delen ska baseras på en utvärdering som rådet ska göra av huruvida den deltagande medlemsstaten har vidtagit effektiva åtgärder.
Om rådet anser att medlemsstaten har vidtagit effektiva åtgärder ska inte någon rörlig del tillämpas.
Beslutet att inte tillämpa den rörliga delen ska antas med kvalificerad majoritet.
2.
Om ytterligare böter beslutas, ska de beräknas på samma sätt som för den rörliga delen av böterna enligt punkt 1.
3.
Inga enskilda bötesbelopp enligt punkterna 1 och 2 får överskrida en övre gräns på 0,2 % av BNP.”
13.
Artikel 13 ska upphävas och hänvisningen till den i artikel 15 ska ersättas med en hänvisning till ”artikel 12”.
14.
Artikel 16 ska ersättas med följande:
”Artikel 16
De böter som indrivits i enlighet med artikel 12 i denna förordning ska utgöra sådana andra inkomster som avses i artikel 311 i EUF-fördraget, och ska föras till en permanent krismekanism för de medlemsstater som har euron som valuta .
Tills denna mekanism har inrättats ska böterna avsättas till finansieringsinstrument med riskdelning för EU-relevanta projekt som finansieras av Europeiska investeringsbanken i enlighet med bestämmelserna i det till fördragen fogade protokollet (nr 5) om Europeiska investeringsbankens stadga.”
14a.
Följande artikel ska införas:
”Artikel 17a
1.
Senast ...
Ü  UT, var vänlig och för in datum: ... år efter den dag då denna förordning träder i kraft Ü och därefter vart tredje år sk a kommissionen offentliggöra en rapport om tillämpningen av denna förordning.
2.
Rapporten och eventuella åtföljande förslag ska överlämnas till Europaparlamentet och rådet.
3.
Om man i rapporten fastställer att det föreligger hinder för genomförandet av de regler och bestämmelser i fördragen som styr den ekonomiska och monetära unionen, ska kommissionen lämna de nödvändiga rekommendationerna till Europeiska rådet.
4.
15.
Alla hänvisningar till ”artikel 104” i förordningen ska ersättas med hänvisningar till ”artikel 126 i EUF-fördraget”.
16.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning .
För en medlemsstat som är föremål för förfarandet vid alltför stora underskott [datum för antagande av denna förordning - ska införas] och under en treårsperiod från korrigeringen av det alltför stora underskottet ska kravet enligt skuldkriteriet anses vara uppfyllt om den berörda medlemsstaten gör tillräckliga framsteg när det gäller att uppfylla det enligt bedömningen i rådets yttranden om dess stabilitets- eller konvergensprogram.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Utfärdad i […].
På rådets vägnar
Ordförande
YTTRANDE FRÅN utskottet för rättsliga frågor
Sharon Bowles
Ordförande
Utskottet för ekonomi och valutafrågor
BRYSSEL
Vid utskottssammanträdet den 12 april 2011 behandlade utskottet detta ärende.
Syftet med lagstiftningspaketet för ekonomisk styrning är att tillgodose behovet av större samordning och närmare övervakning av den ekonomiska politiken i den ekonomiska och monetära unionen.
Paketet består av sex lagstiftningsförslag.
I bilagan återfinns en separat granskning för vart och ett av förslagen.
För enkelhetens skull anges här utskottets slutsatser angående lämpligheten i den rättsliga grunden för varje enskilt fall:
– Förslag till Europaparlamentets och rådets förordning om förebyggande och korrigering av makroekonomiska obalanser ( KOM(2010)0527 – 2010/0281(COD) )
– Förslag till rådets direktiv om krav på medlemsstaternas budgetramverk ( KOM(2010)0523 – 2010/0277(NLE) )
– Förslag till Europaparlamentets och rådets förordning om ändring av förordning (EG) nr 1466/97 om förstärkning av övervakningen av de offentliga finanserna samt övervakningen och samordningen av den ekonomiska politiken ( KOM(2010)0526 – 2010/0280(COD) )
Syftet med detta förslag är att förstärka samordningen av medlemsstaternas ekonomiska politik.
– Förslag till rådets förordning om ändring av förordning (EG) nr 1467/97 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott ( KOM(2010)0522 – 2010/0276(CNS) )
– Förslag till Europaparlamentets och rådets förordning om verkställighetsåtgärder för att korrigera alltför stora makroekonomiska obalanser i euroområdet ( KOM(2010)0525 – 2010/0279(COD) )
Vid utskottssammanträdet den 12 april 2011 antog utskottet för rättsliga frågor enhälligt
Följande ledamöter var närvarande vid slutomröstningen: Klaus-Heiner Lehne (ordförande), Evelyn Regner (vice ordförande), Piotr Borys, Sergio Gaetano Cofferati, Christian Engström, Lidia Joanna Geringer de Oedenberg, Sajjad Karim, Kurt Lechner, Eva Lichtenberger, Antonio López-Istúriz White, Arlene McCarthy, Antonio Masip Hidalgo, Alajos Mészáros, Angelika Niebler, Bernhard Rapkay, Alexandra Thein, Diana Wallis, Rainer Wieland, Cecilia Wikström, Tadeusz Zwiefka. följande rekommendationer.
Med vänlig hälsning
Klaus-Heiner Lehne
Bilaga Bilaga
Ärende: Yttrande över den rättsliga grunden för förslaget till rådets förordning om ändring av förordning (EG) nr 1467/97 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott ( KOM(2010)0522 – 2010/0276(CNS) )
Lagstiftningspaketet för ekonomisk styrning består av sex lagstiftningsförslag som syftar till att förstärka samordningen och övervakningen av den ekonomiska politiken i den ekonomiska och monetära unionen (EMU) i samband med Europa 2020-strategin och den europeiska planeringsterminen, vilka utgör en ny övervakningscykel där processerna inom ramen för stabilitets- och tillväxtpakten och de allmänna riktlinjerna för den ekonomiska politiken sammanförs.
Dessa förslag utgör ett svar på de svagheter som det nuvarande systemet är behäftat med och som uppdagats i samband med den globala ekonomiska och finansiella krisen.
Enligt kommissionen måste systemet stärkas för att ” befästa makroekonomisk stabilitet och hållbara offentliga finanser som en förutsättning för en varaktig produktions- och sysselsättningstillväxt ”
Förslag till rådets förordning (EU) nr …/… om ändring av förordning (EG) nr 1467/97 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott, motiveringen. .
Förslagen följer två meddelanden
”Förstärkt samordning av den ekonomiska politiken” av den 12 maj 2010 och ”Förstärkt samordning av den ekonomiska politiken för stabilitet, tillväxt och nya arbetstillfällen – Verktyg för en kraftfullare ekonomisk styrning” av den 30 juni 2010. från kommissionen och en överenskommelse i Europeiska rådet från juni 2010 om behovet av förstärkt samordning av medlemsstaternas ekonomiska politik.
Lagstiftningspaketet för ekonomisk styrning lades fram den 29 september 2010.
Förslaget till rådets förordning om ändring av förordning (EG) nr 1467/97 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott håller för närvarande på att granskas av utskottet för ekonomi och valutafrågor, med Diogo Feio som föredragande.
Utskottet för sysselsättning och sociala frågor är rådgivande utskott (föredragande: David Casa).
Europaparlamentet medverkar inom ramen för samrådsförfarandet.
Bakgrund
I denna förordning anges bestämmelser för ett påskyndande och förtydligande av förfarandet vid alltför stora underskott, vilket definieras redan i artikel 126 i EUF-fördraget.
Avsikten är att förhindra allvarliga finanspolitiska misstag som kan äventyra de offentliga finansernas hållbarhet och potentiellt även hota EMU.
Medlemsstaterna har därför en skyldighet att undvika alltför stora offentliga underskott, vilka fastställs enligt två huvudkriterier: underskott och skuld.
Enligt kommissionens motivering
Se fotnot 1, motiveringen. är det nödvändigt med en reform av den korrigerande delen av stabilitets- och tillväxtpakten för att bemöta ett antal brister som blivit uppenbara i och med den ekonomiska och finansiella krisen.
Följaktligen är förslaget särskilt inriktat på följande åtgärder:
– ” Skuldkriteriet i förfarandet vid alltför stora underskott måste bli tillämpligt i praktiken […]. ”
Skuldutvecklingen ska följas mer noggrant och jämställas med underskottsutvecklingen.
Den föreslagna rättsliga grunden
Protokollet om förfarandet vid alltför stora underskott, som är fogat till fördragen, innehåller ytterligare bestämmelser om genomförandet av det förfarande som beskrivs i denna artikel.
Rådet ska enhälligt, i enlighet med ett särskilt lagstiftningsförfarande och efter att ha hört Europaparlamentet och Europeiska centralbanken, anta lämpliga bestämmelser som därefter ska ersätta det nämnda protokollet.
Om inte annat följer av övriga bestämmelser i denna punkt ska rådet, på förslag av kommissionen och efter att ha hört Europaparlamentet, fastställa närmare regler och definitioner för tillämpningen av bestämmelserna i det nämnda protokollet.
Artikel 136
1.
a) stärka samordningen och övervakningen av dessa staters budgetdisciplin,
b) för dessa medlemsstater utarbeta riktlinjer för den ekonomiska politiken och se till att de överensstämmer med de riktlinjer som har antagits för hela unionen, samt se till att de övervakas.
2.
När det gäller de åtgärder som avses i punkt 1 får endast de rådsmedlemmar delta i omröstningen som företräder medlemsstater som har euron som valuta.
Domstolens synsätt
Enligt rättspraxis ska en åtgärd, i princip, baseras på bara en rättslig grund.
Om bedömningen av en unionsåtgärd visar att det finns två avsikter med densamma eller att den har två beståndsdelar, och om en av dessa kan identifieras som den huvudsakliga eller avgörande avsikten eller beståndsdelen, medan den andra endast är av underordnad betydelse, måste åtgärden ha en enda rättslig grund, nämligen den som krävs med hänsyn till den huvudsakliga eller avgörande avsikten eller beståndsdelen
Mål C-91/05, kommissionen mot rådet, REG 2008, s.
I-3651. .
Endast om det visas att det finns flera avsikter med den aktuella åtgärden eller att den har flera beståndsdelar, vilka har ett sådant samband att de inte kan åtskiljas, utan att den ena är sekundär och indirekt i förhållande till den andra, ska en sådan rättsakt i undantagsfall antas med stöd av de däremot svarande olika rättsliga grunderna.
I-4829.
Analys av den rättsliga grunden
Artikel 126 är en del av avdelning VIII i kapitel I i EUF-fördraget som handlar om ekonomisk politik.
Däri anges vilka steg som ska följas av kommissionen och rådet när dessa tillämpar förfarandet vid alltför stora underskott (underskottsförfarandet).
Kapitel 4 i avdelning VIII innehåller särskilda bestämmelser för de medlemsstater som har euron som valuta.
Enligt artikel 136 får rådet sålunda besluta om särskilda åtgärder för de medlemsstater som har euron som valuta, närmare bestämt att
– stärka samordningen och övervakningen av dessa staters budgetdisciplin, och
– utarbeta riktlinjer för politiken.
I artikel 136 understryks att dessa åtgärder ska antas ”i enlighet med det tillämpliga förfarandet bland dem som anges i artiklarna 121
För de medlemsstater som har euron som valuta. samt att fastställa närmare bestämmelser för tillämpningen av underskottsförfarandet.
Analys av förslaget.
De föreslagna åtgärdernas syfte och innehåll
Som vi har sett ska en lagstiftningsåtgärd i princip ha en enda rättslig grund.
Endast om det visas att det finns flera avsikter med den aktuella åtgärden eller att den har flera beståndsdelar, vilka har ett sådant samband att de inte kan åtskiljas, utan att den ena är sekundär och indirekt i förhållande till den andra, ska en sådan rättsakt i undantagsfall antas med stöd av de däremot svarande olika rättsliga grunderna.
Mål C-91/05, kommissionen mot rådet, REG 2008, s.
I-3651.
Det föreliggande förslaget syftar till att förändra och förbättra den mekanism som inrättats genom förordning (EG) nr 1467/97 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott.
I sin motivering beskriver kommissionen de viktigaste punkterna för den planerade reformen enligt följande:
b) Det införs en rad nya finansiella sanktioner för medlemsstater i euroområdet, som ska avskräcka från alltför stora underskott i de offentliga finanserna och, i de fall det ändå uppstår sådana, bidra till att de omgående korrigeras.
c) En tydligare och flexiblare ram för kommissionens eventuella rekommendationer.
Av detta framgår att de huvudsakliga ändamålen med förslaget är att avskräcka från och korrigera alltför stora underskott, förhindra allvarliga finanspolitiska misstag samt att fastställa närmare bestämmelser för tillämpningen av förfarandet vid alltför stora underskott.
I skäl 14 i ingressen står det: ” För att säkerställa att deltagande medlemsstater följer unionens ramverk för den finanspolitiska tillsynen, bör regelbaserade sanktioner utformas utifrån artikel 136 i fördraget ”.
Även om det förefaller som att regelbaserade sanktioner är en viktig del av det system som föreslås, och att de bidrar till ett effektivt verkställande av underskottsförfarandet, finns det inget fog för att detta skulle utgöra huvudsyftet med den föreslagna förordningen.
Slutsats
YTTRANDE från utskottet för sysselsättning och sociala frågor
till utskottet för ekonomi och valutafrågor
över förslaget till rådets förordning om ändring av förordning (EG) nr 1467/97 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott
( KOM(2010)0522 – C7-0396/2010 – 2010/0276(CNS) )
Föredragande:
David Casa
KORTFATTAD MOTIVERING
Bakgrund
Den 29 september 2010 presenterade kommissionen ett lagstiftningspaket i syfte att förstärka den ekonomiska styrningen inom EU och euroområdet.
Paketet består av sex förslag: fyra av dem behandlar de offentliga finanserna och innefattar en reform av stabilitets- och tillväxtpakten medan målet med de två nya förordningarna är att kartlägga och ta itu med framväxande makroekonomiska obalanser inom EU och euroområdet.
Kommissionen föreslår att medlemsstaternas efterlevnad av stabilitets- och tillväxtpakten förstärks och att samordningen av finanspolitiken skärps.
I den så kallade preventiva delen av stabilitets- och tillväxtpakten har den nuvarande förordningen (EG) nr 1466/97 om ”förstärkning av övervakningen av de offentliga finanserna samt övervakningen och samordningen av den ekonomiska politiken” ändrats i syfte att se till att medlemsstaterna följer en ”försiktig och ansvarsfull” finanspolitik under ekonomiskt goda tider för att bygga upp en nödvändig buffert inför sämre tider.
I den så kallade korrigerande delen har dessutom ändringsförslag till förordning (EG) nr 1467/97 om ”förfarandet vid alltför stora underskott” lagts fram för att se till att skuldutvecklingen följs mer noggrant och jämställs med underskottsutvecklingen.
Vidare har ett direktiv med krav på medlemsstaternas budgetramar lagts fram för att uppmuntra till ansvar för de offentliga finanserna genom att sätta upp minimikrav för nationella finansramar och se till att de är förenliga med förpliktelserna enligt fördraget.
För att stödja ändringarna i de preventiva och korrigerande delarna av stabilitets- och tillväxtpakten föreslog kommissionen också en skärpning av tillsynsmekanismerna för medlemsstaterna i euroområdet.
Iakttagelser
Detta förslag till yttrande berör kommissionens förslag om ändring av förordning (EG) nr 1467/97 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott, till vilket föredraganden föreslår följande ändringar:
- Förstärkningen av övervakningen av de offentliga finanserna bör alltid lyda under EU:s övergripande mål, och särskilt under kraven i artikel 9 i fördraget om Europeiska unionens funktionssätt, som hör samman med främjandet av en hög sysselsättningsnivå, garantier för ett fullgott socialt skydd och kampen mot social utestängning.
- Vid övervakningen av överensstämmelsen med reglerna om budgetdisciplin och då beslut fattas i detta syfte bör särskild hänsyn tas inte enbart till allvarliga ekonomiska utan också sociala nedgångar som kan påverka regeringarnas finansiella ställning.
- Möjligheten för medlemsstater som genomför strukturreformer att avvika från sina respektive medelfristiga budgetmål bör inte vara kopplad till pensionsreformer som syftar till att främja vissa modeller.
Denna möjlighet bör i stället beviljas för de medlemsstater som genomför strukturreformer som bidrar till att bevara eller skapa arbetstillfällen och till att minska fattigdomen.
- De böter som drivits in från medlemsstater som inte efterlever sina respektive rekommendationer bör användas till att stödja EU:s långsiktiga investeringar och sysselsättningsmål och inte enbart utdelas till medlemsstater som inte omfattas av något förfarande vid alltför stora underskott, såsom kommissionen föreslår.
- Förstärkningen av den ekonomiska styrningen bör gå hand i hand med en skärpning av den demokratiska legitimiteten för den europeiska styrningen.
Europaparlamentets roll bör i detta sammanhang stärkas för hela övervakningsprocessen.
Regelbundna samråd med arbetsmarknadens parter och ett utökat deltagande för de nationella parlamenten är även en förutsättning för en trovärdig och transparent övervakningsram.
ÄNDRINGSFÖRSLAG
Utskottet för sysselsättning och sociala frågor uppmanar utskottet för ekonomi och valutafrågor att som ansvarigt utskott infoga följande ändringsförslag i sitt betänkande:
Ändringsförslag
1
Förslag till förordning – ändringsakt
Skäl 1
Kommissionens förslag
Ändringsförslag
(1) Samordningen av medlemsstaternas ekonomiska politik inom unionen bör enligt fördraget innebära att man följer riktlinjerna om stabila priser, sunda offentliga finanser och monetära förhållanden samt en stabil betalningsbalans.
(1) Samordningen av medlemsstaternas ekonomiska politik inom unionen bör enligt fördraget om Europeiska unionens funktionssätt innebära att man följer riktlinjerna om hög sysselsättningsnivå och social sammanhållning, stabila priser, sunda offentliga finanser och monetära förhållanden samt en stabil betalningsbalans.
Ändringsförslag
2
Förslag till förordning – ändringsakt
Skäl 1a (nytt)
Kommissionens förslag
Ändringsförslag
(1a) I fördraget om Europeiska unionens funktionssätt föreskrivs att unionen, vid fastställandet och genomförandet av sin politik och verksamhet, ska beakta de krav som är förknippade med främjandet av hög sysselsättningsnivå, garantier för ett fullgott socialt skydd och kampen mot social utestängning.
Ändringsförslag
3
Förslag till förordning – ändringsakt
Skäl 1b (nytt)
Kommissionens förslag
Ändringsförslag
Ändringsförslag
4
Förslag till förordning – ändringsakt
Skäl 3
Kommissionens förslag
Ändringsförslag
(3) Stabilitets- och tillväxtpakten grundas på målet om sunda offentliga finanser, som ett sätt att stärka förutsättningarna för prisstabilitet och stark varaktig tillväxt som kan bidra till ökad sysselsättning.
(3) Stabilitets- och tillväxtpakten grundas på målet om sunda offentliga finanser, som ett sätt att stärka förutsättningarna för prisstabilitet och stark varaktig tillväxt som kan bidra till ökad sysselsättning , och den bör därför främja långsiktiga investeringar till förmån för en smart och hållbar tillväxt som inbegriper alla .
Ändringsförslag
5
Förslag till förordning – ändringsakt
Skäl 4a (nytt)
Kommissionens förslag
Ändringsförslag
(4a) Den stärkta övervakningen av de offentliga finanserna bör dock bidra till unionens tillväxt- och sysselsättningsmål och bör vid en allvarlig konjunkturnedgång eller en betydande ökning av arbetslösheten kombineras med insatser för att stimulera ekonomin, skydd och skapande av sysselsättning och social sammanhållning, samtidigt som medlemsstaternas särskilda prioriteringar och behov respekteras.
Ändringsförslag
6
Förslag till förordning – ändringsakt
Skäl 4b (nytt)
Kommissionens förslag
Ändringsförslag
(4b) Förstärkningen av den ekonomiska styrningen bör gå hand i hand med en skärpning av den demokratiska legitimiteten för europeisk styrning, vilket bör uppnås genom att Europaparlamentet och de nationella parlamenten i högre utsträckning och vid rätt tidpunkt deltar under hela förfarandena för samordningen av den ekonomiska politiken, och till fullo utnyttjar de instrument som fastställs i EUF ‑fördraget, särskilt de allmänna riktlinjerna för medlemsstaternas och unionens ekonomiska politik och riktlinjerna för medlemsstaternas sysselsättningspolitik.
Ändringsförslag
7
Förslag till förordning – ändringsakt
Skäl 12
Kommissionens förslag
Ändringsförslag
(12) Vid bedömningen av om tidsfristen bör förlängas för att korrigera ett alltför stort underskott, bör särskild hänsyn tas till omfattande och allvarliga konjunkturnedgångar .
(12) Vid bedömningen av om tidsfristen bör förlängas för att korrigera ett alltför stort underskott, bör särskild hänsyn tas till en allvarlig konjunkturnedgång eller en betydande ökning av arbetslösheten .
Ändringsförslag
8
Förslag till förordning – ändringsakt
Kommissionens förslag
Ändringsförslag
”1.
”1.
Ändringsförslag
9
Förslag till förordning – ändringsakt
Förordning (EG) nr 1467/97
Kommissionens förslag
Ändringsförslag
”1a.
Under en treårsperiod från och med den [date of entering into force of this Regulation - to be inserted] ska denna indikators retroaktiva natur beaktas vid tillämpningen.”
”1a.
Under en treårsperiod från och med den ...* ska denna indikators retroaktiva natur beaktas vid tillämpningen.”
____________
* EUT – för in datumet för denna förordnings ikraftträdande.
Ändringsförslag
10
Förslag till förordning – ändringsakt
Förordning (EG) nr 1467/97
Kommissionens förslag
Ändringsförslag
”3.
Rapporten ska på lämpligt sätt ta upp det ekonomiska lägets utveckling på medellång sikt (särskilt tillväxtpotential, rådande konjunkturförhållanden, inflation, alltför stora makroekonomiska obalanser) samt utvecklingen av de offentliga finanserna på medellång sikt (särskilt ansträngningar att konsolidera finanserna under ”goda tider”, offentliga investeringar, politiskt genomförande av unionens gemensamma tillväxtstrategi och de offentliga finansernas allmänna kvalitet, särskilt då följandet av rådets direktiv […] om krav på medlemsstaternas finanspolitiska ramverk).
Rapporten ska vid behov också innehålla en analys av skuldställningen på medellång sikt (särskilt belysa riskfaktorer adekvat, inklusive skuldernas löptids- och valutastruktur, stock-/flödesjusteringar, ackumulerade reserver och andra offentliga tillgångar; garantier särskilt till finanssektorn; till åldrandet både explicit och implicit relaterade skulder samt privata skulder om de implicit utgör eventualförpliktelser för den offentliga sektorn).
Dessutom ska kommissionen vederbörligen beakta eventuella andra faktorer som enligt den berörda medlemsstaten har betydelse för en samlad kvalitativ bedömning av överskridandet av referensvärdet och som medlemsstaten har förelagt kommissionen och rådet.
I detta sammanhang ska särskild hänsyn tas till budgetmässiga ansträngningar för att främja internationell solidaritet och uppnå unionens politiska mål, inklusive finansiell stabilitet.”
”3.
Rapporten ska på lämpligt sätt ta upp det sociala och ekonomiska lägets utveckling på medellång sikt (särskilt tillväxtpotential, rådande konjunkturförhållanden, fattigdomsnivå, inkomstklyftor, arbetslöshet, inflation, alltför stora makroekonomiska obalanser) samt utvecklingen av de offentliga finanserna på medellång sikt (särskilt ansträngningar att konsolidera finanserna under ”goda tider”, offentliga investeringar, politiskt genomförande av unionens strategi för tillväxt och sysselsättning och de offentliga finansernas allmänna kvalitet, särskilt då följandet av rådets direktiv […] om krav på medlemsstaternas finanspolitiska ramverk).
Rapporten ska vid behov också innehålla en analys av skuldställningen på medellång sikt (särskilt belysa riskfaktorer adekvat, inklusive skuldernas löptids- och valutastruktur, stock-/flödesjusteringar, ackumulerade reserver och andra offentliga tillgångar; garantier särskilt till finanssektorn; till åldrandet både explicit och implicit relaterade skulder samt privata skulder om de implicit utgör eventualförpliktelser för den offentliga sektorn).
Dessutom ska kommissionen vederbörligen beakta eventuella andra faktorer som enligt den berörda medlemsstaten har betydelse för en samlad kvalitativ bedömning av överskridandet av referensvärdet och som medlemsstaten har förelagt kommissionen och rådet.
I detta sammanhang ska särskild hänsyn tas till budgetmässiga ansträngningar för att främja internationell solidaritet och uppnå unionens politiska mål, inklusive finansiell stabilitet.”
Ändringsförslag
11
Förslag till förordning – ändringsakt
Förordning (EG) nr 1467/97
”5.
Vid alla budgetbedömningar inom ramen för förfarandet vid alltför stora underskott och förfarandet vid alltför stora skulder ska kommissionen och rådet vederbörligen beakta genomförandet av genomgripande strukturreformer av pensionssystemen eller de sociala trygghetssystemen, som främjar unionens tillväxtmål, eller reformer som genomförs till följd av rådets rekommendationer i enlighet med artikel 121 i EUF-fördraget.”
Ändringsförslag
12
Förslag till förordning – ändringsakt
Förordning (EG) nr 1467/97
Kommissionens förslag
Ändringsförslag
”7.
Om skuldkvoten överskrider referensvärdet, ska reformens kostnad bara beaktas om underskottet ligger nära referensvärdet.
För detta ändamål ska under fem år från och med reformens ikraftträdande dess nettokostnads påverkan på underskotts- och skuldutvecklingen beaktas enligt en linjär degressiv skala.
Det ska också beaktas om denna nettokostnad minskar genom att ovannämnda pensionsreform helt eller delvis upphävs.”
”7.
Om skuldkvoten överskrider referensvärdet, ska reformens hela kostnad bara beaktas om underskottet ligger nära referensvärdet.
För detta ändamål ska , från och med reformens ikraftträdande , dess nettokostnads påverkan på underskotts- och skuldutvecklingen beaktas enligt en linjär degressiv skala.
Det ska också beaktas om denna nettokostnad minskar genom att ovannämnda pensionsreformer helt eller delvis upphävs.”
Ändringsförslag
13
Förslag till förordning – ändringsakt
Förordning (EG) nr 1467/97
Kommissionens förslag
Ändringsförslag
”4.
I rådets rekommendation ska det även fastställas en tidsfrist för korrigeringen av det alltför stora underskottet, vilken ska slutföras under det år som följer på året då underskottet fastställdes, om inte särskilda omständigheter föreligger.
I rekommendationen ska rådet begära att medlemsstaten uppnår årliga budgetmål som enligt rekommendationens underliggande prognos som ett riktmärke motsvarar en årlig minsta förbättring på minst 0,5 % av BNP av sitt konjunkturrensade saldo, utan engångsåtgärder och tillfälliga åtgärder, för att korrigera det alltför stora underskottet inom tidsfristen i rekommendationen.”
”4.
I rådets rekommendation ska det även fastställas en tidsfrist för korrigeringen av det alltför stora underskottet, vilken ska slutföras under det år som följer på året då underskottet fastställdes, om inte särskilda omständigheter föreligger.
I rekommendationen ska rådet, samtidigt som full hänsyn tas till artikel 9 i EUF ‑fördraget, särskilt när det gäller främjande av hög sysselsättningsnivå, garantier för ett fullgott socialt skydd och kampen mot social utestängning, och till unionens tillväxt- och sysselsättningsmål, begära att medlemsstaten uppnår årliga budgetmål som enligt rekommendationens underliggande prognos som ett riktmärke motsvarar en årlig minsta förbättring på minst 0,5 % av BNP av sitt konjunkturrensade saldo, utan engångsåtgärder och tillfälliga åtgärder, för att korrigera det alltför stora underskottet inom tidsfristen i rekommendationen.”
Ändringsförslag
14
Förslag till förordning – ändringsakt
Förordning (EG) nr 1467/97
Kommissionens förslag
Ändringsförslag
”5.
Rådet ska bedöma om det, jämfört med de ekonomiska prognoserna i sin rekommendation, föreligger oväntade negativa ekonomiska händelser med stora negativa effekter för de offentliga finanserna.
”5.
Rådet ska bedöma om det, jämfört med de ekonomiska prognoserna i sin rekommendation, föreligger oväntade negativa ekonomiska eller sociala händelser med stora negativa effekter för de offentliga finanserna.
Ändringsförslag
15
Förslag till förordning – ändringsakt
Kommissionens förslag
Ändringsförslag
”1.
I föreläggandet ska rådet begära att medlemsstaten uppnår årliga budgetmål som enligt rekommendationens underliggande prognos som ett riktmärke motsvarar en årlig minsta förbättring på minst 0,5 % av BNP av sitt konjunkturrensade saldo, utan engångsåtgärder och tillfälliga åtgärder, för att korrigera det alltför stora underskottet inom tidsfristen i rekommendationen.
Rådet ska också ange åtgärder som främjar att dessa mål uppnås.”
”1.
I föreläggandet ska rådet begära att medlemsstaten uppnår årliga budgetmål som enligt rekommendationens underliggande prognos som ett riktmärke motsvarar en årlig minsta förbättring på minst 0,5 % av BNP av sitt konjunkturrensade saldo, utan engångsåtgärder och tillfälliga åtgärder, för att korrigera det alltför stora underskottet inom tidsfristen i rekommendationen.
Rådet ska också ange åtgärder som främjar att dessa mål uppnås.”
Ändringsförslag
16
Förslag till förordning – ändringsakt
Kommissionens förslag
Ändringsförslag
”2.
”2.
Rådet ska bedöma om det, jämfört med de ekonomiska prognoserna i sitt föreläggande, föreligger oväntade negativa ekonomiska eller sociala händelser med stora negativa effekter för de offentliga finanserna.
Ändringsförslag
17
Förslag till förordning – ändringsakt
Kommissionens förslag
Ändringsförslag
2.
2.
Ändringsförslag
18
Förslag till förordning – ändringsakt
Förordning (EG) nr 1467/97
Artikel 7
Kommissionens förslag
Ändringsförslag
7.
7.
Artikel 7 ska ersättas med följande:
”7.
Ett påskyndat förfarande ska användas om det rör sig om ett avsiktligt planerat underskott som enligt rådets beslut är alltför stort.”
Ändringsförslag
19
Förslag till förordning – ändringsakt
Förordning (EG) nr 1467/97
Artikel 8
Kommissionens förslag
Ändringsförslag
Ändringsförslag
20
Förslag till förordning – ändringsakt
Kommissionens förslag
Ändringsförslag
1a .
Kommissionen och rådet ska rapportera sina resultat i enlighet med punkt 1 till Europaparlamentet.
Ändringsförslag
21
Förslag till förordning – ändringsakt
Förordning (EG) nr 1467/97
Artikel 16
Kommissionens förslag
Ändringsförslag
De böter som anges i artikel 12 i denna förordning ska utgöra andra inkomster enligt artikel 311 i fördraget om Europeiska unionens funktionssätt och ska användas genom en unionsmekanism för finansiell stabilitet till stöd för unionens långsiktiga investerings- och sysselsättningsmål .”
ÄRENDETS GÅNG
Titel
Ändring av rådets förordning (EG) nr 1467/97 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott
Referensnummer
KOM(2010)0522 – C7-0396/2010 – 2010/0276(CNS)
Ansvarigt utskott
ECON
Yttrande
Tillkännagivande i kammaren
EMPL
13.12.2010
Föredragande av yttrande
Utnämning
David Casa
21.10.2010
Behandling i utskott
1.12.2010
25.1.2011
Antagande
16.3.2011
Slutomröstning: resultat
+:
–:
0:
39
4
1
Slutomröstning: närvarande ledamöter
Regina Bastos, Edit Bauer, Jean-Luc Bennahmias, Pervenche Berès, Mara Bizzotto, Philippe Boulland, David Casa, Alejandro Cercas, Marije Cornelissen, Frédéric Daerden, Karima Delli, Proinsias De Rossa, Frank Engel, Sari Essayah, Richard Falbr, Ilda Figueiredo, Nadja Hirsch, Stephen Hughes, Liisa Jaakonsaari, Danuta Jazłowiecka, Martin Kastler, Ádám Kósa, Patrick Le Hyaric, Veronica Lope Fontagné, Olle Ludvigsson, Elizabeth Lynne, Thomas Mann, Elisabeth Morin-Chartier, Csaba Őry, Rovana Plumb, Konstantinos Poupakis, Sylvana Rapti, Licia Ronzulli, Elisabeth Schroedter, Jutta Steinruck, Traian Ungureanu
Slutomröstning: närvarande suppleanter
Georges Bach, Raffaele Baldassarre, Sven Giegold, Thomas Händel, Antigoni Papadopoulou, Evelyn Regner
Slutomröstning: närvarande suppleanter (art.
187.2)
Liam Aylward, Fiona Hall
ÄRENDETS GÅNG
Titel
Ändring av rådets förordning (EG) nr 1467/97 om påskyndande och förtydligande av tillämpningen av förfarandet vid alltför stora underskott
Referensnummer
KOM(2010)0522 – C7-0396/2010 – 2010/0276(CNS)
Begäran om samråd med parlamentet
29.11.2010
Ansvarigt utskott
Tillkännagivande i kammaren
ECON
13.12.2010
Rådgivande utskott
Tillkännagivande i kammaren
BUDG
13.12.2010
EMPL
13.12.2010
Inget yttrande avges
Beslut
BUDG
20.10.2010
Föredragande
Utnämning
Diogo Feio
21.9.2010
Bestridande av den rättsliga grunden
JURI:s yttrande
JURI
12.4.2011
Behandling i utskott
26.10.2010
24.1.2011
22.3.2011
Antagande
19.4.2011
Slutomröstning: resultat
+:
–:
0:
29
7
10
Slutomröstning: närvarande ledamöter
Burkhard Balz, Sharon Bowles, Udo Bullmann, Nikolaos Chountis, George Sabin Cutaş, Rachida Dati, Leonardo Domenici, Derk Jan Eppink, Diogo Feio, Elisa Ferreira, Vicky Ford, Ildikó Gáll-Pelcz, José Manuel García-Margallo y Marfil, Jean-Paul Gauzès, Sven Giegold, Sylvie Goulard, Liem Hoang Ngoc, Wolf Klinz, Jürgen Klute, Rodi Kratsa-Tsagaropoulou, Philippe Lamberts, Astrid Lulling, Arlene McCarthy, Íñigo Méndez de Vigo, Ivari Padar, Alfredo Pallone, Anni Podimata, Antolín Sánchez Presedo, Olle Schmidt, Edward Scicluna, Peter Simon, Theodor Dumitru Stolojan, Ivo Strejček, Kay Swinburne, Marianne Thyssen, Ramon Tremosa i Balcells, Corien Wortmann-Kool
Slutomröstning: närvarande suppleanter
Marta Andreasen, Herbert Dorfmann, Robert Goebbels, Carl Haglund, Krišjānis Kariņš, Barry Madlener, Thomas Mann, Claudio Morganti, Andreas Schwab
Slutomröstning: närvarande suppleanter (art.
187.2)
Karima Delli
Ingivande
2.5.2011
A7-0194/2011
***
REKOMMENDATION
om utkastet till rådets beslut om ingående av protokollet om fastställande av de fiskemöjligheter och den ekonomiska ersättning som föreskrivs i partnerskapsavtalet om fiske mellan Europeiska unionen och Demokratiska Republiken São Tomé e Príncipe
(05371/2011 – – C7‑0119/2011 – 2010/0355(NLE))
Fiskeriutskottet
Föredragande:
Luis Manuel Capoulas Santos
PE 458.638v02-00
Teckenförklaring
* Samrådsförfarandet
*** Besiktningsförfarande
***I Ordinarie lagstiftningsförfarande (första behandlingen)
***II Ordinarie lagstiftningsförfarande (andra behandlingen)
***III Ordinarie lagstiftningsförfarande (tredje behandlingen)
(Det angivna förfarandet baseras på den rättsliga grund som angetts i förslaget till akt.)
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING............................................................................................................................6
YTTRANDE från utskottet för utveckling ........................................................11
YTTRANDE från budgetutskottet ............................................................................15
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................19
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om utkastet till rådets beslut om ingående av protokollet om fastställande av de fiskemöjligheter och den ekonomiska ersättning som föreskrivs i partnerskapsavtalet om fiske mellan Europeiska unionen och Demokratiska Republiken São Tomé e Príncipe .
(05371/2011 – C7-0119/2011 – 2010/0355(NLE) )
(Godkännande)
Europaparlamentet utfärdar denna resolution
– med beaktande av utkastet till rådets beslut (05371/2011),
– med beaktande av fiskeriutskottets rekommendation och yttrandena från utskottet för utveckling och budgetutskottet ( A7-0194/2010 ).
1.
2.
Europaparlamentet uppdrar åt talmannen att översända parlamentets ståndpunkt till rådet och kommissionen samt till regeringarna och parlamenten i medlemsstaterna och i Demokratiska republiken São Tomé och Príncipe.
MOTIVERING
Inledning
Förhandlingar om och ingående av partnerskapsavtal om fiske ingår som en del i det allmänna målet att upprätthålla och bevara EU-flottans fiskeverksamhet, även för fjärrfiskeflottan, och att utveckla partnerskap och samarbete med tredjeländer för att främja ett hållbart utnyttjande av fiskeresurserna utanför EU:s vatten samtidigt som hänsyn tas till miljömässiga, sociala och ekonomiska aspekter.
Därför antog Europeiska rådet den 23 juli 2007 förordning (EG) nr 894/2007 om ingående av ett partnerskapsavtal om fiske mellan Demokratiska republiken São Tomé e Príncipe och Europeiska gemenskapen
EUT´L 205, 7.8.2007, s.
35; rättelse i EUT 330, 15.12.2007, s.
60. .
Detta avtal, som är tillämpligt i perioder om fyra år som förlängs automatiskt om inte någon av parterna säger upp avtalet, upphävde och ersatte det första fiskeavtalet som ingicks 1984 mellan EG och São Tomé och Príncipe.
Till gällande partnerskapsavtal från 2006 lades ett protokoll som fastställde fiskemöjligheter och den ekonomiska ersättningen för perioden mellan den 1 juni 2006 och 31 maj 2010, då detsamma löper ut.
Samtidigt med detta förslag till rådets beslut om ingående av det nya protokollet, inledde kommissionen två andra förfaranden: Ett förslag till rådets beslut om undertecknande på unionens vägnar och provisorisk tillämpning av det nya protokollet
De båda förslagen antogs av rådet den 24 februari 2011.
I enlighet med artikel 13 i det nya protokollet ska detta tillämpas provisoriskt från och med den dag det undertecknas av båda parter.
Det nya protokollet undertecknades den 13 maj 2011, dvs. samma dag som rådet förelade parlamentet sin begäran om godkännande.
Analys av det nya protokollet
Huvudinnehållet i det nya protokollet är följande:
– Årlig ekonomisk ersättning: 682 500 euro (med ett totalt belopp på 2 047 500 euro för hela perioden), fördelat enligt följande:
a) ett årligt belopp för tillträdet till São Tomé och Príncipes exklusiva ekonomiska zon på 455 000 euro motsvarande en referensfångstmängd på 7 000 ton per år, och
b) ett specifikt belopp på 227 500 euro per år till stöd för genomförandet av São Tomé och Príncipes sektoriella fiskeripolitik.
Den ekonomiska ersättningen som EU betalar ska öka med 65 euro per ton om EU-fartygens totala fångst överstiger 7 000 ton per år.
– Fiskemöjligheter: tillstånd ges för fiske med 28 notfartyg för tonfiske och 12 fartyg med ytlångrev.
Dessa fiskemöjligheter kommer att kunna justeras upp eller ned utifrån årliga utvärderingar av beståndens tillstånd, vilket också medför att den ekonomiska ersättningen justeras på lämpligt sätt.
Fördelningen av fiskemöjligheterna mellan de berörda medlemsstaterna, som omfattas av en särskild rådets förordning, är följande: notfartyg för tonfiske: Spanien – 16 fartyg; Frankrike – 12 fartyg; fartyg för fiske med ytlångrev: Spanien – 9 fartyg; Portugal – 3 fartyg.
– Förskott och avgifter från fartygsägarna: 35 euro per ton fångad tonfisk i São Tomé och Príncipes fiskezon.
De årliga förskotten ligger på 6 125 euro per notfartyg för tonfiske, vilket motsvarar avgifterna för en årsfångst på 175 ton, och 2 275 euro för ytlångrevsfartyg, vilket motsvarar avgifterna för en årsfångst på 65 ton.
Nedanstående tabell jämför vissa delar av det gamla och det nya protokollet samt utvecklingen av fiskemöjligheternas fördelning mellan medlemsstaterna.
Protokollets giltighetstid
fyra år
1.6.2006–31.5.2010
tre år
2011–2014
Paraferat
25 maj 2006
15 juli 2010
Årlig ekonomisk ersättning
682 500 euro, 227 500 euro av detta belopp är avsatt för São Tomé och Príncipes sektoriella fiskeripolitik
Avgift som ska betalas av fartygsägarna
35 euro per fångstton
35 euro per fångstton
- Notfartyg för tonfiske: 5 250 euro/år (referensfångster: 150 ton)- Fartyg som bedriver ytfiske med långrev: 1 295 euro/år (referensfångster: 55 ton)
- Notfartyg för tonfiske: 6 125 euro/år (referensfångster: 175 ton)
Referenstonnage per år
8 500 ton/år
7 000 ton/år
Erbjudna fiskemöjligheter
Notfartyg för tonfiske (2006/2010)
Fartyg med ytlångrev
(2006/2010)
Fartyg med ytlångrev
(2011/2014)
SPANIEN
13
16
13
9
FRANKRIKE
12
12
PORTUGAL
5
3
TOTALT
25 fartyg
28 fartyg
18 fartyg
12 fartyg
Enligt den utvärderingsrapport som gjordes av oberoende experter
Utvärdering i efterhand av protokollet för 2006–2010 och förhandsbedömning av det framtida protokollet. under det föregående protokollets giltighetstid, var utnyttjande av fiskemöjligheterna bättre för fartyg som fiskar med snörpvad (med ett medeltal på 79 procent) än fartyg med ytlångrev (med ett medeltal på 42 procent).
Mot bakgrund av denna utnyttjandegrad de senaste åren för ytlångrevsfartyg, har fiskemöjligheterna minskats från 18 till 12 fartyg i förhållande till det tidigare protokollet.
En lätt ökning av antalet tillgängliga licenser för kategorin notfartyg har å andra sidan observerats för att kompensera att vissa aktörer den senaste tiden flyttat sin verksamhet från Indiska oceanen till Atlanten på grund av problemen med sjöröveri.
Den genomsnittliga årliga fångstmängden var 1 252 ton mellan 2006 och 2009, en nivå som ligger betydligt under referensfångstmängden.
I det nya protokollet har man därför kunnat konstatera en följdriktig minskning av referensfångstmängden (från 8 500 till 7 000 ton/år), som återspeglar de senaste årens tendens.
Med hänsyn till behoven inom fiskesektorn i Republiken São Tomé och Príncipe har ändå de årliga anslagen för sektorsstöd ökat i jämförelse med de anslag som ursprungligen föreslogs i det förra protokollet.
Även det nya protokollet innehåller en exklusivitetsklausul, något som fanns redan i avtalstexten, och en bättre specificering av innehållet i översyns- och upphävandeklausulerna för betalningen av den ekonomiska ersättningen och för avbrytande av protokollets tillämpning under vissa omständigheter, framför allt om avgörande delar av de mänskliga rättigheterna enligt artikel 9 i Cotonouavtalet har överträtts (artiklarna 8 och 9 i det nya protokollet).
Liksom i det föregående protokollet är fiskezonerna belägna i vatten som ligger mer än 12 sjömil från baslinjerna.
Enligt protokollet ska minst 20 procent av sjömännen som mönstrar på gemenskapsfartygen vara från São Tomé och Príncipe, eller eventuellt från en AVS-stat, och på begäran av São Tomé och Príncipes behöriga myndigheter ska fartygen ta ombord en observatör utsedd av landets fiskeministerium.
Föredragandens anmärkningar och kommentarer
Förhandsutvärderingen kom fram till att fiskeavtalet med São Tomé och Príncipe tillgodoser EU-flottans behov och skulle kunna bidra till att upprätthålla lönsamheten inom EU:s tonfiske i Atlanten, genom att EU:s fartyg och de verksamheter som är beroende av fisket erbjuds en stabil rättslig ram på mellanlång sikt och bidrar till att upprätthålla kontinuiteten i de fiskeområden som omfattas av avtal i Guineabukten.
Det hör till de minst utvecklade länderna, och São Tomé och Príncipes BNP domineras av jordbruk, förädling av jordbruksprodukter och fiske.
Detta tillsammans med beroendet av livsmedelsimport, leder till ett underskott i handelsbalansen och ett beroende av utländskt stöd.
São Tomé och Príncipes fiske är koncentrerat på kustresurserna och producerar nära 4 000 ton fisk per år.
Omkring 15 procent av den aktiva befolkningen är fortfarande beroende av fisket för sin försörjning.
Denna resurs utgör 74 procent av den animaliska proteinkonsumtionen i São Tomé och Príncipe.
Enligt efterhandsutvärderingen har betydande framsteg gjorts när det gäller kontroll och övervakning av fisket (de första stegen har tagits för att inrätta ett satellitövervakningssystem för fartyg, en ny rättslig grund har skapats för att upprätta ett fartygsregister och förvalta det), och São Tomé och Príncipe deltar och syns i högre grad i regionala eller underregionala organisationer som internationella kommissionen för bevarandet av tonfisk (Iccat) och den regionala kommittén för fiske i Guineabukten (Corep).
Utvärderingen kom också fram till att mer än 50 procent av EU:s ekonomiska ersättning har anslagits till budgeten för São Tomé och Príncipes fiskerimyndighet, vilket ligger i linje med São Tomé och Príncipes myndigheters åtagande i det föregående protokollet.
Alla arter som fiskas av gemenskapsfartygen är migrerande arter.
Avtalet bidrar i allmänhet med nära 0,36 procent av de totala fångstmängderna av de artbestånd som fisket riktas mot, och inga fångster av gemenskapsfartyg inom ramen för avtalet utnyttjar mer än 0,55 procent av den totala fångstmängden av artbestånden i fråga.
Enligt utvärderingsrapporten håller sig utnyttjandet av arter som gulfenad tonfisk, bonit och svärdfisk inom gränserna för hållbarhet.
Det råder en viss osäkerhet om eventuella negativa effekter för vissa arter, men avtalets påverkan på situationen i allmänhet är minimal, och det betraktas som hållbart och i linje med Iccats rekommendationer.
När det gäller förfarandet framhåller föredraganden det negativa i att inget av kommissionens förslag för det nya protokollet antogs förrän den 13 december 2010, nära sex månader efter att det paraferades.
Detta har försenat förfarandets avslutning och dess provisoriska tillämpning vilket har lett till ett förlängt verksamhetsuppehåll för gemenskapsflottan i detta område eftersom också tidsperioden på sex månader, enligt artikel 9 i rådets förordning (EG) nr 1006/2008 av den 29 september 2008, löpt ut
EUT L 286, 29.10.2008, s.
33. .
Slutsatser
Föreliggande förslag gagnar väsentligen båda parter, och föredraganden rekommenderar därför att det antas.
Föredraganden uppmanar emellertid kommissionen att förelägga parlamentet slutsatserna från de möten och överläggningar som hållits i den gemensamma kommitté som avses i avtalet samt det sektorsprogram för fiske som nämns i protokollet tillsammans med resultaten av de årliga utvärderingarna.
till fiskeriutskottet
över förslaget till rådets beslut om ingående av ett nytt protokoll om fastställande av de fiskemöjligheter och den ekonomiska ersättning som föreskrivs i partnerskapsavtalet om fiske mellan Demokratiska Republiken São Tomé e Príncipe och Europeiska gemenskapen
( KOM(2010)0735 – C7‑…/2011 – 2010/0355(NLE) )
Föredragande: Isabella Lövin
KORTFATTAD MOTIVERING
Fiskeavtalet mellan Europeiska gemenskapen och Demokratiska republiken São Tomé e Príncipe löpte ut den 31 maj 2010.
Möjligheten att inte ge sitt godkännande ska ses som en sista utväg och styrkas av bevis för att avtalets tillämpningsområde inte respekteras på vederbörligt sätt, såvida inte parlamentet nekar till ingående av ett protokoll av andra orsaker.
Enligt förslaget till avtal förbinder sig parterna till en partnerskapsram, som underlättar utvecklingen av en hållbar fiskeripolitik och ett ansvarsfullt utnyttjande av fiskeresurserna i Demokratiska republiken São Tomé e Príncipes fiskeområde, vilket är i båda parternas intresse.
Texten till det nya protokollet är förenlig med parternas önskan om att stärka partnerskapet och samarbetet inom fiskerisektorn med hjälp av samtliga tillgängliga finansiella instrument.
Det ekonomiska bidraget uppgår till 2 047 500 euro under de tre år som detta protokoll är giltigt.
Beloppet omfattar
· 455 000 euro per år, vilket motsvarar en referensfångstmängd på 7 000 ton per år för 40 fartyg, och
· 227 500 euro per år, vilket motsvarar EU:s stöd till den sektoriella fiskeripolitiken i Demokratiska republiken São Tomé e Príncipe.
Till detta måste summan som fartygsägarna betalar läggas till – licensavgifter på 6 125 euro för notfartyg och 2 275 euro för fartyg med ytlångrev, samt 35 euro per ton tonfisk som fångats i São Tomé e Príncipes exklusiva ekonomiska zon.
São Tomé e Príncipe får 100 euro per ton fångad tonfisk, med en garanterad utbetalning för minst 7 000 ton per år, samt ytterligare finansiering för att utveckla den nationella fiskerisektorn.
Om EU-fartygens totala fångst i São Tomé e Príncipes vatten överstiger 7 000 ton per år ska den ekonomiska ersättningen som EU betalar ökas med 65 euro per ton, och fartygsägarna ska betala 35 euro per ton.
Om den kvantitet som fångas av EU:s fartyg överstiger den kvantitet som motsvarar det dubbla totala årsbeloppet, ska det utestående beloppet för den överskjutande kvantiteten betalas det påföljande året.
För utvecklingsländer kan detta vara problematiskt av flera anledningar.
En genomläsning av avtalets utvärdering tyder på att följande punkter bör beaktas vid genomförandet av avtalet:
· São Tomé e Príncipe är ett föga utvecklat och ytterst skuldsatt land.
74 procent av det animaliska proteinet utgörs av fisk i den nationella kosten.
· Fiskerimyndigheten och fiskeförvaltningen är fortfarande svaga och utvecklingen av fisket i São Tomé e Príncipe bristfällig, även efter det att landet fått ekonomiskt stöd från det senaste partnerskapsavtalet om fiske, vilket beskrivs i avtalets utvärdering.
· De fartyg som ägs av europeiska aktörer och som är under Ekvatorialguineas och Gabons flagg, har privata licenser i São Tomé e Príncipes vatten.
Detta bör undersökas av kommissionen, eftersom det försvagar exklusivitetsklausulen i partnerskapsavtalet om fiske.
· Fördelarna med avtalet för São Tomé e Príncipe är begränsade till det ekonomiska stödet, eftersom det enligt utvärderingen varken finns landningsplatser, hamnbesök, lokal sysselsättning eller några andra ekonomiska fördelar.
· Inga observatörer har mobiliserats på EU:s fartyg och det finns en viss oro över huruvida EG-fartygen uppfyller rapporteringskraven.
· Vissa av de fångade arterna är särskilt utsatta, särskilt storögd tonfisk och makohaj.
Det finns också anledning till oro över fiske med långrev med stora bifångster av sjöfåglar och sköldpaddor som följd.
Avtalet har dock medfört betydande stöd till budgeten för São Tomé e Príncipes fiskerimyndighet.
En flottförteckning har upprättats och kontrollen har förbättrats.
De första stegen mot ett satellitbaserat kontrollsystem för fartyg har tagits.
I utvärderingen framgår det att även om den övergripande utvärderingen har varit långsam, och många områden kvarstår att behandla, bör avtalets bidrag vid tillhandahållandet av budgetstöd för dessa genomföranden inte underskattas av parterna.
******
Utskottet för utveckling uppmanar fiskeriutskottet att som ansvarigt utskott föreslå att kommissionens förslag godkänns.
Utskottet för utveckling anser att kommissionen på vederbörligt sätt bör ta följande punkter i beaktande vid genomförandet av avtalet:
a) Insynen i förfarandena för att fastställa den totala fångsten bör förbättras, liksom åtgärderna för att bekämpa olagligt, orapporterat och oreglerat fiske (IUU), särskilt genom förbättrad infrastruktur för kontroll och övervakning av fisket i São Tomé e Príncipes exklusiva ekonomiska zon, i syfte att trygga ett ansvarsfullt och hållbart fiske.
b) De europeiska fiskefartygens tillgång till återstoden av den tillåtna fångstmängden av fiskeresurser bör begränsas och vara förenlig med måttet maximalt hållbara avkastning, efter det att lokalbefolkningens näringsbehov mötts.
c) Hållbara fiskemetoder bör främjas genom att det säkerställs att all fiskeverksamhet som omfattas av partnerskapsavtalet om fiske uppfyller samma hållbarhetskriterier som fiskeverksamheten i EU:s farvatten.
d) Det bör, vad gäller korruptionsproblemen, inte finnas några som helst tvivel om ordningens integritet.
e) Den lokala regeringens ansvar bör utökas och måste också garantera förbättrade levnadsvillkor för lokala fiskare, utveckling av lokalt, hållbart, småskaligt fiske och lokala, bärkraftiga beredningsföretag samt efterlevnaden av miljöstandarder.
f) De miniminormer och villkor som fastställts på regional nivå, såsom de avseende bordning av observatörer och rapporteringskrav, ska respekteras.
g) Årliga rapporter om genomförandet av avtalet bör utarbetas och skickas till parlamentet och rådet, i syfte att främja insynen och säkerställa att de extra anslagen för att stödja den sektoriella fiskeripolitiken används för just detta ändamål.
h) Både andemeningen och ordalydelsen i exklusivitetsklausulen bör följas.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
2.5.2011
Slutomröstning: resultat
+:
–:
0:
23
Slutomröstning: närvarande ledamöter
Thijs Berman, Corina Creţu, Leonidas Donskis, Charles Goerens, Catherine Grèze, Eva Joly, Miguel Angel Martínez Martínez, Gay Mitchell, Norbert Neuser, Bill Newton Dunn, Maurice Ponga, Birgit Schnieber-Jastram, Alf Svensson, Eleni Theocharous, Ivo Vajgl
Slutomröstning: närvarande suppleanter
Kriton Arsenis, Proinsias De Rossa, Agustín Díaz de Mera García Consuegra, Enrique Guerrero Salom, Martin Kastler, Krzysztof Lisek, Csaba Őry, Bart Staes
Slutomröstning: närvarande suppleanter (art.
187.2)
Edit Bauer
till fiskeriutskottet
över utkastet till rådets beslut om ingående av ett nytt protokoll om fastställande av de fiskemöjligheter och den ekonomiska ersättning som föreskrivs i partnerskapsavtalet om fiske mellan Demokratiska Republiken São Tomé e Príncipe och Europeiska gemenskapen
( KOM(2010)0735 – C7‑.../2011 – 2010/0355(NLE) )
Föredragande: François Alfonsi
KORTFATTAD MOTIVERING
Fiskeavtalet mellan Europeiska gemenskapen och São Tomé e Príncipe löpte ut den 31 maj 2010 efter att ha varit i kraft i tre år.
Avtalsvillkoren är följande:
Typ av utgifter
2011
2012
2013
TOTALT
Fångstmängd på 7 000 ton/år à 65 €/ton
455 000 €
455 000 €
455 000 €
1 365 000 €
Genomförande av den sektoriella fiskeripolitiken i São Tomé e Príncipe
227 500 €
227 500 €
227 500 €
682 500 €
Summa:
682 500 €
682 500 €
682 500 €
2 047 500 €
Administrativa utgifter
206 000 €
Totalt inklusive administrativa utgifter
682 500 €
682 500 €
682 500 €
2 253 500 €
Efter en gemensam utvärdering av beståndens tillstånd kan det på vissa villkor ges möjlighet att anpassa fiskekvoterna.
EU:s ekonomiska ersättning kommer att omfatta följande delar:
- Ett belopp på 455 000 EUR per år för rätten att fiska 7 000 ton per år (65 euro per ton).
- Ett belopp på 227 500 EUR per år för att stödja och genomföra den sektoriella fiskeripolitiken i São Tomé e Príncipe.
- En finansieringsram på 206 000 EUR för administrativa utgifter för perioden 2011–2013.
Det finns ingen övre gräns för vilka ytterligare mängder av tonfisk som får fångas av EU‑fartyg.
Varje överskjutande ton fångst kommer att kosta 65 EUR.
Om EU-fartygens fångster överskrider en mängd som motsvarar det dubbla totala årsbeloppet kommer betalningen för de fångster som överskrider detta gränsvärde att göras först året därpå.
São Tomé e Príncipe ligger på 101:a plats av 178 länder i Transparency Internationals korruptionsindex 2010.
Kommissionen måste se efter i vad mån pengarna har använts, och kommer att användas, för de ändamål som fastställts i överenskommelsen med São Tomé e Príncipe.
Budgetutskottet anser därför att följande punkter bör beaktas i samband med genomförandet av avtalet:
· Kommissionen ska varje år se efter om de medlemsstater vars fartyg bedriver fiske med stöd av protokollet till avtalet har efterlevt kraven på fångstrapportering.
Om så inte skett ska kommissionen avslå deras ansökningar om fisketillstånd för det kommande året.
· Kommissionen ska årligen rapportera till Europaparlamentet och rådet om resultaten av det fleråriga sektorsprogram som beskrivs i artikel 7 i protokollet samt om hur medlemsstaterna uppfyllt kraven på fångstrapportering.
· Kommissionen ska, innan protokollet löper ut eller förhandlingar om att eventuellt ersätta det inleds, förelägga Europaparlamentet och rådet en utvärdering i efterhand av protokollet, tillsammans med en kostnads-nyttoanalys.
Budgetutskottet uppmanar fiskeriutskottet att som ansvarigt utskott föreslå för parlamentet att det ger sitt godkännande till ingåendet av avtalet, och önskar att följande punkter beaktas på vederbörligt sätt av kommissionen och São Tomé e Príncipe vid genomförandet av avtalet:
a) Kommissionen ska varje år se efter om de medlemsstater vars fartyg bedriver fiske med stöd av protokollet till avtalet har efterlevt kraven på fångstrapportering.
Om så inte skett ska kommissionen avslå deras ansökningar om fisketillstånd för det kommande året.
b) Kommissionen ska årligen rapportera till Europaparlamentet och rådet om resultaten av det fleråriga sektorsprogram som beskrivs i artikel 7 i protokollet samt om hur medlemsstaterna uppfyllt kraven på fångstrapportering.
c) Kommissionen ska, innan protokollet löper ut eller förhandlingar om att eventuellt ersätta det inleds, förelägga Europaparlamentet och rådet en utvärdering i efterhand av protokollet, tillsammans med en kostnads-nyttoanalys.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
2.5.2011
Slutomröstning: resultat
+:
–:
0:
21
1
Slutomröstning: närvarande ledamöter
Slutomröstning: närvarande suppleanter
Jürgen Klute
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
24.5.2011
Slutomröstning: resultat
+:
–:
0:
17
1
1
Slutomröstning: närvarande ledamöter
Josefa Andrés Barea, Kriton Arsenis, Alain Cadec, Carmen Fraga Estévez, Pat the Cope Gallagher, Marek Józef Gróbarczyk, Iliana Malinova Iotova, Isabella Lövin, Guido Milana, Maria do Céu Patrão Neves, Crescenzio Rivellini, Ulrike Rodust, Struan Stevenson, Catherine Trautmann, Jarosław Leszek Wałęsa
Slutomröstning: närvarande suppleanter
Jean-Paul Besset, Izaskun Bilbao Barandica, Ole Christensen, Chris Davies
Slutomröstning: närvarande suppleanter (art.
187.2)
Pablo Arias Echeverría
A7-0255/2011
BETÄNKANDE
om en ny handelspolitik för Europa i samband med Europa 2020-strategin
(2010/2152(INI))
Utskottet för internationell handel
Föredragande:
Daniel Caspary
PE 460.634v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING..........................................................................................................................17
YTTRANDE från utskottet för utveckling ........................................................19
YTTRANDE från utskottet för industrifrågor, forskning och energi 24
YTTRANDE från utskottet för den inre marknaden och konsumentskydd 29
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................33
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om en ny handelspolitik för Europa i samband med Europa 2020-strategin
( 2010/2152(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av meddelandet från kommissionen till Europaparlamentet, rådet, Europeiska ekonomiska och sociala kommittén och Regionkommittén ”Handel, tillväxt och världspolitik, Handelspolitiken – en hörnsten i Europa 2020-strategin” ( KOM(2010)0612 ),
– med beaktande av kommissionens meddelande ”Europa 2020, En strategi för smart och hållbar tillväxt för alla” ( KOM(2010)2020 ),
– med beaktande av kommissionens meddelande ”Ett konkurrenskraftigt Europa i världen – Ett bidrag till EU:s tillväxt- och sysselsättningsstrategi” ( KOM(2006)0567 ),
– med beaktande av sin resolution av den 17 februari 2011 om Europa 2020
Antagna texter, P7_TA(2011)0068 . ,
– med beaktande av sin resolution av den 11 maj 2011 om läget i förhandlingarna om ett frihandelsavtal mellan EU och Indien
Antagna texter, P7_TA-PROV(2011)0224 . ,
– med beaktande av sin resolution av den 11 maj 2011 om handelsförbindelserna mellan EU och Japan
Antagna texter, P7_TA-PROV(2011)0225 . ,
– med beaktande av sin resolution av den 8 juni 2011 om handelsförbindelserna mellan EU och Kanada
Antagna texter, P7_TA-PROV(2011)0257 . ,
– med beaktande av sin resolution av den 6 april 2011 om den framtida EU-politiken för internationella investeringar
Antagna texter, P7_TA-PROV(2011)0141 . ,
– med beaktande av sin resolution av den 17 februari 2011 om frihandelsavtalet mellan EU och Sydkorea
Antagna texter, P7_TA-PROV(2011)0063 . ,
– med beaktande av meddelandet från kommissionen till rådet, Europaparlamentet och Europeiska ekonomiska och sociala kommittén ”Att bidra till en hållbar utveckling: rättvis handel och icke-statliga handelsrelaterade system för hållbar utveckling” av den 5 maj 2009 ( KOM(2009)0215 ),
– med beaktande av sin resolution av den 25 november 2010 om den internationella handelspolitiken inom ramen för de krav som klimatförändringarna medför
Antagna texter, P7_TA(2010)0445 . ,
– med beaktande av sin resolution av den 25 november 2010 om mänskliga rättigheter samt sociala normer och miljönormer i internationella handelsavtal
Antagna texter, P7_TA(2010)0434 . ,
– med beaktande av sin resolution av den 25 november 2010 om företagens sociala ansvar och miljöansvar vid internationella handelsavtal
Antagna texter, P7_T7(2010)0446. ,
– med beaktande av sin resolution av den 21 oktober 2010 om EU:s handelsförbindelser med Latinamerika
Antagna texter, P7_T7(2010)0387. ,
– med beaktande av sin resolution av den 21 september 2010 om handelsförbindelser och ekonomiska förbindelser med Turkiet
Antagna texter, P7_T7(2010)0324. ,
– med beaktande av sin resolution av den 16 juni 2010 om EU 2020
Antagna texter, P7_TA(2010)0223 . ,
– med beaktande av sin resolution av den 26 mars 2009 om ett frihandelsavtal mellan EU och Indien
EUT C 117 E, 6.5.2010, s.
166. ,
– med beaktande av sin resolution av den 5 februari 2009 om handel och ekonomiska förbindelser med Kina
EUT C 67 E, 18.3.2010, s.
132. ,
– med beaktande av sin resolution av den 5 februari 2009 om att förstärka de europeiska små och medelstora företagens roll i den internationella handeln
EUT C 67 E, 18.3.2010, s.
101. ,
– med beaktande av sin resolution av den 18 december 2008 om varumärkesförfalskningens inverkan på den internationella handeln
EUT C 45 E, 23.2.2010, s.
47. ,
– med beaktande av kommissionens meddelande av den 17 oktober 2008 ”De yttersta randområdena: en tillgång för Europa”,
– med beaktande av sin resolution av den 4 september 2008 om handel med tjänster
– med beaktande av sin resolution av den 20 maj 2008 om råvaruhandel
EUT C 279 E, 19.11.2009, s.
5. ,
– med beaktande av sin resolution av den 24 april 2008 om ”Mot en reformerad Världshandelsorganisation”
EUT C 259 E, 29.10.2009, s.
77. ,
– med beaktande av sin resolution av den 19 februari 2008 om EU:s strategi för att få till stånd marknadstillträde för europeiska företag
EUT C 184 E, 6.8.2009, s.
16. ,
– med beaktande av sin resolution av den 13 december 2007 om handel och ekonomiska förbindelser med Korea
EUT C 323 E, 18.12.2008, s.
520. ,
– med beaktande av sin resolution av den 22 maj 2007 om EU i världen – konkurrenskraftens externa aspekter
EUT C 102 E, 24.4.2008, s.
128. ,
– med beaktande av sin resolution av den 12 oktober 2006 om EU:s ekonomiska och kommersiella förbindelser med Mercosur i syfte att ingå ett interregionalt associeringsavtal
EUT C 308 E, 16.12.2006, s.
182. ,
– med beaktande av sin resolution av den 28 september 2006 om EU:s ekonomiska och kommersiella förbindelser med Indien
EUT C 306 E, 15.12.2006, s.
400. ,
– med beaktande av sin resolution av den 1 juni 2006 om transatlantiska förbindelser mellan EU och Förenta staterna
EUT C 298 E, 8.12.2006, s.
235. ,
– med beaktande av ordförandeskapets slutsatser från Europeiska rådets möte den 17-18 juni 2010,
– med beaktande av artikel 48 i arbetsordningen,
– med beaktande av betänkandet från utskottet för internationell handel och yttrandena från utskottet för utveckling, utskottet för industrifrågor, forskning och energi och utskottet för den inre marknaden och konsumentskydd ( A7‑0255/2011 ), och av följande skäl:
EU:s och USA:s andel av världens relativa BNP
”Convergence, Catch Up and Overtaking”, PwC, 2010. minskar samtidigt som tillväxtekonomierna är på snabb frammarsch
Denna relativa minskning av unionens BNP återspeglas i hur handeln har utvecklats
Uppgifter från Eurostat.
D. Unionen stod för 19 procent av världens varuexport 1999 och 17,1 procent av exporten 2009, vilket motsvarar en minskning med 10 procent i relativ export.
E. Unionen stod för 19,5 procent av världens varuimport 1999 och 17,6 procent av importen 2009, vilket motsvarar en minskning med 10 procent i relativ import.
F. Exporten av tjänster ökade från 26,7 procent till 30,2 procent av unionens totala export mellan 1999 och 2009
Eurostat, FN:s databas UN Servicetrade. .
G. 50 länder (30 om EU räknas som en enhet) står för 80 procent av världens handel.
Demografiska förändringar
Europeiska kommissionen, 2009 års åldranderapport; Eurostat/Unece arbetsgrupp 2010. påverkar även den ekonomiska utvecklingen
Unionens ekonomi beror till stor del på deltagandet i den externa tillväxten
I. Målen om tillväxt, välstånd, arbetstillfällen och bevarande av den europeiska sociala modellen är alla sammanlänkade och stöder varandra.
J. Kommissionen beräknar att 90 procent av världens tillväxt år 2015 kommer att skapas utanför unionen.
K. Öppnare marknader leder till högre produktivitet, bidrar till ökad extern konkurrenskraft och skulle omedelbart kunna bidra till över 1,5 procent av den direkta ekonomiska tillväxten och innebära stora fördelar för konsumenterna.
M. Med tanke på unionens demografiska framtidsutsikter och deras negativa effekter för tillväxtpotentialen är det av största vikt att utnyttja tillväxtpotentialen i ökad produktivitet och utrikeshandel.
En framtida europeisk handelspolitisk strategi bör beakta de särdrag som kännetecknar EU:s företag och regioner samt beroendet av extern tillväxt
N. Kommissionen föreslår i sitt meddelande ”Handel, tillväxt och världspolitik” konkreta kortsiktiga åtgärder, men tar inte upp unionens framtida roll i en förändrad värld.
O. Kommissionen har lagt fram ett förslag till Europaparlamentets och rådets förordning om införande av övergångsordningar för bilaterala investeringsavtal mellan medlemsstater och tredjeländer som en del av EU:s investeringspolitik.
Europaparlamentet uppmanar kommissionen att utarbeta en sådan prognos som utgångspunkt och lägga fram en reviderad strategi på medellång och lång sikt före sommaren 2012, eftersom meddelandet om handel, tillväxt och världspolitik inte gör detta.
Europaparlamentet är medvetet om att handelspolitiken inte är ett självändamål
a) mänskliga rättigheter,
b) jobbgarantier och jobbskapande,
c) arbetstagares rättigheter och ILO:s grundläggande arbetsrättsliga normer,
d) företagens sociala ansvar,
e) jordbrukspolitiken,
f) miljöpolitiken,
g) klimatförändringar,
h) kampen mot fattigdom inom och utanför EU,
i) utvecklingspolitiken,
j) skyddet av konsumenternas intressen och rättigheter,
k) tryggad råvaru- och energiförsörjning,
l) utrikespolitiken,
m) grannskapspolitiken,
n) industripolitiken,
o) skyddet av äganderätten, däribland immateriella rättigheter,
p) främjandet av de rättsstatliga principerna.
Antagna texter P7_TA (2010)0434. , om företagens sociala ansvar och miljöansvar vid internationella handelsavtal
Antagna texter P7_TA (2010)0446. och om den internationella handelspolitiken inom ramen för de krav som klimatförändringarna medför
Europaparlamentet framhåller att handelspolitiken är ett viktigt inslag i unionens nya industripolitik och att handeln bör bygga på rättvis global konkurrens och fullständig ömsesidighet för att upprätthålla en sund tillverkningsbas i Europa.
Parlamentet föredrar starkt en multilateral strategi inom WTO
Parlamentet betraktar frihandelsavtal som viktiga instrument för marknadstillträde
Parlamentet efterlyser fler och bättre resultat från dialoger på hög nivå med viktiga handelspartner som Förenta staterna, Kina, Japan och Ryssland.
Huvudprioriteringen är fortfarande öppna marknader och marknadstillträde
Europaparlamentet betonar att det främsta bidraget till EU:s ekonomiska framgång är de olika ekonomiska aktörernas verksamhet, däribland små och medelstora företag och multinationella företag, och uppmanar därför kommissionen att ta hänsyn till de olika ekonomiska aktörernas behov och intressen i samband med alla handelsförhandlingar och nya interna bestämmelser.
EU:s konkurrenskraft och ekonomiska framgång kan inte säkras utan tjänster och väl skyddade utländska direktinvesteringar
Antagna texter, P7_TA(2011)0141 . .
Europaparlamentet efterlyser positiv ömsesidighet på internationella marknader för offentlig upphandling
Europaparlamentet uppmanar kommissionen att arbeta för ett positivt ömsesidigt tillträde inom denna viktiga ekonomiska sektor, och påminner om att man när det gäller ömsesidigt tillträde inte bör sträva efter att stänga våra marknader utan att i stället öppna de utländska marknaderna för offentlig upphandling.
Europaparlamentet efterlyser en ambitiös insats för att begränsa regleringsmässiga hinder i och utanför Europa
Europaparlamentet uppmanar kommissionen att systematiskt utvärdera hur EU:s interna politik och bestämmelser påverkar den globala konkurrensförmågan och att i sina förslag ge företräde åt de alternativ som minst sannolikt kommer att påverka EU-företagens konkurrenskraft negativt i och utanför Europa.
Parlamentet deltar i kampen mot fattigdom i och utanför EU
Europaparlamentet uppmanar kommissionen att i samband med avtal om ekonomiskt partnerskap beakta parlamentets tidigare resolutioner om behovet av att visa flexibilitet i förhandlingarna med våra partner och fullgöra åtagandena om särskild och differentierad behandling för utvecklingsländerna.
Europaparlamentet betonar att utrikeshandelspolitiken ska skydda EU:s förmåga att bevara en stark jordbrukssektor som kan garantera livsmedelstryggheten och livsmedelssuveräniteten för 500 miljoner konsumenter i EU.
Europaparlamentet kräver en hållbar och icke snedvriden råvaruförsörjning
Det krävs ett bättre tullsamarbete i och utanför EU
Europaparlamentet uppmanar kommissionen och medlemsstaterna att allvarligt överväga förslaget att inrätta en gemensam europeisk tullmyndighet som ska säkra en mer effektiv tillämpning av tullbestämmelser och tullförfaranden inom EU:s tullområde.
Europaparlamentet efterlyser ett korrekt skydd av immateriella rättigheter som även tar hänsyn till de fattigaste människornas intressen
o
o o
MOTIVERING
Kommissionens dokument innehåller goda idéer för de kommande månaderna, men ingen riktig framtidsstrategi läggs fram.
Den 9 november 2010 lade Europeiska kommissionen fram sitt meddelande ”Handel, tillväxt och världspolitik” om den framtida handelspolitiken för EU.
Detta meddelande, som ska lägga fram de externa aspekterna av Europa 2020-strategin, är i första hand en fortsättning på strategin Europa i världen från 2006.
I ett betänkande som utarbetades av samma föredragande tog Europaparlamentet 2007 ställning till strategin Europa i världen och välkomnade detta initiativ.
Kommissionen och parlamentet inledde under 2010 en utvärdering av denna strategi.
Av denna utvärdering framgår tydligt att många av de angivna målen för Europa i världen ännu inte har uppnåtts.
Föredraganden uppmanar därför kommissionen, medlemsstaterna och alla deltagare att undersöka varför många mål ännu inte har kunnat uppnås och att dra lämpliga slutsatser av detta.
De flesta av de mål som formulerades då ska fortfarande genomföras, enligt kommissionens senaste dokument.
Argumenten för de åtgärder som angavs i det tidigare kommissionsdokumentet, som finns förklarade i motiveringen till betänkandet ”EU i världen – konkurrenskraftens externa aspekter” (2006/2292), gäller även i dag och upprepas därför inte här.
När det gäller innehållet hänvisar föredraganden till motiveringen i sitt betänkande från 2006 om konkurrenskraftens utrikespolitiska aspekter
Föredraganden välkomnar kommissionens meddelande ”Handel, tillväxt och världspolitik” – vid en tidpunkt då EU genom Lissabonfördragets ikraftträdande även har fått nya befogenheter, t.ex. när det gäller investeringspolitiken.
I samband med detta välkomnas särskilt att kommissionen erkänner att vårt välstånd och vår tillväxt beror på ett fungerande internationellt handelssystem.
Ändå kritiserar föredraganden att meddelandet, som visserligen tar upp många relevanta frågor, underlåter att presentera en framtidsinriktad handels- och investeringsstrategi.
Meddelandet ”Handel, tillväxt och världspolitik” handlar enligt föredraganden snarare om riktlinjer för politiken under de kommande månaderna än om en omfattande handelsstrategi för EU, som står inför utmaningarna från en global ekonomi i snabb förändring och en kraftig förskjutning av den ekonomiska jämvikten.
Världen har förändrats dramatiskt under de senaste åren ...
Världshandeln har tack vare WTO och många multilaterala och bilaterala initiativ fått ett enormt uppsving.
Vid genomförandet av Lissabonstrategin år 2000 hade EU fortfarande 25 procent av det globala mervärdet, men år 2020 räknar man med en andel på 18 procent.
Däremot hade världens två mest folkrika länder, Kina och Indien, under år 2000 endast 10 procent av världshandeln, en andel som år 2020 enligt olika källor kommer att ha ökat till 25 procent.
Bara denna förändring visar att en sådan förändring också måste påverka EU:s politik.
Sedan 1990-talet har allt fler tillväxtekonomier och utvecklingsländer i allt större utsträckning integrerats i världshandeln och utvecklats till en bärande motor i världsekonomin.
Detta visade sig särskilt under krisåren 2008 och 2009, då framför allt tillväxtekonomierna hade en stabiliserande effekt på den globala ekonomin.
EU:s och USA:s exportandel i förhållande till den totala globala exporten låg under 2009 på knappt 29 procent, jämfört med knappt 37 procent 1999.
BRIK-länderna (Brasilien, Ryssland, Indien och Kina) däremot gick från en andel på 9,3 procent av den globala exporten till en andel på 20,4 procent år 2009, med en tendens till ytterligare ökningar.
Många tillväxtekonomier uppvisar handelsöverskott, exporterna och ekonomin ökar kraftigt och skuldsättningen minskar.
Det är framför allt syd-syd-handeln som ökar kraftigt, och beroendet av efterfrågan i industriländerna har sjunkit avsevärt.
EU måste dessutom tänka på att befolkningstillväxten inom EU minskar kraftigt, medan invånarantalet i utvecklingsländerna däremot ökar blixtsnabbt.
Detta kommer att påverka ländernas ekonomiska situation.
Med tanke på att 18 procent respektive 36 miljoner arbetsplatser inom EU redan i dag är beroende av utrikeshandeln och att 90 procent av den globala ekonomiska tillväxten år 2015 troligen kommer att genereras utanför EU, är det särskilt viktigt att utarbeta och genomföra en långsiktig strategi för utrikeshandel, som tar hänsyn till den föränderliga rollen för EU inom den globala ekonomin.
... och därför bör kommissionen snabbt lägga fram en långsiktig strategi för utrikeshandeln
Mot bakgrund av denna utveckling uppmanar föredraganden kommissionen att utarbeta en analys och långtidsplanering som tar hänsyn till de aktuella förutsättningarna för den globala ekonomin och den aktuella situationen för EU samt den sannolika framtida utvecklingen.
YTTRANDE från utskottet för utveckling
till utskottet för internationell handel
över en ny handelspolitik för Europa i samband med Europa 2020-strategin
( 2010/2152(INI) )
Föredragande: Birgit Schnieber-Jastram
FÖRSLAG
Utskottet för utveckling uppmanar utskottet för internationell handel att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet understryker därför att det är extremt viktigt att utforma en handelspolitik som bidrar till att uppfylla millennieutvecklingsmål 8 (utveckla ett globalt partnerskap för utveckling), samtidigt som skillnaderna mellan medelinkomstländer, låginkomstländer och bräckliga stater beaktas.
Europaparlamentet påminner om att EU, för att främja en ekonomisk tillväxt som kommer alla till del och som gynnar de fattiga, inom ramen för sin handelspolitik måste sträva efter att inom två år slutföra Doharundan på ett sätt som främjar utveckling och ytterligare stödja handeln och den regionala integrationen mellan de sydliga länderna.
Europaparlamentet påminner om att Aid for Trade-strategin syftar till att hjälpa utvecklingsländer att förhandla, genomföra och dra fördel av handelsavtal, att utöka sin handel och att påskynda utrotandet av fattigdomen.
Europaparlamentet uppmanar EU att avstå från att utöva onödiga påtryckningar på utvecklingsländerna för att kunna sluta investeringsavtal som begränsar deras möjlighet att införa bestämmelser till förmån för sociala utvecklingsmål.
Europaparlamentet uppmanar EU att respektera den överenskommelse som nåddes under det svenska ordförandeskapet om att lägga fram en konkret plan för genomförandet av FN:s ram för att ”skydda, respektera och åtgärda”.
Punkt 18 i resolutionen om rättvis handel och utveckling ( 2005/2245(INI) ).
A6-0207/2006 .
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
3.3.2011
Slutomröstning: resultat
+:
–:
0:
19
Slutomröstning: närvarande ledamöter
Thijs Berman, Ricardo Cortés Lastra, Nirj Deva, Leonidas Donskis, Charles Goerens, András Gyürk, Eva Joly, Franziska Keller, Gay Mitchell, Norbert Neuser, Birgit Schnieber-Jastram, Michèle Striffler, Alf Svensson, Eleni Theocharous, Iva Zanicchi, Gabriele Zimmer
Slutomröstning: närvarande suppleanter
Fiona Hall, Cristian Dan Preda
Slutomröstning: närvarande suppleanter (art.
187.2)
Jolanta Emilia Hibner
YTTRANDE från utskottet för industrifrågor, forskning och energi
till utskottet för internationell handel
över en ny handelspolitik för Europa inom ramen för Europa 2020-strategin
( 2010/2152(INI) )
Föredragande: Andrzej Grzyb
FÖRSLAG
Utskottet för industrifrågor, forskning och energi uppmanar utskottet för internationell handel att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
– ta hänsyn till alla aspekter när det gäller konkurrenskraften hos den europeiska industrin, små och medelstora företag, jordbrukssektorn och livsmedelsindustrin, med tanke på det växande handelsunderskottet när det gäller jordbruksprodukter och den höga standard som måste hållas av EU-industrin,
– främja sådant samarbete med utvecklingsländer som är fördelaktigt för båda parter,
– försöka bekämpa tredjeländers handelssnedvridande åtgärder, t.ex. exportavgifter och orättvist offentligt stöd till inhemsk produktion.
Parlamentet efterlyser en starkare koppling mellan regelverken för den externa marknaden och den inre marknaden för att minska onödiga kostnader för företag och undanröja regleringshinder, och snabba på innovation och tillgång till handel.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
12.4.2011
Slutomröstning: resultat
+:
–:
0:
44
2
1
Slutomröstning: närvarande ledamöter
Slutomröstning: närvarande suppleanter
Antonio Cancian, António Fernando Correia De Campos, Francesco De Angelis, Ilda Figueiredo, Matthias Groote, Andrzej Grzyb, Satu Hassi, Yannick Jadot, Silvana Koch-Mehrin, Bernd Lange, Werner Langen, Mario Pirillo, Algirdas Saudargas, Catherine Trautmann
till utskottet för internationell handel
över en ny handelspolitik för Europa i samband med Europa 2020-strategin
( 2010/2152(INI) )
Föredragande:
Malcolm Harbour
FÖRSLAG
Utskottet för den inre marknaden och konsumentskydd uppmanar utskottet för internationell handel att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet framhåller åter att det mellan Europeiska unionen och dess handelsparter behövs balanserade handelsavtal, som ingås i en anda av ömsesidighet och som är till nytta för båda parter.
Europaparlamentet anser att EU samtidigt bör överväga att delta i en dialog för att uppmuntra dessa länder att förstärka sina regionala handelsförbindelser med upprättande av en gemensam tullunion som slutmål.
Europaparlamentet anser med tanke på den åldrande befolkningen att den äldre arbetskraften är en värdefull tillgång till handeln, och att hinder bör avskaffas för att uppmuntra och stimulera de äldre att fortsätta arbeta.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att ta vederbörlig hänsyn till betydelsen av innovation för en stark och hållbar tillväxt genom att se till att innovationerna får ordentlig finansiering, nämligen genom inrättande av EU‑projektobligationer och lagstiftning som tillåter riskkapitalfonder att investera fritt i hela EU.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
13.4.2011
Slutomröstning: resultat
+:
–:
0:
33
3
Slutomröstning: närvarande ledamöter
Pablo Arias Echeverría, Adam Bielan, Lara Comi, Anna Maria Corazza Bildt, António Fernando Correia De Campos, Jürgen Creutzmann, Christian Engström, Evelyne Gebhardt, Louis Grech, Małgorzata Handzlik, Iliana Ivanova, Philippe Juvin, Sandra Kalniete, Eija-Riitta Korhola, Edvard Kožušník, Kurt Lechner, Toine Manders, Mitro Repo, Robert Rochefort, Zuzana Roithová, Heide Rühle, Matteo Salvini, Christel Schaldemose, Andreas Schwab, Eva-Britt Svensson, Róża Gräfin von Thun und Hohenstein, Kyriacos Triantaphyllides, Emilie Turunen, Bernadette Vergnaud, Barbara Weiler
Slutomröstning: närvarande suppleanter
Ashley Fox, María Irigoyen Pérez, Constance Le Grip, Konstantinos Poupakis, Olle Schmidt, Marc Tarabella
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
21.6.2011
Slutomröstning: resultat
+:
–:
0:
23
4
1
Slutomröstning: närvarande ledamöter
William (The Earl of) Dartmouth, Laima Liucija Andrikienė, Kader Arif, David Campbell Bannerman, Daniel Caspary, Marielle De Sarnez, Christofer Fjellner, Yannick Jadot, Metin Kazak, Bernd Lange, David Martin, Emilio Menéndez del Valle, Vital Moreira, Paul Murphy, Cristiana Muscardini, Godelieve Quisthoudt-Rowohl, Niccolò Rinaldi, Tokia Saïfi, Helmut Scholz, Peter Šťastný, Robert Sturdy, Keith Taylor, Iuliu Winkler, Pablo Zalba Bidegain, Paweł Zalewski
Slutomröstning: närvarande suppleanter
Catherine Bearder, George Sabin Cutaş, Mário David, Syed Kamall, Maria Eleni Koppa, Elisabeth Köstinger, Jörg Leichtfried, Inese Vaidere, Jarosław Leszek Wałęsa
A7-0276/2011
***
REKOMMENDATION
om förslaget till rådets beslut om ingående av avtalet genom skriftväxling mellan Europeiska unionen och Konungariket Norge om ytterligare handelsförmåner för jordbruksprodukter, uppnådda på grundval av artikel 19 i avtalet om Europeiska ekonomiska samarbetsområdet
(14206/2010 – C7‑0101/2011 – 2010/0243(NLE))
Utskottet för internationell handel
Föredragande: Helmut Scholz
PE 456.787v02-00
Teckenförklaring
* Samrådsförfarande
*** Godkännandeförfarande
***I Ordinarie lagstiftningsförfarande (första behandlingen)
***II Ordinarie lagstiftningsförfarande (andra behandlingen)
***III Ordinarie lagstiftningsförfarande (tredje behandlingen)
(Det angivna förfarandet baseras på den rättsliga grund som angetts i förslaget till akt.)
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION...................5
MOTIVERING............................................................................................................................6
YTTRANDE från utskottet för jordbruk och landsbygdens utveckling 8
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................11
FÖRSLAG TILL EUROPAPARLAMENTETS LAGSTIFTNINGSRESOLUTION
om förslaget till rådets beslut om ingående av avtalet genom skriftväxling mellan Europeiska unionen och Konungariket Norge om ytterligare handelsförmåner för jordbruksprodukter, uppnådda på grundval av artikel 19 i avtalet om Europeiska ekonomiska samarbetsområdet
(14206/2010 – C7‑0101/2011 – 2010/0243(NLE) )
(Godkännande)
Europaparlamentet utfärdar denna resolution
– med beaktande av förslaget till rådets beslut (14206/2010),
– med beaktande av avtalet genom skriftväxling mellan Europeiska unionen och Konungariket Norge om ytterligare handelsförmåner för jordbruksprodukter, uppnådda på grundval av artikel 19 i avtalet om Europeiska ekonomiska samarbetsområdet (14372/2010),
– med beaktande av begäran om godkännande som rådet har lagt fram i enlighet med artiklarna 207.4 första stycket och 218.6 andra stycket led a i fördraget om Europeiska unionens funktionssätt ( C7‑0101/2011 ),
1.
Europaparlamentet godkänner att avtalet ingås.
2.
MOTIVERING
Som medlem av Europeiska ekonomiska samarbetsområdet (EES) drar Norge nytta av den inre marknadens fördelar, men jordbruk och fiske är undantagna från fri omsättning i EES‑avtalet från 1992.
Det senaste avtalet mellan Konungariket Norge och Europeiska gemenskapen på grundval av artikel 19 i EES-avtalet trädde i kraft i juli 2003.
Det innehöll en ordning för handel med ost mellan parterna och ömsesidiga medgivanden för ett antal olika jordbruksprodukter inklusive tullkvoter.
Från mars 2008 till januari 2010 hölls nya förhandlingar som resulterade i det föreliggande förslaget till avtal som innehåller följande bestämmelser.
Medgivanden som Norge beviljat EU:
Ytterligare full liberalisering av grovt räknat cirka 20 procent av EU:s export till Norge, eller 250 miljoner euro.
Sammanlagt kommer cirka 60 procent (räknat i värdet av handeln) av jordbrukshandeln mellan Konungariket Norge och Europeiska unionen att vara helt fri.
För mer känsliga produkter som kött, mjölkprodukter, frukt, grönsaker och prydnadsväxter kommer Norge att bevilja följande tullkvoter och nedsatta tullavgifter:
· Nya tullkvoter, i köttsektorn (600 ton för fläskkött, 800 ton för fjäderfäkött och 900 ton för nötkött) på villkor att dessa kvantiteter omvandlas till MGN-kvoter inom ramen för WTO när ett framtida WTO-avtal ska genomföras.
Medgivanden som EU beviljat Norge:
Fullständig liberalisering för produkter där Norge erbjuder fullständig liberalisering , och tilläggskvoter för ost (3 200 ton), färska hallon (400 ton), potatischips (200 ton) o ch foder till sällskapsdjur (13 000 ton).
Norge har en positiv handelsbalans gentemot EU totalt sett , men när det gäller handeln på jordbruksområdet har EU en positiv balans gentemot Norge.
EU:s export av jordbruksprodukter fördubblades mellan 2000 och 2007 till 1,6 miljarder euro.
YTTRANDE från utskottet för jordbruk och landsbygdens utveckling
till utskottet för internationell handel
över utkastet till rådets beslut om ingående av avtalet genom skriftväxling mellan Europeiska unionen och Konungariket Norge om ytterligare handelsförmåner för jordbruksprodukter, uppnådda på grundval av artikel 19 i avtalet om Europeiska ekonomiska samarbetsområdet
(14206/2010 – C7‑0101/2011 – 2010/0243(NLE) )
Föredragande:
Richard Ashworth
KORTFATTAD MOTIVERING
Det senaste avtalet genom skriftväxling mellan Europeiska unionen (då Europeiska gemenskapen) och Konungariket Norge på grundval av artikel 19 i EES-avtalet trädde i kraft i juli 2003.
Det innehöll en ordning för handel med ost mellan parterna och ömsesidiga medgivanden för ett antal olika jordbruksprodukter inklusive tullkvoter.
I artikel 19 i avtalet om Europeiska ekonomiska samarbetsområdet (EES) föreskrivs en successiv liberalisering av handeln med jordbruksprodukter mellan de avtalsslutande parterna.
För det ändamålet bör parterna vartannat år se över handelsvillkoren för jordbruksprodukter och inom ramen för avtalet, på basis av förmånsbehandling, bilateralt eller multilateralt och till ömsesidig nytta, fatta beslut om ytterligare minskningar av varje slag av handelshinder inom jordbrukssektorn.
Detta förslag, i vilket föreskrivs ytterligare liberalisering av handeln med jordbruksprodukter, är resultatet av de bilaterala förhandlingar om handel med jordbruksprodukter som ägde rum mellan mars 2008 och januari 2010.
De nya förmånerna kommer att bestå av ytterligare fullständig liberalisering för vissa känsliga produkter och därmed kommer cirka 60 procent av handeln med jordbruksprodukter mellan Konungariket Norge och Europeiska unionen att vara helt fri.
För mer känsliga produkter som kött, mjölkprodukter, frukt, grönsaker och prydnadsväxter har man enats om tullkvoter eller nedsatta tullar.
Särskilda bestämmelser har fastställts för förvaltningen av tullkvoterna för ost.
Budgetkonsekvenser: Förlusten av tullintäkter uppskattas till cirka 4,96 miljoner euro (netto efter avdrag för uppbördskostnader).
På grundval av ovannämnda synpunkter anser utskottet för jordbruk och landsbygdens utveckling att ifrågavarande avtal, som ska ingås på basis av det föreslagna rådsbeslutet, är i linje med ansträngningarna att uppnå en successiv liberalisering av handeln med jordbruksprodukter mellan Europeiska unionen och Konungariket Norge.
Utskottet anser vidare att man i avtalet på vederbörligt sätt har beaktat ovannämnda känsliga produkter och föreskrivit lämpliga lösningar i fråga om tullkvoter eller nedsatta tullar.
******
Utskottet för jordbruk och landsbygdens utveckling uppmanar utskottet för internationell handel att som ansvarigt utskott föreslå att parlamentet ger sitt godkännande.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
24.5.2011
Slutomröstning: resultat
+:
–:
0:
35
1
2
Slutomröstning: närvarande ledamöter
John Stuart Agnew, Richard Ashworth, Liam Aylward, José Bové, Luis Manuel Capoulas Santos, Vasilica Viorica Dăncilă, Michel Dantin, Paolo De Castro, Albert Deß, Herbert Dorfmann, Hynek Fajmon, Lorenzo Fontana, Béla Glattfelder, Martin Häusling, Esther Herranz García, Peter Jahr, Elisabeth Jeggle, Jarosław Kalinowski, Elisabeth Köstinger, Agnès Le Brun, George Lyon, Mairead McGuinness, Krisztina Morvai, Mariya Nedelcheva, James Nicholson, Rareş-Lucian Niculescu, Wojciech Michał Olejniczak, Georgios Papastamkos, Marit Paulsen, Britta Reimers, Alfreds Rubiks, Giancarlo Scottà, Czesław Adam Siekierski, Sergio Paolo Francesco Silvestris, Csaba Sándor Tabajdi, Marc Tarabella
Slutomröstning: närvarande suppleanter
Luís Paulo Alves, Salvatore Caronna, Esther de Lange
Slutomröstning: närvarande suppleanter (art.
187.2)
Pablo Zalba Bidegain
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
13.7.2011
Slutomröstning: resultat
+:
–:
0:
24
1
1
Slutomröstning: närvarande ledamöter
William (The Earl of) Dartmouth, Laima Liucija Andrikienė, Kader Arif, David Campbell Bannerman, Daniel Caspary, Marielle De Sarnez, Christofer Fjellner, Metin Kazak, David Martin, Vital Moreira, Paul Murphy, Cristiana Muscardini, Franck Proust, Godelieve Quisthoudt-Rowohl, Niccolò Rinaldi, Helmut Scholz, Peter Šťastný, Keith Taylor, Paweł Zalewski
Slutomröstning: närvarande suppleanter
Josefa Andrés Barea, George Sabin Cutaş, Norbert Glante, Syed Kamall, Elisabeth Köstinger
Slutomröstning: närvarande suppleanter (art.
187.2)
Rosa Estaràs Ferragut, Vicky Ford
A7-0304/2011
BETÄNKANDE
om förslaget till Europaparlamentets och rådets beslut om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning (ansökan EGF/2010/027 NL/Noord-Brabant huvudgrupp 18 från Nederländerna)
(KOM(2011)0386 – C7‑0173/2011 – 2011/2137(BUD))
Budgetutskottet
Föredragande: Barbara Matera
PE 469.713v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
BILAGA: EUROPAPARLAMENTETS OCH RÅDETS BESLUT..............................................6
MOTIVERING............................................................................................................................8
BILAGA: SKRIVELSE FRÅN UTSKOTTET FÖR SYSSELSÄTTNING OCH SOCIALA FRÅGOR 12
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om förslaget till Europaparlamentets och rådets beslut om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning (ansökan EGF/2010/027 NL/Noord-Brabant huvudgrupp 18 från Nederländerna)
( KOM(2011)0386 – C7‑0173/2011 – 2011/2137(BUD) )
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2011)0386 – C7‑0173/2011 ),
– med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
EUT C 139, 14.6.2006, s.
1. , särskilt punkt 28,
EUT L 406, 30.12.2006, s.
1. ,
– med beaktande av trepartsförfarandet i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006,
– med beaktande av skrivelsen från utskottet för sysselsättning och social frågor,
– med beaktande av betänkandet från budgetutskottet ( A7‑0304/2011 ), och av följande skäl:
A. Europeiska fonden för justering för globaliseringseffekter (nedan kallad ”fonden”) inrättades för att ge kompletterande stöd till arbetstagare som blivit arbetslösa till följd av de genomgripande strukturförändringar som skett inom världshandeln på grund av globaliseringen och för att underlätta deras återinträde på arbetsmarknaden.
B. Tillämpningsområdet för fonden har utvidgats, och från och med den 1 maj 2009 är det möjligt att söka stöd för åtgärder som riktas till arbetstagare som har blivit uppsagda som en direkt följd av den globala finansiella och ekonomiska krisen.
C. Unionens ekonomiska stöd till arbetstagare som har blivit uppsagda bör vara dynamiskt och ges så snabbt och effektivt som möjligt, i enlighet med Europaparlamentets, rådets och kommissionens gemensamma uttalande, som antogs vid förlikningsmötet den 17 juli 2008, och med vederbörlig hänsyn till bestämmelserna i det interinstitutionella avtalet av den 17 maj 2006 när det gäller antagandet av beslut om utnyttjande av fonden.
E. Ansökan uppfyller kriterierna för berättigande till stöd enligt förordningen om Europeiska fonden för justering för globaliseringseffekter.
BILAGA: EUROPAPARLAMENTETS OCH RÅDETS BESLUT
om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning (ansökan EGF/2010/027 NL/Noord-Brabant huvudgrupp 18 från Nederländerna)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA BESLUT
med beaktande av fördraget om Europeiska unionens funktionssätt,
med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
EUT C 139, 14.6.2006, s.
1. , särskilt punkt 28,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1927/2006 av den 20 december 2006 om upprättande av Europeiska fonden för justering för globaliseringseffekter
EUT L 406, 30.12.2006, s.
1. , särskilt artikel 12.3,
EUT C […], […], s. […]. , och
av följande skäl:
(2) Tillämpningsområdet för fonden har utvidgats, och från och med den 1 maj 2009 är det möjligt att söka stöd för åtgärder som riktas till arbetstagare som har blivit uppsagda som en direkt följd av den globala finansiella och ekonomiska krisen.
(3) Det interinstitutionella avtalet av den 17 maj 2006 gör det möjligt att använda medel från fonden upp till ett belopp på högst 500 miljoner euro per år.
Ansökan uppfyller villkoren för fastställande av det ekonomiska stödet enligt artikel 10 i förordning (EG) nr 1927/2006.
Kommissionen föreslår därför att ett belopp på 667 823 euro ska anslås.
(5) Fonden bör därför utnyttjas för att bevilja det ekonomiska stöd som Nederländerna ansökt om.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Europeiska fonden för justering för globaliseringseffekter ska belastas med 667 823 euro i åtagande- och betalningsbemyndiganden ur Europeiska unionens allmänna budget för 2011.
Artikel 2
Detta beslut ska offentliggöras i Europeiska unionens officiella tidning .
Utfärdat i [Bryssel/Strasbourg] den
På Europaparlamentets vägnar På rådets vägnar
Ordförande Ordförande
MOTIVERING
Europeiska fonden för justering för globaliseringseffekter inrättades för att ge kompletterande stöd till arbetstagare som blivit arbetslösa till följd av genomgripande strukturförändringar i världshandelsmönstret.
Enligt bestämmelserna i punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 om budgetdisciplin och sund ekonomisk förvaltning
EUT C 139, 14.6.2006, s.
1. och artikel 12 i förordning (EG) nr 1927/2006
EUT L 406, 30.12.2006, s.
1. får det årliga belopp som avdelas för fonden inte överstiga 500 miljoner euro som tas från eventuella marginaler under det samlade utgiftstaket för det föregående året och/eller från annullerade åtagandebemyndiganden under de två senaste åren, med undantag för sådana som ingår under rubrik 1b.
Anslagen förs in i budgeten i form av en avsättning så snart kommissionen har funnit tillräckliga marginaler och/eller frigjort åtaganden.
För att kunna ta fonden i anspråk ska kommissionen, efter en positiv prövning av ansökan, lägga fram ett förslag till budgetmyndigheten om utnyttjande av fonden tillsammans med en begäran om överföring.
Parallellt med detta kan ett trepartsmöte ordnas för att komma överens om användning av fonden och vilka belopp som behövs.
Trepartsmötet kan vara i förenklad form.
II.
Lägesrapport: kommissionens förslag
Den 28 juni 2011 antog kommissionen ett nytt förslag till beslut om utnyttjande av Europeiska fonden för globaliseringseffekter till förmån för Nederländerna för att stödja återintegrering på arbetsmarknaden av arbetstagare som har blivit uppsagda som en följd av den globala finansiella och ekonomiska krisen.
Detta är den nionde ansökan som ska behandlas inom ramen för budgeten för 2011 och avser utnyttjande av ett totalbelopp på 667 823 euro från fonden till förmån för Nederländerna.
Denna ansökan, ärende EGF/2010/027 NL/ Noord-Brabant huvudgrupp 18 från Nederländerna, lämnades in till kommissionen den 20 december 2010 och kompletterades med ytterligare uppgifter fram till den 7 mars 2011.
Ett av kriterierna för kommissionens bedömning var utvärderingen av kopplingen mellan uppsägningarna och stora strukturella förändringar i världshandelsmönstren eller finanskrisen, vilket i just detta fall hör samman med det globala efterfrågetappet för den grafiska branschen, som 2009 var - 8,6 procent för Nederländerna.
Dessutom minskade övriga branschers beställningar på tryckt reklammaterial kraftigt, på grund av budgetnedskärningar inom tryckeri- och förlagsverksamhet.
När det gäller att belägga antalet uppsägningar uppfyller fallet Noord-Brabant helt och hållet villkoren i artikel 2 c i förordning (EG) nr 1927/2006, där det anges att på mindre arbetsmarknader eller vid särskilda omständigheter kan en ansökan om bidrag från EGF godtas även om de interventionskriterier som fastställts i artikel 2 a eller 2 b inte till fullo uppfylls, om uppsägningarna har allvarliga följder för sysselsättningen och den lokala ekonomin.
Nederländerna begär i denna ansökan undantag från artikel 2 b, enligt vilken minst 500 arbetstagare ska ha sagts upp under en referensperiod på nio månader vid företag som är verksamma inom en huvudgrupp enligt Nace rev.
2 i en region eller två regioner som gränsar till varandra på Nuts II-nivå i en medlemsstat.
Ansökan avser 199 uppsägningar i 14 företag i sektorn Nace rev.
2 huvudgrupp 18 (Grafisk produktion och reproduktion av inspelningar) inom Nuts II-regionen Noord-Brabant (NL41), under referensperioden på nio månader från den 16 januari till den 16 oktober 2010.
De nederländska myndigheterna anser att ansökan uppfyller kraven i artikel 2 c i förordning (EG) nr 1927/2006 på grund av de särskilda omständigheter som råder.
De uppsägningar som ansökan gäller har skett i samma huvudgrupp enligt Nace rev.
Noord-Brabant gränsar dessutom till Zuid‑Holland på Nuts II-nivån.
Det exceptionella är kombinationen av dessa faktorer vilka sammantaget försätter arbetstagarna och den berörda regionen i en ovanlig och svår situation.
Enligt Nederländerna är situationen i Noord-Brabant mycket ansträngd.
I denna provins ökade arbetslösheten från 3,1 procent det tredje kvartalet 2008 till 5 procent det tredje kvartalet 2010.
I Veghel och Uden, det nästa största centret för den grafiska sektorn i Noordosst-Brabant var arbetslösheten inom den grafiska branschen 88 procent högre i oktober 2010 än i oktober 2008.
Enligt prognosen kommer arbetsmarknaden i Noord-Brabant dessutom att försämras ytterligare på grund av krisen inom teknisk industri och bygg- och anläggningssektorn, vilket kommer att kraftigt försämra de arbetslösas möjligheter att hitta ett nytt arbete.
Under 2009 beviljades Nederländerna dessutom samfinansiering från fonden för att stödja arbetstagare som sagts upp inom samma sektor och i samma Nuts II-region.
Kommissionen anser därför att uppsägningarna har allvarliga följder för sysselsättningen och den lokala ekonomin, och att dels den svåra ekonomiska situationen och osäkerheten på arbetsmarknaden i Noord-Brabant, dels de övriga uppsägningar som skett av samma orsaker och under samma tidsperiod inom samma huvudgrupp enligt Nace rev.
2 i andra nederländska Nuts II-regioner gör att ansökan uppfyller kriterierna i artikel 2 c i förordning (EG) nr 1927/2006.
Enligt de nederländska myndigheterna var det dessutom omöjligt att förutse den finansiella och ekonomiska krisen och vilka följder den skulle få för sektorn.
Kommissionens bedömning var också grundad på en beskrivning av regionen och de berörda myndigheterna och intressenterna.
Det samordnade paketet med personliga tjänster som ska finansieras, inbegripet dess förenlighet med de åtgärder som finansieras genom strukturfonderna, omfattar åtgärder för att på nytt integrera de berörda 199 arbetstagarna i anställning, exempelvis föreberedande åtgärder, rådgivning och utbildning.
Dessa personliga tjänster inleddes den 16 januari 2010.
De nederländska myndigheterna beaktade i sin ansökan och kompletterande information kriterierna i artikel 6 i förordning (EG) nr 1927/2006 genom att
• intyga att det ekonomiska bidraget från Europeiska fonden för justering för globaliseringseffekter inte ersätter åtgärder som företagen är skyldiga att vidta till följd av den nationella lagstiftningen eller kollektivavtal,
• visa att åtgärderna ger stöd till enskilda arbetstagare och inte ska användas för omstrukturering av företag eller sektorer,
• bekräfta att de aktuella åtgärder som avses ovan inte får stöd från andra finansiella EU-instrument.
När det gäller förvaltnings- och kontrollsystem har Nederländerna meddelat kommissionen att det ekonomiska stödet kommer att förvaltas och kontrolleras av samma organ som förvaltar och kontrollerar stödet från Europeiska socialfonden i Nederländerna.
Byrån för sociala frågor och sysselsättning kommer att vara förvaltningsmyndighetens förmedlande organ.
Kommissionen bedömer att ansökan uppfyller kriterierna för berättigande till stöd enligt förordningen om Europeiska fonden för justering för globaliseringseffekter och rekommenderar att budgetmyndigheterna bifaller ansökan.
För att utnyttja fonden har kommissionen överlämnat en begäran om överföring till budgetmyndigheten om ett sammanlagt belopp på 667 823 euro från reserven för Europeiska fonden för justering för globaliseringseffekter (40 02 43) för åtagandebemyndiganden till budgetpost 04 05 01.
Föredraganden välkomnar det faktum att 2011 års budget, efter upprepade uppmaningar från parlamentet, för första gången fastställer betalningsbemyndigandena (47 608 950 euro) under fondens budgetrubrik.
Föredraganden påminner om att fonden skapades som ett separat särskilt instrument med egna mål och tidsfrister och som sådant förtjänar ett målinriktat anslag, som innebär att man undviker överföringar från andra budgetposter, något som inträffade tidigare, och som kunde inverka negativt på uppfyllandet av de olika målen.
Enligt det interinstitutionella avtalet får fonden utnyttjas upp till det årliga taket på 500 miljoner euro.
Detta är det fjärde förslaget om utnyttjande av fonden som lämnats in till budgetmyndigheten under 2011.
Om man drar ifrån det aktuella begärda beloppet (667 823 euro) från de anslag som finns tillgängliga återstår därför ett tillgängligt belopp på 458 415 504 euro till slutet av 2011.
III.
Förfarandet
Kommissionen har lagt fram en begäran om överföring för att få med ett särskilt åtagandebemyndigande i 2011 års budget så som föreskrivs i punkt 28 i det interinstitutionella avtalet av den 17 maj 2006.
Enligt en intern överenskommelse ska utskottet för sysselsättning och sociala frågor delta i processen för att kunna ge konstruktivt stöd och bidra till bedömningen av ansökningar ur fonden.
Efter utvärdering ska Europaparlamentets utskott för sysselsättning och sociala frågor ge sin syn på användningen av fonden i en skrivelse som kommer att bifogas rapporten.
I Europaparlamentets, rådets och kommissionens gemensamma uttalande, som antogs under medlingsmötet den 17 juli 2008, bekräftades vikten av att säkerställa ett snabbt förfarande, med vederbörlig hänsyn till det interinstitutionella avtalet, för att anta beslut om utnyttjande av fonden.
BILAGA: SKRIVELSE FRÅN UTSKOTTET FÖR SYSSELSÄTTNING OCH SOCIALA FRÅGOR
ES/jm
D(2011)34759
Alain Lamassoure
Ordförande för budgetutskottet
ASP 13E158
Ärende: Yttrande om utnyttjandet av Europeiska fonden för justering för globaliseringseffekter i ärendet EGF/2010/027 NL/Noord-Brabant huvudgrupp 18 ( KOM(2011)0386 )
Till ordföranden
Utskottet för sysselsättning och sociala frågor (EMPL) och dess arbetsgrupp för Europeiska fonden för justering för globaliseringseffekter granskade utnyttjandet av fonden för ärende EGF/2010/027 NL/Noord-Brabant huvudgrupp 18 och antog följande yttrande.
EMPL-utskottet och arbetsgruppen för Europeiska fonden för justering för globaliseringseffekter är positiva till att fonden utnyttjas för denna ansökan.
I detta sammanhang vill EMPL-utskottet framföra vissa synpunkter, utan att därför ifrågasätta betalningsöverföringarna.
Enligt förordning (EEG) nr 1893/2006. som sades upp i Nuts II‑regionen Noord-Brabant i Nederländerna mellan den 16 januari och den 16 oktober 2010.
C) Kommissionen bekräftade i samband med bedömningen 2010 av andra ansökningar från samma sektor och regioner att den grafiska sektorn hade drabbats av den ekonomiska krisen.
D) Ansökan utgör en del av ett paket med fyra ansökningar som samtliga avser uppsägningar i sex olika Nuts II-regioner i Nederländerna med verksamhet i den grafiska sektorn.
Denna ansökan är främst kopplad till ansökningarna EGF/2010/029 NL/Zuid-Holland och Utrecht huvudgrupp 18, som lämnades in på grundval av artikel 2 b och EGF/2009/027 Noord-Brabant och Zuid Holland huvudgrupp 18 inom samma sektor och den angränsande Nuts II-regionen.
2.
F) De nederländska myndigheterna hävdar att trots en dyrbar omstrukturering av sektorn och insatserna för att förbereda arbetstagarna inför de nya arbetsmetoderna i en utbudsstyrd bransch, förlorade de nederländska företagen gentemot sina konkurrenter utanför EU samt att krisens negativa konsekvenser för sektorn inte kunde ha förutsetts.
G) Enligt de statistiska prognoserna kommer dessutom arbetsmarknaden för teknisk industri och bygg- och anläggningssektorn ytterligare att försämras, vilket kommer att kraftigt försämra de arbetslösas möjligheter att hitta ett nytt arbete.
I) 27,6 procent av de uppsagda arbetstagarna var process- och maskinoperatörer och montörer och 41,2 procent var fackmän och tekniker.
J) EU-budgeten för 2011 omfattar för första gången anslag till betalningar till EGF-fondens budgetpost 04 05 01 som också i detta fall överstiger överföringen av betalningar från andra oanvända budgetposter.
Utskottet för sysselsättning och sociala frågor uppmanar därför budgetutskottet att som ansvarigt utskott infoga följande förslag i sitt resolutionsförslag avseende Noord-Brabants ansökan:
1.
2.
Europaparlamentet gläder sig över att fondens bidrag är planerat att enbart stödja aktiva arbetsmarknadsåtgärder (utbildning och rådgivning) och inte kommer att användas för bidrag.
Med vänlig hälsning
Pervenche Berès
R ESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
8.9.2011
Slutomröstning: resultat
+:
–:
0:
26
1
Slutomröstning: närvarande ledamöter
Slutomröstning: närvarande suppleanter
Derk Jan Eppink, Roberto Gualtieri, Peter Šťastný, Georgios Stavrakakis
A7-0311/2011
BETÄNKANDE
om förslaget till Europaparlamentets och rådets beslut om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning (ansökan EGF/2011/003 DE/Arnsberg and Düsseldorf automotive från Tyskland)
(KOM(2011)0447 – C7‑0209/2011 – 2011/2163(BUD))
Budgetutskottet
Föredragande: Barbara Matera
PE 470.070v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
BILAGA: EUROPAPARLAMENTETS OCH RÅDETS BESLUT..............................................6
MOTIVERING............................................................................................................................8
BILAGA: SKRIVELSE FRÅN UTSKOTTET FÖR SYSSELSÄTTNING OCH SOCIALA FRÅGOR 12
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om förslaget till Europaparlamentets och rådets beslut om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning (ansökan EGF/2011/003 DE/Arnsberg and Düsseldorf automotive från Tyskland)
( KOM(2011)0447 – C7‑0209/2011 – 2011/2163(BUD) )
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2011)0447 – C7‑0209/2011 ),
– med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
EUT C 139, 14.6.2006, s.
1. , särskilt punkt 28,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1927/2006 av den 20 december 2006 om upprättande av Europeiska fonden för justering för globaliseringseffekter
EUT L 406, 30.12.2006, s.
1. ,
– med beaktande av trepartsförfarandet enligt punkt 28 i det interinstitutionella avtalet av den 17 maj 2006,
– med beaktande av skrivelsen från utskottet för sysselsättning och sociala frågor,
– med beaktande av betänkandet från budgetutskottet ( A7‑0311/2011 ), och av följande skäl:
A. Europeiska unionen har inrättat lagstiftningsinstrument och budgetinstrument för att ge extra stöd till arbetstagare som drabbats av konsekvenserna av de genomgripande strukturförändringar som skett inom världshandeln och för att underlätta deras återinträde på arbetsmarknaden.
B. Tillämpningsområdet för fonden har utvidgats, och från och med den 1 maj 2009 är det möjligt att söka stöd för åtgärder som riktas till arbetstagare som har blivit uppsagda som en direkt följd av den globala finansiella och ekonomiska krisen.
C. Unionens ekonomiska stöd till arbetstagare som har blivit uppsagda bör vara dynamiskt och ges så snabbt och effektivt som möjligt, i enlighet med Europaparlamentets, rådets och kommissionens gemensamma uttalande, som antogs vid förlikningsmötet den 17 juli 2008, och med vederbörlig hänsyn till det interinstitutionella avtalet av den 17 maj 2006 när det gäller antagandet av beslut om utnyttjande av fonden.
D. Tyskland har ansökt om medel från fonden med anledning av 778 uppsägningar, som alla omfattas av stödet, vid fem företag verksamma inom huvudgrupp 29 enligt Nace rev 2 (tillverkning av motorfordon, släpfordon och påhängsvagnar) i Nuts II-regionerna Arnsberg (DEA5) och Düsseldorf (DEA1) i Tyskland.
Europaparlamentet välkomnar den planerade förstärkningen av budgetposten för Europeiska fonden för justering för globaliseringseffekter 04 05 01 med 50 000 000 euro genom ändringsbudget 3/2011, som kommer att användas för att täcka det belopp som behövs för denna ansökan.
BILAGA: EUROPAPARLAMENTETS OCH RÅDETS BESLUT
av den ...
om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning (ansökan EGF/2011/003 DE/Arnsberg and Düsseldorf automotive från Tyskland)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA BESLUT
med beaktande av fördraget om Europeiska unionens funktionssätt,
med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
EUT C 139, 14.6.2006, s.
1. , särskilt punkt 28,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1927/2006 av den 20 december 2006 om upprättande av Europeiska fonden för justering för globaliseringseffekter
EUT L 406, 30.12.2006, s.
1. , särskilt artikel 12.3,
EUT C […], […], s. […]. , och
av följande skäl:
(2) Tillämpningsområdet för fonden har utvidgats, och från och med den 1 maj 2009 är det möjligt att söka stöd för åtgärder som riktas till arbetstagare som har blivit uppsagda som en direkt följd av den globala finansiella och ekonomiska krisen.
(3) Det interinstitutionella avtalet av den 17 maj 2006 gör det möjligt att använda medel från fonden upp till ett belopp på högst 500 miljoner euro per år.
(4) Tyskland lämnade den 9 februari 2011 in en ansökan om medel från fonden med anledning av uppsägningar vid fem företag som är verksamma inom huvudgrupp 29 (tillverkning av motorfordon, släpfordon och påhängsvagnar) enligt Nace rev 2, i Nuts 2-regionerna Arnberg (DEA5) och Düsseldorf (DEA1), och kompletterade ansökan med ytterligare uppgifter fram till den 28 april 2011.
Ansökan uppfyller villkoren för fastställande av det ekonomiska stödet enligt artikel 10 i förordning (EG) nr 1927/2006.
Kommissionen föreslår därför att ett belopp på 4 347 868 euro ska anslås.
(5) Fonden bör därför utnyttjas för att bevilja det ekonomiska stöd Tyskland ansökt om.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Europeiska fonden för justering för globaliseringseffekter ska belastas med 4 347 868 euro i åtagande- och betalningsbemyndiganden ur Europeiska unionens allmänna budget för 2011.
Artikel 2
Detta beslut ska offentliggöras i Europeiska unionens officiella tidning .
Utfärdat i [Bryssel/Strasbourg] den
På Europaparlamentets vägnar På rådets vägnar
Ordförande Ordförande
MOTIVERING
Europeiska fonden för justering för globaliseringseffekter inrättades för att ge kompletterande stöd till arbetstagare som blivit arbetslösa till följd av genomgripande strukturförändringar i världshandelsmönstret.
Enligt bestämmelserna i punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 om budgetdisciplin och sund ekonomisk förvaltning
EUT C 139, 14.6.2006, s.
1. samt i artikel 12 i förordning (EG) nr 1927/2006
EUT L 406, 30.12.2006, s.
1. , får det årliga belopp som avdelas för fonden inte överstiga 500 miljoner euro, och detta belopp får tas från outnyttjade marginaler under utgiftstaken för det föregående året samt från outnyttjade åtagandebemyndiganden som frigjorts under de två senaste åren, med undantag för sådana som ingår under rubrik 1b i budgetramen.
Anslagen förs in i budgeten i form av en avsättning så snart kommissionen har funnit tillräckliga marginaler och/eller frigjort åtaganden.
För att kunna ta fonden i anspråk ska kommissionen, efter en positiv prövning av ansökan, lägga fram ett förslag till budgetmyndigheten om utnyttjande av fonden tillsammans med en begäran om överföring.
Parallellt kan ett trepartsförfarande anordnas för att nå en överenskommelse om utnyttjande av fonden och de belopp som krävs.
Trepartsförfarandet kan ske i förenklad form.
II.
Aktuellt läge: Kommissionens förslag
Den 20 juli 2011 antog kommissionen ett nytt förslag till beslut om utnyttjande av Europeiska fonden för globaliseringseffekter till förmån för Tyskland för att stödja återintegrering på arbetsmarknaden av arbetstagare som har blivit uppsagda som en följd av den globala finansiella och ekonomiska krisen.
Detta är den femtonde ansökan som behandlas under budgetåret 2011 och den innebär en användning av totalt 4 347 868 euro ur fonden för Tysklands del.
Det gäller 778 uppsägningar, som alla omfattas av stödet, i fem företag verksamma inom huvudgrupp 29 (tillverkning av motorfordon, släpfordon och påhängsvagnar) enligt Nace rev 2 i Nuts 2‑regionerna Arnsberg (DEA5) och Düsseldorf (DEA1) i Tyskland, under referensperioden på nio månader från den 1 mars 2010 till den 1 december 2010.
Denna ansökan, ärende EGF/2011/003 DE/Arnsberg och Düsseldorf automotive från Tyskland, lämnades in till kommissionen den 9 februari 2011 och kompletterades med ytterligare uppgifter fram till den 28 april 2011.
Ansökan grundades på interventionskriteriet i artikel 2 b i förordningen om Europeiska fonden för justering för globaliseringseffekter enligt vilka minst 500 arbetstagare ska ha sagts upp under en referensperiod på nio månader vid företag som är verksamma inom en Nace rev.
2-sektor i en region eller två regioner som gränsar till varandra på Nuts II-nivå i en medlemsstat.
Ett av kriterierna för kommissionens bedömning var utvärderingen av kopplingen mellan uppsägningarna och stora strukturella förändringar i världshandelsmönstren eller finanskrisen, vilket i just detta fall hör samman med den minskade efterfrågan på nya motorfordon i Europeiska unionen till följd av den finansiella och ekonomiska krisen.
Som ett resultat av denna minskade produktionen av motorfordon i Tyskland med 13,8 % under 2009 jämfört med 2008 och med 14 % under 2010 jämfört med 2008.
Denna plötsliga drastiska krisrelaterade minskning i efterfrågan på motorfordon, som inte kunde förutses, ledde, enligt de tyska myndigheterna, dessutom till en betydande minskning av utnyttjandet av produktionskapaciteten och till en kraftig minskning av intäkterna för leverantörerna inom motorfordonsindustrin.
Enligt de tyska myndigheterna kommer de 778 uppsägningar som omfattas av denna ansökan att ytterligare bidra till en ökning av arbetslösheten i regionerna Arnsberg och Düsseldorf, som redan allvarligt drabbats genom avskedandena hos Nokia i Bochum och stängningen av General Motors.
Det samordnade paket med individanpassade tjänster som ska finansieras, inbegripet dess komplementaritet med åtgärder som finansieras genom strukturfonderna, omfattar följande åtgärder:
– Kortfristigt understöd till arbetssökande - under den tid som arbetstagarna deltar i aktiva arbetsmarknadspolitiska åtgärder.
– Fortbildning - riktad till friställda arbetstagare som saknar erkända yrkeskvalifikationer eller vars kvalifikationer behöver uppdateras, men också till industriarbetare.
– Rådgivning om företagsetablering - vägledning och stöd för genomförande och finansiering av företagsetableringar.
– Seminarier och gruppdiskussioner - handledning och erfarenhetsutbyte i små grupper av arbetstagare med liknande yrkesbakgrund.
– Vägledning på den internationella och nationella arbetsmarknaden - förbereda ett antal arbetstagare för jobb utanför regionen, och även utanför Tyskland.
– Aktiveringstillägg - incitament för arbetstagare som tar ett nytt jobb med lägre lön.
– Platssökning - särskilda personer kommer att hålla kontakt med potentiella arbetsgivare och söka efter de lämpligaste kandidaterna för de lediga platser som finns samt kartlägga de yrkesspecifika utbildningsbehov kandidaterna har.
– Handledning och stöd för arbetstagare som hittat ett nytt arbete och till arbetslösa arbetstagare - att hjälpa arbetstagare att anpassa sig till det nya jobbet och stödja arbetstagare som befinner sig i arbetslöshet.
När det gäller kriterierna i artikel 6 i förordning (EG) nr 1927/2006 intygade eller meddelade de tyska myndigheterna följande i sin ansökan och kompletterande information:
• Det ekonomiska bidraget från Europeiska fonden för justering för globaliseringseffekter ersätter inte åtgärder som företagen är skyldiga att vidta till följd av den nationella lagstiftningen eller kollektivavtal.
• Åtgärderna ger stöd till enskilda arbetstagare och ska inte användas för omstrukturering av företag eller sektorer.
• De bidragsberättigande åtgärder som avses ovan får inte stöd från något annat av EU:s finansieringsinstrument.
När det gäller förvaltnings- och kontrollsystemen har Tyskland meddelat kommissionen att det ekonomiska stödet kommer att förvaltas och kontrolleras av samma organ som förvaltar och kontrollerar stödet från Europeiska socialfonden.
Kommissionens bedömer att ansökan uppfyller kriterierna för berättigande till stöd enligt förordningen om Europeiska fonden för justering för globaliseringseffekter och rekommenderar att budgetmyndigheterna bifaller ansökan.
För att utnyttja fonden har kommissionen överlämnat en begäran om överföring till budgetmyndigheten av ett sammanlagt belopp på 4 347 868 euro från reserven för Europeiska fonden för justering för globaliseringseffekter (40 02 43) i åtagandebemyndiganden till fondens budgetpost 04 05 01.
Föredraganden välkomnar det faktum att 2011 års budget, efter upprepade uppmaningar från parlamentet, för första gången visar betalningsbemyndigandena (47 608 950 euro) under fondens budgetpost och välkomnar förstärkningen av budgetpost 04 05 01 med 50 000 000 euro såsom förutses genom ÄB 3/2011.
Föredraganden påminner om att fonden skapades som ett separat särskilt instrument med egna mål och tidsfrister och som sådant förtjänar ett eget anslag, vilket innebär att man undviker överföringar från andra budgetposter, något som inträffade tidigare och som kunde inverka negativt på uppfyllandet av de olika målen.
Enligt det interinstitutionella avtalet får fonden utnyttjas upp till det årliga taket på 500 miljoner euro.
Detta är det femtonde förslaget om utnyttjande av fonden som lämnats in till budgetmyndigheten under 2011.
Om man drar ifrån det aktuella begärda beloppet (4 347 868 euro) från de anslag som finns tillgängliga återstår därför ett tillgängligt belopp på 420 413 131 euro till slutet av 2011.
III.
Förfarandet
Kommissionen har lagt fram en begäran om överföring för att införa specifika åtagandebemyndiganden i 2011 års budget, såsom föreskrivs i punkt 28 i det interinstitutionella avtalet av den 17 maj 2006.
Enligt en intern överenskommelse ska utskottet för sysselsättning och sociala frågor delta i processen för att konstruktivt stödja och bidra till bedömningen av ansökningarna om medel ur fonden.
Efter sin bedömning kommer Europaparlamentets utskott för sysselsättning och sociala frågor att lägga fram sina synpunkter på utnyttjandet av fonden, vilka kommer att bifogas som en skrivelse till detta betänkande.
I Europaparlamentets, rådets och kommissionens gemensamma uttalande, som antogs under förlikningsmötet den 17 juli 2008, bekräftades vikten av att säkerställa ett snabbt förfarande, med vederbörlig hänsyn till det interinstitutionella avtalet, för att anta beslut om utnyttjande av fonden.
BILAGA: SKRIVELSE FRÅN UTSKOTTET FÖR SYSSELSÄTTNING OCH SOCIALA FRÅGOR
EK/jm
D(2011)44589
Alain Lamassoure
Ordförande för budgetutskottet
ASP 13E158
Ärende: Yttrande över utnyttjande av Europeiska fonden för justering för globaliseringseffekter för ansökan EGF/2011/003 DE/Arnsberg and Düsseldorf automotive från Tyskland ( KOM(2011)0447 )
EMPL-utskottet och arbetsgruppen för Europeiska fonden för justering för globaliseringseffekter är positiva till att fonden utnyttjas för denna ansökan.
I detta sammanhang vill EMPL-utskottet framföra vissa synpunkter, utan att därför ifrågasätta betalningsöverföringarna.
EMPL-utskottets synpunkter grundar sig på följande överväganden:
A) Denna ansökan bygger på artikel 2b i förordningen för Europeiska fonden för justering för globaliseringseffekter och gäller 778 arbetstagare i huvudgrupp 29 Nace rev.
2 i Nuts II‑regionerna Arnsberg och Düsseldorf som sades upp under referensperioden mellan den 1 mars 2010 och den 1 december 2010.
C) Denna ansökan avser främst uppsägningar hos underleverantörer, där omsättningen minskade med 26 procent mellan 2008 och 2009.
D) De tyska myndigheterna anför vidare att underleverantörerna under en tid hade verkat under press från fordonstillverkarna för att minska sina marginaler och därför drabbades särskilt hårt av den plötsliga och svåra kris som ledde till en kraftig minskning av produktionskapacitetsutnyttjandet och ett kraftigt inkomstbortfall för underleverantörerna i fordonsindustrin med ett stort antal konkurser som följd vilka alla medförde personalminskningar.
E) Kommissionen har redan i tidigare ansökningar rörande fordonsindustrin bekräftat att den finansiella och ekonomiska krisen i synnerhet drabbat biltillverkarna och deras underleverantörer mot bakgrund av att 60 till 80 procent av all nya bilar som säljs i Europa köps på kredit.
G) 66,5 procent av de uppsagda arbetstagarna tillhör antingen kategorin arbetare inom hantverksarbete, byggverksamhet och tillverkning eller process- och maskinoperatörer samt montörer och 11,3 procent av dem hade varit anställda i lågkvalificerade yrken.
H) Kommissionen informerade EMPL-utskottet om att ändringsbudget nr 3
Utskottet för sysselsättning och sociala frågor uppmanar därför budgetutskottet att som ansvarigt utskott infoga följande förslag i sitt resolutionsförslag avseende Tysklands ansökan:
1.
Europaparlamentet instämmer med kommissionen att villkoren för ekonomiskt stöd enligt artikel 2b i förordningen om Europeiska fonden för justering för globaliseringseffekter (1927/2006) är uppfyllda och att Tyskland därför är berättigat till stöd enligt förordningen.
3.
Europaparlamentet noterar denna första tyska ansökan baserad på artikel 2b och det faktum att varje företag har inrättat sitt eget övergångsföretag för att förverkliga det samordnade paketet med individanpassade tjänster.
Europaparlamentet välkomnar möjligheten för arbetstagare utan erkänd utbildning eller med föråldrade kvalifikationer att delta i intensivutbildning i syfte att förvärva kompetens som motsvarar den enskildes önskemål och förutsättningar och arbetsmarknadens behov.
Med vänlig hälsning
R ESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
22.9.2011
Slutomröstning: resultat
+:
–:
0:
17
3
2
Slutomröstning: närvarande ledamöter
Slutomröstning: närvarande suppleanter
Maria Da Graça Carvalho, Jan Mulder
Slutomröstning: närvarande suppleanter (art.
187.2)
Kinga Gál
A7-0342/2011
Föredragande: Jürgen Creutzmann
PE 467.028v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING..........................................................................................................................14
YTTRANDE från utskottet för ekonomi och valutafrågor ....................17
YTTRANDE från utskottet för rättsliga frågor ...........................................22
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................27
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om hasardspel online på den inre marknaden
( 2011/2084(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens meddelande av den 24 mars 2011 med titeln ”Grönbok om onlinespel på den inre marknaden” ( KOM(2011)0128 ),
– med beaktande av artiklarna 51, 52 och 56 i fördraget om Europeiska unionens funktionssätt,
– med beaktande av protokollet om tillämpning av subsidiaritets- och proportionalitetsprinciperna, fogat till fördraget om Europeiska unionens funktionssätt,
– med beaktande av EU-domstolens relevanta rättspraxis
2010 (C-316/07, C-358/07, C-359/07, C-360/07, C-409/07 och C-410/07), Carmen Media 2010 (C-46/08) och Engelmann 2010 (C-64/08). ,
– med beaktande av rådets slutsatser av den 10 december 2010 och lägesrapporterna från de franska, svenska, spanska och ungerska rådsordförandeskapen om ramen för spel och vadhållning i EU‑medlemsstaterna,
– med beaktande av sin resolution av den 10 mars 2009 om integriteten för hasardspel online
EUT C 87 E, 1.4.2010, s.
30. ,
– med beaktande av sin resolution av den 8 maj 2008 om vitboken om idrott
EUT C 271 E, 12.11.2009, s.
51. ,
– med beaktande av Europaparlamentets och rådets direktiv 2010/13/EU av den 10 mars 2010 om samordning av vissa bestämmelser som fastställs i medlemsstaternas lagar och andra författningar om tillhandahållande av audiovisuella medietjänster
EUT L 95, 15.4.2010, s.
1. ,
– med beaktande av Europaparlamentets och rådets direktiv 2005/29/EG av den 11 maj 2005 om otillbörliga affärsmetoder som tillämpas av näringsidkare gentemot konsumenter på den inre marknaden och om ändring av rådets direktiv 84/450/EEG och Europaparlamentets och rådets direktiv 97/7/EG, 98/27/EG och 2002/65/EG samt Europaparlamentets och rådets förordning (EG) nr 2006/2004
EUT L 149, 11.6.2005, s.
22. ,
– med beaktande av Europaparlamentets och rådets direktiv 97/7/EG av den 20 maj 1997 om konsumentskydd vid distansavtal
EGT L 144, 4.6.1997, s.
19. ,
– med beaktande av Europaparlamentets och rådets direktiv 2005/60/EG av den 26 oktober 2005 om åtgärder för att förhindra att det finansiella systemet används för penningtvätt och finansiering av terrorism
EUT L 309, 25.11.2005, s.
15. ,
– med beaktande av kommissionens meddelande av den 6 juni 2011 med titeln ”Insatser mot korruption på EU:s territorium”,
– med beaktande av Europaparlamentets och rådets direktiv 95/46/EG av den 24 oktober 1995 om skydd för enskilda personer med avseende på behandling av personuppgifter och om det fria flödet av sådana uppgifter
EGT L 281, 23.11.1995, s.
31. ,
– med beaktande av Europaparlamentets och rådets direktiv 2002/58/EG av den 12 juli 2002 om behandling av personuppgifter och integritetsskydd inom sektorn för elektronisk kommunikation
EGT L 201, 31.7.2002, s.
37. ,
– med beaktande av kommissionens meddelande av den 18 januari 2011 med titeln ”Utveckling av idrottens europeiska dimension”,
– med beaktande av rådets direktiv 2006/112/EG av den 28 november 2006 om ett gemensamt system för mervärdesskatt
EUT L 347, 11.12.2006, s.
1. ,
– med beaktande av Europaparlamentets och rådets direktiv 2006/123/EG av den 12 december 2006 om tjänster på den inre marknaden
EUT L 376, 27.12.2006, s.
36. ,
– med beaktande av Europaparlamentets och rådets direktiv 2000/31/EG av den 8 juni 2000 om vissa rättsliga aspekter på informationssamhällets tjänster, särskilt elektronisk handel, på den inre marknaden
EGT L 178, 17.7.2000, s.
1. ,
– med beaktande av artikel 48 i arbetsordningen,
– med beaktande av betänkandet från utskottet för den inre marknaden och konsumentskydd och yttrandena från utskottet för ekonomi och valutafrågor samt utskottet för rättsliga frågor (A7‑.../2011), och av följande skäl:
B. Tillämpningen av subsidiaritetsprincipen gör att det inte finns någon särskild europeisk lagstiftningsakt för reglering av hasardspel online.
C. Speltjänster omfattas av ett antal EU-rättsakter, såsom direktivet om audiovisuella medietjänster, direktivet om otillbörliga affärsmetoder, direktivet om konsumentskydd vid distansavtal, direktivet om åtgärder för att förhindra penningtvätt, dataskyddsdirektivet, direktivet om integritet och elektronisk kommunikation och direktivet om ett gemensamt system för mervärdesskatt.
D. Sektorn för hasardspel regleras på olika sätt i olika medlemsstater, vilket inte bara gör det svårt för reglerade aktörer att erbjuda lagliga gränsöverskridande speltjänster, utan också gör det svårt för tillsynsmyndigheterna att skydda konsumenterna och bekämpa olagliga hasardspel online och eventuella brott som har samband med sådana spel på EU-nivå.
E. Det finns ett mycket stort mervärde i att agera på EU-nivå för att bekämpa brottslighet och bedrägerier och i synnerhet för att slå vakt om idrottens integritet och skydda spelare och konsumenter.
F. I artikel 56 i EUF-fördraget garanteras friheten att tillhandahålla tjänster.
I. Konsumenterna måste informeras om de eventuellt skadliga effekterna av hasardspel online och skyddas mot faror på detta område, särskilt beroende, bedrägerier, svindel och minderårigas spel.
J. Hasardspel utgör en betydande inkomstkälla som de flesta medlemsstater använder för allmännyttiga och välgörande ändamål, till exempel idrott.
K. Idrottens integritet måste ovillkorligen garanteras genom att man förstärker kampen mot korruption och riggade matcher.
Europaparlamentet välkomnar kommissionens klargörande att den politiska process som inletts i och med grönboken absolut inte syftar till en avreglering/liberalisering av hasardspel online, och gläder sig över att kommissionen i sin grönbok tar hänsyn till parlamentets tydliga och konsekventa ståndpunkt om hasardspel.
1) styra människors naturliga drift att spela genom att begränsa marknadsföringen till vad som är absolut nödvändigt för att informera potentiella spelare om var de kan spela lagligt och genom att kräva att all marknadsföring av hasardspel online systematiskt ska åtföljas av en varning för överdrivet eller patologiskt spelande,
2) bekämpa den olagliga sektorn för hasardspel genom att stärka de tekniska och rättsliga möjligheterna att upptäcka och straffa olagliga aktörer och genom att verka för ett utbud av lagliga speltjänster av hög kvalitet,
3) säkerställa ett effektivt skydd för spelare, i synnerhet för minderåriga och andra sårbara grupper,
4) förebygga riskerna för beroende vid hasardspel,
5) säkerställa att hasardspel genomförs under korrekta, rättvisa, ansvarsfulla och öppna former,
6) verka för konkreta åtgärder som garanterar idrottstävlingarnas integritet,
7) säkerställa att en del av de pengar som satsas går till idrotten och hästsporten,
8) säkerställa att en betydande del av de offentliga intäkterna från hasardspel används för att främja allmännyttiga eller välgörande ändamål, och
9) säkerställa att spelmarknaden är fri från brott, bedrägerier och alla former av penningtvätt.
Subsidiaritetsprincipen och EU:s mervärde
Europaparlamentet betonar att medlemsstaterna har rätt att reglera och kontrollera sina spelmarknader i enlighet med EU:s lagstiftning om den inre marknaden, sina traditioner och sin kultur.
Europaparlamentet betonar vikten av att få spelare att avstå från olagliga hasardspel, vilket förutsätter att det finns ett lagligt utbud inom ramen för ett system som är enhetligt i EU, särskilt när det gäller beskattning, och som tillämpar gemensamma minimistandarder för ansvarsskyldighet och integritet.
Europaparlamentet påpekar att EU-domstolen i ett flertal domar har godtagit att beviljandet av exklusiva rättigheter till en enskild aktör som står under strikt offentlig övervakning kan vara ett sätt att bättre skydda konsumenterna mot bedrägerier och att mer effektivt bekämpa brottslighet inom sektorn för hasardspel online.
Europaparlamentet understryker att leverantörer av hasardspel online alltid måste följa den nationella lagstiftningen i de länder där spelet bedrivs samt att medlemsstaterna alltjämt bör ha exklusiv rätt att införa alla åtgärder de anser nödvändiga för att bekämpa olagliga hasardspel online i syfte att tillämpa den nationella lagstiftningen och strypa tillgången till marknaden för olagliga leverantörer.
Samarbete mellan tillsynsmyndigheter
Europaparlamentet betonar särskilt att ”spread betting”, en form av hasardspel som huvudsakligen sker online och där konsumenterna potentiellt kan förlora många gånger sin ursprungliga insats, måste vara föremål för mycket strikta villkor för konsumenttillgång och bör vara reglerat, vilket redan är fallet i många medlemsstater, i likhet med vad som gäller för finansiella derivat.
Europaparlamentet uppmanar kommissionen att initiera bildandet av ett nätverk med nationella organisationer som tar hand om spelberoende för att möjliggöra utbyte av erfarenheter och bästa praxis.
”Cross-Border Alternative Dispute Resolution in the European Union”, 2011,
Hasardspel och idrott – behovet av att garantera integriteten
46.
MOTIVERING
Sektorn för hasardspel online ökar stadigt.
Enligt aktuella uppgifter äger i dag 10 procent av alla hasardspel i Europa rum på internet eller via liknande förmedlingskanaler, såsom mobiltelefoner eller interaktiva TV-plattformar.
Denna andel blir allt större och marknadsvolymen överstiger nu 10 miljarder euro.
Marknaden för platsbaserade hasardspel och marknaden för onlinespel kännetecknas av ett brett produktutbud: å ena sidan klassiska lottospel och lotterier, men också sportvadslagning, poker, bingospel och vadslagning vid häst- och hundkapplöpningar enligt totalisatormetoden.
Internet är till sin natur ett gränsöverskridande medium.
Hasardspel online låter sig därför inte stoppas av gränser.
Men eftersom utbudet och antalet spelare hela tiden ökar blir också den rådande fragmenteringen av marknaden i Europa på detta område allt tydligare.
I många medlemsstater råder totalförbud eller förbud med möjlighet att bevilja tillstånd, andra har en helt öppen och liberaliserad marknad.
Som EU-domstolen har konstaterat i flera domar är hasardspel inte standardtjänster.
Därför har de uttryckligen uteslutits ur tjänstedirektivet även om det fria tillhandahållandet av tjänster enligt artikel 56 i EUF-fördraget naturligtvis även gäller för hasardspel.
Medlemsstaterna kan bland annat på grundval av artiklarna 51 och 52 i EUF-fördraget i stor utsträckning själva reglera sina marknader så länge dessa bestämmelser är förenliga med de mål som ska uppnås, till exempel att bekämpa spelberoende.
På grund av att traditionerna skiljer sig avsevärt åt är subsidiaritetsprincipen av särskilt stor betydelse inom denna sektor.
Medlemsstaterna beslutar i stor utsträckning själva hur de vill reglera sin spelmarknad.
Men dessa starkt varierande bestämmelser medför också att marknaden på internet snedvrids.
Hasardspelsaktörer i medlemsstater med öppna marknader och låga skatter kan också nås i länder där hasardspel online är förbjudet eller så konkurrerar de med onlineaktörer som har tillstånd.
Dessa aktörer och aktörer med platsbaserade hasardspel i dessa länder har svårt att hävda sig i konkurrensen.
Dessutom finns det en oreglerad svart marknad på internet av betydande omfattning.
Därför måste det centrala målet vara att avsevärt begränsa denna svarta och gråa marknad.
Medlemsstaterna kan på grundval av subsidiaritetsprincipen besluta sig för detta alternativ.
Ett bättre alternativ vore att skapa ett lagligt utbud av hasardspel online.
Detta får dock under inga omständigheter leda till att det skapas ett (statligt) monopol för hasardspel online eftersom monopol endast sällan säkerställer ett tillräckligt utbud.
Följaktligen bör marknaden öppnas upp och tillräckliga incitament skapas för företag att erbjuda ett lagligt utbud.
För att uppnå detta är en modell med tillstånd det bästa sättet, under förutsättning att den bygger på principen om konkurrens utan diskriminering.
I detta system, som med framgång redan har införts i några medlemsstater, som Frankrike och Italien, fastställer nationella tillsynsmyndigheter villkoren för att bevilja tillstånd.
Sedan systemet med tillstånd infördes har andelen aktörer med tillstånd i till exempel Frankrike ökat snabbt: aktörer med tillstånd svarar nu för mer än 80 procent av den franska marknaden för hasardspel online.
En förutsättning för en öppen och ordnad marknad för hasardspel online är en oberoende och stark nationell tillsynsmyndighet.
Den måste fastställa ramvillkoren för hasardspel och framför allt även kunna genomdriva dem.
Nationella tillsynsmyndigheter måste således få erforderlig behörighet för att beivra överträdelser och vidta åtgärder mot aktörer utan tillstånd.
Eftersom internet till sin natur är gränsöverskridande kan inte medlemsstaterna på egen hand reglera alla områden av hasardspel online.
Därför krävs ett starkt utökat samarbete mellan de nationella tillsynsmyndigheterna.
Hittills förekommer samarbete endast i liten omfattning, till exempel i form av bilaterala förfaranden.
Men det skulle behövas institutionaliserat samarbete, till exempel på grundval av informationssystemet för den inre marknaden, för att snabbt och effektivt utbyta information.
Även ett utbyggt nätverk av tillsynsmyndigheter som samordnas av kommissionen är tänkbart.
Endast med en gemensam europeisk strategi går det att förhindra att aktörer utan tillstånd utnyttjar luckor i regelverket och spelar ut nationella tillsynsmyndigheter mot varandra.
Därför krävs att kommissionen och medlemsstaterna handlar snabbt för att skydda konsumenterna i EU mot oseriösa aktörer.
Hasardspel medför en risk för beroende.
Studier visar att sedan hasardspel online introducerades för ungefär 10 år sedan har antalet människor som vänder sig till stödcenter för spelberoende ökat markant.
Det finns redan åtskilliga initiativ, både från tillsynsmyndigheter och i form av uppförandekoder och frivilliga åtaganden, som försöker begränsa problemspelande och spelberoende på internet.
Men det leder knappast till några resultat om varje medlemsstat tillämpar olika standarder.
Till exempel krävs i en del medlemsstater en elektronisk legitimation för identitetskontroll på internet.
Utlänningar har ofta inte en sådan legitimation och är därför uteslutna från hasardspel online, även om de är varaktigt bosatta i denna medlemsstat.
Därför är det viktigt med europeiska tekniska standarder som kan utarbetas gemensamt av branschen, konsumentskyddsorganisationer och kommissionen.
De minskar också hindren för marknadstillträde för hasardspelsaktörer från andra europeiska länder.
Låga hinder för marknadstillträde är en viktig åtgärd för att skapa en laglig och reglerad spelmarknad.
Skydd av minderåriga mot hasardspel är ett annat generellt mål som inte är beroende av olika traditioner eller kulturer.
Det ligger därför nära till hands att på EU-nivå fastställa minimistandarder för att skydda minderåriga, förhindra spelberoende men även bekämpa penningtvätt och annan brottslighet relaterad till hasardspel.
Detta skulle kunna ske i form av ett förslag till direktiv från kommissionen där det fastställs minimistandarder som gäller i hela EU och som är bindande för alla leverantörer av hasardspel online som har tillstånd.
Därutöver skulle det stå medlemsstaterna fritt att fastställa ytterligare kriterier.
Beslutsamt handlande från kommissionens och medlemsstaternas sida är viktigt för att i hela EU säkerställa en enhetlig och hög minimiskyddsnivå för konsumenterna.
I de flesta medlemsstater bidrar intäkterna från hasardspel till välgörande eller allmännyttiga ändamål och till att främja idrotten.
Men detta gäller endast för lagliga spelaktörer med tillstånd.
Aktörer utan tillstånd betalar ingen skatt och lämnar följaktligen inte heller några bidrag till samhället.
En marknad som regleras på nationell nivå skulle medföra att leverantörerna av hasardspel online blev tvungna att betala en stor del av skatterna på spel i spelarens land.
Detta är viktigt för att de offentliga intäkterna från hasardspel i hela Europa ska kunna användas för att främja idrott och andra allmännyttiga ändamål.
Vid till exempel hästkapplöpningar kan det på detta sätt säkerställas att uppfödarna får en del av intäkterna från vadslagning som behövs för fortsatt finansiering av uppfödningen.
Tyvärr har det tidigare gång på gång förekommit vadslagningsbedrägerier inom idrotten som äventyrar idrottens integritet.
Alla berörda parter – det vill säga idrottsföreningarna, supportrarna, spelaktörerna och spelarna – har ett direkt intresse av att trygga idrottens integritet och stoppa vadslagningsbedrägerier.
Vadslagningsbedrägerier kan bäst förebyggas på EU-nivå.
Därför bör kommissionen gemensamt med medlemsstaterna utveckla ett system som effektivt förhindrar vadslagningsbedrägerier.
Ett gemensamt agerande mot vadslagningsbedrägerier får också större tyngd gentemot utomeuropeiska kriminella vadslagningsbedragare.
För att bevara idrottens integritet måste intressekonflikter mellan aktörer inom sportvadslagning och idrottsföreningar undvikas.
Men enbart reklam för hasardspel eller sponsring av en idrottsförening utgör i sig inte en intressekonflikt.
YTTRANDE från utskottet för ekonomi och valutafrågor
till utskottet för den inre marknaden och konsumentskydd
över hasardspel online på den inre marknaden
( 2011/2084(INI) )
Föredragande: Sophie Auconie
FÖRSLAG
Utskottet för ekonomi och valutafrågor uppmanar utskottet för den inre marknaden och konsumentskydd att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet betonar särskilt att spread betting, en form av hasardspel som huvudsakligen sker online och där konsumenterna potentiellt kan förlora många gånger sin ursprungliga insats, måste vara föremål för mycket strikta villkor för konsumenttillgång och bör vara reglerad, vilket redan är fallet i många medlemsstater, i likhet med vad som gäller för finansiella derivat.
Europaparlamentet är positivt till en rättslig definition av minimistandarder för konsumentskydd, särskilt för de mest sårbara konsumenterna, utan att detta påverkar medlemsstaternas rätt att anta en strängare lagstiftning.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
31.8.2011
Slutomröstning: resultat
+:
–:
0:
38
2
Slutomröstning: närvarande ledamöter
Burkhard Balz, Sharon Bowles, Udo Bullmann, Pascal Canfin, Nikolaos Chountis, Rachida Dati, Leonardo Domenici, Diogo Feio, Markus Ferber, Ildikó Gáll-Pelcz, José Manuel García-Margallo y Marfil, Jean-Paul Gauzès, Sven Giegold, Liem Hoang Ngoc, Jürgen Klute, Philippe Lamberts, Astrid Lulling, Arlene McCarthy, Sławomir Witold Nitras, Ivari Padar, Alfredo Pallone, Antolín Sánchez Presedo, Olle Schmidt, Edward Scicluna, Theodor Dumitru Stolojan, Ivo Strejček, Marianne Thyssen, Corien Wortmann-Kool,
Slutomröstning: närvarande suppleant(er)
Sophie Auconie, Pervenche Berès, Herbert Dorfmann, Sari Essayah, Vicky Ford, Ashley Fox, Olle Ludvigsson, Thomas Mann, Sirpa Pietikäinen, Andreas Schwab, Theodoros Skylakakis, Catherine Stihler
Slutomröstning: närvarande suppleant(er) (art.
187.2)
Kriton Arsenis (S&D), Knut Fleckenstein (S&D), Bill Newton Dunn (ALDE)
13.7.2011
över hasardspel online på den inre marknaden
Föredragande:
Sajjad Karim
FÖRSLAG
Utskottet för rättsliga frågor uppmanar utskottet för den inre marknaden och konsumentskydd att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
De förenade målen C–316/07, C–358/07, C–359/07, C–360/07, C–409/07 och C–410/07, Markus Stoß, ännu ej offentliggjorda. har klargjort att medlemsstaternas lagstiftningsmässiga begränsningar måste vara motiverade och sammanhängande och måste överensstämma med de rättsliga mål som eftersträvas i syfte att skydda konsumenterna, förhindra bedrägerier och skydda den allmänna ordningen.
6.
Europaparlamentet konstaterar att det hade kunnat göras fler framsteg i de överträdelseförfaranden som pågår sedan 2008 och att det aldrig har inletts något ärende i EU-domstolen mot en enskild medlemsstat.
Europaparlamentet bekräftar sin ståndpunkt att vadslagning om idrott är ett slags kommersiell användning av idrottstävlingar, och rekommenderar att kommissionen och medlemsstaterna ska skydda idrottstävlingar från otillåten kommersiell användning, framför allt genom att erkänna idrottsorganens äganderätt till tävlingar som de anordnar, detta inte bara för att garantera en skälig ekonomisk vinst på alla nivåer av professionell idrott och amatöridrott, utan också för att stärka kampen mot uppgjorda matcher.
Europaparlamentet uppmanar kommissionen att lägga fram meningsfulla lagstiftningsförslag som kan utgöra en rättslig ram som ger de europeiska företagen säkerhet beträffande rättsläget och skyddar konsumenterna.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
11.7.2011
Slutomröstning: resultat
+:
–:
0:
22
Slutomröstning: närvarande ledamöter
Raffaele Baldassarre, Luigi Berlinguer, Sebastian Valentin Bodu, Françoise Castex, Christian Engström, Marielle Gallo, Klaus-Heiner Lehne, Antonio Masip Hidalgo, Bernhard Rapkay, Evelyn Regner, Francesco Enrico Speroni, Dimitar Stoyanov, Alexandra Thein, Rainer Wieland, Cecilia Wikström, Tadeusz Zwiefka
Slutomröstning: närvarande suppleanter
Kurt Lechner, Eva Lichtenberger, Toine Manders, Paulo Rangel, Dagmar Roth-Behrendt
Slutomröstning: närvarande suppleanter (art.
187.2)
Giuseppe Gargani
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
6.10.2011
Slutomröstning: resultat
+:
–:
0:
30
1
3
Slutomröstning: närvarande ledamöter
Adam Bielan, Lara Comi, Anna Maria Corazza Bildt, António Fernando Correia De Campos, Jürgen Creutzmann, Christian Engström, Evelyne Gebhardt, Louis Grech, Małgorzata Handzlik, Iliana Ivanova, Edvard Kožušník, Kurt Lechner, Toine Manders, Hans-Peter Mayer, Phil Prendergast, Mitro Repo, Robert Rochefort, Zuzana Roithová, Christel Schaldemose, Andreas Schwab, Emilie Turunen, Bernadette Vergnaud, Barbara Weiler
Slutomröstning: närvarande suppleanter
Marielle Gallo, Anna Hedh, Constance Le Grip, Emma McClarkin, Sylvana Rapti, Oreste Rossi, Wim van de Camp
Slutomröstning: närvarande suppleanter (art.
187.2)
Alexander Alvaro, Monika Hohlmeier, Axel Voss, Pablo Zalba Bidegain
A7-0371/2011
24.10.2011
BETÄNKANDE
om reform av EU:s regler om statligt stöd avseende tjänster av allmänt ekonomiskt intresse
(2011/2146(INI))
Utskottet för ekonomi och valutafrågor
Föredragande: Peter Simon
PE 469.843v03-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING..........................................................................................................................11
YTTRANDE från utskottet för industrifrågor, forskning och energi 14
YTTRANDE från utskottet för den inre marknaden och konsumentskydd 17
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................20
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om reform av EU:s regler om statligt stöd avseende tjänster av allmänt ekonomiskt intresse
( 2011/2146(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av artiklarna 14 och 16 i fördraget om Europeiska unionens funktionssätt samt protokoll nr 26 till detta,
– med beaktande av meddelandet från kommissionen av den 23 mars 2011: Reform av EU:s regler om statligt stöd avseende tjänster av allmänt ekonomiskt intresse ( KOM(2011)0146 ),
– med beaktande av kommissionens arbetsdokument av den 23 mars 2011 som behandlar tillämpningen av EU:s statsstödsregler på tjänster av allmänt ekonomiskt intresse sedan 2005 och resultaten från det offentliga samrådet ( SEK(2011)0397 ),
– med beaktande av det offentliga samråd som kommissionen anordnade 2010 om regler om statligt stöd avseende tjänster av allmänt ekonomiskt intresse,
– med beaktande av ”Vägledning om hur Europeiska unionens bestämmelser om statligt stöd, offentlig upphandling och den inre marknaden ska tillämpas på tjänster av allmänt ekonomiskt intresse, särskilt sociala tjänster av allmänt intresse” av den 7 december 2010 ( SEK(2010)1545 ),
– med beaktande av kommissionens direktiv 2006/111/EG av den 16 november 2006 om insyn i de finansiella förbindelserna mellan medlemsstater och offentliga företag samt i vissa företags ekonomiska verksamhet
EUT L 318, 17.11.2006, s.
17. ,
– med beaktande av kommissionens beslut 2005/842/EG av den 28 november 2005 om tillämpningen av artikel 86.2 i EG-fördraget på statligt stöd i form av ersättning för offentliga tjänster som beviljas vissa företag som fått i uppdrag att tillhandahålla tjänster av allmänt ekonomiskt intresse
– med beaktande av gemenskapens rambestämmelser för statligt stöd i form av ersättning för offentliga tjänster
EUT C 297, 29.11.2005, s.
4. ,
– med beaktande av kommissionens meddelande av den 19 januari 2001 – Tjänster i allmänhetens intresse i Europa
EGT C 17, 19.1.2001, s.
4. ,
– med beaktande av kommissionens meddelande av den 26 september 1996: Tjänster i allmänhetens intresse i Europa
EGT C 281, 26.9.1996 s.
3. ,
– med beaktande av Regionkommitténs yttrande av den 1 juli 2011: Reform av EU:s regler om statligt stöd avseende tjänster av allmänt ekonomiskt intresse
EUT C 259, 2.9.2011, s.
40. ,
– med beaktande av yttrandet av den 15 juni 2011 från Europeiska ekonomiska och sociala kommittén om ”Meddelande från kommissionen till Europaparlamentet, rådet, Europeiska ekonomiska och sociala kommittén och Regionkommittén – Reform av EU:s regler om statligt stöd avseende tjänster av allmänt ekonomiskt intresse”
EUT C 248, 25.8.2011, s.
149. .
– med beaktande av domstolens dom av den 24 juli 2003, Altmark Trans GmbH och Regierungspräsidium Magdeburg mot Nahverkehrsgesellschaft Altmark GmbH
– med beaktande av sina resolutioner av den 5 juli 2011 om framtiden för sociala tjänster av allmänt intresse
Antagna texter, P7_TA(2011)0319 . , av den 14 mars 2007 om sociala tjänster av allmänt intresse i Europeiska unionen
EUT C 301 E, 13.12.2007, s.
140. , av den 27 september 2006 om kommissionens vitbok om tjänster av allmänt intresse
EUT C 306 E, 15.12.2006, s.
277. , av den 14 januari 2004 om grönboken ”Tjänster i allmänhetens intresse”
EUT C 92 E, 16.4.2004, s.
126. , av den 17 oktober 2001 om kommissionens meddelande ”Tjänster i allmänhetens intresse”
EGT C 140 E, 13.6.2002, s.
27. och av den 7 november 1997 om kommissionens meddelande ”Tjänster i allmänhetens intresse i Europa”
EGT C 371 E, 8.12.1997, s.
4. ,
– med beaktande av artikel 48 i arbetsordningen,
– med beaktande av betänkandet från utskottet för ekonomi och valutafrågor och yttrandena från utskottet för industrifrågor, forskning och energi och utskottet för den inre marknaden och konsumentskydd ( A7‑0371/2011 ), och av följande skäl:
A. Tjänster av allmänt ekonomiskt intresse har en viktig plats bland unionens gemensamma värden och främjar grundläggande rättigheter och den sociala, ekonomiska och territoriella sammanhållningen, och är således avgörande för kampen mot ojämlikhet i samhället och i allt högre grad också för en hållbar utveckling.
B. Tjänster av allmänt ekonomiskt intresse ger ett viktigt bidrag till medlemsstaternas ekonomiska styrka och konkurrenskraft och därmed inte bara till att förebygga och övervinna ekonomiska kriser utan också till att skapa allmänt välstånd.
C. Tillhandahållandet av tjänster av allmänt ekonomiskt intresse främjar ett framgångsrikt genomförande av Europa 2020-strategin, och dessa tjänster kan bidra till att uppnå tillväxtmål inom särskilt sysselsättning, utbildning och social integration, så att man i slutändan kan uppnå de satta målsättningarna för produktivitet, sysselsättning och social sammanhållning.
D. Kostnadseffektiva lösningar genom konkurrerande privata företag ligger i medborgarnas intresse och är avgörande med tanke på budgetsituationen.
E. Tjänster av allmänt ekonomiskt intresse är tjänster som inte alltid skulle kunna erbjudas utan statligt ingripande, i alla fall inte i tillräcklig omfattning.
F. Sociala tjänster av allmänt intresse spelar en viktig roll för att säkerställa grundläggande rättigheter och de bidrar på ett avgörande sätt till lika möjligheter.
G. I den nuvarande EU-lagstiftningen fastställs undantag från anmälningsplikten för sjukhus och offentligt subventionerade bostäder, dvs. tjänster av allmänt ekonomiskt intresse som tillgodoser grundläggande sociala behov.
H. Artiklarna 106 och 107 i EUF-fördraget utgör den rättsliga grunden för reformen av statsstödsregler för tjänster av allmänt ekonomiskt intresse, och artikel 14 i EUF-fördraget gör det möjligt för Europaparlamentet och rådet, genom förordningar i enlighet med det ordinarie lagstiftningsförfarandet, att fastställa de principer och villkor, särskilt ekonomiska och finansiella, på grundval av vilka sådana tjänster utförs, utan att detta påverkar medlemsstaternas befogenheter.
I. I protokoll nr 26 till EUF-fördraget fastställs att tjänster av allmänt ekonomiskt intresse ska utmärkas av en hög nivå på kvalitet, säkerhet och överkomlighet, likabehandling och främjande av allmän tillgång och användarnas rättigheter, samtidigt som deras avgörande roll erkänns uttryckligen.
Europaparlamentet noterar de mål som kommissionen har med förslaget till reform, dvs. att skapa klarhet kring tillämpningen av reglerna om statligt stöd avseende tjänster av allmänt ekonomiskt intresse med beaktande av deras mångfald.
Parlamentet föreslår att kommissionen i detta sammanhang inte begränsar sig till att enbart åberopa EU-domstolens beslut utan att utforma avgörande kriterier för att hjälpa till att förstå och tillämpa de begrepp som används.
Europaparlamentet framhåller de särdrag som kännetecknar tjänster av allmänt ekonomiskt intresse på regional och lokal nivå, vilka inte påverkar konkurrensen på den inre marknaden, och där ett förenklat och transparent förfarande borde vara möjligt för att främja innovation och medverkan från små och medelstora företag.
13.
14.
Europaparlamentet anser att det kommande kommissionsförslaget om EU 2020‑projektobligationer skulle kunna och bör vara en avgörande drivkraft för utvecklingen av tjänster av allmänt ekonomiskt intresse i medlemsstaterna och på EU‑nivå.
Europaparlamentet önskar i detta sammanhang understryka att ett vidareutvecklat samarbete mellan offentliga myndigheter, genom gemensamt resursutnyttjande, innebär en stor potential när det gäller att öka effektiviteten vid användningen av offentliga medel och att modernisera de allmännyttiga tjänsterna i syfte att tillmötesgå medborgarnas nya behov på lokal nivå.
Förenkling/Proportionalitet
Kommissionen uppmanas att i detta sammanhang göra det enklare att förstå reglerna och föreskriva skyldigheterna när det gäller de offentliga ersättningarna för tjänster av allmänt ekonomiskt intresse och därmed uppnå större rättssäkerhet för offentliga myndigheter och tjänsteleverantörer.
Sociala tjänster
Lokala tjänster
Kvalitets- och effektivitetsaspekter
°
° °
MOTIVERING
1.
Betydelsen av tjänster av allmänt ekonomiskt intresse
Tjänster av allmänt ekonomiskt intresse spelar inte bara en avgörande roll för enskilda medborgare utan är också av enorm betydelse för hela samhällets välstånd.
Mångfalden av sådana tjänster är stor, och att avgöra vad som är en allmännyttig tjänst, dvs. vilka tjänster som bör erbjudas i allmänhetens intresse, är inom EU en uppgift för nationella, regionala och lokala myndigheter.
Genom de statliga interventionerna ska det säkerställas att alla medborgare får tillgång till dessa tjänster och att tjänsterna kan erbjudas alla medborgare till ett överkomligt pris och med en hög kvalitet.
De erbjudna tjänsterna ger ett avgörande bidrag till den ekonomiska kapaciteten och konkurrenskraften och främjar den sociala, ekonomiska och territoriella sammanhållningen i EU.
Ett framgångsrikt genomförande av tillväxtstrategin Europa 2020, inte minst på områdena sysselsättning, utbildning och social integration, främjas genom tillhandahållandet av tjänster av allmänt ekonomiskt intresse.
En särskild betydelse har de sociala tjänsterna av allmänt intresse som spelar en viktig roll för att säkerställa grundläggande rättigheter och att avgörande bidra till lika möjligheter.
2.
Reform av regl erna om statligt stöd till tjänster av allmänt ekonomiskt intresse
Enligt artikel 14 i EUF-fördraget fastställs dessutom att unionen och medlemsstaterna, inom ramen för sina respektive befogenheter och inom fördragens tillämpningsområde, ska sörja för att sådana tjänster utförs på grundval av principer och villkor, särskilt ekonomiska och finansiella, som gör det möjligt för dem att fullgöra sina uppgifter.
Vid reformen av EU:s statsstödsregler måste därför båda artiklarna beaktas och det måste säkerställas att reglerna inte skapar hinder för en rimlig ersättning till de företag som anförtrotts att tillhandahålla tjänster av allmänt ekonomiskt intresse.
Den konkreta tillämpningen av reglerna om förbud mot och kontroll av statligt stöd förklarades av kommissionen 2005 i rambestämmelserna och beslutet om tjänster av allmänt ekonomiskt intresse som löper ut i slutet av året och därför måste ses över.
Med rambestämmelserna, beslutet och ”Vägledning[en] om hur Europeiska unionens bestämmelser om statligt stöd […] på tjänster av allmänt ekonomiskt intresse” kunde betydande förbättringar när det gäller tillämpning och begriplighet uppnås.
Det samråd om det nu gällande paketet som kommissionen inledde 2010 har dock visat att de rättsliga instrumenten måste bli ännu klarare samt enklare, effektivare och mer proportionella.
Samråden gav också vid handen att inte bara de administrativa kostnaderna utan också osäkerheter och missförstånd när det gäller centrala begrepp i dessa regler såsom uppdragsbeskrivning, rimlig vinst, företag, ekonomiska och icke-ekonomiska tjänster eller relevans för den inre marknaden, kan ha lett till att reglerna inte tillämpats.
Ett grundläggande problem är att finansieringen och organisationen av offentliga tjänster i EU hänger på enskilda domar och rättsliga tolkningar.
Utan en klar rättslig ram kan osäkerhetsmomenten och missförstånden inte undanröjas.
Eftersom det med artikel 14 i EUF‑fördraget skapades en ny rättslig grund för en ny övergripande rättslig ram som bestämmer de principer och villkor, särskilt ekonomiska och finansiella, för offentliga tjänster, kan den nödvändiga rättssäkerheten och klarheten äntligen skapas på denna grund.
Det är därför av högsta prioritet att kommissionen lägger fram en sådan horisontell rättlig ram före utgången av 2011.
Man bör dock beakta att reformen av EU:s statsstödsregler för tjänster av allmänt ekonomiskt intresse endast utgör en del av denna i högsta grad nödvändiga ram.
Man måste också beakta behovet av en särskild, sektorsspecifik lagstiftning för vissa tjänster.
3.
Centrala faktorer
3.1 Förenkling, klarhet och proportionalitet
De mål som kommissionen har med reformen, dvs. att skapa större klarhet kring reglerna om statligt stöd för tjänster av allmänt ekonomiskt intresse och att vilja säkerställa en diversifierad och proportionerlig behandling som motsvarar mångfalden av de olika typerna av tjänster av allmänt ekonomiskt intresse, välkomnas.
Också strävan att förenkla tillämpningen av statsstödsreglerna så att myndigheternas administrativa kostnader står i rimlig proportion till åtgärdens effekter på konkurrensen på den inre marknaden, skulle kunna leda till ett bättre genomförande av reglerna.
I detta sammanhang bör reglerna om förbudet mot och kontrollen av statligt stöd till de företag som fått i uppdrag att tillhandahålla offentliga tjänster utformas i enlighet med de administrativa instansernas kapacitet så att en korrekt tillämpning av reglerna kan säkerställas och i synnerhet så att de företag som fått i uppdrag att tillhandahålla offentliga tjänster kan uppfylla de uppgifter de anförtrotts.
Tröskelvärdena för befrielse från anmälningsplikten för ersättning för tjänster av allmänt ekonomiskt intresse är ett sätt att minska den administrativa bördan.
En allmän höjning av de nu gällande tröskelvärdena som bestäms genom tillämpningen av beslutet om tjänster av allmänt ekonomiskt intresse bör därför beaktas för att ytterligare minska den administrativa bördan.
En ytterligare förenkling skulle kunna bestå i att införa en de minimis-regel för statsstöd till företag som fått i uppdrag att tillhandahålla tjänster av allmänt ekonomiskt intresse och som på grund av sitt lokalt begränsat verksamhetsområde förmodligen endast får försumbara effekter på handeln mellan medlemsstaterna.
Här måste det säkerställas att ersättningen endast används till den aktuella tjänsten av allmänt ekonomiskt intresse.
En metod baserad på kombinerade index för storleken på kommunen, beloppet för ersättningen och omsättningen för det företag som fått i uppdrag att tillhandahålla tjänster av allmänt ekonomiskt intresse skulle kunna vara ett lämpligt alternativ.
3.2 Sociala tjänster
För sociala tjänster av allmänt ekonomiskt intresse som till sin natur är lokalt begränsade bör man överväga särskilda förhöjda tröskelvärden för storleken på ersättningen när man kan anta att det inte kan bli fråga om några följder för handeln mellan medlemsstaterna så länge tröskelvärdena inte överskrids.
Att utvidga det allmänna undantaget från anmälningsplikten till andra typer av sociala tjänster av allmänt ekonomiskt intresse, såsom äldrevård och handikappomsorg eller hälsovård, bör övervägas.
Offentliga tjänster måste vara av hög kvalitet och tillgängliga för alla befolkningsgrupper.
De särskilda uppgifterna för och arten på sociala tjänster av allmänt intresse bör inte bara skyddas utan klart definieras inom ramen för sektorsspecifika regler.
Det är oroande att vissa medlemsstater är så pass återhållsamma med att klassificera statsstöd till allmännyttiga bostadsföretag som sociala tjänster av allmänt ekonomiskt intresse att de gör det först när tjänsterna uteslutande är avsedda för missgynnade och socialt svaga grupper.
En sådan restriktiv tolkning går stick i stäv med det övergripande målet om social mångfald.
För att de sociala tjänsterna av allmänt ekonomiskt intresse ska kunna fylla sin särskilda funktion, måste de vara tillgängliga för alla medborgare, oavsett inkomst och förmögenhet.
3.3 Det stora handlingsutrymmet för nationella, regionala och lokala myndigheter
Tjänster av allmänt ekonomiskt intresse måste vara av hög kvalitet och den allmänna tillgången måste främjas.
Det primära ansvaret för att skapa förutsättningar för att beställa, tillhandahålla, finansiera och organisera tjänster av allmänt ekonomiskt intresse ligger hos medlemsstaterna och är förankrat i protokoll nr 26 till Lissabonfördraget.
Det stora handlingsutrymme som nationella, regionala och lokala myndigheter i EU har för tjänster av allmänt ekonomiskt intresse poängteras därmed särskilt i fördragen.
Reformen av EU:s statsstödsregler kan därför endast ske under strikt beaktande av subsidiaritetsprincipen.
I enlighet med konkurrensreglerna i EUF-fördraget är också kommissionens befogenhet begränsad till att enbart kontrollera statsstödet till tillhandahållandet av tjänster av allmänt ekonomiskt intresse, och fastställandet av kvalitets- och effektivitetskriterier kan på europeisk nivå endast ske på grundval av artikel 14 i EUF-fördraget med beaktande av subsidiaritetsprincipen.
YTTRANDE från utskottet för industrifrågor, forskning och energi
till utskottet för ekonomi och valutafrågor
över reformen av EU:s regler om statligt stöd avseende tjänster av allmänt ekonomiskt intresse
( 2011/2146(INI) )
Föredragande:
Gunnar Hökmark
FÖRSLAG
Utskottet för industrifrågor, forskning och energi uppmanar utskottet för ekonomi och valutafrågor att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet anser att statligt stöd ska bidra till att stimulera lokal företagaranda och den lokala ekonomin, skapa lokala arbetstillfällen och främja konkurrensen på bland annat telekommunikationsmarknaden.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
26.9.2011
Slutomröstning: resultat
+:
–:
0:
33
6
Slutomröstning: närvarande ledamöter
Slutomröstning: närvarande suppleanter
YTTRANDE från utskottet för den inre marknaden och konsumentskydd
till utskottet för ekonomi och valutafrågor
över reformen av EU:s regler om statligt stöd avseende tjänster av allmänt ekonomiskt intresse
( 2011/2146(INI) )
Föredragande: António Fernando Correia De Campos
FÖRSLAG
Europaparlamentet välkomnar kommissionens meddelande om reformen av EU-reglerna för statligt stöd avseende tjänster av allmänt ekonomiskt intresse.
2.
Europaparlamentet välkomnar kommissionens avsikt att avge ytterligare förklaringar och fastställa ytterligare kriterier när det gäller skillnaden mellan icke-ekonomiska och ekonomiska verksamheter för att undvika klagomål till EU‑domstolen och överträdelseförfaranden från kommissionens sida.
Europaparlamentet framhåller de särdrag som kännetecknar tjänster av allmänt ekonomiskt intresse på regional och lokal nivå, vilka inte påverkar konkurrensen på den inre marknaden, och menar att ett förenklat och öppet förfarande borde vara möjligt för att främja innovation och medverkan från små och medelstora företag.
Europaparlamentet erinrar om att reglerna för statligt stöd strikt bör följa subsidiaritetsprincipen och garantera de lokala och regionala myndigheternas frihet att själva avgöra hur de vill organisera, finansiera och utföra uppdraget att tillhandahålla offentliga tjänster.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
26.9.2011
Slutomröstning: resultat
+:
–:
0:
27
8
Slutomröstning: närvarande ledamöter
Pablo Arias Echeverría, Adam Bielan, Lara Comi, Anna Maria Corazza Bildt, António Fernando Correia De Campos, Jürgen Creutzmann, Cornelis de Jong, Evelyne Gebhardt, Małgorzata Handzlik, Malcolm Harbour, Philippe Juvin, Sandra Kalniete, Edvard Kožušník, Toine Manders, Phil Prendergast, Mitro Repo, Heide Rühle, Matteo Salvini, Christel Schaldemose, Andreas Schwab, Emilie Turunen, Bernadette Vergnaud, Barbara Weiler
Slutomröstning: närvarande suppleanter
Pascal Canfin, Frank Engel, Marielle Gallo, Anna Hedh, María Irigoyen Pérez, Othmar Karas, Constance Le Grip, Antonyia Parvanova, Sylvana Rapti, Olle Schmidt, Kyriacos Triantaphyllides, Anja Weisgerber
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
17.10.2011
Slutomröstning: resultat
+:
–:
0:
27
8
1
Slutomröstning: närvarande ledamöter
Burkhard Balz, Udo Bullmann, Pascal Canfin, Nikolaos Chountis, George Sabin Cutaş, Leonardo Domenici, Derk Jan Eppink, Diogo Feio, Ildikó Gáll-Pelcz, Jean-Paul Gauzès, Sven Giegold, Sylvie Goulard, Liem Hoang Ngoc, Gunnar Hökmark, Wolf Klinz, Jürgen Klute, Philippe Lamberts, Werner Langen, Astrid Lulling, Arlene McCarthy, Alfredo Pallone, Anni Podimata, Antolín Sánchez Presedo, Peter Simon, Peter Skinner, Ivo Strejček, Kay Swinburne, Marianne Thyssen
Slutomröstning: närvarande suppleanter
Sophie Auconie, Philippe De Backer, Saïd El Khadraoui, Ashley Fox, Olle Ludvigsson, Thomas Mann, Andreas Schwab, Theodoros Skylakakis
Slutomröstning: närvarande suppleanter (art.
187.2)
Diana Wallis
A7-0385/2011
Föredragande: Santiago Fisas Ayxela
PE 466.981v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
MOTIVERING..........................................................................................................................21
YTTRANDE från utskottet för ekonomi och valutafrågor ....................26
YTTRANDE från utskottet för miljö, folkhälsa och livsmedelssäkerhet 31
YTTRANDE från utskottet för den inre marknaden och konsumentskydd 35
YTTRANDE från utskottet för rättsliga frågor ...........................................40
YTTRANDE från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor 43
YTTRANDE från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män 47
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................52
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om idrottens europeiska dimension
( 2011/2087(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens meddelande av den 18 januari 2011 ”Utveckling av idrottens europeiska dimension” ( KOM(2011)0012 ),
– med beaktande av kommissionens vitbok om idrott ( KOM(2007)0391 ),
– med beaktande av kommissionens meddelande ”Insatser mot korruption på EU:s territorium” ( KOM(2011)0308 ),
– med beaktande av Europarådets två konventioner, konventionen om läktarvåld och olämpligt uppträdande vid idrottsevenemang av den 19 augusti 1985, och konventionen mot dopning av den 19 augusti 1990,
– med beaktande av sin resolution av den 5 juni 2003 om kvinnor och idrott
EUT
– med beaktande av sin resolution av den 21 april 2004 om respekt för centrala arbetsnormer i produktionen av sportartiklar för de olympiska spelen
EUT C 104 E, 30.4.2004, s.
757. ,
– med beaktande av sin resolution av den 14 april 2005 om dopning inom idrotten
EUT C 33 E, 9.2.2006, s.
590. ,
– med beaktande av sin förklaring av den 14 mars 2006 om bekämpning av rasism inom fotbollen
EUT C 291 E, 30.11.2006, s.
143. ,
– med beaktande av sin resolution av den 15 mars 2006 om tvångsprostitution i samband med internationella idrottsevenemang
EUT
C 291 E, 30.11.2006, s 292. ,
– med beaktande av sin resolution av den 29 mars 2007 om framtiden för professionell fotboll i Europa
EUT C 27 E, 31.1.2008, s.
232. ,
– med beaktande av sin resolution av den 13 november 2007 om idrottens roll i utbildningen
EUT C 282 E, 6.11.2008, s.
131. ,
– med beaktande av sin resolution av den 8 maj 2008 om vitboken om idrott
EUT C 271 E, 12.11.2009, s.
51. ,
– med beaktande av sin resolution av den 19 februari 2009 om den sociala ekonomin
EUT C 76 E, 25.3.2010, s.
16. ,
– med beaktande av sin resolution av den 10 mars 2009 om integriteten för hasardspel online
EUT C 87 E, 1.4.2010, s.
30. ,
– med beaktande av sin resolution av den 5 juli 2011 om kommissionens femte sammanhållningsrapport och strategin för sammanhållningspolitiken efter 2013
P7_TA(2011)0316 . ,
– med beaktande av sin skriftliga förklaring 62/2010 av den 16 december 2010 om ökat EU-stöd till idrott på gräsrotsnivå,
– med beaktande av rådets beslut 2010/37/EG av den 27 november 2009 i anslutning till Europeiska frivilligåret för främjandet av aktivt medborgarskap (2011),
– med beaktande av rådets slutsatser av den 18 november 2010 om idrottens roll som upphov till och pådrivande faktor för aktiv social integration
EUT C 326, 3.12.2010, s.
5. ,
– med beaktande av rådets slutsatser av den 17 juni 2010 om den nya strategin för sysselsättning och tillväxt,
– med beaktande av rådets resolution av den 1 juni 2011 om en EU-arbetsplan för idrott för 2011–2014
EUT C 162, 1.6.2011, s.
1. ,
– med beaktande av Punta del Este-deklarationen från december 1999 och Unescos rundabordsmöte om traditionella idrotter och spel (TSG – traditional sports and games)
Almaty, Kazakstan, 5–6 november 2006. , som handlar om erkännande av traditionella idrotter och spel som en del av ett immateriellt kulturarv och en symbol för kulturell mångfald,
– med beaktande av EU-domstolens och tribunalens rättspraxis, liksom även beslut från kommissionen i idrottsfrågor,
– med beaktande av stadgan för insatser för att undanröja diskriminering av hbt-personer inom idrotten,
– med beaktande av artiklarna 6, 19 och 165 i fördraget om Europeiska unionens funktionssätt,
– med beaktande av artikel 48 i arbetsordningen,
– med beaktande av Regionkommitténs yttrande
CdR 66/2011 slutlig. av den 11–12 oktober 2011 och yttrandet från Europeiska ekonomiska och sociala kommittén av den 26–27 oktober 2011 ”Utveckling av idrottens europeiska dimension”
CESE 1594/2011 – SOC/413. ,
– med beaktande av betänkandet från utskottet för kultur och utbildning och yttrandena från utskottet för ekonomi och valutafrågor, utskottet för miljö, folkhälsa och livsmedelssäkerhet, utskottet för den inre marknaden och konsumentskydd, utskottet för rättsliga frågor, utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor och utskottet för kvinnors rättigheter och jämställdhet ( A7‑0385/2010 ), och av följande skäl:
B. Idrottens särdrag bör ges företräde i Europeiska domstolens domar om idrottsfrågor samt i kommissionens beslut om dessa.
C. Alla intressenter, också de politiskt ansvariga, måste ta hänsyn till idrottens särdrag samt till dess strukturer baserade på frivilligarbete och dess sociala och fostrande funktioner.
E. EU bör i sina åtgärder på idrottens område alltid ta hänsyn till idrottens särdrag och respektera dess sociala, fostrande och kulturella aspekter.
I. EU:s idrottspolitik måste utvecklas så den inriktar sig på och stöder både den professionella idrottens och amatöridrottens syften och mål.
J. EU bör ha som prioritet att stödja och främja idrott för personer med intellektuella eller fysiska funktionshinder, eftersom idrotten är så viktig för social integration, folkhälsa och gränsöverskridande frivilligarbete.
K. Frivilligarbetet är hörnstenen för största delen av amatöridrotten i Europa.
L. 35 miljoner frivilligarbetare gör det möjligt att utveckla idrott för alla och sprida idrottens ideal, vilket även idrottsklubbar och idrottsföreningar utan vinstsyfte gör.
N. Främjande av fysisk aktivitet och idrott bidrar till omfattande besparingar inom den offentliga hälso- och sjukvården.
O. Idrottens bidrag till bättre hälsa och välbefinnande är en avgörande faktor för att motivera medborgarna att delta i idrott och fysisk aktivitet.
P. Dopning står i strid med idrottens värderingar och utsätter idrottsmänniskor för allvarliga faror samt medför allvarliga och bestående skador för hälsan.
Q. Elitidrott förhöjer vissa av idrottens mest grundläggande värden, sprider dem i samhället och främjar där ett aktivt idrottsutövande.
R. Många toppidrottare befinner sig i en osäker situation efter att de avslutat sin idrottskarriär.
S. Det är av grundläggande betydelse att sådana idrottare förbereds på livet efter idrottskarriären genom att erbjudas allmän eller yrkesinriktad utbildning parallellt med idrottsutbildningen.
T. Idrottarnas grundläggande rättigheter måste garanteras och skyddas.
U. Verbalt och fysiskt våld samt diskriminerande beteenden riskerar att utvecklas i samband med idrottstävlingar.
V. Idrott för kvinnor är inte är tillräckligt värderat och att kvinnor är underrepresenterade i idrottsorganisationernas beslutsorgan.
Y. Intrång i idrottsorganisationernas immateriella rättigheter och framväxten av digital piratkopiering, särskilt genom otillåtna direktsändningar från idrottsevenemang, är ett hot mot ekonomin i hela idrottssektorn.
Z. Idrotten fungerar inte som en typisk näringsgren på grund av motståndarnas ömsesidiga beroende av varandra och på grund av den tävlingsbalans som måste finnas för att resultaten även i fortsättningen ska vara ovissa.
Idrotten är viktig och utgör en källa till glädje för många medborgare, oavsett om de är deltagare, supportrar eller åskådare.
Ökad insyn och demokratisk redovisningsskyldighet kan åstadkommas i idrottsklubbarna genom att supportrarna får vara med i sina klubbars ägande- och styrelsestrukturer.
Finansieringen av gräsrotsidrotten kan endast tryggas om innehavarna av de nödvändiga nationella spellicenserna, som betalar skatter och avgifter och finansierar andra aktiviteter av allmänt intresse i medlemsstaterna, i lag åläggas att betala till allmännyttiga ändamål och effektivt skyddas från olaglig konkurrens.
Idrotten kan spela en roll inom olika områden för unionens externa förbindelser, bland annat som ett diplomatiskt verktyg.
Europaparlamentet uppmanar med kraft kommissionen att inom den kommande fleråriga budgetramen föreslå en särskild och ambitiös budget för idrottspolitiken, mot bakgrund av vilken nytta idrotten för med sig för folkhälsan samt ur social, kulturell och ekonomisk synvinkel.
Europaparlamentet uppmanar med kraft medlemsstaterna att fastställa klara riktlinjer för hur idrott och fysisk aktivitet ska tas med på alla utbildningsstadier runtom i medlemsstaterna.
Europaparlamentet rekommenderar kommissionen att uppmuntra idrottsutövande bland äldre, eftersom detta är ett bra sätt att umgås och behålla en god hälsa.
Europaparlamentet understryker att idrotten måste göras tillgänglig för alla medborgare i många olika sammanhang: i skolan, på arbetsplatsen, såsom fritidsverksamhet eller genom klubbar och föreningar.
Europaparlamentet framhåller idrottens enorma samhällsintegrerande kraft på många områden, på områden såsom medborgarengagemang och demokratiförståelse, hälsofrämjande åtgärder, stadsutveckling, social integration, arbetsmarknad, sysselsättning, kompetensutveckling och utbildning.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att stödja och uppmuntra europeisk forskning om damidrottens särart, om orsakerna till att kvinnor och flickor slutar idrotta och om den fortsatta ojämlikheten i fråga om kvinnors tillgång till idrott.
Europaparlamentet anser att EU:s anslutning till Europarådets antidopningkonvention är ett nödvändigt steg på väg mot en samordning av ett mera enhetligt genomförande av Världsantidopningskoden i medlemsstaterna.
Europaparlamentet ställer sig positivt till att medlemsstaterna i samverkan med europeiska idrottsförbund tar fram minimistandarder för säkerheten på idrottsarenor och vidtar alla lämpliga åtgärder för att garantera största möjliga säkerhet för idrottare och åskådare.
Idrottens ekonomiska dimension
Europaparlamentet uppmanar kommissionen och medlemsstaterna att inrätta ett system för erkännande av kvalifikationer som förvärvats av frivilliga och av kvalifikationer som krävs för utövandet av reglerade yrken med anknytning till idrotten.
Europaparlamentet uppmanar medlemsstaterna att se till att idrottare kan få högre utbildning samt tillförsäkra ett harmoniskt erkännande av deras kvalifikationer inom idrott och utbildning för att förbättra den yrkesmässiga rörligheten.
47.
Europaparlamentet understryker att det är viktigt att det kommersiella utnyttjandet av audiovisuella rättigheter till idrottsarrangemang sker på ett centraliserat sätt, med exklusiva rättigheter och enligt territoriella principer, för att garantera att inkomster fördelas rättvist mellan elitidrott och breddidrott.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att skydda de immateriella rättigheterna till idrottsligt innehåll och att samtidigt respektera allmänhetens rätt till information.
Europaparlamentet upprepar sin begäran till kommissionen att fastställa riktlinjer för statligt stöd genom att precisera vilken typ av offentligt stöd som är berättigat för att idrotten ska kunna fylla sin sociala, kulturella och fostrande funktion.
59.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att på ett konkret sätt främja utbyte av bästa praxis och ett tätt samarbete inom teknik och forskning på idrottsområdet.
Organisationen av idrott
64.
Europaparlamentet uppmanar idrottens styrande organ att förbättra insynen i spelaragenternas verksamhet och att samarbeta med medlemsstaternas myndigheter för att få bort korruptionen.
Europaparlamentet uttrycker sin åsikt om att system som införts av idrottens styrande organ för att öka insynen i samband med internationella spelarövergångar är ett steg i rätt riktning eftersom de tjänar principen om god ledning och syftar till att garantera idrottstävlingarnas integritet.
Europaparlamentet uppmanar kommissionen att genom att till fullo beakta artikel 165 i EUF-fördraget senast 2012 lägga fram ett förslag i syfte att skapa bättre förståelse för idrottens särskilda behov och vidta konkreta åtgärder för att tillmötesgå dessa.
Samarbetet med tredjeländer och internationella organisationer
En europeisk identitet genom idrott
- att årligen organisera en ”Europeisk idrottsdag” till förmån för såväl amatöridrottens och den professionella idrottens sociala och kulturella roll som för nyttan med idrott ur folkhälsosynvinkel,
- att stödja en årlig utnämning av en ”europeisk idrottshuvudstad” under ledning av ACES (Association des capitales européennes du sport – Organisationen av europeiska idrottshuvudstäder), med finansiellt stöd och nödvändiga kontroller,
- att stödja lokala, traditionella, ursprungliga idrotter, vilka ingår i EU:s rika kulturella och historiska mångfald och symboliserar dess valspråk ”Förenade i mångfalden”, genom att öka medvetenheten om dessa idrotter, bland annat genom en europeisk idrottskarta och europeiska festivaler,
- att upprätta ett utbytesprogram och relevanta åtgärder för unga amatöridrottare och tränare så att de kan lära sig nya träningsmetoder, ta fram bästa metoder och med idrottens hjälp utveckla europeiska värden såsom rent spel, respekt och social integration samt främja interkulturell dialog,
- att bidra till att inrätta ett utbytesprogram för idrottstränare,
- att samarbeta med medlemsstaterna och idrottsorganisationerna för att slå vakt om den grundläggande integriteten för idrott på gräsrotsnivå,
- att stödja medlemsstaternas arbete med uppgiftsinsamling och forskning för att utbyta exempel på bästa praxis.
o
o o
MOTIVERING
Artikel 165 i fördraget om Europeiska unionens funktionssätt (EUF-fördraget) ger EU en ny behörighet för idrott, manar EU att bidra till att främja idrottsfrågor och anger att EU-åtgärder bör inriktas mot att utveckla idrottens europeiska dimension.
Meddelandet från kommissionen är det första policydokument som har utfärdats på idrottsområdet efter att Lissabonfördraget har trätt i kraft, vilket ger EU ett mandat att stödja, samordna, och komplettera policyåtgärder som vidtas av medlemsstaterna på idrottsområdet.
Under förra perioden utarbetade Europaparlamentet, som en återspegling av vikten av detta, andra resolutionsförslag, nämligen om framtiden för professionell fotboll i Europa
Antagna texter, P6_TA(2007) 0100. , om idrottens roll i utbildningen”
Antagna texter, P6_TA(2007) 0503. och om vitboken om idrott
Antagna texter, P6_TA(2008) 0198. (genomförd av kommissionen under 2007).
– Varför idrott är viktigt för samhället
Idrott utgör i sig ett viktigt socialt fenomen och en allmännytta.
För många är det den viktigaste formen av rekreation, oavsett om de deltar själva, eller om de är åskådare.
När den är som bäst för idrotten människor samman, oavsett deras härkomst, bakgrund, religiösa trosåskådning eller ekonomiska status.
Idrott främjar europeiska medborgares aktiva bidrag till samhället och hjälper till att bygga upp en känsla av social integration.
– Förbättra hälsan genom idrott
Fysisk aktivitet är en av de viktigaste faktorerna som avgör människans hälsotillstånd i det moderna samhället.
Brist på fysisk aktivitet har en negativ effekt på europeiska medborgares hälsa, eftersom det ökar risken för att utveckla fetma, bli överviktig och ådra sig olika sjukdomar.
Dessa negativa följder är en börda för medlemsstaternas hälsovårdsbudget och allmänna ekonomi.
– Dopning, våld och intolerans
Dopning kvarstår som ett viktigt hot mot idrott.
Många aktörer efterlyser en mer aktiv strategi från EU i kampen mot dopning genom att unionen ansluter sig till Europarådets konvention mot dopning, i den mån unionens behörighet inom detta område berättigar till detta.
Åskådarvåld och oroligheter kvarstår även som ett alleuropeiskt fenomen och det finns ett behov av en europeisk strategi med åtgärder för att minska de medföljande riskerna.
– Idrotten och ekonomin
Idrott utgör en stor och snabbt växande del av ekonomin och är ett viktigt bidrag till tillväxt och arbeten, med mervärden och anställningseffekter som överstiger genomsnittliga tillväxtsiffror.
Hållbar finansiering av idrott är dock en fråga som behöver studeras närmare.
– Organisering av idrott
God ledning inom idrott är ett villkor för att möta utmaningar med idrottens och EU:s rättsliga ramverk.
Sådana utmaningar inkluderar: medborgarnas fria rörlighet och idrottarnas nationalitet, spelarövergångar (problem avseende handlingarnas legalitet och transparens i finansflöden), idrottstävlingars integritet och en europeisk dialog inom idrottssektorn.
Kommissionens meddelande:
Den 18 januari 2011 antog Europeiska kommissionen meddelandet ”Utveckling av idrottens europeiska dimension”.
Det fastslår kommissionens idéer om insatser på EU-nivå inom idrotten.
Det föreslår konkreta åtgärder för kommissionen och/eller medlemsstaterna inom tre breda kapitel: idrottens sociala roll, idrottens ekonomiska dimension och organisationen av idrott.
Meddelandets huvudbudskap:
– Nyckelutmaningar med avseende på idrott (t.ex. dopning av amatöridrottare och våld med anknytning till idrott) identifieras.
– Autonomin hos strukturer som styr idrott respekteras och behörigheterna för medlemsstaterna inom organisationen av idrott erkänns.
– Det hävdas emellertid att åtgärder på EU-nivå vad gäller organisering av idrott kan tillhandahålla betydande mervärde.
– Varje kapitel avslutas med en lista över möjliga uppföljningsåtgärder som kommissionen och medlemsstaterna kan vidta.
– Förslagens komplexitet på idrottsområdet erkänns.
– Ett fortsatt informellt samarbete mellan medlemsstater föreslås för att säkerställa fortsatt utbyte av bästa praxis och vidarespridning av resultat.
I meddelandet fastställs att EU-åtgärder bidrar till de allmänna målen i Europa 2020-strategin genom att förbättra anställningsbarhet och rörlighet genom åtgärder som främjar social integration i, och genom, idrott, utbildning och träning och europeiska riktlinjer för fysisk aktivitet.
Syftet med de åtgärder som föreslås i meddelandet är att uppmuntra till debatt mellan intressenter, bemöta utmaningar inom idrotten och hjälpa sektorn att utvecklas.
Idrottsutövare, idrottsorganisationer och EU-medborgare förväntas dra nytta av planerna som utmynnar ur EU:s nya roll vilken i enlighet med Lissabonfördraget ska vara att stödja och koordinera idrottspolicy i medlemsstaterna.
För närvarande tillhandahåller kommissionen stöd till projekt och nätverk på idrottsområdet, antingen genom idrottsspecifika stimulansåtgärder, i synnerhet de förberedande åtgärderna på idrottsområdet, eller genom existerande program på olika relevanta områden.
Dessa inkluderar livslångt lärande, folkhälsa, ungdom, medborgarskap, forskning och teknologisk utveckling, social integration, kampen mot rasism, miljöskydd och andra områden.
Föredragandens kommentarer och framtida utmaningar:
Angående idrottens värde:
– Föredraganden tror starkt på att idrott, med dess utbildningsmässiga och kulturella värde, kan bidra till Europeiska unionens strategiska mål.
– Idrott bidrar till integration, eftersom den är öppen för alla medborgare, oavsett kön, etnicitet, religion, ålder, nationalitet och social status.
– Föredraganden är medveten om att idrott bland kvinnor inte är tillräckligt värderat och att kvinnor är underrepresenterade i idrottsorganisationernas beslutsfattande organ.
– Föredraganden uppmuntrar medlemsstaterna att beakta äldre idrottares erfarenhet när de söker tillträde till tränaryrket och att etablera speciella vägar för idrottsutövare som önskar bedriva högre utbildning, samt att se till att det finns handledare som följer upp dem.
– Frivilligarbetare möjliggör att många idrottsevenemang kan förflyta smidigt.
Föredraganden skulle vilja understryka vikten av deras bidrag.
Om att bemöta de stora frågorna:
– Föredraganden är av åsikten att det bör vara medlemsstaternas ansvar att främja hälsofördelarna med idrott.
På EU-nivå bör fokus ligga på större frågor som dopning, människohandel, idrottsutövares rörlighet, rasism, och våld inom idrott.
– Det bör göras varje möjlig ansträngning för att förebygga kriminella handlingar som utgör ett hot mot idrott, t.ex. penningtvätt, uppgjorda matcher, människohandel och utnyttjande av minderåriga.
– Föredraganden uppmanar medlemsstaterna att förbjuda tillträde till idrottsstadion för supportrar som har uppvisat våldsamt eller diskriminerande beteende.
Föredraganden föreslår ett europeiskt register för personer som har förbjudits tillträde till idrottsevenemang.
Om god ledning:
– Standarder för idrottsledning genom utbyte av bästa praxis bör främjas.
– Medlemsstaternas lagstiftning om försäljning av medierättigheter bör harmoniseras för att förhindra en situation där endast stora organisationer drar nytta av försäljningen.
– Föredraganden vidkänner vikten av rättvis fördelning av inkomst mellan idrottsklubbar av olika storlekar och mellan professionella idrotter och amatöridrotter.
– Även vikten av utbildningsbidrag betonas, eftersom de är en effektiv skyddsmekanism för utbildningscentrum och för en rimlig avkastning på investering.
Om rättvisa idrottstävlingar:
– Idrottsevenemangens integritet är viktig.
Medlemsstater bör anta regleringsåtgärder för att säkerställa att idrott skyddas mot olämpliga influenser som vadslagning eller uppgjorda matcher.
– Föredraganden uppmanar medlemsstaterna att göra det brottsligt att attackera tävlingars integritet.
– Idrottstävlingars rättvisa och öppenhet är avgörande för att skydda idrottsmäns och idrottskvinnors integritet.
– Idrottsförbund har inte de strukturella och rättsliga medlen för att agera effektivt mot uppgjorda tävlingar.
– Föredraganden stöder licensieringssystemen och finansiell fair play.
– Föredraganden erkänner idrottsdomstolars legitima rätt att lösa tvister på idrottsområdet och efterfrågar därför bildandet av en europeisk kammare vid Idrottens skiljedomstol (CAS).
Angående budgeten:
– Det behövs lämplig budgettäckning för idrott för att den förberedande åtgärden ska övergå i ett specifikt program som tillägnas den nya behörigheten.
Angående möjligheter och arbetstillfällen:
– Medlemsstaternas utbildningsprogram bör vara koordinerade på ett sätt som tillåter unga idrottsutövare att kombinera utbildning med idrottsträning.
– Det bör finnas kurser för unga människor som vill göra en idrottskarriär och kombinera den med studier.
– Idrott bör främjas i skolor med tanke på dess fördelar med att bryta ned sociala barriärer och integrera marginaliserade grupper.
– Idrott har potentialen att bidra till jobbskapande och en smart, hållbar och integrerande tillväxt.
Angående turism:
– Synergier mellan idrott och turism behöver identifieras, i synnerhet genom uppgradering av kollektiva infrastrukturer.
– Föredraganden noterar att stora evenemang och idrott erbjuder utmärkta möjligheter för att utnyttja utvecklingen av turismpotentialen i Europa.
Angående traditionella idrotter och spel:
– Föredraganden anser starkt att vi bör bevara lokala, traditionella idrotter, eftersom dessa utgör en del av vårt kulturarv och förstärker känslan av europeiskt medborgarskap.
Detta är en sann symbol för den kulturella mångfalden i våra samhällen.
– Föredraganden noterar att en del traditionella spel och idrotter redan har försvunnit och att de som har överlevt löper en förestående risk att försvinna.
– Föredraganden uppmanar kommissionen att utarbeta en stadga för inhemska idrotter och att stödja dess spridning.
Europeisk identitet genom idrott:
– Föredraganden uppmanar kommissionen att organisera en årligt förekommande ”Europeisk idrottsdag” för att höja den allmänna medvetenheten om idrottens fördelar.
– Möjliga initiativ inkluderar konferenser och debatter om idrott, rabatt på idrottsartiklar i butiker och främjandet av en hälsosam livsstil.
– Föredraganden uppmuntrar kommissionen att stödja den årliga utnämningen av en ”Europeisk idrottshuvudstad” under ledning av ACES, med finansiellt stöd och nödvändiga kontroller.
– Föredraganden föreslår att den europeiska flaggan ska vaja vid stora idrottsevenemang i Europa och föreslår att den ska framträda på sporttröjor tillhörande medlemsstaternas idrottsutövare.
Träning och rörlighet inom idrott:
– Betonar att träning av spelare på lokal nivå behövs för en hållbar utveckling av idrott i Europa.
– Föredraganden föreslår att ett utbytesprogram för unga idrottare ska skapas för att ge idrottare möjlighet att träna med utländska lag.
– Studenter och skolelever bör vara berättigade att delta i dessa utbyten.
Studenterna skulle ha möjlighet att lära sig nya träningsmetoder och utveckla sin europeiska medvetenhet.
Programmet skulle förstärka interkulturell dialog.
Om samarbetet med tredjeländer och internationella organisationer:
– Föredraganden uppmanar kommissionen och medlemsstaterna att i samband med samarbetet med tredjeländer ta upp problem såsom internationell överföring av spelare, utnyttjande av minderåriga spelare, piratkopieringsverksamhet och illegal vadslagning.
– Idrottsklubbarna bör vara tvungna att efterleva migrationslagstiftning vad gäller rekrytering av ungdomar från tredjeländer.
Detta kommer att säkerställa att idrottsutövarna behandlas väl tills det att de återvänder till sina ursprungsländer.
Om idrottsagenter:
YTTRANDE från utskottet för ekonomi och valutafrågor
till utskottet för kultur och utbildning
över idrottens europeiska dimension
( 2011/2087(INI) )
Föredragande: Burkhard Balz
FÖRSLAG
Utskottet för ekonomi och valutafrågor uppmanar utskottet för kultur och utbildning att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
– med beaktande av sin resolution av den 19 februari 2009 om den sociala ekonomin ( 2008/2250(INI) ),
– med beaktande av att idrott är ett socialt och kulturellt fenomen, men att den också kan ses som en ekonomisk dynamisk sektor och generera betydande indirekta intäkter och bidra till Europa 2020-strategin,
– med beaktande av att idrott inte är som annan ekonomisk verksamhet, utan en unik företeelse som organisationsmässigt är uppbyggt kring förbund, som inte fungerar som affärsdrivande företag, och att skillnad måste göras mellan de idrottsliga aspekterna och de kommersiella intressena,
Europaparlamentet välkomnar artikel 165 i EUF-fördraget, som för första gången ger EU en rättslig bas för åtgärder på idrottsområdet och således för ekonomiska stödprogram på EU‑nivå.
Europaparlamentet betonar att det ömsesidiga erkännandet av kurser och specialistutbildningar inom en gemensam europeisk ram för personer som har specialyrken inom idrotten (domare, tränare) är särskilt viktigt eftersom det bidrar till att öka konkurrenskraften på lång sikt, vilket i sin tur innebär att intäktsförluster kan undvikas.
Europaparlamentet uppmanar kommissionen att lägga fram konkreta förslag för att åtgärda de brister och skillnader som finns i bestämmelserna för den till sin natur gränsöverskridande verksamhet som bedrivs av idrottsagenter, och som synliggjordes i den oberoende studie som 2009 gjordes på uppdrag av kommissionen.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
22.9.2011
Slutomröstning: resultat
+:
–:
0:
29
Slutomröstning: närvarande ledamöter
Udo Bullmann, Pascal Canfin, George Sabin Cutaş, Rachida Dati, Derk Jan Eppink, Diogo Feio, Elisa Ferreira, Ildikó Gáll-Pelcz, Jean-Paul Gauzès, Sven Giegold, Sylvie Goulard, Liem Hoang Ngoc, Othmar Karas, Wolf Klinz, Philippe Lamberts, Astrid Lulling, Hans-Peter Martin, Ivari Padar, Olle Schmidt, Marianne Thyssen
Slutomröstning: närvarande suppleanter
Pervenche Berès, David Casa, Herbert Dorfmann, Saïd El Khadraoui, Sari Essayah, Mojca Kleva, Thomas Mann, Gianni Pittella, Andreas Schwab
14.9.2011
över idrottens europeiska dimension
( 2011/2087(INI) )
Föredragande: Sophie Auconie
FÖRSLAG
Utskottet för miljö, folkhälsa och livsmedelssäkerhet uppmanar utskottet för kultur och utbildning att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
– med beaktande av att enligt artikel 165 i Lissabonfördraget (FEUF) ska EU:s insatser syfta till att utveckla idrottens europeiska dimension genom att främja rättvisa och öppenhet i idrottstävlingar och samarbete mellan organisationer och myndigheter med ansvar för idrott samt genom att skydda idrottsutövarnas fysiska och moraliska integritet, särskilt när det gäller de yngsta utövarna.
Europaparlamentet uppmanar medlemsstaterna och de lokala myndigheterna att inte bara använda sig av privata idrottsanläggningar, eftersom detta kan leda till bristande jämlikhet, utan också öppna de offentliga idrottsanläggningarna för ett brett deltagande på jämlik basis och utbyta exempel på god praxis i detta hänseende.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att mer kraftfullt stödja hälso- och sjukvårdspersonalens roll i främjandet av idrottsdeltagande och att undersöka hur sjukförsäkringsbolag kan erbjuda incitament som uppmuntrar personer att börja idrotta.
R ESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
12.9.2011
Slutomröstning: resultat
+:
–:
0:
41
1
Slutomröstning: närvarande ledamöter
János Áder, Kriton Arsenis, Sophie Auconie, Pilar Ayuso, Paolo Bartolozzi, Sandrine Bélier, Sergio Berlato, Milan Cabrnoch, Martin Callanan, Nessa Childers, Chris Davies, Bairbre de Brún, Anne Delvaux, Edite Estrela, Julie Girling, Françoise Grossetête, Jolanta Emilia Hibner, Karin Kadenbach, Christa Klaß, Jo Leinen, Peter Liese, Kartika Tamara Liotard, Linda McAvan, Radvilė Morkūnaitė-Mikulėnienė, Miroslav Ouzký, Antonyia Parvanova, Mario Pirillo, Pavel Poc, Anna Rosbach, Oreste Rossi, Daciana Octavia Sârbu, Carl Schlyter, Richard Seeber, Theodoros Skylakakis, Salvatore Tatarella, Anja Weisgerber, Marina Yannakoudakis
Slutomröstning: närvarande suppleanter
YTTRANDE från utskottet för den inre marknaden och konsumentskydd
till utskottet för kultur och utbildning
över idrottens europeiska dimension
( 2011/2087(INI) )
Föredragande:
Eija-Riitta Korhola
FÖRSLAG
Utskottet för den inre marknaden och konsumentskydd uppmanar utskottet för kultur och utbildning att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
A. Idrott är en dynamisk tillväxtsektor och ett redskap för social sammanhållning i ordets sanna bemärkelse, och den har en mycket viktig social, hälsorelaterad och ekonomisk betydelse i EU och dess regioner, där den kan bidra mycket till lokal utveckling av både infrastruktur och ekonomi, och fungera som en stor turistattraktion.
B. På grund av sina särdrag omfattas speltjänster varken av tjänstedirektivet (2006/123/EG) eller det nya direktivet om konsumenters rättigheter (som godkändes av Europaparlamentet den 23 juni 2011).
C. För att trygga finansieringen inom gräsrotsidrotten måste innehavarna av de nödvändiga nationella spellicenserna, som betalar skatter och avgifter och finansierar andra aktiviteter av allmänt intresse i medlemsstaterna, i lag åläggas betala till allmännyttiga ändamål och effektivt skyddas från olaglig konkurrens.
D. Kränkningar av immateriella rättigheter utgör ett verkligt hot mot finansieringen av europeisk idrott på lång sikt.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att inrätta ett system för erkännande av kvalifikationer som förvärvats av frivilliga och av kvalifikationer som krävs för utövandet av reglerade yrken med anknytning till idrotten.
Europaparlamentet insisterar på att rätten att ge ensamrätt på lotterier och andra sifferspel ska ligga kvar hos medlemsstaterna, med tanke på att de europeiska paraplyorganisationerna inom idrott anser att de nationella lotteriernas ekonomiska bidrag till idrotten och framför allt till gräsrotsidrotten är oumbärligt.
Europaparlamentet understryker idrottens fostrande betydelse och uppmuntrar de initiativ som tagits av idrottsorganisationerna och spelarrangörerna för att fostra idrottsutövarna till god praxis vid vadslagning i samband med idrott.
10.
14.
Europaparlamentet stöder kommissionens tillvägagångssätt att undersöka de ekonomiska och juridiska aspekterna på spelarövergångar samt vilken inverkan dessa har på idrottstävlingarna och framför allt på politiken för utbildning av unga spelare inom föreningarna.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
26.9.2011
Slutomröstning: resultat
+:
–:
0:
33
2
Slutomröstning: närvarande ledamöter
Pablo Arias Echeverría, Adam Bielan, Lara Comi, Anna Maria Corazza Bildt, António Fernando Correia De Campos, Jürgen Creutzmann, Cornelis de Jong, Evelyne Gebhardt, Mikael Gustafsson, Małgorzata Handzlik, Malcolm Harbour, Philippe Juvin, Sandra Kalniete, Edvard Kožušník, Kurt Lechner, Toine Manders, Phil Prendergast, Mitro Repo, Heide Rühle, Christel Schaldemose, Andreas Schwab, Emilie Turunen, Bernadette Vergnaud, Barbara Weiler
Slutomröstning: närvarande suppleanter
Frank Engel, Marielle Gallo, Anna Hedh, María Irigoyen Pérez, Othmar Karas, Constance Le Grip, Antonyia Parvanova, Sylvana Rapti, Olle Schmidt, Kyriacos Triantaphyllides, Anja Weisgerber
Föredragande:
Toine Manders
FÖRSLAG
Utskottet för rättsliga frågor uppmanar utskottet för kultur och utbildning att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
A. De värden som idrotten förkroppsligar utsätts för överdrivet kommersiellt tryck som utövas mot bakgrund av ett oklart rättsläge och tar sig uttryck till exempel i form av uppgjorda matcher.
B. Kränkningar av immateriella rättigheter utgör ett allvarligt hot mot finansieringen av europeisk idrott på lång sikt.
C. Det är endast idrottens ekonomiska dimension som omfattas av unionslagstiftningen och reglerna för hur idrottstävlingar organiseras måste förbli utanför dennas tillämpningsområde.
1.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
10.10.2011
Slutomröstning: resultat
+:
–:
0:
14
3
1
Slutomröstning: närvarande ledamöter
Raffaele Baldassarre, Luigi Berlinguer, Sebastian Valentin Bodu, Françoise Castex, Christian Engström, Marielle Gallo, Sajjad Karim, Antonio Masip Hidalgo, Jiří Maštálka, Bernhard Rapkay, Evelyn Regner, Francesco Enrico Speroni, Dimitar Stoyanov, Diana Wallis
Slutomröstning: närvarande suppleanter
Kurt Lechner, Toine Manders, Paulo Rangel
Slutomröstning: närvarande suppleanter (art.
187.2)
Pablo Zalba Bidegain
( 2011/2087(INI) )
Föredragande:
Emine Bozkurt
FÖRSLAG
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor uppmanar utskottet för kultur och utbildning att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet framhåller behovet av insatser mot aktörer som bedriver otillåten spelverksamhet inom EU samt aktörer som bedriver spelverksamhet utanför EU, eftersom dessa kan kringgå övervakningssystemen mot oegentligheter inom idrotten.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
29.9.2011
Slutomröstning: resultat
+:
–:
0:
48
Slutomröstning: närvarande ledamöter
Jan Philipp Albrecht, Sonia Alfano, Alexander Alvaro, Roberta Angelilli, Vilija Blinkevičiūtė, Rita Borsellino, Emine Bozkurt, Simon Busuttil, Carlos Coelho, Rosario Crocetta, Tanja Fajon, Hélène Flautre, Kinga Gál, Kinga Göncz, Nathalie Griesbeck, Sylvie Guillaume, Salvatore Iacolino, Lívia Járóka, Juan Fernando López Aguilar, Monica Luisa Macovei, Clemente Mastella, Véronique Mathieu, Louis Michel, Jan Mulder, Antigoni Papadopoulou, Georgios Papanikolaou, Carmen Romero López, Birgit Sippel, Csaba Sógor, Renate Sommer, Valdemar Tomaševski, Kyriacos Triantaphyllides, Wim van de Camp, Axel Voss, Renate Weber, Tatjana Ždanoka
Slutomröstning: närvarande suppleanter
Edit Bauer, Anna Maria Corazza Bildt, Cornelis de Jong, Ioan Enciu, Monika Hohlmeier, Franziska Keller, Jean Lambert, Mariya Nedelcheva, Hubert Pirker, Debora Serracchiani, Gianni Vattimo
Slutomröstning: närvarande suppleanter (art.
187.2)
Anna Rosbach
YTTRANDE från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män
till utskottet för kultur och utbildning
över idrottens europeiska dimension
( 2011/2087(INI) )
Föredragande: Joanna Senyszyn
FÖRSLAG
Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män uppmanar utskottet för kultur och utbildning att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
– med beaktande av sin resolution av den 21 april 2004 om respekt för centrala arbetsnormer i produktionen av sportartiklar för de olympiska spelen
EUT C 104 E, 30.4.2004, s.
757. ,
– med beaktande av sin resolution av den 5 juni 2003 om kvinnor och idrott
EUT
– med beaktande av sin resolution av den 15 mars 2006 om tvångsprostitution i samband med internationella idrottsevenemang
EUT
C 291 E, 30.11.2006, s 292. ,
– med beaktande av den europeiska stadgan om kvinnors rättigheter inom idrotten (”European Chart of Women’s rights in Sports – Jump in Olympia.
Strong(er) Women through Sport”),
Europaparlamentet uppmanar kommissionen och medlemsstaterna samt relevanta aktörer, idrottsorganisationer och idrottsförbund att garantera män och kvinnor lika tillgång till beslutsfattande positioner inom idrotten och lika tillgång till tränarjobb och till administrativa tjänster inom idrottsorganisationerna.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att överväga mixade idrottsprogram för att utmana och skingra missuppfattningar om kvinnors förmåga, motverka diskriminering och könsstereotypa föreställningar samt stärka kvinnans roll.
11 Europaparlamentet anser att kvinnliga elitidrottare är positiva förebilder för unga, och påpekar därför att medierna spelar en viktig roll för att öka de kvinnliga idrottarnas synlighet.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att höja medvetenheten om vikten av åldersanpassad och barnvänlig idrottsundervisning av god kvalitet för flickor och pojkar redan från förskolan, och föreslår därför att lämpliga strategier och riktlinjer utarbetas.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att göra allt för att främja och garantera en jämn könsfördelning inom skolidrotten och vid offentliga idrottsanläggningar.
17.
Europaparlamentet uppmuntrar till barnpassningsverksamhet vid idrottsanläggningar och idrottshallar, så att mammor och pappor som har hand om små barn kan få lika möjligheter att utöva idrott.
R ESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
15.9.2011
Slutomröstning: resultat
+:
–:
0:
31
1
Slutomröstning: närvarande ledamöter
Regina Bastos, Edit Bauer, Andrea Češková, Tadeusz Cymański, Edite Estrela, Ilda Figueiredo, Iratxe García Pérez, Zita Gurmai, Mary Honeyball, Teresa Jiménez-Becerril Barrio, Nicole Kiil-Nielsen, Rodi Kratsa-Tsagaropoulou, Constance Le Grip, Barbara Matera, Elisabeth Morin-Chartier, Siiri Oviir, Antonyia Parvanova, Raül Romeva i Rueda, Nicole Sinclaire, Joanna Katarzyna Skrzydlewska, Britta Thomsen, Marina Yannakoudakis, Anna Záborská
Slutomröstning: närvarande suppleanter
Izaskun Bilbao Barandica, Jill Evans, Christa Klaß, Kartika Tamara Liotard, Mariya Nedelcheva, Katarína Neveďalová, Norica Nicolai, Antigoni Papadopoulou, Joanna Senyszyn
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
10.11.2011
Slutomröstning: resultat
+:
–:
0:
28
2
Slutomröstning: närvarande ledamöter
Magdi Cristiano Allam, Zoltán Bagó, Malika Benarab-Attou, Lothar Bisky, Piotr Borys, Silvia Costa, Santiago Fisas Ayxela, Mary Honeyball, Cătălin Sorin Ivan, Petra Kammerevert, Morten Løkkegaard, Marek Henryk Migalski, Katarína Neveďalová, Doris Pack, Chrysoula Paliadeli, Marco Scurria, Joanna Senyszyn, Emil Stoyanov, Hannu Takkula, Sampo Terho, Helga Trüpel, Gianni Vattimo, Sabine Verheyen
Slutomröstning: närvarande suppleanter
Slutomröstning: närvarande suppleanter (art.
187.2)
Pablo Zalba Bidegain
A7-0400/2011
Utskottet för utrikesfrågor
Föredragande:
Marek Siwiec och Mário David
PE 469.805v02-00
INNEHÅLL
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION.................................................3
YTTRANDE från utskottet för utveckling ........................................................28
YTTRANDE från budgetutskottet ............................................................................32
YTTRANDE från utskottet för sysselsättning och sociala frågor ...36
YTTRANDE från utskottet för industrifrågor, forskning och energi 41
YTTRANDE från utskottet för regional utveckling ...................................46
YTTRANDE från utskottet för kultur och utbildning ...............................50
YTTRANDE från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor 55
YTTRANDE från utskottet för konstitutionella frågor ..........................59
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET.....................................................62
FÖRSLAG TILL EUROPAPARLAMENTETS RESOLUTION
om översynen av den europeiska grannskapspolitiken
( 2011/2157(INI) )
Europaparlamentet utfärdar denna resolution
– med beaktande av de gemensamma meddelandena från kommissionen och unionens höga representant för utrikes frågor och säkerhetspolitik av den 25 maj 2011 om ny respons på ett grannskap i förändring ( KOM(2011)0303 ) och av den 8 mars 2011 om ett partnerskap för demokrati och delat välstånd med södra Medelhavsområdet ( KOM(2011)0200 ),
– med beaktande av kommissionens meddelanden av den 11 mars 2003 om ett utvidgat europeiskt grannskap: En ny ram för förbindelserna med våra grannländer i öster och söder ( KOM(2003)0104 ), av den 12 maj 2004 om europeiska grannskapspolitiken –strategidokument ( KOM(2004)0373 ), av den 4 december 2006 om stärkande av den europeiska grannskapspolitiken ( KOM(2006)0726 ), av den 5 december 2007 om en stark europeisk grannskapspolitik ( KOM(2007)0774 ), av den 3 december 2008 om ett östligt partnerskap ( KOM(2008)0823 ), av den 20 maj 2008 om Barcelonaprocessen: en union för Medelhavsområdet ( KOM(2008)0319 ), av den 12 maj 2010 om utvärdering av den europeiska grannskapspolitiken ( KOM(2010)0207 ) och av den 24 maj 2011 om en dialog om migration, rörlighet och säkerhet med länderna i södra Medelhavsområdet ( KOM(2011)0292 ),
– med beaktande av utvecklingen av den europeiska grannskapspolitiken sedan 2004, och i synnerhet kommissionens lägesrapporter om dess genomförande,
– med beaktande av de handlingsplaner som antagits gemensamt med Egypten, Israel, Jordanien, Libanon, Marocko, den palestinska myndigheten och Tunisien, samt med Armenien, Azerbajdzjan, Georgien och Moldavien, och av associeringsagendan med Ukraina,
– med beaktande av rådets (utrikes frågor) slutsatser om den europeiska grannskapspolitiken av den 26 juli 2010 och 20 juni 2011 och rådets (utrikes frågor/handel) slutsatser av den 26 september 2011,
– med beaktande av slutsatserna från mötet den 13 december 2010 med utrikesministrarna i de länder som omfattas av det östliga partnerskapet,
– med beaktande av de gemensamma förklaringarna från toppmötena i Prag den 7 maj 2009 respektive Warszawa den 29–30 september 2011 om det östliga partnerskapet,
– med beaktande av Barcelonaförklaringen om upprättandet av ett partnerskap mellan Europa och Medelhavsområdet, vilken antogs vid utrikesministrarnas konferens om Europa-Medelhavsområdet den 27–28 november 1995,
– med beaktande av att Europeiska rådet vid sitt möte i Bryssel den 13–14 mars 2008 godkände Barcelonaprocessen: en union för Medelhavsområdet,
– med beaktande av förklaringen från det Medelhavstoppmöte som hölls i Paris den 13 juli 2008,
– med beaktande av slutsatserna från associeringsrådet EU–Marocko av den 13 oktober 2008, som gav Marocko en framskjuten ställning,
– med beaktande av slutsatserna från associeringsrådet EU–Jordanien av den 26 oktober 2010, som gav Jordanien en framskjuten ställning,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1638/2006 av den 24 oktober 2006 om fastställande av allmänna bestämmelser för upprättandet av ett europeiskt grannskaps- och partnerskapsinstrument
EUT L 310, 9.11.2006, s.
1. ,
– med beaktande av sin skriftliga förklaring nr 15/2011 av den 27 september 2011 om inrättandet av Erasmus- och Leonardo da Vinci-program för Europa‑Medelhavsområdet,
– med beaktande av Europeiska revisionsrättens särskilda rapport nr 13/2010 med titeln ”Har det nya europeiska grannskaps- och partnerskapsinstrumentet införts på ett bra sätt och leder det till att resultat uppnås i Södra Kaukasien (Armenien, Azerbajdzjan och Georgien)?”,
EUT L 211, 27.8.2011. ,
– med beaktande av sina resolutioner om översynen av den europeiska grannskapspolitiken – den östliga dimensionen och om översynen av den europeiska grannskapspolitiken – den sydliga dimensionen av den 7 april 2011 ( B7‑0198/2011 och B7-0199/2011 ),
– med beaktande av sina resolutioner av den 19 januari 2006 om den europeiska grannskapspolitiken
EUT C 287 E, 19.1.2006, s.
312. , av den 15 november 2007 om stärkande av den europeiska grannskapspolitiken
EUT C 282 E, 6.11.2008, s.
443. , av den 6 juli 2006 om det europeiska grannskaps- och partnerskapsinstrumentet (ENPI)
EUT C 303 E, 13.12.2006, s.
760. , av den 5 juni 2008 om rådets årliga rapport till Europaparlamentet om de viktigaste aspekterna och de grundläggande vägvalen när det gäller den gemensamma utrikes- och säkerhetspolitiken (Gusp)
EUT C 285 E, 26.11.2009, s.
11. , av den 19 februari 2009 om översynen av det europeiska grannskaps- och partnerskapsinstrumentet
EUT C 76 E, 25.3.2010, s.
83. , av den 19 februari 2009 om Barcelonaprocessen: union för Medelhavsområdet
EUT C 76 E, 25.3.2010, s.
76. , av den 17 januari 2008 om en strategi för regionalpolitiken vid Svarta havet
EUT C 41 E, 19.2.2009, s.
64. , av den 20 januari 2011 om en EU-strategi för Svarta havet
Antagna texter, P7_TA(2011)0025 . , av den 20 maj 2010 om en union för Medelhavsområdet
Antagna texter, P7_TA(2010)0192 . , av den 20 maj 2010 om behovet av en EU-strategi för Sydkaukasien
Antagna texter, P7_TA(2010)0193 . , av den 9 september 2010 om situationen i Jordanfloden, särskilt det nedre flodområdet
Antagna texter, P7_TA(2010)0314 . , av den 3 februari 2011 om situationen i Tunisien
Antagna texter, P7_TA(2011)0038 . , av den 17 februari 2011 om situationen i Egypten
Antagna texter, P7_TA(2011)0064 . , av den 10 mars 2011 om det södra grannskapet och särskilt Libyen, inklusive humanitära aspekter
Antagna texter, P7_TA(2011)0095 . , av den 7 juli 2011 om Syrien, Jemen och Bahrain mot bakgrund av situationen i arabvärlden och Nordafrika, av den 15 september 2011 och 20 januari 2011 om situationen i Vitryssland och alla sina tidigare resolutioner om Vitryssland och av den 15 september 2011 om situationen i Libyen
Antagna texter, P7_TA(2011)0386 . respektive Syrien
Antagna texter, P7_TA(2011)0387 . ,
– med beaktande av de rekommendationer som antogs av kommittéerna i den parlamentariska församlingen för unionen för Medelhavsområdet vid dess sjunde sammanträdesperiod som hölls i Rom den 3 och 4 mars 2011,
– med beaktande av den konstituerande akten för den parlamentariska församlingen Euronest av den 3 maj 2011,
– med beaktande av slutsatserna från det inledande mötet för församlingen för regionala och lokala myndigheter i Europa–Medelhavsområdet (Arlem), vilket hölls i Barcelona den 21 januari 2010,
– med beaktande av sin resolution om de kulturella aspekterna i EU:s yttre åtgärder ( 2010/2161(INI) )1,
– med beaktande av artiklarna 8 och 21 i fördraget om Europeiska unionen,
– med beaktande av artikel 48 i arbetsordningen,
– med beaktande av betänkandet från utskottet för utrikesfrågor och yttrandena från utskottet för utveckling, budgetutskottet, utskottet för sysselsättning och sociala frågor, utskottet för industrifrågor, forskning och energi, utskottet för regional utveckling, utskottet för kultur och utbildning, utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor och utskottet för konstitutionella frågor ( A7-0400/2011 ), och av följande skäl:
A. Respekt för och främjande av demokrati och mänskliga rättigheter, i synnerhet kvinnors, barns och minoriteters rättigheter; rättvisa och rättssäkerhet, grundläggande friheter, bland annat yttrandefrihet, samvetsfrihet, religions- eller trosfrihet, frihet att vara öppen med sin sexuella läggning, mötes- och föreningsfrihet och mediefrihet, inklusive obegränsad tillgång till information, kommunikation och internet; en förstärkning av det civila samhället, säkerhet, bland annat fredlig konfliktlösning och goda grannförbindelser; demokratisk stabilitet, välstånd, en rättvis fördelning av inkomster, rikedomar och möjligheter; social sammanhållning, korruptionsbekämpning och främjande av en god samhällsstyrning och hållbar utveckling tillhör EU:s grundläggande principer och mål och måste utgöra de gemensamma värden som ligger till grund för översynen av den europeiska grannskapspolitiken.
B. Det ligger i högsta grad i EU:s intresse att vara ambitiöst i det ekonomiska samarbetet och anta en ömsesidigt gynnsam, ansvarsfull och flexibel strategi som bygger på stöd till demokratiseringsprocesser och försvar av de mänskliga rättigheterna.
E. Samarbetet inom den parlamentariska församlingen Euronest syftar till att skapa positiva effekter genom att tjäna som ett forum för att utbyta åsikter, skapa gemensamma synsätt kring vår tids globala utmaningar när det gäller demokrati, politik, ekonomi, energitrygghet och sociala frågor samt stärka banden mellan länderna i regionen och EU.
F. I artikel 49 i EU-fördraget står det att varje europeisk stat som respekterar de värden som unionen bygger på – det vill säga demokrati, rättsstatsprincipen och respekt för de mänskliga rättigheterna och de grundläggande friheterna – och som förbinder sig att främja dem, får ansöka om att bli medlem av unionen.
G. Starkare förbindelser kräver en tydlig och konstaterad reformvilja med målet att göra konkreta framsteg som uppfyller de förutbestämda riktmärkena.
J. Europaparlamentet har genom sin skriftliga förklaring nr 15/2011 av den 27 september 2011 gett sitt stöd till inrättandet av Erasmus- och Leonardo da Vinci-program för Europa–Medelhavsområdet.
2.
Europaparlamentet anser att en fullständig och effektiv respekt för religionsfriheten (individuellt, kollektivt, offentligt, privat och institutionellt) bör fastställas som en prioritet, särskilt för alla religiösa minoriteter i området, tillsammans med behovet av konkret hjälp för dessa grupper.
Europaparlamentet uppmanar kommissionen att göra projekten inom det östliga partnerskapet och unionen för Medelhavsområdet synligare i partnerländerna och lättare att förstå för medborgarna i dessa länder, bland annat genom att tydliggöra det mervärde som det innebär att samarbeta med EU.
Hållbar ekonomisk och social utveckling
Europaparlamentet uppmanar med kraft kommissionen att stödja uppbyggnaden av administrativ kapacitet i sysselsättningsfrågor och sociala frågor, med särskild tonvikt på kapacitetsbyggande inom juridiska tjänster, vilket kommer att säkerställa bättre förberedelser för genomförandet av reformer.
Europaparlamentet uppmanar kommissionen att ta till sig strategidokumenten för fattigdomsminskning och låta dessa vara den vägledande politiska ramen för en ekonomisk tillväxt på medellång sikt som gynnar de fattiga, och för en rättvisare resursfördelning utifrån landets behov.
Associeringsavtal
Sektor iellt samarbete
Europaparlamentet hänvisar också till den understödjande roll som EU kan spela för att åtgärda miljöproblem i våra grannländer, särskilt när det gäller att eliminera omfattande lager av gamla bekämpningsmedel som kan medföra kemiska föroreningar i stor skala.
Parlamentet uppmanar därför kommissionen att stärka och öka Taiex1 och programmen för partnersamverkan med lokala myndigheter i EU och partnerskapsländer.
Rörlighet
Europaparlamentet påpekar i detta sammanhang att medlemsstaterna måste respektera principen om icke-avvisning (”non-refoulement”) och göra allt för att underlätta uppbyggnaden av ett tillgängligt och rättvist europeiskt asylsystem som tillhandahåller skydd.
Europaparlamentet uppmanar rådet och kommissionen att inleda en strukturerad dialog med myndigheter i tredjeländer i syfte att utarbeta en rörlighetsstrategi som gynnar alla parter, underlätta viseringsförfaranden, i ökad utsträckning använda de möjligheter som erbjuds genom EU:s viseringskodex och förbättra och harmonisera tillämpningen av denna för att garantera lika och rättvisa villkor för sökande i alla medlemsstater, med särskilt fokus på effekterna av det ömsesidiga beroendet mellan utvecklingsbistånd, säkerhet, reguljär migration och irreguljär migration enligt definitionerna i den övergripande strategin för migration.
Den regionala dimensionen
Europaparlamentet framhåller euroregionernas mycket viktiga bidrag till uppnåendet av de sammanhållningspolitiska målen, och uppmuntrar kommissionen att främja och stödja dessa regioners utveckling, särskilt i gränsområden, i syfte att stärka euroregionernas roll i den europeiska grannskapspolitiken.
Europaparlamentet påminner om att den europeiska grannskapspolitiken i sina multilaterala aspekter bör stödja ett snabbt och effektivt igångsättande av konkreta projekt som fastställts av unionen för Medelhavsområdet och som är avsedda att möjliggöra en gemensam utvecklings- och integrationsprocess, inte minst genom samfinansiering av genomförbarhetsstudier och stöd till en ökning av koncessionslånen.
EU och konfliktlösning
Så här efter revolutionerna i Nordafrika betonar Europaparlamentet vikten av stöd till rättsväsendet i övergångsskedet och vädjar till alla partnerländer att samarbeta med den internationella rättskipningen, särskilt Internationella brottmålsdomstolen.
Den parlamentariska dimensionen
Europaparlamentet bekräftar sin beredvillighet att välkomna företrädare från det vitryska parlamentet till Euronest så snart som parlamentsvalen i Vitryssland betraktas som demokratiska av världssamfundet, inklusive OSSE.
Finansiering
Europaparlamentet anser att översynen av det europeiska grannskapsinstrumentet måste vara förenlig med, och genomföras inom ramen för, den pågående utvärderingen av den fleråriga budgetramen för 2007–2013 och förhandlingarna om perioden efter 2013, så att man slipper inleda nya förhandlingar om finansieringen av grannskapspolitiken under 2012 och 2013.
Europaparlamentet understryker att den omfördelning av anslagen som behövs för en ökad finansiering av den europeiska grannskapspolitiken bör utgå från tydliga prioriteringar och därför inte ske på bekostnad av EU:s enda verktyg för krishantering och fredsskapande, nämligen stabilitetsinstrumentet, så som kommissionen har föreslagit.
*
* *
114.Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik, Europeiska utrikestjänsten, regeringarna och parlamenten i medlemsstaterna och länderna i den europeiska grannskapspolitiken samt till generalsekreteraren för unionen för Medelhavsområdet.
Föredragande: Michèle Striffler
FÖRSLAG
Utskottet för utveckling uppmanar utskottet för utrikesfrågor att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Därför uppmanar parlamentet kommissionen och Europeiska utrikestjänsten att alltid ha dessa mål, nämligen att minska och på sikt utrota fattigdomen, för ögonen när de genomför den europeiska grannskapspolitiken, oavsett om det handlar om partnerländerna i det östra grannskapet eller om dem i det södra grannskapet.
2.
Europaparlamentet begär att mandatet för EU:s särskilde representant i södra Medelhavsområdet ska omfatta utvecklingsfrågor, eftersom representanten kan spela en avgörande roll för att se till att de demokratiska framstegen åtföljs av bestående framsteg på utvecklingsområdet, särskilt en förbättring av de sociala och ekonomiska villkoren i de berörda länderna.
Europaparlamentet understryker att det är särskilt viktigt att EU:s program för utveckling och mänskliga rättigheter stöder det civila samhället, där de verkliga aktörerna i processerna finns, i synnerhet kvinno- och ungdomsorganisationer.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
7.11.2011
Slutomröstning: resultat
+:
–:
0:
21
Slutomröstning: närvarande ledamöter
Thijs Berman, Leonidas Donskis, Charles Goerens, András Gyürk, Eva Joly, Franziska Keller, Miguel Angel Martínez Martínez, Norbert Neuser, Birgit Schnieber-Jastram, Michèle Striffler, Alf Svensson, Patrice Tirolien, Ivo Vajgl, Anna Záborská
Slutomröstning: närvarande suppleanter
Santiago Fisas Ayxela, Fiona Hall, Krzysztof Lisek, Isabella Lövin, Horst Schnellhardt, Giancarlo Scottà, Jan Zahradil
Slutomröstning: närvarande suppleanter (art.
187.2)
Föredragande:
Göran Färm
FÖRSLAG
Europaparlamentet anser att en konstruktiv långsiktig grannskapspolitik inte bara är av avgörande betydelse för partnerskapsländerna när det gäller att främja framsteg mot fred, demokrati, stabilitet och välstånd, utan också av strategisk betydelse för EU med tanke på hur viktiga partnerländerna i både öster och söder är för vår gemensamma säkerhet, miljö och ekonomiska utveckling.
Europaparlamentet anser att översynen av det europeiska grannskapsinstrumentet måste vara förenlig med, och genomföras inom ramen för, den pågående utvärderingen av den fleråriga budgetramen för 2007–2013 och förhandlingarna om perioden efter 2013, detta för att slippa inleda nya förhandlingar om finansieringen av grannskapspolitiken under 2012 och 2013.
Parlamentet anser att det är nödvändigt att det reviderade europeiska grannskapsinstrumentet inte försummar denna dimension och att det har möjlighet att snabbt stödja och samverka med andra finansieringsinstrument som rör flyktingar, till exempel Europeiska flyktingfonden, Europeiska återvändandefonden och Europeiska fonden för de yttre gränserna.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
7.11.2011
Slutomröstning: resultat
+:
–:
0:
25
2
Slutomröstning: närvarande ledamöter
Marta Andreasen, Francesca Balzani, Reimer Böge, Lajos Bokros, Isabelle Durant, James Elles, José Manuel Fernandes, Eider Gardiazábal Rubial, Salvador Garriga Polledo, Carl Haglund, Lucas Hartong, Jutta Haug, Sidonia Elżbieta Jędrzejewska, Ivailo Kalfin, Jan Kozłowski, Alain Lamassoure, Vladimír Maňka, Barbara Matera, Nadezhda Neynsky, Dominique Riquet, László Surján, Derek Vaughan
Slutomröstning: närvarande suppleanter
François Alfonsi, Frédéric Daerden, Jürgen Klute, Georgios Stavrakakis
Slutomröstning: närvarande suppleanter (art.
187.2)
Marisa Matias
Föredragande: Sylvana Rapti
FÖRSLAG
Utskottet för sysselsättning och sociala frågor uppmanar utskottet för utrikesfrågor att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
A. En hållbar ekonomisk tillväxt förutsätter en helhetssyn till förmån för sysselsättning och socialt skydd.
B. Den europeiska grannskapspolitiken är avgörande för stabiliteten i EU:s grannländer och bidrar till säkerhet och utveckling för alla och det finns ett gemensamt intresse av att ett större område runt Europa är demokratiskt, stabilt, välmående och fredligt.
C. EU tjänar globalt som en modell för social utveckling och kan erbjuda värdefull expertis om ansvarsfull tillväxt.
D. Den nya europeiska grannskapspolitiken omprövas och måste ständigt omprövas, i förhållande såväl till den utveckling som sker i grannländerna som till frågor av gemensamt intresse och bör omformas och inrättas för att kunna hantera de historiska utmaningarna samt prioritera akuta situationer.
E. Initiativtagandet till de demokratiska förändringarna i Nordafrika kom från invånare, huvudsakligen bland den unga generationen, i samhällen med ojämlik förmögenhetsfördelning, stor arbetslöshet, bristande social trygghet och avsaknad av utbildning och framtidsutsikter – invånare som till och med lever under fattigdomsgränsen och överlever endast tack vare den informella ekonomin.
F. Regionen med partnerländerna i södra Medelhavsområdet har en av världens lägsta förvärvsfrekvenser och händelserna i början av 2011 har i vissa partnerländer öppnat nya möjligheter att ta sig an de utmaningar som sysselsättningsskapandet innebär.
G. Den europeiska grannskapspolitiken kräver att problemen i den östliga respektive den sydliga dimensionen behandlas lika, med hänsyn till såväl demokratin som till ekonomiska och sociala frågor.
H. Befolkningsutvecklingen i olika regioner som omfattas av den europeiska grannskapspolitiken varierar kraftigt.
Europaparlamentet uppmanar med kraft grannskapsländerna att ratificera alla ILO:s grundläggande arbetskonventioner och anpassa den nationella lagstiftningen därefter.
Europaparlamentet framhåller att den europeiska grannskapspolitiken bör utgöra grunden för effektivt samarbete mot illegal invandring, eftersom partnerländerna är både ursprungs- och genomgångsländer för illegala invandrare, tillsammans med effektiv gränskontroll, bekämpande av organiserad brottslighet och således främjande av de mänskliga rättigheterna.
Europaparlamentet välkomnar initiativ för studentutbyte och utbyte inom yrkesutbildningen, såsom den nyligen antagna skriftliga förklaringen om inrättandet av Erasmus- och Leonardo da Vinci-program i Europa–Medelhavsområdet.
Europaparlamentet understryker vikten av att samordna politiken mellan EU och medlemsstaterna för att få bättre resultat på områden av ömsesidigt intresse, men också för att fastställa standardiserade villkor.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
7.11.2011
Slutomröstning: resultat
+:
–:
0:
31
3
Slutomröstning: närvarande ledamöter
Edit Bauer, Jean-Luc Bennahmias, Pervenche Berès, Philippe Boulland, Milan Cabrnoch, Alejandro Cercas, Ole Christensen, Frédéric Daerden, Karima Delli, Frank Engel, Richard Falbr, Marian Harkin, Roger Helmer, Liisa Jaakonsaari, Ádám Kósa, Veronica Lope Fontagné, Elizabeth Lynne, Thomas Mann, Elisabeth Morin-Chartier, Siiri Oviir, Konstantinos Poupakis, Sylvana Rapti, Elisabeth Schroedter, Jutta Steinruck, Traian Ungureanu, Andrea Zanoni
Slutomröstning: närvarande suppleanter
Georges Bach, Raffaele Baldassarre, Edite Estrela, Julie Girling, Richard Howitt, Ria Oomen-Ruijten, Emilie Turunen
Slutomröstning: närvarande suppleanter (art.
187.2)
Catherine Bearder
Föredragande: Bogdan Kazimierz Marcinkiewicz
FÖRSLAG
Europaparlamentet välkomnar förslaget om att skapa en europeisk energigemenskap, och anser att detta skulle kunna utgöra ett viktigt steg mot ett samarbete med våra grannländer.
Europaparlamentet uppmanar kommissionen att vidareutveckla EU:s Svartahavsstrategi, eftersom den utgör en viktig del av EU:s energistrategi gentemot omvärlden med tanke på dess geostrategiska roll, som gör att den i hög grad kan bidra till energitrygghet och diversifiering av energikällor.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
20.10.2011
Slutomröstning: resultat
+:
–:
0:
35
4
Slutomröstning: närvarande ledamöter
Slutomröstning: närvarande suppleanter
Maria Badia i Cutchet, Jolanta Emilia Hibner, Sajjad Karim, Bernd Lange, Markus Pieper, Hannu Takkula, Silvia-Adriana Ţicău, Catherine Trautmann, Hermann Winkler
Slutomröstning: närvarande suppleanter (art.
187.2)
Judith Sargentini
Föredragande: Lena Kolarska-Bobińska
FÖRSLAG
Utskottet för regional utveckling uppmanar utskottet för utrikesfrågor att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
6.10.2011
Slutomröstning: resultat
+:
–:
0:
40
2
1
Slutomröstning: närvarande ledamöter
François Alfonsi, Luís Paulo Alves, Charalampos Angourakis, Catherine Bearder, Jean-Paul Besset, Victor Boştinaru, Philip Bradbourn, Zuzana Brzobohatá, John Bufton, Alain Cadec, Salvatore Caronna, Tamás Deutsch, Rosa Estaràs Ferragut, Brice Hortefeux, Danuta Maria Hübner, Filiz Hakaeva Hyusmenova, Juozas Imbrasas, María Irigoyen Pérez, Seán Kelly, Mojca Kleva, Elżbieta Katarzyna Łukacijewska, Ramona Nicole Mănescu, Riikka Manner, Iosif Matula, Erminia Mazzoni, Lambert van Nistelrooij, Jan Olbrycht, Monika Smolková, Georgios Stavrakakis, Nuno Teixeira, Michail Tremopoulos, Viktor Uspaskich, Oldřich Vlasák, Kerstin Westphal, Joachim Zeller
Slutomröstning: närvarande suppleanter
Jens Geier, Lena Kolarska-Bobińska, Maurice Ponga, Elisabeth Schroedter, Patrice Tirolien, Giommaria Uggias, Derek Vaughan, Sabine Verheyen
Föredragande: Marek Henryk Migalski
FÖRSLAG
Utskottet för kultur och utbildning uppmanar utskottet för utrikesfrågor att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet uppskattar den effekt som Europa-Medelhavsuniversitetet har haft och anser att denna framgång bör spridas och att ett liknande initiativ bör inledas för den östliga partnerskapsregionen.
Europaparlamentet påpekar dessutom att kultur- och rörlighetsprogrammen även bör beakta rörligheten för konstnärer och personer som bedriver konstnärsstudier, eftersom det underlättar ett kreativt och kulturellt berikande utbyte.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
5.10.2011
Slutomröstning: resultat
+:
–:
0:
26
2
Slutomröstning: närvarande ledamöter
Magdi Cristiano Allam, Maria Badia i Cutchet, Malika Benarab-Attou, Lothar Bisky, Jean-Marie Cavada, Santiago Fisas Ayxela, Mary Honeyball, Cătălin Sorin Ivan, Petra Kammerevert, Morten Løkkegaard, Marek Henryk Migalski, Katarína Neveďalová, Doris Pack, Chrysoula Paliadeli, Marie-Thérèse Sanchez-Schmid, Marietje Schaake, Marco Scurria, Hannu Takkula, Sampo Terho, László Tőkés, Helga Trüpel, Sabine Verheyen, Milan Zver
Slutomröstning: närvarande suppleanter
Slutomröstning: närvarande suppleanter (art.
187.2)
Jacky Hénin
( 2011/2157(INI) )
Föredragande:
Hélène Flautre
FÖRSLAG
Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor uppmanar utskottet för utrikesfrågor att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
Europaparlamentet anser att översynen av den europeiska grannskapspolitiken ger EU en möjlighet att effektivt uppnå sina mål och följa sina värderingar enligt artiklarna 2, 3, 6, 8 och 21 i EU-fördraget.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
17.10.2011
Slutomröstning: resultat
+:
–:
0:
35
2
Slutomröstning: närvarande ledamöter
Jan Philipp Albrecht, Rita Borsellino, Simon Busuttil, Philip Claeys, Carlos Coelho, Tanja Fajon, Hélène Flautre, Kinga Gál, Kinga Göncz, Ágnes Hankiss, Anna Hedh, Salvatore Iacolino, Sophia in ‘t Veld, Lívia Járóka, Teresa Jiménez-Becerril Barrio, Juan Fernando López Aguilar, Baroness Sarah Ludford, Monica Luisa Macovei, Véronique Mathieu, Claude Moraes, Jan Mulder, Georgios Papanikolaou, Carmen Romero López, Judith Sargentini, Birgit Sippel, Csaba Sógor, Rui Tavares, Kyriacos Triantaphyllides, Axel Voss, Auke Zijlstra
Slutomröstning: närvarande suppleanter
Edit Bauer, Anna Maria Corazza Bildt, Dimitrios Droutsas, Ana Gomes
Slutomröstning: närvarande suppleanter (art.
187.2)
Albert Deß, Mikael Gustafsson, Gabriele Zimmer
FÖRSLAG
Utskottet för konstitutionella frågor uppmanar utskottet för utrikesfrågor att som ansvarigt utskott infoga följande i sitt resolutionsförslag:
För att denna dimension ska fungera väl bör en systematisk utvärdering göras av hur Euronest och den parlamentariska församlingen för unionen för Medelhavsområdet fungerar i praktiken i syfte att förbättra dem där det är möjligt.
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
24.10.2011
Slutomröstning: resultat
+:
–:
0:
15
1
1
Slutomröstning: närvarande ledamöter
Andrew Henry William Brons, Carlo Casini, Andrew Duff, Roberto Gualtieri, Zita Gurmai, Stanimir Ilchev, Constance Le Grip, David Martin, Paulo Rangel, György Schöpflin, József Szájer, Rafał Trzaskowski
Slutomröstning: närvarande suppleanter
Sandrine Bélier, Zuzana Brzobohatá, Marietta Giannakou, Helmut Scholz, Alexandra Thein
RESULTAT AV SLUTOMRÖSTNINGEN I UTSKOTTET
Antagande
17.11.2011
Slutomröstning: resultat
+:
–:
0:
57
5
Slutomröstning: närvarande ledamöter
Gabriele Albertini, Pino Arlacchi, Bastiaan Belder, Elmar Brok, Arnaud Danjean, Mário David, Michael Gahler, Ana Gomes, Andrzej Grzyb, Takis Hadjigeorgiou, Anna Ibrisagic, Anneli Jäätteenmäki, Jelko Kacin, Othmar Karas, Ioannis Kasoulides, Nicole Kiil-Nielsen, Maria Eleni Koppa, Andrey Kovatchev, Eduard Kukan, Vytautas Landsbergis, Krzysztof Lisek, Sabine Lösing, Ulrike Lunacek, Mario Mauro, Kyriakos Mavronikolas, Francisco José Millán Mon, Alexander Mirsky, María Muñiz De Urquiza, Annemie Neyts-Uyttebroeck, Norica Nicolai, Raimon Obiols, Pier Antonio Panzeri, Ioan Mircea Paşcu, Alojz Peterle, Bernd Posselt, Hans-Gert Pöttering, Cristian Dan Preda, Fiorello Provera, Tokia Saïfi, José Ignacio Salafranca Sánchez-Neyra, Nikolaos Salavrakos, Jacek Saryusz-Wolski, Werner Schulz, Marek Siwiec, Hannes Swoboda, Kristian Vigenin, Boris Zala
Slutomröstning: närvarande suppleanter
Charalampos Angourakis, Véronique De Keyser, Andrew Duff, Göran Färm, Hélène Flautre, Roberto Gualtieri, Doris Pack, Helmut Scholz, György Schöpflin, Alf Svensson, Traian Ungureanu, Ivo Vajgl
Slutomröstning: närvarande suppleanter (art.
187.2)
Marije Cornelissen, Rui Tavares, Ramon Tremosa i Balcells
30.5.2005
FÖRSLAG TILL RESOLUTION
till följd av uttalandena av rådet och kommissionen
från Armin Laschet
för utskottet för utrikesfrågor
om en reform av Förenta Nationerna
Europaparlamentets resolution om en reform av Förenta Nationerna
Europaparlamentet utfärdar denna resolution
–
med beaktande av sin resolution av den 29 januari 2004 om förbindelserna mellan EU och FN, EUT C 96 E, 21.4.2004, s.
75.
–
med beaktande av rapporten ”A more secure world: our shared responsibility” (”En säkrare värld: vårt delade ansvar”) från FN:s högnivåpanel om hot, utmaningar och förändringar, offentliggjord den 1 december 2004.
–
med beaktanden av översynsrapporten om FN:s millenieprojekt och handlingsplanen för att uppnå millennieutvecklingsmålen inom 2015,
–
med beaktande av rapporten ”In larger freedom: towards development, security and human rights for all” (”I större frihet: på väg mot utveckling, säkerhet och mänskliga rättigheter för alla”) från FN:s generalsekreterare, offentliggjord den 21 mars 2005,
–
A.
Högnivåpanelens rapport innehåller mer än hundra rekommendationer om ändringar och behovet att reformera FN för att kunna möta olika utmaningar och hot, från fattigdom, infektionssjukdomar, miljöskador och civilt våld till terrorism, massförstörelsevapen och ickespridning av kärnvapen, och generalsekreterarens rapport understryker och stöder de flesta av dessa rekommendationer.
B.
Högnivåpanelen presenterar i sin rapport en ny syn på kollektiv säkerhet, och uppmärksammar alla de allvarliga hot mot internationell fred och säkerhet som aktualiserats runt om i världen.
C.
D.
I högnivåpanelens rapport anges klart och tydligt att våld, i den mån det är nödvändigt, endast får tillgripas som sista utväg, och att FN:s säkerhetsråd bör slå fast detta i en resolution om principerna för användning av våld, och den ger tveklöst stöd åt den ”framväxande norm” enligt vilken det finns ett kollektivt internationellt ansvar att erbjuda skydd i händelse av folkmord och andra former av storskaligt dödande, etniska rensningar eller allvarliga kränkningar av internationell folkrätt som enskilda regeringar har visat sig maktlösa mot eller ovilliga att förhindra.
E.
Att införa verklig multilateralism är det lämpligaste sättet att lösa de problem och hot som det internationella samfundet står inför, under förutsättning att det bygger på välanpassade institutioner och effektiva förfaranden för att fatta beslut och se till att de genomförs.
F.
Generalsekreteraren understryker i sin rapport nödvändigheten att vidta åtgärder och omgående genomföra en reform, och presenterar en rad konkreta åtgärder som utan vidare kan vidtas efter beslut av stats- och regeringscheferna i september 2005.
G.
EU:s medlemsstater måste gå i spetsen när det gäller ansträngningar att få till stånd universellt anslutning till multilaterala konventioner.
Kollektiv säkerhet i det tjugoförsta århundradet: förebyggande, medvetandegörande och delat ansvar
1.
Europaparlamentet välkomnar varmt generalsekreterarens rapport som följde rapporten från högnivåpanelen om hot, utmaningar och förändringar, och den beslutsamhet som ligger till grund för denna om att genomföra en konsekvent och genomgående reform av FN för att anpassa organisationen till de nya förhållanden som råder runt om i världen samt se till att den tillhandahåller kollektiv säkerhet i det tjugoförsta århundradet på ett sätt som är effektivt, rättvist och långsiktigt samt garanterar den demokratiska insynen.
2.
Europaparlamentet uppmanar rådet att fullt ut stödja Kofi Annans rapport om reformen, och uppmanar det luxemburgska ordförandeskapet att försöka få rådet att anta ett beslut om en gemensam hållning från EU:s sida i förhållande till konkreta FN-reformer.
3.
4.
5.
6.
7.
Europaparlamentet stöder garantier för leveranser av det bränsle som krävs för att utveckla fredliga användningsområden, t.ex. en lösning där IAEA skulle garantera leveranser till marknadspriser av klyvbart material till civila kärnenergianvändare för de stater som frivilligt avstår från att utveckla nationella anläggningar för anrikning av uran och separering av plutonium.
8.
Europaparlamentet stöder tanken att FN utvecklar en strategi för att bekämpa terrorism som kännetecknas av respekt för de mänskliga rättigheterna och rättsstatsprincipen, som inbegriper det civila samhället och som bygger på de fem pelarna att avskräcka potentiella terrorister från att begå eller stödja terroristhandlingar, blockera terroristers tillgång till finansiering och materiella resurser, avskräcka stater från att stödja terrorism, utveckla staters förmåga att bekämpa terrorism samt skydda de mänskliga rättigheterna.
9.
Europaparlamentet ser fram emot att FN:s generalförsamling avslutar arbetet med en heltäckande konvention om terrorism som utgår från en tydlig och accepterad definition som beaktar de mänskliga rättigheterna och demokratiska friheterna, och som bland annat innehåller hänvisningar till begreppsdefinitionerna i den internationella överenskommelsen från 1999 om bekämpning av terrorismfinansiering och i FN:s säkerhetsråds resolution 1566, och i vilken det på nytt fastslås att sådana handlingar som omfattas av de tolv tidigare överenskommelserna om bekämpning av terrorism utgör terrorism samt förklaras att sådana handlingar uppfyller brottsrekvisitet för brott mot folkrätten.
10.
En värld utan nöd: en gemensam och balanserad syn på en ny utvecklingspolitik för FN
11.
12.
13.
Europaparlamentet framhåller behovet av att ytterligare främja vetenskaplig forskning och utveckling för att garantera en hållbar miljö, bekämpa klimatförändringarna och tillgodose utvecklingsländernas särskilda behov när det gäller jordbruk, naturresurser och miljöförvaltning.
14.
Europaparlamentet erinrar om att ett framgångsrikt partnerskap måste baseras på en tvåvägsprocess där utvecklingsländerna måste stärka sin förvaltning, bekämpa korruptionen och maximera de inhemska resurserna för att finansiera nationella utvecklingsstrategier, samtidigt som industriländerna måste understödja dessa ansträngningar genom att bli effektivare i sin tilldelning av utvecklingsstöd, underlätta tillgången till sina marknader och bevilja skuldlättnader.
15.
16.
Parlamentet stöder fullt ut generalsekreterarens särskilda uppmaningar inom detta område, inklusive att fastställa en tydlig tidsplan för när de utvecklade länderna skall uppnå målet att avsätta 0,7 procent av BNI till offentligt utvecklingsbistånd, att erkänna Afrikas särskilda behov, att inleda en rad snabba initiativ för att göra större omedelbara framsteg mot millennieutvecklingsmålen, inklusive avskaffande av användarnas avgifter för grundläggande hälsovård och utbildning.
17.
Parlamentet bekräftar att FN:s beslutsfattande organ bör ha behörigheten – och ansvaret – att både fastställa gemensamma nyttigheter och införa normer för att garantera och anta bestämmelser för bevarande och skydd av dessa gemensamma nyttigheter, och att bl.a. fastställa internationella regler som syftar till att klargöra förhållandet mellan handel och miljö i syfte att skydda de multilaterala miljöavtalen från handelsbestämmelserna.
Förnyade institutioner för större representativitet och effektivitet
18.
19.
20.
21.
22.
Europaparlamentet stöder till fullo högnivåpanelens förslag att införa en mekanism för vägledande omröstning i säkerhetsrådet, genom vilken medlemmarna kunde uppmana till offentlig tillkännagivande av ståndpunkterna rörande en föreslagen insats, och där nej‑röster inte har vetoeffekt och den slutliga omröstningen inte är juridiskt bindande, men i stället skulle ansvaret i förhållande till vetomöjligheten öka.
23.
24.
25.
26.
27.
28.
29.
30.
31.
32.
33.
34.
35.
36.
37.
38.
Europaparlamentet uppmanar medlemsstaterna att stödja och stärka FN:s ”demokratiska rådslag” som främjar demokratin i FN:s medlemsstater och stödjer utvecklingen av demokratiska strukturer inom FN-systemet genom att vara en modell för demokratier i sin linda, och samtidigt hindra att FN-organ har sina säten i icke-demokratiska, auktoritära stater, vilket kan skada FN:s trovärdighet.
39.
40.
41.
42.
Europaparlamentet uppmanar enträget EU:s medlemsstater att utan dröjsmål stödja reformförslaget i generalsekreterarens rapport som följer på rapporten från högnivåpanelen, och göra allt man kan för att genomföra dessa reformer i lämpliga områden och att i samarbete med EU:s institutioner se till att få fram nödvändiga resurser för detta syfte.
43.
Europaparlamentet uppmanar presidiet att ge en grupp experter i uppdrag att utarbeta en skiss över hur den totala reformen av FN-systemet skulle inverka dels på FN-stadgan, dels på verksamheten vid EU:s institutioner.
44.
Europaparlamentet beslutar att en genomföra en serie informationskampanjer riktade till allmänheten såväl inom som utom Europa för att informera om FN-reformens historiska betydelse om och de konsekvenser denna kommer att få för det institutionella systemet i Europa.
45.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, EU:s medlemsstater, FN:s generalsekreterare, ordföranden för FN:s säkerhetsråd, ordföranden för FN:s generalförsamling, ordföranden för FN:s ekonomiska och sociala råd, medlemmarna i högnivåpanel för en reform av FN samt EU‑medlemsstaternas parlament, Förenta staternas kongress, interparlamentariska unionen och Europarådets parlamentariska församling.
22.6.2005
FÖRSLAG TILL RESOLUTION
i enlighet med artikel 81 i arbetsordningen
från utskottet för miljö, folkhälsa och livsmedelssäkerhet
om kommissionens förslag till rådets beslut om anpassning till den tekniska utvecklingen av bilagan till Europaparlamentets och rådets direktiv 2002/95/EG av den 27 januari 2003 om begränsning av användningen av vissa farliga ämnen i elektriska och elektroniska produkter
Europaparlamentets resolution om kommissionens förslag till rådets beslut om anpassning till den tekniska utvecklingen av bilagan till Europaparlamentets och rådets direktiv 2002/95/EG av den 27 januari 2003 om begränsning av användningen av vissa farliga ämnen i elektriska och elektroniska produkter
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till rådets beslut om anpassning till den tekniska utvecklingen av bilagan till EUT L 37, 13.2.2003, s.
19. av den 27 januari 2003 om begränsning av användningen av vissa farliga ämnen i elektriska och elektroniska produkter (KOM-AC_DR(2005)CMT-2005-1948-2),
–
–
–
med beaktande av artikel 81 i arbetsordningen, och av följande skäl:
A.
I artikel 4.1 i direktiv 2002/95/EG begränsas användningen av vissa farliga ämnen i nya elektriska och elektroniska produkter som släpps ut på marknaden från och med den 1 juli 2006, om inte undantag medges i bilagan.
B.
C.
23. .
D.
E.
Kommissionen hävdar i skäl 2 i förslaget till beslut att vissa material och komponenter som innehåller vissa farliga ämnen bör undantas från förbudet, eftersom ”det fortfarande inte är praktiskt möjligt att bortskaffa eller ersätta nämnda farliga ämnen i dessa material och komponenter”.
F.
Kommissionen hävdar i skäl 3 att eftersom ”riskbedömningen av dekabromdifenyleter (...) har visat att det i dagsläget inte behövs några fler åtgärder för att minska riskerna för konsumenterna (...) kan dekaBDE undantas från bestämmelserna i artikel 4.1 i direktiv 2002/95/EG”.
Ändringar av detta slag kräver ett lagstiftningsförslag i den bemärkelse som avses i artikel 251 i fördraget.
G.
H.
I.
1.
2.
Europaparlamentet uppmanar rådet att motsätta sig förslaget, såvida inte kommissionen ändrar det genom att dra tillbaka inslaget om dekaBDE.
3.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet och kommissionen och till medlemsstaternas regeringar och parlament.
i enlighet med artikel 113 i arbetsordningen
från Cristiana Muscardini
om EU:s energipolitik
Europaparlamentet utfärdar denna resolution
–
med beaktande av artikel 113 i arbetsordningen,
A.
B.
Det är omöjligt att styra klimatförändringarna.
C.
D.
1.
Europaparlamentet uppmanar kommissionen och rådet att se till att medlemsstaterna blir skyldiga att snarast möjligt ta alla tänkbara initiativ för att öka den europeiska energiproduktionen.
2.
Europaparlamentet uppmanar kommissionen och rådet att införa sanktionsåtgärder mot de stater som inte agerar i tid.
3.
Europaparlamentet uppmanar kommissionen och rådet att se till att även finansministrarna deltar i sammanträden om energi och klimatförändringar.
7.6.2006
FÖRSLAG TILL RESOLUTION
till följd av fråga för muntligt besvarande B6‑…/…
från Raül Romeva i Rueda
för utskottet för utrikesfrågor
om eldhandvapen och lätta vapen, inför konferensen 2006 för översyn av Förenta nationernas handlingsprogram för att förebygga, motverka och avskaffa olaglig handel med eldhandvapen och lätta vapen i alla avseenden, och i riktning mot att utarbeta ett internationellt vapenhandelsfördrag
Europaparlamentets resolution om eldhandvapen och lätta vapen, inför konferensen 2006 för översyn av Förenta nationernas handlingsprogram för att förebygga, motverka och avskaffa olaglig handel med eldhandvapen och lätta vapen i alla avseenden, och i riktning mot att utarbeta ett internationellt vapenhandelsfördrag
Europaparlamentet utfärdar denna resolution
–
med beaktande av sina resolutioner av den 15 mars 2001 EGT C 343, 5.12.2001, s.
–
med beaktande av sin tidigare resolution av den 17 november 2005 P6_TA(2005)0436 . om rådets sjätte årliga rapport enligt tillämpningsbestämmelse 8 i Europeiska unionens uppförandekod för vapenexport (2005/2013(INI)),
–
–
med beaktande av slutsatserna från mötet med rådet för allmänna frågor och yttre förbindelser den 3 oktober 2005, där man gav uttryck för EU:s stöd för att internationell vapenhandel skall ske inom FN:s ramar, vilket skulle medföra bindande gemensamma normer för den världsomspännande handeln med konventionella vapen Europeiska unionens råd, 2678:e mötet med rådet (allmänna frågor) i Luxemburg den 3 oktober 2005. ,
–
med beaktande av Förenta nationernas handlingsprogram för att förebygga, motverka och avskaffa olaglig handel med SALW i alla avseenden, som antogs i juli 2001,
–
med beaktande av FN:s andra mellanstatliga tvåårsmöte för överläggningar om genomförandet av FN:s handlingsprogram för att förebygga, motverka och avskaffa olaglig handel med SALW i alla avseenden, som hölls den 11-15 juli 2005,
–
med beaktande av att FN:s generalförsamling i december 2005 antog ett internationellt instrument som skall ge staterna möjlighet att i rätt tid och pålitligt upptäcka och spåra olagliga SALW Beslut A/60/463 (L.55), den 8 december 2005. ,
–
med beaktande av att protokollet från 2001 om olaglig tillverkning av och handel med skjutvapen, delar och komponenter till dessa och ammunition trädde i kraft den 6 juli 2005 Protokollet är känt under benämningen ”FN:s protokoll om skjutvapen” och antogs i maj 2001 genom generalförsamlingens resolution 55/255. ,
–
med beaktande av FN:s översynskonferens om organisationens handlingsprogram, som enligt planerna skall äga rum mellan den 26 juni och den 7 juli 2006, och behovet av att se till att denna konferens och dess uppföljning blir lyckade,
–
A.
Det är välkommet att det internationella stödet ökar för ett rättsligt bindande internationellt vapenhandelsfördrag som förbjuder transaktioner som riskerar att undergräva de mänskliga rättigheterna eller den internationella humanitära rätten eller som hotar stabiliteten i länder eller regioner som sannolikt kommer att bidra till att väpnade konflikter bryter ut eller trappas upp.
B.
C.
D.
E.
Tiden är mogen för att det internationella samfundet skall ta itu med spridning och missbruk av SALW med hjälp av bindande internationella normer som grundas på allomfattande respekt för internationell rätt, inklusive mänskliga rättigheter och internationell humanitär rätt.
F.
G.
Det är beklagligt att FN:s breda samråd om att bekämpa olaglig förmedlingsverksamhet med SALW gjort så få framsteg samt att det saknas vilja att förhandla om ett rättsligt bindande internationellt instrument om vapenförmedling.
H.
FN:s handlingsprogram ålägger staterna att bedöma ansökningar om exporttillstånd i enlighet med stränga nationella bestämmelser och förfaranden som täcker alla SALW och överensstämmer med staternas befintliga ansvar och berörd internationell rätt och som särskilt beaktar risken för att dessa vapen skall dirigeras om till den olagliga handeln.
I.
Strategier för minskning och kontroll av SALW måste på ett lämpligt sätt integreras och bli en väsentlig del av internationella program för konfliktförebyggande verksamhet och fredsbyggande efter konflikter.
J.
De pågående kampanjinsatserna från civilsamhällets sida välkomnas och stöds.
1.
Europaparlamentet uppmanar de stater som är parter i konferensen 2006 om översyn av FN:s handlingsprogram att komma överens om en uppsättning övergripande principer om vapentransaktioner, i överensstämmelse med deras befintliga ansvar i enlighet med internationell, regional och nationell lagstiftning, inbegripet ett krav på att inte sända vapen som sannolikt kommer att bidra till kränkningar av de mänskliga rättigheterna och brott mot mänskligheten eller som främjar regional eller nationell instabilitet och väpnade konflikter.
2.
Europaparlamentet uppmanar det internationella samfundet att påbörja förhandlingar om ett internationellt fördrag om vapenhandel inom FN:s ramar omedelbart efter översynskonferensen 2006 om FN:s handlingsprogram, i syfte att upprätta ett rättsligt bindande instrument för att reglera vapentransaktioner i enlighet med definitionen i föregående punkt.
3.
4.
Europaparlamentet betonar att de skyldigheter som redan existerar i enlighet med internationell rätt när det gäller vapentransaktioner, särskilt sådana som omfattar kriterier för mänskliga rättigheter och humanitär rätt, bör kodifieras.
5.
Europaparlamentet uppmanar alla stater som undertecknat FN-protokollet om skjutvapen att utan dröjsmål ratificera protokollet och införliva det med nationell lagstiftning.
6.
Europaparlamentet uppmanar alla stater att se till att brott mot vapenembargon (inklusive ekonomiskt eller logistiskt stöd) definieras som brott i nationell lagstiftning.
7.
Europaparlamentet understryker att reformer som syftar till att förbättra de väpnade styrkornas funktionssätt, öppenhet och ansvarsskyldighet, och även brottsbekämpande myndigheter och straffrättsliga system, kan bidra till en trygg miljö där medborgarna inte längre känner behov av att äga vapen.
8.
9.
Europaparlamentet uppmanar alla stater att med sin nationella lagstiftning införliva uppförandekoden för personal vid brottsbekämpande myndigheter Uppförandekod för personal vid brottsbekämpande myndigheter, antagen genom generalförsamlingens resolution 34/169 av den 17 december 1979. och de grundläggande principerna för sådan personals användning av våld och skjutvapen Grundläggande principer för användning av våld och skjutvapen genom personal vid brottsbekämpande myndigheter, antagna av FN:s åttonde kongress om förebyggande av brott och behandling av gärningsmän i Havanna på Kuba den 27 augusti – 7 september 1990. .
10.
Europaparlamentet rekommenderar mycket starkt att regeringarna
a) bör förbjuda att civilpersoner utan tillstånd innehar och använder SALW och automatiska och halvautomatiska gevär och kulsprutor,
b) bör utveckla program för information och utbyte mellan stater som önskar samarbeta i frågor som rör kontroll av civilpersoners innehav av SALW,
c) bör ta upp frågan om att minska den överdrivna och inte önskvärda efterfrågan efter SALW i samhället och att de därför bör främja program och åtgärder för att minska denna efterfrågan och förebygga eller minska våld och osäkerhet i städerna och på landsbygden samt koncentrera sig på grupper som är särskilt utsatta för våld som hänger samman med SALW.
11.
Europaparlamentet uppmanar särskilt staterna att utveckla nationell lagstiftning för systematisk genomgång och licensiering av SALW och automatiska och halvautomatiska kulsprutor och att förhindra att vapen skaffas av personer som har ett våldsamt förflutet, särskilt våld i hemmet, eller har begått vapenhandelsbrott eller brott mot bestämmelser för vapenkontroll.
12.
Europaparlamentet uppmanar de stater som är parter i FN:s handlingsprogram och som kommer att bli parter i det framtida vapenhandelsfördraget att utveckla program för tekniskt stöd för att hjälpa tredjelandsorganisationer eller regionala organisationer som önskar utveckla lagstiftningskontroll för att reglera vapenhandeln.
13.
Europaparlamentet uppmanar de stater som är parter i FN:s handlingsprogram och som kommer att bli parter i det framtida vapenhandelsfördraget att inrätta rapporterings- och övervakningsförfaranden för att stödja staterna när de genomför sina åtaganden.
14.
Europaparlamentet uppmanar EU:s delegation att försvara principerna och rekommendationerna i denna resolution vid FN:s översynskonferens om organisationens handlingsprogram, som enligt planernas skall hållas mellan den 26 juni och den 7 juli 2006.
15.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, regeringarna och parlamenten i medlemsstaterna, FN:s generalsekreterare, det parlamentariska forumet om SALW och Interparlamentariska unionens församling.
i enlighet med artikel 174 i arbetsordningen
från talmanskonferensen
om antal ledamöter i utskotten
Beslut om antal ledamöter i utskotten
Europaparlamentet fattar detta beslut
–
med beaktande av artikel 174 i arbetsordningen,
–
med beaktande av sitt beslut av den 21 juli 2004 om antal ledamöter i utskotten Antagna texter av den 21 juli 2004, P6_TA(2004)0001 . .
1.
Europaparlamentet beslutar att från och med den 1 januari 2007 ändra antalet ledamöter i utskotten enligt följande:
CO1 – Utskottet för utrikesfrågor: 86 ledamöter
CO2 – Utskottet för utveckling: 36 ledamöter
CO3 – Utskottet för internationell handel: 33 ledamöter
CO4 – Budgetutskottet: 50 ledamöter
CO5 – Budgetkontrollutskottet: 40 ledamöter
CO6 – Utskottet för ekonomi och valutafrågor: 51 ledamöter
CO7 – Utskottet för sysselsättning och sociala frågor: 52 ledamöter
CO8 – Utskottet för miljö, folkhälsa och livsmedelssäkerhet: 68 ledamöter
CO9 – Utskottet för industrifrågor, forskning och energi: 54 ledamöter
C10 – Utskottet för den inre marknaden och konsumentskydd: 44 ledamöter
C11 – Utskottet för transport och turism: 52 ledamöter
C12 – Utskottet för regional utveckling: 57 ledamöter
C13 – Utskottet för jordbruk och landsbygdens utveckling: 47 ledamöter
C14 – Fiskeriutskottet: 40 ledamöter
C15 – Utskottet för kultur och utbildning: 38 ledamöter
C16 – Utskottet för rättsliga frågor: 28 ledamöter
C17 – Utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor: 60 ledamöter
C18 – Utskottet för konstitutionella frågor: 28 ledamöter
C19 – Utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män: 40 ledamöter
C20 – Utskottet för framställningar: 40 ledamöter
2.
Europaparlamentet beslutar att från och med den 1 januari 2007 ändra antalet ledamöter i underutskotten enligt följande:
SCO1A – Underutskottet för mänskliga rättigheter: 36 ledamöter
SCO1B – Underutskottet för säkerhet och försvar: 36 ledamöter
FÖRSLAG TILL RESOLUTION
till följd av uttalandena av rådet och kommissionen
från Marco Pannella och Marco Cappato
för ALDE-gruppen
om initiativet för ett allmänt moratorium för dödsstraff
Europaparlamentet utfärdar denna resolution
–
med beaktande av sina tidigare resolutioner om ett allmänt moratorium för dödsstraff och framför allt den resolution som antogs den 23 oktober 2003,
–
med beaktande av de resolutioner om ett moratorium för avrättningar som antagits av olika FN-organ, bland annat kommissionen för mänskliga rättigheter,
–
med beaktande av EU:s uttalanden till stöd för ett allmänt moratorium för dödsstraff,
–
med beaktande av sin skriftliga förklaring om dödsstraffet: om ett allmänt moratorium för avrättningar i syfte att uppnå ett totalt avskaffande,
–
A.
EU beslutade i sina riktlinjer för politiken gentemot tredje land i fråga om dödsstraff som Europeiska rådet antog i Luxemburg den 6 juni 1998 att inom internationella organisationer verka för ett allmänt moratorium för dödsstraff och inom rimlig tid ett avskaffande av dödsstraffet.
B.
C.
Den 27 juli 2006 antog den italienska deputeradekammaren enhälligt ett förslag där man krävde att den italienska regeringen, efter samråd med sina samarbetspartner i EU men utan krav på enhällighet, vid FN:s nästa generalförsamling lägger fram ett förslag till resolution om ett allmänt moratorium för dödsstraff i syfte att uppnå att dödsstraffet helt avskaffas i världen.
D.
Den 9 januari 2007 beslutade den italienska regeringen och Europarådet att gemensamt försöka samla så mycket stöd som möjligt för ett initiativ i FN:s generalförsamling för ett allmänt moratorium för dödsstraff i syfte att helt avskaffa dödsstraffet.
E.
Den 22 januari 2007 beslutade rådet (allmänna frågor och yttre förbindelser) att Tyskland som ordförandeland för EU i New York skulle undersöka möjligheterna för en förnyad debatt och förutsättningarna för förhandlingar om förslaget om ett allmänt moratorium för dödsstraff.
1.
Europaparlamentet stöder aktivt den italienska deputeradekammaren och regeringens initiativ som även har rådets, kommissionens och Europarådets stöd.
2.
Europaparlamentet upprepar sin uppmaning till rådets ordförandeskap att snarast börja arbeta med ett resolutionsförslag om ett allmänt moratorium för avrättningar som skall läggas fram för FN:s generalförsamling.
3.
Europaparlamentet uppmanar alla EU:s institutioner och medlemsstaterna att politiskt och diplomatiskt göra allt för att denna resolution skall antas av den pågående generalförsamlingen.
4.
Europaparlamentet uppmanar rådets ordförandeskap och kommissionen att för parlamentet redovisa de resultat som uppnås under den pågående generalförsamlingen.
5.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådets ordförandeskap, kommissionen, medlemsstaternas parlament, FN:s generalsekreterare samt alla länder som har företrädare i FN:s generalförsamling.
till följd av uttalandena av rådet och kommissionen
från Thierry Cornillet, Philippe Morillon, Marielle De Sarnez och Marios Matsakis
för ALDE-gruppen
om den humanitära situationen i Darfur
Europaparlamentets resolution om den humanitära situationen i Darfur
Europaparlamentet utfärdar denna resolution
-
med beaktande av sina tidigare resolutioner om situationen i Darfur, särskilt resolutionerna antagna den 16 september 2004, 23 juni 2005, 6 april 2006 och 28 september 2006,
-
med beaktande av begreppet ”ansvar att skydda” som FN har beslutat att tillämpa, vilket innebär att när nationella myndigheter uppenbarligen underlåter att skydda sin befolkning mot folkmord, krigsförbrytelser, etnisk rensning och brott mot mänskligheten kan FN:s säkerhetsråd besluta att skicka militära styrkor i enlighet med kapitel VII i FN-stadgan,
-
med beaktande av säkerhetsrådets resolutioner om Sudan, särskilt resolution 1706 om att placera en ny fredsbevarande styrka i Darfur,
-
med beaktande av FN:s konvention om barnets rättigheter som är bindande och inte medger några undantag,
-
med beaktande av att Desmond Tutu, 1983 års mottagare av Nobels fredspris, krävt en betydande FN-styrka med ett effektivt mandat för att skydda civilbefolkningen i Darfur, och av följande skäl:
A.
Det är oerhört tragiskt att konflikten i Darfurregionen mellan reguljära styrkor, regeringsstödd milis och rebeller har krävt minst 400 000 dödsoffer och drivit över 2,5 miljoner människor på flykt de senaste tre åren, trots att ett fredsavtal för Darfur undertecknades i Abuja i Nigeria den 5 maj 2006.
B.
Enligt FN:s observatörer har de 2,5 miljonerna flyktingar och fördrivna inte längre tillgång till hjälp från internationella organisationer och dör av undernäring och sjukdomar.
C.
Många hjälporganisationer har tvingats lämna Darfur därför att biståndsarbetarnas personliga säkerhet är hotad.
D.
Den rådande situationen i Darfur destabiliserar allvarligt hela regionen och leder till humanitära katastrofer i Tchad och Centralafrikanska republiken.
E.
Antalet offer ökar för varje dag och en internationell insats blir alltmer nödvändig.
1.
Europaparlamentet kräver att regeringarna i EU:s medlemsstater, rådet och kommissionen tar sitt ansvar och gör allt för att verkligen skydda befolkningen i Darfur från en humanitär katastrof.
2.
3.
Europaparlamentet kräver att ett flygförbud införs över hela Darfur, med undantag endast för flyg med hjälpsändningar.
4.
Europaparlamentet uppmanar rådet och kommissionen att arbeta för att skapa förutsättningar för att politiska förhandlingar återupptas mellan alla parter i konflikten, något som kan göra det möjligt för flyktingar och fördrivna att återvända till sina byar och hemtrakter på ett säkert sätt.
5.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, medlemsstaternas regeringar och parlament, Afrikanska unionens generalsekreterare, Arabförbundets generalsekreterare, FN:s generalsekreterare och FN:s säkerhetsråd.
från Martine Roure
för PSE-gruppen
om bekämpande av rasism och främlingsfientlighet
Europaparlamentets rekommendation till rådet om bekämpande av rasism och främlingsfientlighet
Europaparlamentet utfärdar denna rekommendation
–
med beaktande av sitt betänkande av den 4 juli 2002 Betänkande Ceyhun – T5-363/2002, EUT C 271 E, 12.11.2003, s.
379. ,
–
med beaktande av den gemensamma åtgärden 96/443/RIF om åtgärder mot rasism och främlingsfientlighet,
–
med beaktande av rådets rambeslut om kommissionens bekämpande av rasism och främlingsfientlighet (KOM(2001)0664) EGT C 75 E, 26.3.2002, s.
269. ,
–
A.
B.
C.
Trots flera års förhandlingar inom rådet har man ännu inte lyckats nå någon överenskommelse om detta förslag till rambeslut.
D.
Det tyska ordförandeskapet har markerat att det avser att återuppta förhandlingarna om rambeslutet om bekämpande av rasism och att det betraktar antagandet av detta rambeslut som en prioriterad fråga.
E.
Den text som nu diskuteras är resultatet av flera års förhandlingar och bör ligga till grund för utarbetandet av en mer omfattande europeisk lagstiftning på detta område.
F.
G.
1.
Europaparlamentet riktar följande rekommendation till rådet:
a) avge ett starkt politiskt budskap för ett medborgarnas Europa och säkerställa ett gott skydd för de grundläggande rättigheterna genom att anta detta rambeslut,
b) säkerställa att rambeslutet ger ett europeiskt mervärde i förhållande till den gemensamma åtgärden från 1996,
c) tydligare definiera undantagen och möjligheterna att undanta vissa gärningar från straffrättsligt ansvar,
d) bibehålla möjligheten till undantag från principen om dubbel straffbarhet i syfte att möjliggöra ömsesidig rättslig hjälp mellan medlemsstater i samband med väckandet av åtal på grund av rasistiska och främlingsfientliga gärningar,
e) inbegripa en bestämmelse om icke-försämring, så att genomförandet av rambeslutet inte kan leda till att det befintliga skyddet försvagas,
f) inrätta en komplett rättslig ram för bekämpandet av rasism och främlingsfientlighet genom att möjliggöra ett snabbt antagande av ett områdesöverskridande direktiv om bekämpande av diskriminering i enlighet med artikel 13 i EG-fördraget samt besluta om effektiva, proportionerliga och avskräckande straffrättsliga påföljder.
2.
Europaparlamentet uppdrar åt talmannen att översända denna rekommendation till rådet och, för kännedom, till kommissionen och till medlemsstaternas parlament och regeringar.
till följd av uttalandena av Europeiska rådet och kommissionen
från Jan Marinus Wiersma, Hannes Swoboda, Reino Paasilinna och Panagiotis Beglitis
för PSE-gruppen
om toppmötet mellan EU och Ryssland
Europaparlamentets resolution om toppmötet mellan EU och Ryssland
Europaparlamentet utfärdar denna resolution
–
med beaktande av partnerskaps- och samarbetsavtalet mellan Europeiska gemenskaperna och deras medlemsstater som den ena parten och Ryska federationen som den andra parten, vilket trädde i kraft 1997 och upphör att gälla 2007,
–
med beaktande av människorättsdialogen mellan EU och Ryssland,
–
med beaktande av sina tidigare resolutioner om Ryssland och särskilt resolutionen av den 26 maj 2005 om förbindelserna mellan EU och Ryssland EUT C 117 E, 18.5.2006, s.
235. ,
–
med beaktande av sin resolution av 13 december 2006 om toppmötet mellan EU och Ryssland Antagna texter, P6_TA(2006)0566 . ,
–
A.
Förbindelserna mellan EU och Ryssland har vuxit sig allt starkare under de senaste åren och lett till en djup och omfattande ekonomisk integration och ett ömsesidigt beroende som kommer att öka ännu mer under den närmaste framtiden.
B.
Ett ökat samarbete och goda grannförbindelser mellan EU och Ryssland är av avgörande betydelse för stabiliteten, säkerheten och välfärden i hela Europa och dess grannländer.
C.
Ett avtal om strategiskt partnerskap mellan EU och Ryska federationen är avgörande för detta ökade samarbete, särskilt när det gäller att vidareutveckla de ekonomiska förbindelserna i en anda av jämlikhet, öppenhet och respekt för internationellt erkända förfaranden, att stärka säkerheten och stabiliteten i Europa genom att hitta fredliga politiska lösningar på regionala konflikter i det gemensamma grannskapet samt att ytterligare stärka respekten för mänskliga rättigheter och rättsstatsprincipen liksom den demokratiska ramen för dessa förbindelser.
D.
Ett skyndsamt genomförande av de fyra gemensamma områdena, dvs. ett gemensamt ekonomiskt område, ett område för frihet, säkerhet och rättvisa, ett område för yttre säkerhet och ett område för forskning, utbildning och kultur bör stå i centrum i förhandlingarna om det nya strategiska partnerskapsavtalet.
E.
Ett framtida avtal mellan EU och Ryska federationen bör innehålla de principer i energistadgan som syftar till att stärka banden och minska EU:s oro för att Ryssland använder sina stora energitillgångar som ett politiskt vapen.
F.
Litauen hotar att blockera ett energiavtal mellan EU och Ryska federationen på grund av att den ryska oljeledningen Druzhbas anknytning till Litauens raffinaderi Mazeikiu Nafta varit stängd sedan juni 2006 efter det att Rysslands oljeledningsoperatör Transneft anklagats för att avsiktligt fördröja reparationer av oljeläckor.
G.
H.
EU och Ryssland diskuterar att inrätta en jourtelefon vid energikriser som skall göra det möjligt för befattningshavare i Bryssel och Moskva att genast kontakta varandra för att förhindra eventuella avbrott i olje- och gasförsörjningen till följd av politiska eller tekniska problem.
I.
Ett nytt ramavtal mellan EU och Ryssland, som skall ersätta partnerskaps- och samarbetsavtalet som löper ut 2007 och som skall omfatta Bulgarien och Rumänien, skulle vara ett positivt bevis på att både EU och Ryssland vill ha en grund för ett fortsatt intensivt samarbete, i synnerhet när det gäller gemensamma intressen som energi och säkerhet.
J.
K.
Efter flera månaders förhandlingar mellan kommissionen, det tyska ordförandeskapet och Polen å ena sidan och Ryssland å andra sidan, förefaller Ryssland villigt att försöka bryta det politiska dödläget och nå fram till en kompromiss med EU, vilket gör att båda sidorna kan inleda förhandlingar om det nya ramavtalet.
L.
Det internationella samfundet hyser en ökad oro över hur mänskliga rättigheter och rättsstatsprincipen respekteras i Ryssland, framför allt yttrandefriheten och mötesfriheten.
M.
Både EU-medborgare som reser till Ryssland och ryska medborgare som försöker komma in i EU möts i dag av omfattande visumkontroller.
N.
USA:s planer på att placera ut ett antirobotsystem på europeisk mark i Polen och Tjeckien har upprört Ryssland och gett upphov till en het debatt om maktbalansen och en eventuell kapprustning.
1.
2.
3.
4.
5.
Europaparlamentet uppmanar Ryssland, som är medlem i FN, OSSE och Europarådet, att fullgöra sina skyldigheter när det gäller att fullt ut iaktta och respektera mänskliga rättigheter, församlingsfriheten och yttrandefriheten.
6.
Europaparlamentet uppmanar eftertryckligen kommissionen och rådet att även i fortsättningen övervaka den rådande situationen och utvecklingen framöver i Ryssland, och påminner om att en bredare debatt om situationen i Ryssland bör vara en prioriterad fråga hos rådet.
7.
Europaparlamentet understryker vikten av att samarbeta med Ryssland som en nödvändig strategisk partner för att trygga freden, stabiliteten och säkerheten och för att bekämpa internationell terrorism och våldsbenägen extremism samt att behandla andra säkerhetsproblem som rör miljö- och kärnkraftshot, narkotika, vapen- och människohandel och gränsöverskridande organiserad brottslighet inom det europeiska grannskapet i samarbete med OSSE och andra aktörer i internationella fora.
8.
9.
10.
11.
12.
13.
14.
15.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, medlemsstaternas regeringar och parlament samt Ryska federationens regering och parlament.
till följd av ett uttalande av kommissionen
från Cristiana Muscardini, Brian Crowley, Roberta Angelilli, Adam Bielan, Gintaras Didžiokas och Ryszard Czarnecki
för UEN-gruppen
om kampen mot den ökande extremismen i Europa
Europaparlamentets resolution om kampen mot den ökande extremismen i Europa
Europaparlamentet utfärdar denna resolution
–
med beaktande av de internationella människorättsinstrumenten, särskilt den internationella konventionen om avskaffande av alla former av rasdiskriminering och europeiska konventionen om skydd för de mänskliga rättigheterna och de grundläggande friheterna, som båda undertecknats av samtliga EU-medlemsstater och av ett stort antal tredjeländer,
–
med beaktande av artiklarna 6 och 7 i EU-fördraget och artikel 13 i EG-fördraget,
–
med beaktande av stadgan om de grundläggande rättigheterna och arbetsordningen för Europeiska unionens byrå för grundläggande rättigheter ,
–
med beaktande av sin lagstiftningsresolution av den 29 november 2007 om förslaget till rådets rambeslut om bekämpande av vissa former av och uttryck för rasism och främlingsfientlighet enligt strafflagstiftningen, Antagna texter: P6_TA-PROV(2007)0552 .
–
med beaktande av sina tidigare resolutioner om rasism, främlingsfientlighet och extremism,
–
A.
Rekryteringen av islamistiska fundamentalister och den våldsamma propagandakampanj som genomförs i form av bland annat terroristattacker i Europeiska unionen och som grundar sig på antisemitism och hat mot de europeiska värdena, är djupt oroväckande.
B.
Extremistiska rörelser och partier som grundar sin ideologi och sina politiska uttalanden, metoder och ageranden på intolerans, rasism och antisemitism håller återigen på att öka i antal, vilket är också oroväckande.
C.
Även den våldsamma verksamhet och de terroristattacker som genomförs av vänsterextremistiska rörelser som grundar sig på spridning av hat och klasskrig är oroväckande.
D.
Sådana ideologier är oförenliga med demokrati och mänskliga rättigheter och med de principer och värden som EU grundar sig på.
E.
Ingen medlemsstat kan bortse från de faktiska hot som extremismen utgör mot demokratin, och därför är det en utmaning för hela Europa att bekämpa spridningen av främlingsfientlighet och andra extremistiska politiska yttringar.
F.
Information om de rörelser och grupper som uppmuntrar till hat, attacker mot demokratiska institutioner, terroristattacker och annat våld kan framför allt hittas i vissa medier och på ett stort antal hemsidor på Internet.
1.
Europaparlamentet fördömer bestämt alla hatattacker, uppmanar de nationella myndigheterna att göra sitt yttersta för att straffa de skyldiga och för att bekämpa straffriheten i samband med sådana attacker, och uttalar sitt fulla stöd för alla som fallit offer för sådana attacker liksom deras familjer.
2.
Europaparlamentet påpekar att extremiströrelser som uppmuntrar till våld i vissa fall missbrukar föreningsfriheten ur politisk synvinkel.
Åtgärder som är avsedda att begränsa dessa rörelsers handlingsförmåga bör stå i proportion till den fara de utgör och med likställdhet och frihet för alla som klara målsättningar.
3.
Europaparlamentet uppmanar medlemsstaterna att ta itu med de sociala och ekonomiska problemen såsom arbetslöshet, invandring och säkerhet, som de extremistiska rörelserna drar nytta av, och att utveckla strategier för utbildning om ett demokratiskt medborgarskap som grundar sig på medborgerliga rättigheter och skyldigheter.
4.
Europaparlamentet uppmanar kommissionen och rådet att leda arbetet med att finna framför allt förebyggande politiska och juridiska lösningar och inte glömma bort viktiga frågor rörande utbildning för ungdomar och information till allmänheten, utbildning om totalitarism och kunskapsspridning om de mänskliga rättigheterna och de grundläggande friheterna för att se till att de handlingar och händelser som faktiskt har inträffat i Europa inte glöms bort.
5.
Europaparlamentet uppmanar kommissionen att kontrollera att gällande lagstiftning som är avsedd att förhindra uppmuntran till politiskt och religiöst våld verkligen tillämpas.
6.
Europaparlamentet uppmanar medierna att genom sin verksamhet främja och sprida principer och värden såsom demokrati, liberalism och tolerans.
7.
Europaparlamentet betonar behovet av en lösning på den skadliga Internetanvändningen och betonar att den Internetövervakning som avser att förhindra terroristattacker måste förhindra att Internet kan användas för att uppmuntra till terroristattacker.
8.
Europaparlamentet uppmanar kommissionen att stödja de icke-statliga organisationer och organisationer inom det civila samhället som arbetar för att främja demokratiska värderingar, solidaritet, social integrering, interkulturell dialog och social medvetenhet för att på sätt bekämpa radikalisering och våldsam extremism.
9.
Europaparlamentet uppmanar rådet och kommissionen att intensifiera de gemenskapsprogram som syftar till att främja social integrering och utbildning om ett demokratiskt medborgarskap och ta itu med sociala och ekonomiska problem som otrygghet, arbetslöshet och utslagning.
10.
21.4.2008
FÖRSLAG TILL RESOLUTION
till följd av uttalandena av rådet och kommissionen
från Frithjof Schmidt, Raül Romeva i Rueda och Hélène Flautre
för Verts/ALE-gruppen
om situationen i Burma
Europaparlamentets resolution om situationen i Burma
Europaparlamentet utfärdar denna resolution
–
med beaktande av sina resolutioner av den 14 december 2006 och den 21 juni 2007 om Burma,
–
med beaktande av rådets slutsatser av den 19 november 2007 om antagande av ytterligare restriktiva åtgärder mot Burma,
–
med beaktande av rådets förordning (EG) nr 194/2008 av den 25 februari 2008 om förlängning och skärpning av de restriktiva åtgärderna mot Burma och om upphävande av förordning (EG) nr 817/2006,
–
A.
Den burmesiska statens råd för fred och utveckling (SPDC) har efter fjorton års arbete förklarat att en folkomröstning om den nya konstitutionen kommer att hållas den 10 maj 2008 och följas upp av flerpartival 2010.
B.
Burmas regering har förkastat de förslag som lades fram av FN:s sändebud Ibrahim Gambari för att garantera ett fritt och rättvist genomförande av folkomröstningen i närvaro av internationella observatörer.
C.
D.
Sedan folkomröstningen tillkännagavs har regeringen i Burma antagit lag nr 1/2008, som förvägrar medlemmar av religiösa ordnar rösträtt samtidigt som den vidtagit olika åtgärder för att försäkra sig om att få majoriteten av rösterna i valet.
E.
Den största delen av den burmesiska oppositionen har beslutat att bojkotta folkomröstningen.
F.
De sanktioner som EU antagit gentemot den burmesiska regeringen har fram tills nu varit verkningslösa.
1.
Europaparlamentet beklagar djupt den totala avsaknaden av demokratisk legitimitet i samband med folkomröstningen om den nya konstitutionen, eftersom den burmesiska befolkningen har fråntagits alla grundläggande demokratiska rättigheter som skulle göra det möjligt att hålla en öppen debatt om konstitutionen, ändra den och därefter att fritt uttala sig genom folkomröstningen.
2.
Europaparlamentet fördömer den burmesiska regeringens förkastande av de förslag som lagts fram av FN:s särskilda sändebud Ibrahim Gambari för att möjliggöra en öppen och övergripande kampanj inför folkomröstningen om konstitutionen.
3.
Europaparlamentet anser att en hållbar utveckling i Burma, som skapar ett stabilt klimat på lång sikt, enbart kan åstadkommas genom en övergripande process med nationell försoning och dialog samt respekt för de demokratiska värderingarna, mänskliga rättigheter och rättsstatsprincipen.
4.
Europaparlamentet uppmanar regeringen i Burma att tillsätta en oberoende valkommission, se till att ett korrekt röstregister upprättas, häva de långvariga restriktionerna för medierna, tillåta förenings-, yttrande- och mötesfrihet i Burma, annullera de nya förordningarna som kriminaliserar legitima debatter om folkomröstningen och acceptera internationella observatörers närvaro.
5.
Europaparlamentet kräver ett omedelbart och ovillkorligt frisläppande av politiska motståndare till regimen och mer än 1 800 politiska fångar, bland annat Aung San Suu Kyi, ledarna för 88-generationens studentrörelse och ledarna för shanfolkens förbund för demokrati (Shan Nationalities League for Democracy), som fängslades 2005.
6.
Europaparlamentet kräver att man utreder alla dödsfall och fall av personer som saknas sedan kraftåtgärderna i september 2007 mot demonstrerande buddhistiska munkar och demokratiaktivister, och kartlägger var saknade munkar och nunnor befinner sig.
7.
8.
Europaparlamentet uppmanar rådet, kommissionen och medlemsstaterna att engagera Kina, i dess egenskap av medlem av FN:s säkerhetsråd och part i det frivilliga protokollet till FN:s konvention om barnets rättigheter om barns indragning i väpnade konflikter, i att säkerställa att Burma gör verkliga framsteg när det gäller att förhindra brott mot barns rättigheter i samband med väpnade konflikter.
9.
10.
Europaparlamentet stödjer ett aktivt engagemang i och tillträde till Burma genom den särskilde rapportören och andra företrädare för berörda människorättsmekanismer.
11.
12.
13.
14.
Europaparlamentet uppmanar rådet att se till att riktade sanktioner tillämpas på ett effektivt sätt och att ingående utreda vem sanktionerna ska riktas mot samt möjliggöra omprövning av beslut och pågående övervakning samt säkerställa att åtgärder som beslutats även tillämpas.
15.
Europaparlamentet uppmanar rådet att fortsätta att se över sanktionerna med utgångspunkt i specifika riktmärken för mänskliga rättigheter som måste omfatta följande punkter: frigivandet av politiska fångar och alla andra personer som godtyckligt fängslats för att de utövat sina grundläggande mänskliga rättigheter, med andra ord yttrande-, mötes- och föreningsfrihet, en korrekt officiell rapport om antalet personer som dödats, arresterats och häktats av säkerhetsstyrkorna (bland annat under den senaste tidens kraftåtgärder), var och i vilken situation dessa personer befinner sig; upphörande av militära angrepp mot civila, och en övergång till demokrati.
16.
17.
18.
Europaparlamentet uppmanar EU och övriga västländer att erbjuda incitament för reformer som en motvikt till hotet och/eller införandet av sanktioner som på ett positivt sätt kan motivera militären att införa förändringar.
19.
20.
Europaparlamentet uppmanar rådet och kommissionen att stärka stödet till människorättsaktivister och medlemmar av oppositionen i Burma.
21.
22.
Europaparlamentet uppmanar kommissionen att upprätta och utvidga biståndsprogram som syftar till att stärka grupper, såsom kvinnor och etniska och religiösa minoriteter, som har berövats sin rösträtt, och att avhjälpa politiska, etniska, religiösa och andra splittringar.
23.
Europaparlamentet uppmanar kommissionen att öka stödet för burmeser som lever utomlands genom programmet för fördrivna personer inom ramen för instrumentet för utvecklingssamarbete, och att överväga andra stödmöjligheter.
24.
Europaparlamentet betonar att det stöd som ges måste vara kopplat till riktmärken och tidsfrister för att bl.a. bättre kontrollera korruptionsriskerna.
25.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, medlemsstaternas regeringar och parlament, Aseanländernas regeringar och parlament, Nationella demokratiförbundet (NLD) i Burma, Statens råd för fred och utveckling (SPDC) i Burma, Kinas, Indiens och Rysslands regeringar och parlament och FN:s generalsekreterare.
till följd av uttalandena av rådet och kommissionen
från Vittorio Agnoletto
för GUE/NGL-gruppen
om det nionde toppmötet mellan EU och Indien (i Marseille den 29 september 2008)
Europaparlamentets resolution om det nionde toppmötet mellan EU och Indien (i Marseille den 29 september 2008)
Europaparlamentet utfärdar denna resolution
–
med beaktande av det nionde toppmötet mellan EU och Indien som kommer att hållas i Marseille den 29 september 2008,
–
med beaktande av avtalet från 2004 om ett strategiskt partnerskap mellan EU och Indien (KOM(2004)0430),
–
med beaktande av EU:s och Indiens gemensamma handlingsplan som antogs vid det sjätte toppmötet mellan EU och Indien i New Delhi den 7 september 2005,
–
med beaktande av förslaget om att förhandla om ett partnerskaps- och samarbetsavtal med Indien,
–
A.
Dagordningen för det kommande ”Marseilletoppmötet” mellan EU och Indien kommer sannolikt att domineras av översynen av den gemensamma handlingsplanen från 2005, klimatförändringarna, fred och säkerhet, utbildning, hälsa och livsmedelssäkerhet.
B.
Detta toppmöte bör inleda en ny fas i förbindelserna mellan EU och Indien och underlätta diskussionen om regionala frågor som är av gemensamt intresse för EU och Indien.
1.
2.
3.
4.
Europaparlamentet oroar sig över det för närvarande ostadiga politiska läget i Pakistan och det alltmer osäkra läget i Afghanistan och Sri Lanka och uttrycker sin förhoppning om att Indien som det dominerande landet i regionen kommer att främja stabilitet och fred.
5.
6.
7.
Europaparlamentet uppmanar med kraft Indiens regering att fortsätta samarbetet med relevanta FN-människorättsorgan i syfte att effektivt utrota diskriminering på grundval av kast, ett samarbete som bör omfatta kommittén för avskaffande av rasdiskriminering och FN:s särskilda rapportörer med uppdrag att utveckla principer och riktlinjer för att avskaffa diskriminering på grundval av arbete och ursprung.
8.
9.
Europaparlamentet uppmanar Indiens regering att vara särskilt vaksam mot uppkomsten av etniska, religiösa och kulturella spänningar mellan olika grupper, som skulle äventyra landets sekulära arv som präglas av tolerans och samlevnad.
10.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till kommissionen, rådet och Indiens regering och parlament.
till följd av ett uttalande av kommissionen
från Cristiana Muscardini, Adam Bielan, Roberta Angelilli, Mario Borghezio och Antonio Mussa
för UEN-gruppen
om bilindustrins framtid
Europaparlamentets resolution om bilindustrins framtid
Europaparlamentet utfärdar denna resolution
–
med beaktande av slutsatserna från högnivågruppen CARS 21 av den 12 december 2005,
–
med beaktande av sin resolution av den 15 januari 2008 om CARS 21: Ett konkurrenskraftigt motorfordonsregelverk (2007/2120(INI)),
–
med beaktande av ordförandeskapets slutsatser från Europeiska rådet i Bryssel den 15‑16 oktober 2008,
–
med beaktande av kommissionens meddelande av den 29 oktober 2008 med titeln ”Från finanskris till återhämtning: ram för åtgärder på EU-nivå” (KOM(2008)0706),
–
med beaktande av kommissionens meddelande av den 26 november 2008 till Europeiska rådet med titeln ”En ekonomisk återhämtningsplan för Europa” (KOM(2008)0800),
–
med beaktande av rådets (konkurrenskraft) slutsatser av den 5 och 6 mars 2009 om bilindustrin,
–
A.
B.
C.
Bilindustrin är också en mycket viktig arbetsgivare i fråga om kvalificerad arbetskraft, och en central drivkraft för kunskap och innovation, i det att den varje år investerar mer än 20 miljarder euro i forskning och utveckling.
D.
E.
Bilindustrin har nära kopplingar till många andra industrisektorer, och ett stort antal underentreprenörer och leverantörer utgörs av små och medelstora företag, vilka drabbas av finanskrisen i lika hög grad, det vill säga mycket hårt, och med en mycket högre arbetslöshetsrisk.
F.
I en marknadsekonomi är det de enskilda företagen som i första hand måste hantera en kris, men i vissa specifika undantagsfall är ett ingripande av den offentliga sektorn i enlighet med befintliga stadsstödsregler motiverat och till och med nödvändigt, när det gäller en sektor som före finanskrisen var en mycket viktig del av EU:s ekonomi och samhälle.
G.
Vissa medlemsstater har börjat vidta nationella åtgärder för att stödja industrin, vilket har påverkat efterfrågan på bilar positivt.
H.
Medlemsstaternas åtgärdsprogram har granskats av kommissionen, som kunnat konstatera att de är fullständigt förenliga med motsvarande åtgärder som vidtagits på gemenskapsnivå och överensstämmer med bestämmelserna om statligt stöd.
I.
Kommissionen förhandlar just nu om ytterligare avregleringar av handeln inom ramen för Doharundan och i form av nya frihandelsavtal, särskilt i form av det nya frihandelsavtalet med Sydkorea som har direkt inverkan på bilsektorn.
J.
En återgång till kraftiga protektionistiska åtgärder är inte det bästa sättet att lösa den nuvarande finansiella och ekonomiska krisen, eftersom det skulle leda till motåtgärder från konkurrenterna på världsmarknaden och därmed till en destruktiv uppbromsning av världshandeln.
1.
Europaparlamentet anser att det enda sättet att ta itu med och komma till rätta med bilsektorns problem är att man på gemenskapsnivå vidtar samordnade politiska åtgärder med fullt deltagande av sektorns största aktörer på både utbuds- och efterfrågesidan.
2.
Europaparlamentet anser att ett sådant ekonomiskt stödprogram bör baseras på
a) att tillgången till krediter säkras för biltillverkare och leverantörer, varvid Europeiska investeringsbanken kan spela en viktig roll i nya återhämtningsprojekt,
b) att efterfrågan på bilar stimuleras, bland annat genom uppmuntran till att skrota gamla bilar och köpa miljövänliga bilar,
c) att samhällseffekterna av en eventuell omstrukturering dämpas och att kvalificerad arbetskraft bevaras genom att Europeiska fonden för justering av globaliseringseffekter och Europeiska specialfonden används fullt ut,
d) att särskilt stöd för forskning och investeringar tillhandahålls.
3.
4.
5.
Europaparlamentet understryker att bilindustrin också har ett ansvar för att vidta åtgärder för att lösa den pågående krisen och måste göra betydande insatser för att bidra till återhämtningen, samtidigt som man bör ta särskild hänsyn till arbetskraftens intressen och förväntningar i samband med användningen av statligt ekonomiskt stöd.
6.
Europaparlamentet betonar att det statliga ekonomiska stödet alltid måste överensstämma med EU:s bestämmelser om statligt stöd och principerna för den inre marknaden, vars fullständiga och effektiva funktion är en förutsättning för Europas återhämtning och framtida tillväxt.
7.
Europaparlamentet bekräftar ånyo att man måste fortsätta att göra omfattande investeringar i forskning och utveckling, i synnerhet på området för ren teknik som skulle kunna förbättra den europeiska industrins konkurrenskraft och bidra till att bekämpa klimatförändringar.
8.
9.
Europaparlamentet understryker att eftersom den globala krisen påverkar andra globala aktörer inom bilsektorn, särskilt Förenta staterna, måste en kontinuerlig dialog föras med tredjeländer och EU:s huvudsakliga handelspartner på multilateral och bilateral nivå för att man ska kunna komma fram till en övergripande lösning och undvika att protektionistiska och diskriminerande åtgärder som vidtas av tredjeländer drabbar EU:s industri på ett oförsvarligt sätt.
10.
Europaparlamentet uppmanar kommissionen att skjuta upp ingåendet av frihandelsavtalet mellan Europeiska unionen och Sydkorea till dess att man hittat en välbalanserad lösning beträffande konsekvenserna för bilsektorn.
11.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen och medlemsstaternas regeringar och parlament.
25.3.2009
FÖRSLAG TILL RESOLUTION
i enlighet med artikel 113 i arbetsordningen
från Cristiana Muscardini
om kriser, miljö och livskvalitet
Förslag till Europaparlamentets resolution om kriser, miljö och livskvalitet
Europaparlamentet utfärdar denna resolution
–
med beaktande av artikel 113 i arbetsordningen, och av följande skäl:
A.
Samtidigt med den allvarliga ekonomiska krisen, som leder till att miljontals arbetstillfällen går förlorade enbart inom EU, pågår en miljökris och en energikris.
B.
Det måste till nya produktionsmodeller som främjar utvecklingen men som inte skadar miljön eller utarmar planeten.
C.
Med den ökande urbaniseringen blir det allt viktigare att se till att återstående grönområden inte förstörs ytterligare, av omsorg för den ekologiska balansen.
D.
Många grönområden har gått förlorade på grund av bränder som varje år ödelägger miljontals hektar av vår mark och som samtidigt skadar klimatet.
E.
Dessvärre blir det allt vanligare med byggnader som respektlöst bryter mot omgivningens kulturella sammanhang och dess specifika landskapsbild.
F.
En överdriven urbanisering får omedelbara följder för livskvaliteten.
1.
Europaparlamentet uppmanar kommissionen och rådet att bedöma möjligheten att införa bestämmelser om att
a) begränsa markåtgången genom att utnyttja såväl obebyggda som övergivna områden på ett bättre sätt,
b) skydda miljön och landskapet av omsorg för människors fysiska och psykiska hälsa,
c) återplantera brandskadade skogar,
d) skapa nya grönområden nära städerna, och
e) främja en hållbar och ansvarsfull urbanisering.
till följd av uttalandena av rådet och kommissionen
från Gunnar Hökmark
för PPE-DE-gruppen
om resultatet av G20-mötet i London den 2 april 2009
Europaparlamentets resolution om resultatet av G20-mötet i London den 2 april 2009
Europaparlamentet utfärdar denna resolution
–
med beaktande av förklaringen om en global plan för återhämtning och reform från G20‑mötet den 2 april 2009,
–
med beaktande av förklaringen om stärkandet av det finansiella systemet från G20-mötet den 2 april 2009,
–
med beaktande av den handlingsplan som fastställdes i New York vid G20-mötet i september 2008,
–
med beaktande av OECD:s lista över länder som inte uppfyller de internationella standarderna för utbyte av skatteinformation som publicerades den 2 april 2009,
–
med beaktande av Eurogruppens stats- och regeringschefers möte den 12 oktober 2008, vars syfte var att anta en samordnad räddningsplan för att bekämpa den ekonomiska krisen,
–
med beaktande av den rapport från högnivåexpertgruppen för den finansiella tillsynen i EU, med Jacques de Larosières som ordförande, som lämnades till kommissionen den 25 februari 2009 inför Europeiska rådets vårmöte 2009,
–
med beaktande av sin resolution av den 11 mars 2009 om en europeisk återhämtningsplan Antagna texter, P6_TA(2009)0123 . ,
–
med beaktande av resultatet av Europeiska rådets vårmöte,
–
A.
Världsekonomin går snabbt tillbaka under 2009 och även de mest optimistiska prognoserna förutspår endast en svag återhämtning under 2010, vilket således för oss närmare en djup social och politisk kris.
B.
C.
D.
Flera medlemsstater har haft allvarliga problem med betalningsbalansen och några har tvingats söka hjälp från Internationella valutafonden.
E.
Den globala planen för återhämtning och reform omfattar följande mål: 1) återställa förtroende, tillväxt och sysselsättning, 2) åtgärda finanssystemet för att återställa utlåningen, 3) stärka finansregleringarna och bygga upp tilliten, 4) reformera de internationella finansiella institutionerna och ge dem ekonomiskt stöd för att överbrygga krisen och undvika kriser i framtiden, 5) främja världshandeln och globala investeringar och motverka protektionism, i syfte att värna om välfärden, och 6) åstadkomma en inkluderande, miljövänlig och hållbar återhämtning.
1.
2.
Europaparlamentet lovordar den ledande roll som EU spelade vid toppmötet genom att ge vägledning och utforma praktiska lösningar.
3.
4.
Europaparlamentet uppmanar det nyinrättade FSB (Financial Stability Board) och Internationella valutafonden att förelägga parlamentet sin rapport om hur handlingsplanen för att stärka finanssektorn genomförs i praktiken.
5.
Europaparlamentet uppmärksammar att de ofta kraftfulla åtgärder som vidtagits i finanssektorn inte är avsedda att förebygga nedläggningen av vissa företag, utan att förebygga en kollaps i sektorn, vilket skulle få en katastrofal dominoeffekt i resten av finanssektorn samt i den reala ekonomin.
6.
Europaparlamentet föreslår en fördubbling av EU:s system för medelfristigt ekonomiskt stöd till medlemsstater som inte har infört euron från 25 till 50 miljarder euro.
7.
Europaparlamentet uppmanar med eftertryck alla medlemsstater som inte har fått undantag och inte har infört euron att koncentrera sig på att uppfylla Maastrichtkriterierna och att planera för att införa euron så snart som möjligt för att vara bättre skyddade mot framtida kriser.
8.
Europaparlamentet välkomnar ECB:s upprepade räntesänkningar för att främja tillväxten, och dess snabba agerande för att tillhandahålla kortfristiga finansiella medel för att återupprätta utlåningen mellan bankerna.
9.
10.
11.
Europaparlamentet lovordar G20-gruppen för att framför allt ha valt lösningar som bygger på långivning och garantier, vilket kommer att maximera de ekonomiska effekterna och samtidigt bidra till att minska den långsiktiga påverkan på de statliga finanserna som program på mer än en biljon dollar medför.
12.
Europaparlamentet är oroat över de skilda produktionsnivåerna inom euroområdet och efterlyser korrigerande åtgärder på nationell nivå där så behövs.
13.
14.
Europaparlamentet välkomnar den avsevärda ökningen av Internationella valutafondens resurser eftersom fonden är den viktigaste givaren av ekonomiskt stöd till länder som har problem med betalningsbalansen, däribland EU-medlemsstater, och även verkar för att stödja tillväxten på tillväxtmarknader och i utvecklingsländer.
15.
Europaparlamentet uppmanar kommissionen att bedöma hur mycket extra medel som kan komma att behövas för Internationella valutafondens särskilda dragningsrätter och uppmanar ECB att göra en bedömning av vilka effekter dessa extra medel kan få på den globala prisstabiliteten.
16.
Europaparlamentet välkomnar att alla de fyra länder som stod kvar på OECD:s svarta lista över skatteparadis har tagits bort efter att länderna godkände reglerna om skattetransparens strax efter G20-mötet.
17.
18.
Europaparlamentet betonar behovet av att effektivt genomföra klimat- och energipaket och att investera ytterligare i förnyelsebar energi, energikällor med låg koldioxidproduktion och energieffektivitet, vilket bör utgöra en central del av energihandlingsplanen för 2010–2014.
19.
Europaparlamentet betonar behovet av att integrera miljöinnovation i all relevant politik för att i stor skala snabbt främja sådan innovation, och uppmanar kommissionen att undersöka lagstiftningsramar samt rättsliga hinder och marknadsmisslyckanden som kan hindra tillämpningen av miljöteknik och ytterligare innovation.
20.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, Europeiska centralbanken, medlemsstaternas regeringar och parlament samt G20-gruppens medlemmar och IMF.
om G20-toppmötet i Pittsburgh den 24–25 september 2009
Kay Swinburne
för ECR-gruppen
PE428.685v01-00 B7‑0081/2009 Europaparlamentets resolution om G20-toppmötet i Pittsburgh den 24‑25 september 2009
– med beaktande av ledarnas uttalande vid G20-toppmötet i Pittsburgh den 24‑25 september 2009,
– med beaktande av rådets och kommissionens uttalanden om G20-toppmötet i Pittsburgh den 24–25 september 2009,
2.
Europaparlamentet noterar bekymrat att statsskulderna och budgetunderskotten blir allt större.
Parlamentet understryker hur viktigt det är att trygga sunda statsfinanser och övervaka dem på ett lämpligt sätt så att man undviker att skapa alltför stora bördor för kommande generationer.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, Europeiska centralbanken, medlemsstaternas parlament och regeringar samt G20-gruppens och Internationella valutafondens medlemmar.
om främjande av demokrati i EU:s yttre förbindelser
Charles Tannock
,
Adam Bielan
,
Ryszard Antoni Legutko
,
Tomasz Piotr Poręba
för ECR-gruppen
PE428.727v01-00 B7‑0119/2009 Europaparlamentets resolution om främjande av demokrati i EU:s yttre förbindelser
Europaparlamentet utfärdar denna resolution
– med beaktande av den allmänna förklaringen om de mänskliga rättigheterna, särskilt artikel 21 i denna, och den internationella konventionen om medborgerliga och politiska rättigheter,
– med beaktande av artiklarna 3, 6, 11 och 19 i fördraget om Europeiska unionen och artiklarna 177, 300 och 310 i EG-fördraget,
– med beaktande av alla avtal mellan EU och tredjeländer samt de klausuler om mänskliga rättigheter och demokrati som ingår i dessa avtal,
– med beaktande av Europeiska unionens stadga om de grundläggande rättigheterna, som kungjordes i Strasbourg den 12 december 2007,
– med beaktande av FN:s generalförsamlings resolution, ”FN:s millenniedeklaration”, av den 8 september 2000 (A/RES/55/2),
– med beaktande av FN:s generalförsamlings resolution av den 4 december 2000 om att främja och befästa demokratin (A/RES/55/96),
– med beaktande av FN:s generalförsamlings resolution av den 15 september 2005 om resultaten från 2005 års världstoppmöte (A/RES/60/1),
– med beaktande av FN:s generalförsamlings resolution av den 23 mars 2005 om att stärka rollen för regionala, subregionala och andra organisationer och arrangemang när det gäller att främja och befästa demokratin (A/RES/59/201),
– med beaktande av kommissionens meddelande om EU:s stöd till och övervakning av val KOM(2000)0191 .
,
– med beaktande av sin resolution av den 15 mars 2001 om kommissionens meddelande om EU:s stöd till och övervakning av val,
– med beaktande av kommissionens meddelande om Europeiska unionens roll i arbetet för att främja mänskliga rättigheter och demokratisering i tredje land KOM(2001)0252 .
,
– med beaktande av sin resolution av den 25 april 2002 om kommissionens meddelande om Europeiska unionens roll i arbetet för att främja mänskliga rättigheter och demokratisering i tredje land,
– med beaktande av den europeiska säkerhetsstrategin av den 12 december 2003,
– med beaktande av kommissionens meddelande om styre och utveckling KOM(2003)0615 .
,
– med beaktande av Europeiska unionens samförstånd om utveckling från 2005,
– med beaktande av Parisdeklarationen om biståndseffektivitet från 2005 och handlingsprogrammet från Accra från 2008,
– med beaktande av kommissionens meddelande ”Samhällsstyrning och det europeiska samförståndet om utveckling – Mot ett harmoniserat tillvägagångssätt i Europeiska unionen” KOM(2006)0421 .
,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1889/2006 av den 20 december 2006 om inrättande av ett finansieringsinstrument för främjande av demokrati och mänskliga rättigheter i hela världen,
– med beaktande av sitt presidiebeslut av den 18 juni 2007 om inrättande av byrån för främjande av parlamentarisk demokrati,
– med beaktande av sin resolution av den 8 maj 2008 om EU:s valobservatörsuppdrag: mål, tillvägagångssätt och framtida utmaningar,
– med beaktande av rådets slutsatser från maj 2009 ”Stöd till demokratisk samhällsstyrning – Mot förbättrade EU-ramar”,
– med beaktande av frågan av den 30 september 2009 till kommissionen om främjande av demokrati inom ramen för de yttre förbindelserna ( O-0093/2009 - B7-0213/2009 ).
,
B. I Europeiska unionens grundfördrag görs ett beslutsamt åtagande till förmån för demokrati och mänskliga rättigheter.
De politiska Köpenhamnskriterierna om stabila institutioner som garanterar demokrati, rättsstatsprincipen, mänskliga rättigheter samt respekt för och skydd av minoriteter har utgjort nyckelprinciper i utvidgningsprocessen.
C. En bred förståelse för demokrati har bidragit till att politiska, sociala och ekonomiska rättigheter kunnat integreras i EU och spelat en väsentlig roll i världshistorien när det gäller att åstadkomma stabilitet och välstånd.
D. Enligt artikel 11 i EU-fördraget är ett av de främsta målen med den gemensamma utrikes- och säkerhetspolitiken att ”utveckla och befästa demokratin och rättsstatsprincipen samt respekten för de mänskliga rättigheterna och de grundläggande friheterna”.
• Respekt för de mänskliga rättigheterna och de grundläggande friheterna, bland annat föreningsfrihet och frihet att delta i fredliga sammankomster samt yttrande- och åsiktsfrihet.
• Rätt att delta i utövandet av offentliga uppdrag, direkt eller via fritt valda företrädare, rätt att rösta och låta sig väljas i fria, hemliga och regelbundet anordnade val på grundval av allmän och lika rösträtt som garanterar befolkningen rätt att fritt uttrycka sin vilja.
• Ett pluralistiskt system med politiska partier och organisationer.
• Respekt för rättssäkerheten.
• Maktdelning och domstolsväsendets oberoende.
• Öppenhet och ansvar i offentlig förvaltning.
• Fria, oberoende och pluralistiska medier.
F. I enlighet med Millenniedeklarationen är ett demokratiskt samhällsstyre som gör medborgarna delaktiga och som är grundat på folkets vilja den bästa garantin för den rätt män och kvinnor har att leva sina liv och fostra sina barn i värdighet, fria från hunger och från fruktan för våld, förtryck och orättvisor.
G. Mäns och kvinnors förmåga att delta på lika villkor i det politiska livet och i beslutsfattandet är en grundläggande förutsättning för en verklig demokrati.
H. Demokrati, utveckling och respekt för alla mänskliga rättigheter, inbegripet ekonomiska, sociala och kulturella rättigheter, är sinsemellan förbundna och ömsesidigt förstärkande.
I. Demokrati är också tydligt kopplat till säkerhet, vilket bekräftas i den europeiska säkerhetsstrategin, där det står att det bästa sättet att stärka den internationella ordningen är att sprida normer för goda styrelseformer, stödja sociala och politiska reformer, ta itu med korruption och maktmissbruk, etablera rättsstatsprincipen och skydda mänskliga rättigheter.
J. Europeiska unionen förfogar över ett stort antal instrument och verktyg, allt från politisk dialog och diplomatiska initiativ till specifika instrument för finansiering och tekniskt samarbete, för att stödja demokratin över hela världen.
K. Europeiska unionens externa finansieringsinstrument, såsom instrumentet för utvecklingssamarbete, Europeiska grannskaps- och partnerskapsinstrumentet och stabilitetsinstrumentet, ger alla stora möjligheter till demokratiskt styre och stöd till institutionell och kapacitetsmässig uppbyggnad.
N. I parlamentets betänkande från 2004 om kommissionens meddelande om styre och utveckling betonades “vikten av att fortsätta valsystemsreformer och parlamentariska reformer bortom inrättandet av flerpartisystem för att säkerställa mer omfattande och effektivare politisk aktivitet bland befolkningen” A5-0219/2004
.
Europaparlamentet rekommenderar rådet att i sina slutsatser inbegripa konkreta och praktiska förslag till förbättring av samordningen av demokratistödet inom ramen för EU:s instrument på området för utrikespolitik, mänskliga rättigheter och utvecklingspolitik.
Europaparlamentet rekommenderar EU att, i syfte att stärka de samordnade åtgärderna över hela världen till förmån för demokrati, offentligt anta FN:s generalförsamlings definition av demokrati som utgångspunkt för sitt eget demokratiseringsarbete.
Europaparlamentet föreslår att rådet och kommissionen ska fortsätta arbetet med en omfattande och detaljerad analys av allt det demokratistöd EU ger i ett urval av partnerländer, så att det blir möjligt att utfärda praktiska rekommendationer.
Europaparlamentet understryker att EU:s demokratistöd måste vara omfattande och inbegripa alla frågor som tas upp i FN:s generalförsamlings resolution från 2005, och att EU måste anta ett långsiktigt perspektiv i sina insatser.
Europaparlamentet betonar att EU:s insatser för att främja demokratin mer systematiskt bör innebära att man särskilt uppmärksammar de förtroendevaldas, de politiska partiernas och de oberoende mediernas roll.
19.
om insynen och läget i Acta-förhandlingarna
Carl Schlyter
,
Eva Lichtenberger
,
Christian Engström
,
Jan Philipp Albrecht
,
Franziska Keller
för Verts/ALE-gruppen
PE433.016v01-00 B7‑0154/2010 Europaparlamentets resolution om insynen och läget i Acta-förhandlingarna
Europaparlamentet utfärdar denna resolution
– med beaktande av artikel 218 i EUF-fördraget,
– med beaktande av sin resolution av den 9 februari 2010 om en översyn av ramavtalet mellan Europaparlamentet och Europeiska kommissionen under den aktuella valperioden ( B7–0091/2010 ),
– med beaktande av sin resolution av den 11 mars 2009 om allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar (omarbetning), som ska betraktas som parlamentets ståndpunkt vid den första behandlingen ( KOM(2008)0229 − C6-0184/2008 – 2008/0090(COD) ),
– med beaktande av sin resolution av den 18 december 2008 om varumärkesförfalskningens inverkan på den internationella handeln ( 2008/2133(INI) ),
– med beaktande av Europeiska datatillsynsmannens yttrande av den 22 februari 2010 om EU:s pågående förhandlingar om ett handelsavtal för bekämpning av varumärkesförfalskning (Acta),
– med beaktande av Europeiska unionens stadga om de grundläggande rättigheterna, särskilt artikel 8,
– med beaktande av Europaparlamentets och rådets direktiv 2002/58/EG om behandling av personuppgifter och integritetsskydd inom sektorn för elektronisk kommunikation, senast ändrat genom Europaparlamentets och rådets direktiv 2009/136/EG av den 25 november 2009,
– med beaktande av Europaparlamentets och rådets direktiv 2000/31/EG av den 8 juni 2000 om vissa rättsliga aspekter på informationssamhällets tjänster, särskilt elektronisk handel, på den inre marknaden (”direktiv om elektronisk handel”),
B. År 2008 inledde EU och andra OECD-länder förhandlingar om ett nytt plurilateralt avtal för att skärpa tillämpningen av immaterialrätten och bekämpa förfalskningar och piratkopiering (handelsavtalet för bekämpning av varumärkesförfalskning – Acta).
C. I sitt betänkande av den 11 mars 2009 uppmanade parlamentet kommissionen att ”omgående ge allmänheten tillgång till alla handlingar som rör de pågående internationella förhandlingarna om handelsavtalet för bekämpning av varumärkesförfalskning (Acta)”.
E. Som fördragens väktare är kommissionen skyldig att försvara unionens regelverk när den förhandlar om internationella avtal som påverkar lagstiftningen inom EU.
F. Enligt de dokument som läckt ut berör Acta-förhandlingarna bland annat kommande EU‑lagstiftning om tillämpning av materialrätten (COD/2005/0127, straffrättsliga åtgärder till skydd för immateriella rättigheter (IPRED-II)) och det så kallade Telekompaketet, samt befintlig EU-lagstiftning om e-handel och uppgiftsskydd.
G. EU:s pågående ansträngningar att harmonisera åtgärderna för tillämpning av materialrätten bör inte kringgås genom handelsförhandlingar som ligger utanför EU:s normala beslutsprocess.
I. Varje eventuellt Acta-avtal som ingås av EU måste vara förenligt med de rättsliga skyldigheter som ålagts EU avseende respekt för lagstiftning om integritetsskydd, yttrandefrihet och uppgiftsskydd, såsom särskilt fastställts i direktiv 95/46/EG och direktiv 2002/58/EG och i Europadomstolen och EU-domstolens rättspraxis.
Europaparlamentet är ytterst bekymrat över bristen på insyn under Acta-förhandlingarna, vilket står i strid med andan och bokstaven i EUF-fördraget.
Europaparlamentet beklagar parternas utstuderade val att inte förhandla via väletablerade internationella organ, som WIPO och Världshandelsorganisationen, som har etablerade ramar för offentlig information och offentliga samråd.
Europaparlamentet påminner kommissionen om att om den inte ger parlamentet omedelbar och fullständig information om förhandlingarna i enlighet med artikel 218 i EUF-fördraget före nästa förhandlingsomgång i april kommer parlamentet inte att ha något annat val än att väcka talan hos EU-domstolen i enlighet med artikel 263 i EUF‑fördraget för överträdelse av fördragen.
Europaparlamentet framhåller att integritets- och uppgiftsskydd är grundläggande värderingar för EU och erkänns som sådana i artikel 8 i Europeiska konventionen om de mänskliga rättigheterna och i artiklarna 7 och 8 i EU:s stadga om de grundläggande rättigheterna.
8.3.2010 B7-0200/2010 FÖRSLAG TILL RESOLUTION i enlighet med artikel 120 i arbetsordningen
om jämställdhet och våld mot kvinnor
Cristiana Muscardini
PE439.716v01-00 B7‑0200/2010 Europaparlamentets resolution om jämställdhet och våld mot kvinnor
Europaparlamentet utfärdar denna resolution
– med beaktande av sina tidigare resolutioner om lika möjligheter,
– med beaktande av sin resolution av den 26 november 2009 om avskaffande av våld mot kvinnor Antagna texter, P7_TA-PROV(2009)0098 .
,
– med beaktande av artikel 120 i arbetsordningen, och av följande skäl:
A. Andelen kvinnor inom institutionerna har visserligen ökat något, men fortfarande är det lång väg kvar till en jämn balans mellan könen.
B. Kvinnor är kraftigt underrepresenterade även i det civila samhället, både när det gäller ansvarsuppdrag (styrelser och chefspositioner) och representationsuppdrag.
Europaparlamentet uppmanar rådet och kommissionen att rekommendera medlemsstaterna att främja kvinnors deltagande i styrelser för företag som har anknytning till den offentliga sektorn, på både nationell och lokal nivå.
Europaparlamentet uppmanar rådet och kommissionen att, mot bakgrund av de negativa resultaten från den enkät som gjorts för att bedöma kvinnors intresse för EU, vidta åtgärder för att se till att kvinnors verkliga intressen beaktas i EU-politiken.
om situationen i Kirgizistan
Heidi Hautala
,
Bart Staes
,
Nicole Kiil-Nielsen
för Verts/ALE-gruppen
PE442.017v01-00 B7‑0419/2010 Europaparlamentets resolution om situationen i Kirgizistan
Europaparlamentet utfärdar denna resolution
– med beaktande av sina tidigare resolutioner om Kirgizistan och Centralasien, särskilt resolutionen av den 6 maj 2010,
– med beaktande av parlamentets resolution av den 20 februari 2008 om en EU-strategi för Centralasien,
– med beaktande av uttalandena av vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik Catherine Ashton om de nya sammandrabbningarna i Kirgizistan den 11 juni 2010 och om folkomröstningen om konstitutionen den 28 juni 2010,
– med beaktande av rådets (utrikes frågor) slutsatser av den 14 juni 2010,
– med beaktande av EU:s strategi för ett nytt partnerskap med Centralasien, som antogs av Europeiska rådet den 21–22 juni 2007,
– med beaktande av partnerskaps- och samarbetsavtalet mellan EU och Kirgizistan, som trädde i kraft 1999,
A. Den 11 juni 2010 utbröt våldsamma sammandrabbningar i städerna Osh och Jalalabad i södra Kirgizistan vilka fortsatte att eskalera fram till den 14 juni, då hundratals beväpnade män rapporterades storma stadens gator, skjuta civila och sätta affärer i brand, varvid de valde sina mål utifrån etniska kriterier.
E. Enligt den nationella säkerhetstjänstens utredning av händelserna den 11–14 juni anstiftades sammandrabbningarna av medlemmar ur samma klan som den fördrivne presidenten Bakijev i samarbete med radikala islamister, militanta grupper från norra Tadzjikistan och talibaner .
J. EU måste alltid stå fast vid sitt åtagande att mänskliga rättigheter, demokrati och rättsstatliga principer ska ingå i unionens avtal med tredje länder och främja demokratiska reformer genom en konsekvent politik som ökar dess trovärdighet som regional aktör.
Europaparlamentet betonar att de värden som Europeiska unionen bekänner sig till tvingar unionen att agera på alla nivåer med anledning av detta lidande, inklusive genom att anslå mer än de 5 miljoner EUR som hittills har uppbringats; stöd som bör stå i proportion till FN:s begäran om 71 miljoner USD för omedelbar humanitär hjälp.
Europaparlamentet uppmanar enträget rådet att ta ledningen och arrangera en internationell givarkonferens för Kirgizistan, för att behandla de humanitära problemen och de grundläggande behoven i Kirgizistan och tillhandahålla det bistånd som krävs för en hållbar utveckling i landet.
Europaparlamentet uppmanar vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik och medlemsstaterna att stödja och aktivt bidra till en snabb polisiär insats från OSSE för att förhindra att nya våldsamheter bryter ut, för att stabilisera situationen i de städer där sammandrabbningar ägt rum samt för att skydda offren och de mest sårbara personerna och underlätta för flyktingar och internflyktingar att återvända.
Europaparlamentet uttrycker sin oro över rapporterna om gripandet av vissa människorättsaktivister i Kirgizistan, och uppmanar de kirgiziska myndigheterna att vidta alla nödvändiga åtgärder för att garantera att människorättsaktivister obehindrat kan bedriva sitt arbete för att främja och slå vakt om de mänskliga rättigheterna.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik, rådet, kommissionen och OSSE.
om situationen för romerna i Europa
Cornelia Ernst
,
Marie-Christine Vergiat
,
Rui Tavares
,
Willy Meyer
,
Nikolaos Chountis
,
Patrick Le Hyaric
,
Miguel Portas
,
Jacky Hénin
,
Kyriacos Triantaphyllides
för GUE/NGL-gruppen
PE446.583v01-00 B7‑0500/2010 Europaparlamentets resolution om situationen för romerna i Europa
Europaparlamentet utfärdar denna resolution
– med beaktande av internationella och europeiska konventioner om skydd av mänskliga rättigheter och grundläggande friheter, Europeiska konventionen om skydd för de mänskliga rättigheterna och de grundläggande friheterna och därtill hörande rättspraxis från Europeiska domstolen för de mänskliga rättigheterna
samt Europeiska unionens stadga om de grundläggande rättigheterna,
– med beaktande av stadgan om de grundläggande rättigheterna, särskilt artiklarna 21 (icke‑diskriminering) och 45 (rörelse- och uppehållsfrihet),
– med beaktande av artiklarna 2, 6 och 7 i fördraget om Europeiska unionen samt artiklarna 13 (åtgärder mot diskriminering på grund bland annat av ras eller etniskt ursprung), 12 (förbud mot diskriminering på grund av nationalitet) och 18 (fri rörlighet),
– med beaktande av rådets direktiv 2000/43/EG om genomförandet av principen om likabehandling av personer oavsett deras ras eller etniska ursprung
och framför allt av definitionerna av direkt och indirekt diskriminering, samt av Europaparlamentets och rådets direktiv 2004/38/EG om unionsmedborgares och deras familjemedlemmars rätt att fritt röra sig och uppehålla sig inom medlemsstaternas territorier
,
– med beaktande av kommissionens meddelande om integreringen av romerna i samhället och i näringslivet ( KOM(2010)0133 ) samt rapporterna från Europeiska unionens byrå för grundläggande rättigheter,
– med beaktande av sina tidigare resolutioner om bland annat romer, rasism och främlingsfientlighet, åtgärder mot diskriminering samt om fri rörlighet, nämligen resolutionerna av den 31 januari 2008 om en europeisk strategi för romer
, av den 10 juli 2008 om folkräkningen av romerna i Italien på grundval av etniskt ursprung samt av den 25 mars 2010 om det andra europeiska toppmötet om romer,
– med beaktande av sin resolution av den 14 januari 2009 om situationen för de grundläggande rättigheterna i Europeiska unionen 2004–2008,
– med beaktande av rekommendationerna från FN:s kommitté för avskaffande av rasdiskriminering vid dess 77:e session (den 2–27 augusti 2010) med avseende på Danmark, Estland, Frankrike, Rumänien och Slovenien,
E. Den 19 augusti 2010 återsändes 86 romer till Rumänien och Bulgarien, följda av omkring 130 den 20 augusti och omkring 300 den 26 augusti, och regeringen tillkännagav att omkring 800 romer skulle återsändas före utgången av augusti.
I. Djup oro och allvarliga farhågor har uttryckts av Europarådets kommission mot rasism och intolerans, FN:s kommitté för avskaffande av rasdiskriminering, Europarådets kommissarie för mänskliga rättigheter och talmannen i Europarådets parlamentariska församling.
M. Rätten till fri rörlighet är en grundläggande rättighet som inskrivits i EU-fördragen och regleras av bestämmelser i direktiv 2004/38/EG, som blivit föremål både för en rapport från kommissionen och för riktlinjer för hur medlemsstaterna korrekt ska tillämpa direktivet.
N. I sin gemensamma förklaring om det andra europeiska toppmötet om romer, vilket hölls i Cordoba den 8–9 april 2010, åtog sig EU:s trio att
– arbeta för att frågor som berör romerna ska tas med i all europeisk och nationell politik för grundläggande rättigheter och skydd mot rasism, fattigdom och socialt utanförskap,
– förbättra färdplanen för den integrerade plattformen för romers integrering och prioritera de huvudsakliga målen och resultaten,
– se till att Europeiska unionens nuvarande former för ekonomiskt stöd, framför allt strukturfonderna, görs tillgängliga för romer.
O. Utvisningarna av romer är redan i sig allvarliga brott mot de europeiska värderingarna när det gäller mänskliga rättigheter och grundläggande friheter och bryter också mot EU‑medlemsstaternas åtaganden att stärka romernas integrering, i den form dessa åtaganden antagits vid det andra toppmötet om romer.
P. Kommissionen är skyldig att se till att EU-fördragen och unionslagstiftningen följs samt att de mänskliga rättigheterna och de grundläggande friheterna respekteras, skyddas och främjas i EU, och kommissionen ska genast ingripa med kraft så fort det förekommer uppenbara brott i detta hänseende.
Europaparlamentet understryker att dessa åtgärder strider mot EU:s fördrag och lagstiftning, mot direktiv 2000/43/EG, eftersom de är liktydiga med diskriminering på grundval av ras och etnisk tillhörighet, och mot direktiv 2004/38/EG om fri rörlighet för medborgare och deras familjer i EU, och eftersom kollektiva utvisningar är förbjudna enligt stadgan om de grundläggande rättigheterna och Europeiska konventionen om skydd för de mänskliga rättigheterna och de grundläggande friheterna.
Europaparlamentet uppmanar med kraft medlemsstaterna att strikt fullgöra sina skyldigheter och att få bort inkonsekvenserna i sin tillämpning av kraven i direktivet om fri rörlighet.
Europaparlamentet fördömer provocerande uttalanden som kopplar samman minoriteter och invandrare med kriminalitet, eftersom detta cementerar negativa stereotyper som bidrar till stigmatisering och diskriminering av romer.
Europaparlamentet uppmanar medlemsstaterna, däribland särskilt Frankrike, att avhjälpa bristerna i skyddet för minoriteter på sitt territorium genom att underteckna och ratificera Europarådets ramkonvention för skydd av nationella minoriteter.
Parlamentet upprepar också sin uppmaning till rådet och kommissionen om att de bör övervaka hur medlemsstaterna tillämpar fördragen och direktiven om åtgärder mot diskriminering samt fri rörlighet, särskilt i förbindelse med romer, och att nödvändiga åtgärder bör vidtas om så inte är fallet.
28.9.2010 B7-0537/2010 FÖRSLAG TILL RESOLUTION i enlighet med artikel 120 i arbetsordningen
om ersättning av beteckningen ”romer”
Sebastian Valentin Bodu
PE446.628v01-00 B7‑0537/2010 Förslag till Europaparlamentets resolution om ersättning av beteckningen ”romer”
Europaparlamentet utfärdar denna resolution
– med beaktande av att beteckningen ”romer” skapar förvirring och leder till sammanblandning både med beteckningen ”rumäner” (som syftar på invånare i Rumänien) och namnet ”Rom” eller ”Roma” (som syftar på Italiens huvudstad),
– med beaktande av artikel 120 i arbetsordningen, och av följande skäl:
A. En sådan sammanblandning kan få oönskade följder för såväl invånare i Rumänien som invånare i Rom vad beträffar hur dessa invånare uppfattas av medborgare i och utanför EU, liksom för den romska minoritetens etniska identitet.
B. Det finns ett land (Makedonien) som vill ändra sitt namn för att uppfylla EU:s anslutningskrav.
om värphönsindustrin i EU: förbudet mot användning av burar från och med 2012
George Lyon
,
Chris Davies
för ALDE-gruppen
PE450.537v01-00 B7‑0706/2010 Europaparlamentets resolution om värphönsindustrin i EU: förbudet mot användning av burar från och med 2012
Europaparlamentet utfärdar denna resolution
– med beaktande av rådets direktiv 1999/74/EG som trädde i kraft den 3 augusti 1999 och innebar att ett förbud infördes mot användning av burar för uppfödning av värphöns, men även att en övergångsperiod på mer än 12 år beviljades under vilken producenterna skulle ändra sina uppfödningssystem,
– med beaktande av kommissionens förordning 589/2008/EG om tillämpningsföreskrifter för handelsnormerna för ägg,
– med beaktande av rådets förordning (EG) nr 1234/2007 av den 22 oktober 2007 om upprättande av en gemensam organisation av jordbruksmarknaderna och om särskilda bestämmelser för vissa jordbruksprodukter (förordningen om en samlad marknadsordning),
– med beaktande av kommissionens meddelande från 2008 om de olika uppfödningssystemen för värphönor, särskilt de som omfattas av rådets direktiv 1999/74/EG,
A. Direktivet om värphöns välbefinnande (1999/74/EG) innebär ett förbud mot uppfödning av värphöns i icke inredda burar från och med den 1 januari 2012, och medlemsstaterna och producenterna kommer då att ha haft mer än 12 år på sig att se till att de iakttar villkoren i lagstiftningen.
C. Ägg som inte produceras i enlighet med direktiv 1999/74/EG får enligt lag inte säljas i Europeiska unionen.
E. Medlemsstaterna ansvarar för att det införs sanktionssystem som är proportionella, effektiva och avskräckande för att garantera att direktivet genomförs, medan kommissionen, i egenskap av fördragets väktare, övervakar läget för genomförandet i EU och vid behov vidtar åtgärder.
F. Rapporter från GD Jordbruk om det nuvarande läget och uppskattningar som gjorts av sektorn för de kommande åren visar att ett betydande antal medlemsstater och 30 procent av äggproducenterna inte förväntas iaktta förbudet mot burar senast den 1 januari 2012.
G. Direktiv 1999/74/EG omfattar inte några eventuella påföljder som medlemsstaterna kan införa mot andra medlemsstater som har underlåtit att genomföra direktiv 1999/74/EG fullständigt före 2012.
H. Ägg- och fjäderfäproduktionssektorn får inget direktstöd inom ramen för den gemensamma jordbrukspolitiken samtidigt som den måste iaktta EU-standarder för djurhälsa och djurskydd som är bland de högsta i världen.
Europaparlamentet är allvarligt oroat över det stora antal medlemsstater och äggproducenter som ligger efter i tidsschemat när det gäller att iaktta tidsfristen.
Europaparlamentet uppmanar kommissionen att omedelbart skapa klarhet och senast den 1 mars 2011 tala om vilka åtgärder man har för avsikt att vidta för att se till att direktivet iakttas.
Europaparlamentet insisterar på att kommissionen inte ska vidta någon åtgärd mot en medlemsstat som hindrar saluföring och import av ägg som inte har producerats i enlighet med EU:s lagstiftning.
12.
FÖRSLAG TILL RESOLUTION till följd av frågan för muntligt besvarande B7‑0670/2010
om internationella adoptioner i Europeiska unionen
Roberta Angelilli
,
Manfred Weber
,
Simon Busuttil
,
Edit Bauer
för PPE-gruppen
Lorenzo Fontana
,
Fiorello Provera
,
Oreste Rossi
Claudio Morganti
PE455.856/rev/v02-00 B7‑0029/2011 Europaparlamentets resolution om internationella adoptioner i Europeiska unionen
Europaparlamentet utfärdar denna resolution
– med beaktande av FN:s konvention om barnets rättigheter, som antogs av FN:s generalförsamling den 20 november 1989, särskilt artikel 21,
– med beaktande av konventionen om skydd av barn och samarbete vid internationella adoptioner (som undertecknades i Haag 1993) och av Europeiska konventionen av den 25 januari 1996 om utövandet av barns rättigheter (ETS nr 160),
– med beaktande av sin resolution om förbättrad lagstiftning och förbättrat samarbete mellan medlemsstaterna beträffande adoption av minderåriga ( A4-0392/1996 ),
– med beaktande av sin resolution av den 16 januari 2008 om en EU-strategi för barnets rättigheter ( 2007/2093(INI) ),
– med beaktande av den muntliga frågan av den 16 december 2010 till kommissionen om internationella adoptioner i Europeiska unionen ( O-0193/2010 – B7-0670/2010 ),
A. Medlemsstaterna har olika åsikter om vilka principer som bör ligga till grund för adoptioner av barn, adoptionsförfaranden och de rättsliga följderna av adoptioner.
B. De problem som orsakas av skillnaderna i nationell lagstiftning skulle kunna minskas om gemensamma reviderade principer och metoder antogs i fråga om barnadoptioner, vilket även skulle främja adoptivbarnens intressen.
C. Problemet med övergivna barn inom Europa blir allt allvarligare och allt mer brådskande, och för att möta denna kris är det viktigt att barns rätt att adopteras skyddas också på internationell nivå, så att man förhindrar att barn tvingas leva på barnhem.
D. Det finns gällande konventioner om skyddet av barn och föräldrars ansvar, närmare bestämt Europeiska konventionen från 1967 om adoption av minderåriga, som syftar till tillnärmning av medlemsstaternas lagstiftning i fall där adoptionen innebär att barnet flyttas från ett land till ett annat, och konventionen om skydd av barn och samarbete vid internationella adoptioner från 1993.
F. Kränkningar av barns rättigheter, våld mot barn och människohandel med barn för syften som olagliga adoptioner, prostitution, olagligt arbete, tvångsäktenskap, gatutiggeri eller andra olagliga syften är fortfarande ett problem inom EU.
G. Det är ytterst viktigt att barnens intressen sätts i främsta rummet.
Europaparlamentet uppmanar medlemsstaterna och kommissionen att i samarbete med Haagkonferensen, Europarådet och barnorganisationer ta fram en ram för att garantera insyn i och effektiv övervakning av vad som händer med övergivna och adopterade barn samt att samordna sina insatser så att människohandel med barn förhindras.
om stigande livsmedelspriser
Nirj Deva
,
James Nicholson
,
Jan Zahradil
,
Janusz Wojciechowski
,
Michał Tomasz Kamiński
för ECR-gruppen
PE459.651v01-00 B7‑0119/2011 Europaparlamentets resolution om stigande livsmedelspriser
Europaparlamentet utfärdar denna resolution
– med beaktande av artikel 39 i fördraget om Europeiska unionens funktionssätt,
– med beaktande av Parisdeklarationen om biståndseffektivitet från 2005 och handlingsprogrammet från Accra från 2008,
– med beaktande av rekommendationerna från den internationella bedömningen av kunskaper, vetenskap och teknik inom jordbruket i ett utvecklingsperspektiv (IAASTD) från april 2008,
– med beaktande av jordbruksutsikterna för 2008–2017 från FN:s livsmedels- och jordbruksorganisation (FAO) och Organisationen för ekonomiskt samarbete och utveckling (OECD),
– med beaktande av slutsatserna och förklaringen från FAO:s världstoppmöte om livsmedelstrygghet i Rom den 16–18 november 2009,
– med beaktande av FN:s generalsekreterares rapport från 2010 om genomförandet av millenniedeklarationen,
– med beaktande av rapporten från FN:s utvecklingsprogram (UNDP), ”Beyond the Midpoint: Achieving the Millennium Development Goals (MDGs)”, som offentliggjordes i januari 2010,
– med beaktande av resultaten av ”hälsokontrollreformen” av EU:s gemensamma jordbrukspolitik av den 20 november 2008,
– med beaktande av resultaten av FN:s högnivåplenarmöte om millennieutvecklingsmålen i New York den 20–22 september 2010,
– med beaktande av Europaparlamentets och rådets förordning (EG) nr 1337/2008 av den 16 december 2008 om inrättande av en snabbinsatsmekanism för att hantera de kraftigt stigande livsmedelspriserna i utvecklingsländerna,
– med beaktande av sin resolution av den 25 oktober 2007 om stigande priser på foder och livsmedel och sin resolution av den 22 maj 2008 om stigande livsmedelspriser i EU och i utvecklingsländerna,
– med beaktande av sin resolution av den 13 januari 2009 om den gemensamma jordbrukspolitiken och global livsmedelsförsörjning,
– med beaktande av sin resolution av den 26 november 2009 om FAO-toppmötet och tryggad livsmedelsförsörjning,
A. Europeiska unionen som helhet, inklusive dess medlemsstater, är fortfarande den ledande givaren av utvecklingsbistånd.
D. Den globala ekonomiska nedgången och de stigande livsmedels- och bränslepriserna har förvärrat livsmedelsläget i många utvecklingsländer, särskilt i de minst utvecklade länderna, vilket delvis hejdat de framsteg som gjorts inom fattigdomsbekämpningen under det senaste årtiondet.
G. Många utvecklingsländer inser inte sin potential i fråga om livsmedelsproduktion.
I. Klimatförändringens följder för jordbruket, särskilt den minskade avkastningen av grödor på grund av upprepad vattenbrist, torka eller – som en kontrast – översvämningar och jordskred, ligger som en tung börda över jordbruksverksamheten i EU och utvecklingsländerna, eftersom ingendera på långa vägar är självförsörjande när det gäller ett flertal jordbruksråvaror.
J. Jordbruksverksamhet som inte är hållbar, till exempel okontrollerad avskogning, bidrar direkt till bristen på högkvalitativ odlingsbar mark för produktion av sunda livsmedel.
Utmaningar och EU:s utvecklingspolitik
Europaparlamentet understryker behovet av att småskaliga jordbrukare i utvecklingsländerna ges ökad tillgång till äganderätt, mikrokrediter – inklusive icke vinstdrivande mikrokreditsystem som fungerar i nära anslutning till behoven hos lokala livsmedelsproducenter – samt inköp av gödningsmedel, särskilt i de fattigare utvecklingsländerna.
Europaparlamentet uppmanar med eftertryck EU:s medlemsstater och det internationella samfundet att stödja Världslivsmedelsprogrammet när det ska möta nya utmaningar i kampen mot svält till följd av snabbt stigande livsmedels- och oljepriser, chockartade väderförhållanden och minskande livsmedelsförråd.
Hållbar livsmedelsproduktion och internationell handel
Europaparlamentet beaktar att jordbruksproduktionen, för att kunna försörja en världsbefolkning som förväntas uppgå till över 9 miljarder människor 2050, kommer att behöva öka med 70 procent fram till dess, samtidigt som man använder mindre mark, vatten och bekämpningsmedel.
om partnerskapsavtalet om fiske mellan Europeiska unionen och Mauretanien
João Ferreira
för GUE/NGL-gruppen
PE459.743v01-00 B7‑0197/2011/rev.
A. Partnerskapsavtalen om fiske bör bygga på en strävan att uppfylla ekonomiska och sociala mål genom ett nära vetenskapligt och tekniskt samarbete enligt villkor som garanterar ett hållbart utnyttjande av fiskeresurserna.
B. Samarbetet bör grundas på ömsesidigt intresse och åtgärder som genomförs gemensamt eller av de enskilda parterna och kompletterar varandra, samtidigt som förenlighet med den fastställda politiken garanteras.
C. Fiskesektorn, inbegripet närstående industrier, spelar en viktig roll i den ekonomiska och sociala utvecklingen i både tredjeländer och medlemsstaterna.
G. Fiskeavtalet mellan EU och Mauretanien är i ekonomiska termer det viktigaste avtalet av alla de avtal som EU undertecknat.
H. De olika stödmöjligheter som fastställts i olika fiskeavtal mellan EU och Mauretanien har i mycket liten utsträckning konkretiserats.
I. Med undantag för hamnen i Nouadhibou i norra delen av landet finns det ingen fiskehamn längs den 700 kilometer långa Atlantkusten.
J. Eftersom fisket är svagt utvecklat i Mauretanien kommer landet inte i åtnjutande av det mervärde som skulle skapas om det själv skulle exploatera sina fiskeresurser (inbegripet beredningsprocesserna och saluföringen av fisk).
K. En sådan utveckling inom fiskesektorn skulle bidra till en ekonomisk och social utveckling i Mauretanien, och leda till ökad sysselsättning, autonomi, suveränitet och självständighet.
L. Europeiska kommissionen har ännu inte lagt fram efterhandsutvärderingen av avtalet om fiske med Mauretanien.
Europaparlamentet försvarar stöd från EU till byggandet – snarast möjligt – av lämpliga anläggningar för landning av fångst längs den centrala och sydliga delen av Mauretaniens kustremsa så att den fisk som fångas i de mauretanska fiskevattnen landas i inhemska hamnar och inte utanför landet, såsom för närvarande ofta sker.
Europaparlamentet anser att det utnyttjande av ett tredjelands resurser som utländska fartygsägare, inbegripet fartygsägare från EU, står för bör begränsas till sådana resurser som inte utnyttjas av landets egna befolkning.
Europaparlamentet uppmanar Europeiska kommissionen att utan dröjsmål lägga fram efterhandsutvärderingen av partnerskapsavtalet om fiske mellan EU och Mauretanien, samt även efterhandsutvärderingarna av övriga partnerskapsavtal.
Europaparlamentet stöder mer rättvisa ekonomiska förbindelser som upprättas på jämbördig fot och som främjar bekämpningen av grundläggande orättvisor och sociala klyftor, hungersnöd, sjukdomar och fattigdom.
om förslaget till ILO:s konvention som kompletteras med en rekommendation om hushållsarbetare
Pervenche Berès
för utskottet för sysselsättning och sociala frågor
PE456.602v01-00 B7‑0296/2011 Europaparlamentets resolution om förslaget till ILO:s konvention som kompletteras med en rekommendation om hushållsarbetare
Europaparlamentet utfärdar denna resolution
– med beaktande av frågan av den 24 februari 2011 till kommissionen om ILO:s konvention om hushållsarbetare ( O-00092/2011 – B7-0305/2011 ),
– med beaktande av sin resolution av den 23 mars 2006 om demografiska utmaningar och solidaritet mellan generationerna EUT C 292 E, 1.12.2006, s.
131.
,
– med beaktande av sin resolution av den 15 januari 2008 om gemenskapens arbetsmiljöstrategi 2007–2012 EUT C 41 E, 19.2.2009, s.
14.
,
– med beaktande av sin resolution av den 19 oktober 2010 om kvinnor med otrygga anställningsförhållanden Antagna texter, P7_TA(2010)0365 .
,
– med beaktande av sin resolution av den 20 oktober 2010 om vikten av ett system med minimiinkomst för att bekämpa fattigdom och främja ett samhälle som är öppet för alla i Europa Antagna texter, P7_TA(2010)0375 .
,
– med beaktande av sin resolution av den 6 juli 2010 om atypiska anställningsformer, säkra yrkesgångar samt nya former för social dialog Antagna texter, P7_TA(2010)0263 .
,
– med beaktande av rådets direktiv 89/391/EEG av den 12 juni 1989 om åtgärder för att främja förbättringar av arbetstagarnas säkerhet och hälsa i arbetet (ramdirektiv) EGT L 183, 29.6.1989, s.
1.
och dess särdirektiv,
– med beaktande av kommissionens meddelande av den 24 maj 2006 ”Anständigt arbete för alla – EU:s bidrag till agendan för anständigt arbete i världen” ( KOM(2006)0249 ) och sin resolution av den 23 maj 2007 EUT C 102 E, 24.4.2008, s.
321.
om anständigt arbete för alla,
– med beaktande av ILO:s rapporter IV.1 och IV.2 om anständigt arbete för hushållsarbetare, som utarbetades inför Internationella arbetskonferensens 99:e sammanträde i juni 2010 samt rapporterna IV.1 (”Brown Report”) och IV.2 (”Blue Report”, utgiven i två volymer) om anständigt arbete för hushållsarbetare, som utarbetades inför Internationella arbetskonferensens 100:e sammanträde i juni 2011,
– med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande över professionaliseringen av hushållsarbetare EESK, SOC/372, 26 maj 2010.
,
– med beaktande av den europeiska konventionen om migrerande arbetstagares ställning (1977),
– med beaktande av det europeiska avtalet om au pair-anställning (1969),
– med beaktande av rekommendation 1663 i den europeiska stadgan om hushållsarbetares rättigheter (2004),
– med beaktande av artiklarna 115.5 och 110.2 i arbetsordningen, och av följande skäl:
2.
5.
Parlamentet anser också att fokus bör ligga på att skapa anständigt arbete för hushållsarbetare och stöder den definition av hushållsarbetare som anges i konventionen.
Parlamentet ser positivt på att man i konventionen tydligt anger att alla arbetstagare som omfattas av denna definition har rätt att behandlas på ett sätt som är förenligt med grundläggande arbetsnormer, social trygghet, icke-diskriminering och likabehandling medan de söker eller har arbete, skydd mot kränkande metoder av arbetsförmedlingar, fortbildning och karriärsutveckling, hälso- och säkerhetsskydd, mödraskydd och bestämmelser om arbetstid/vilotid, skydd mot kränkningar och trakasserier, förenings- och representationsfrihet, kollektivförhandlingar, kollektivåtgärder och livslångt lärande.
Europaparlamentet vill att tillgången till lättillgänglig barnomsorg av hög kvalitet och till ett överkomligt pris utökas, vilket skulle hjälpa till att garantera att arbetstagare inte tvingas att utföra sådant arbete på informell basis.
Dessutom måste man se till att otryggt hushållsarbete där det är möjligt omvandlas till anständiga, välbetalda hållbara arbetstillfällen.
Europaparlamentet anser att man genom att använda bästa praxis från vissa regioner eller medlemsstater, till exempel standardkontrakt, skulle kunna skapa mer stabila anställningsformer för hushållsarbetare som arbetar hemma hos en familj.
Europaparlamentet anser att konventionen bör innehålla strategier som gör att alla människor, däribland de svagaste och mest utsatta, får effektiv tillgång till den formella arbetsmarknaden och lika möjligheter.
.
9.5.2011 B7-0322/2011 FÖRSLAG TILL RESOLUTION till följd av frågorna för muntligt besvarande B7‑0306/2011 , B7-0307/2011 , B7-0308/2011 , B7-0310/2011 , B7-0311/2011 och B7‑0313/2011
om krisen i den europeiska fiskerisektorn till följd av det stigande priset på olja
Ulrike Rodust
för S&D-gruppen
PE465.610v01-00 B7‑0322/2011 Europaparlamentets resolution om krisen i den europeiska fiskerisektorn till följd av det stigande priset på olja
Europaparlamentet utfärdar denna resolution
– med beaktande av kommissionens förordning (EG) nr 1998/2006 om tillämpningen av artiklarna 87 och 88 i fördraget på stöd av mindre betydelse och med beaktande av förordning (EG) nr 875/2007,
1.
Europaparlamentet uttrycker sin oro över den svåra ekonomiska situation som många europeiska yrkesfiskare står inför, vilken har förvärrats ytterligare av de snabbt stigande bränslepriserna.
2.
Europaparlamentet uppmanar kommissionen att undersöka vilka möjligheter som finns och vidta lämpliga åtgärder för att underlätta den svåra ekonomiska situationen för de europeiska yrkesfiskarna, och då även beakta de finansiella svårigheter som flera länder med stora fiskeflottor står inför för närvarande.
3.
Europaparlamentet uppmanar dessutom kommissionen att undersöka om en höjning av det nuvarande taket på 30 000 euro skulle kunna bidra till att förbättra de europeiska yrkesfiskarnas ekonomiska situation, utan att för den delen snedvrida konkurrensen, skada den miljömässiga och sociala hållbarheten eller äventyra EU:s och medlemsstaternas möjligheter att leva upp till sina åtaganden i ramdirektivet om en marin strategi och Europa 2020-strategin.
Parlamentet uppmanar kommissionen att se till att alla former av stöd till fisket med anledning av det stigande oljepriset även ges med fokus på yrkesfiskare som tillämpar hållbara fiskemetoder.
Europaparlamentet stöder de europeiska yrkesfiskarna och upprepar sin begäran till kommissionen om att den bör försöka göra mer tillförlitliga och korrekta bedömningar av vilken inverkan import av fiskeri- och vattenbruksprodukter har på EU:s marknad och vidta åtgärder för att inte bara förhindra en fortsatt urholkning av tullskyddet utan eventuellt även öka det.
Europaparlamentet stöder kommissionens ansträngningar för att förbättra situationen för de europeiska yrkesfiskarna och framför allt för den småskaliga och kustnära fiskeflottan genom en omfattande reform av den gemensamma fiskeripolitiken.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen och medlemsstaternas regeringar och parlament samt till producentorganisationer och den europeiska bearbetningsindustrin.
15.6.2011 B7-0376/2011 FÖRSLAG TILL RESOLUTION i enlighet med artikel 120 i arbetsordningen
om främjande av energiproduktion genom användning av solpaneler på taken till industrianläggningar
Cristiana Muscardini
PE465.689v01-00 B7‑0376/2011 Förslag till Europaparlamentets resolution om främjande av energiproduktion genom användning av solpaneler på taken till industrianläggningar
Europaparlamentet utfärdar denna resolution
– med beaktande av rådets beslut nr 2002/358/EG av den 25 april 2002 om godkännande, på Europeiska gemenskapens vägnar, av Kyotoprotokollet,
– med beaktande av EU:s medlemsstaters åtagande att tillsammans minska sina växthusgasutsläpp under perioden 2008–2012, så att man uppnår en minskning av utvecklingsländernas totala utsläpp med minst 5 procent jämfört med 1990 års nivåer,
– med beaktande av artikel 120 i arbetsordningen, och av följande skäl:
A. I syfte att uppnå dessa mål föreslås det i Kyotoprotokollet ett antal åtgärder såsom stärkande eller införande av nationella strategier för utsläppningsminskning, t.ex. genom bättre energieffektivitet och utveckling av förnybara energikällor.
om situationen i Syrien
Marietje Schaake
,
,
Louis Michel
,
Charles Goerens
,
Sonia Alfano
,
Kristiina Ojuland
,
Izaskun Bilbao Barandica
,
Ramon Tremosa i Balcells
,
Niccolò Rinaldi
för ALDE-gruppen
PE472.668v01-00 B7‑0487/2011 Europaparlamentets resolution om situationen i Syrien
Europaparlamentet utfärdar denna resolution
– med beaktande av sina tidigare resolutioner om Syrien, särskilt resolutionen av den 7 juli 2011 om situationen i Syrien, Jemen och Bahrain mot bakgrund av situationen i arabvärlden och Nordafrika,
– med beaktande av rådet beslut om Syrien av den 12 april, 9 och 23 maj, 20 och 25 juni samt den 2 september 2011 och av uttalandena från unionens höga representant av den 9, 23 och 29 april, 9 maj, 6, 9 och 11 juni, 9 och 31 juli, 1, 4, 18 och 30 augusti samt den 2 september 2011 om en utvidgning av de restriktiva åtgärderna mot den syriska regimen,
– med beaktande av rådets slutsatser om Syrien av den 12 april, 23 maj, 20 juni och den 18 juli 2011,
– med beaktande av Araförbundets uttalande av den 27 augusti 2011 om situationen i Syrien,
– med beaktande av uttalandet av den 19 augusti 2011 från Europaparlamentets talman om Syrien och reaktionen från det internationella samfundet,
– med beaktande av rapporten från informationsuppdraget till Syrien i enlighet med FN:s människorättsråds resolution S-16/1 av den 17 augusti 2011,
– med beaktande av uttalandet av den 3 augusti 2011 från ordföranden i FN:s säkerhetsråd,
– med beaktande av den resolution om människorättssituationen i Syrien som antogs den 23 augusti 2011 av FN:s råd för mänskliga rättigheter vid dess sjuttonde extra möte,
– med beaktande av det gemensamma meddelandet av den 25 maj 2011 om ny respons på ett grannskap i förändring, vilket kompletterar det gemensamma meddelandet av den 8 mars 2011 om ett partnerskap för demokrati och delat välstånd med södra Medelhavsområdet,
– med beaktande av Romstadgan, som Syrien har undertecknat,
– med beaktande av FN:s internationella konvention om medborgerliga och politiska rättigheter från 1966, som Syrien har anslutit sig till,
– med beaktande av den allmänna förklaringen om de mänskliga rättigheterna från 1948,
– med beaktande av FN:s konvention mot tortyr och annan grym, omänsklig eller förnedrande behandling eller bestraffning från 1975, som Syrien har anslutit sig till,
– med beaktande av EU:s riktlinjer om människorättsförsvarare från 2004, som ändrades 2008,
D. Ett informationsuppdrag från FN har kommit fram till att statliga säkerhetsstyrkor i Syrien kan ha begått brott mot mänskligheten under de våldsamma attackerna mot civila.
E. Städerna Hama, Hums och Latakia har utsatts för storskaliga militära anfall som omfattat både flygbombningar och angrepp från flottan.
F. Den syriska regeringen har stängt av vatten- och elförsörjningen och stoppat tillförseln av livsmedel och läkemedel till hela städer i ett försök att tysta sina egna medborgare.
Rapporter från syriska människorättsaktivister och bilder från mobiltelefoner är det enda sättet att få kännedom om de omfattande människorättsbrotten och systematiska angreppen, som ibland är målinriktade och ibland helt slumpmässiga, mot de fredliga demonstranterna och allmänheten i Syrien.
K. Syriska advokater har i allt större utsträckning blivit utsatta för angrepp under samlingar i solidaritet med offer för det våldsamma förtrycket, där de har krävt ett slut på de godtyckliga frihetsberövandena och tortyren samt ett frigivande av alla personer som hålls orättmätigt fängslade, i synnerhet advokater.
L. Läkare har attackerats medan de har utfört sitt arbete och vårdat sårade oavsett deras åsikter.
N. Distriktsåklagaren i Hama, Muhammad Adnan al-Bakkour, avgick den 1 september i protest mot det pågående brutala våldet mot civila demonstranter.
P. Trots upprepade utfästelser och löften om politiska och demokratiska reformer i Syrien har myndigheterna inte vidtagit några trovärdiga åtgärder för att infria dem, och regeringen har förlorat sin legitimitet.
Q. EU är Syriens viktigaste handelspartner.
S. Den nya strategi som föreslås av kommissionen och den höga representanten som respons på ett grannskap i förändring bygger på ömsesidig ansvarsskyldighet och ett gemensamt åtagande kring de universella värdena mänskliga rättigheter, demokrati och rättstatliga principer.
T. Ledamöter av Europaparlamentet har fört diskussioner med företrädare för den syriska oppositionen i exil vid ett flertal tillfällen under de senaste månaderna.
Europaparlamentet uppmanar de syriska myndigheterna att bevilja oberoende internationella observatörer, människorättsövervakare, humanitära biståndsarbetare och internationella journalister omedelbart tillträde.
Europaparlamentet gläder sig över att rådet den 2 september 2011 antog nya restriktiva åtgärder mot den syriska regimen, inklusive ett förbud mot import av syrisk råolja till EU samt ett reseförbud och ett beslut om frysta tillgångar avseende ytterligare fyra syriska medborgare och tre enheter, bland annat den iranska Quds-styrkan.
Europaparlamentet upprepar sitt starka stöd för de diplomatiska ansträngningar från EU:s medlemsstater i FN:s säkerhetsråd och i andra internationella forum som är inriktade på att få fram lämpliga reaktioner från det internationella samfundet på den rådande krisen i Syrien.
om situationen i Egypten och Syrien, särskilt för de kristna samfunden
Elmar Brok
,
Mario Mauro
,
Ioannis Kasoulides
,
Cristian Dan Preda
Tokia Saïfi
,
Magdi Cristiano Allam
,
Othmar Karas
,
Ria Oomen-Ruijten
,
Gabriele Albertini
,
Inese Vaidere
,
Elena Băsescu
,
Elisabeth Jeggle
,
Monica Luisa Macovei
,
Zuzana Roithová
,
Nadezhda Neynsky
,
Roberta Angelilli
,
Thomas Mann
,
Constance Le Grip
,
Salvatore Iacolino
,
Bernd Posselt
,
Elżbieta Katarzyna Łukacijewska
,
Sari Essayah
,
Anne Delvaux
för PPE-gruppen
PE472.752v02-00 B7‑0555/2011 Europaparlamentets resolution om situationen i Egypten och Syrien, särskilt för de kristna samfunden
Europaparlamentet utfärdar denna resolution
– med beaktande av sina tidigare resolutioner om Egypten och Syrien,
– med beaktande av de uttalanden som vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik gjorde om Syrien den 8 och 31 juli, den 1, 4, 18, 19, 23 och 30 augusti, den 2, 12, och 23 september och den 8 oktober 2011,
– med beaktande av sin resolution av den 20 januari 2011 om situationen för kristna när det gäller religionsfrihet, i vilken Europaparlamentet uppmanade den höga representanten att inrätta en permanent kapacitet inom Europeiska utrikestjänstens direktorat för mänskliga rättigheter för att övervaka situationen vad gäller regeringars och samhällens begränsningar av religionsfriheten och därmed sammanhängande friheter, och att varje år avlägga rapport för Europaparlamentet,
– med beaktande av rådets (utrikes frågor) slutsatser av den 20 februari 2011, i vilka Catherine Ashton (den höga representanten) uppmanades att avlägga rapport om antagna åtgärder och konkreta förslag när det gäller att ytterligare stärka Europeiska unionens insatser för främjande av och respekt för religiösa frågor och religionsfrihet,
– med beaktande av rådets (utrikes frågor) slutsatser av den 10 oktober 2011 om Syrien,
– med beaktande av den internationella konventionen om medborgerliga och politiska rättigheter från 1966, som Egypten och Syrien har anslutit sig till,
Egypten
A. Minst 28 egyptiska medborgare dödades och mer än 350 sårades när militära styrkor den 9 oktober 2011 angrep kopter i Kairo efter en protestaktion mot en attack riktad mot en kyrka i Aswanprovinsen.
B. Sedan början av den arabiska våren har cirka 100 000 kopter lämnat Egypten.
Syrien
Egypten
Europaparlamentet uppmanar de egyptiska myndigheterna att frige de 28 kristna som greps i Maspero.
Europaparlamentet uppmanar eftertryckligen de egyptiska myndigheterna att sätta stopp för diskrimineringen av kopterna, till exempel genom att stryka religiösa hänvisningar i alla officiella handlingar.
Europaparlamentet uppmanar eftertryckligen vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik, Catherine Ashton, att se till att dessa krav genomförs och efterlevs.
10.
Syrien
Europaparlamentet uttrycker sitt djupa deltagande med offrens familjer och berömmer det syriska folket för dess mod och beslutsamhet samt stöder helhjärtat dess strävan att uppnå full respekt för rättsstaten, de mänskliga rättigheterna och de grundläggande friheterna liksom garantier för bättre ekonomiska och sociala villkor.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik, medlemsstaternas regeringar och parlament, Ryska federationens regering och parlament, Folkrepubliken Kinas regering och parlament, Förenta staternas regering och kongress, Arabförbundets generalsekreterare, Arabrepubliken Egyptens regering och Arabrepubliken Syriens regering och parlament.
om Europeiska rådets möte den 8–9 december 2011 ( 2011/2546(RSP) )
Roberto Gualtieri
,
Stephen Hughes
,
Enrique Guerrero Salom
,
Udo Bullmann
för S&D-gruppen
PE479.441v01-00 B7‑0004/2012 Europaparlamentets resolution om Europeiska rådets möte den 8–9 december 2011 ( 2011/2546(RSP) )
Europaparlamentet utfärdar denna resolution
– med beaktande av Europeiska rådets slutsatser av den 8−9 december 2011,
– med beaktande av uttalandet av den 9 december 2011 från euroområdets stats- och regeringschefer,
– med beaktande av paketet med sex lagstiftningsförslag om ekonomisk styrning och de två förslagen från kommissionen om att ytterligare skärpa budgetdisciplinen Förordning om skärpning av den ekonomiska övervakningen och övervakningen av de offentliga finanserna i medlemsstater, COM(2011)0819 , och förordning om gemensamma bestämmelser för övervakning och bedömning av utkast till budgetplaner, COM(2011)0821 .
,
– med beaktande av läget i förhandlingarna om utkastet till internationellt avtal om en starkare ekonomisk union,
– med beaktande av artikel 110.2 i arbetsordningen.
Europaparlamentet bekräftar sitt stöd för det förslag som lades fram i ad hoc‑arbetsgruppen av de ledamöter som utsetts av talmanskonferensen till att företräda parlamentet.
– det i det nya avtalet uttryckligen ska fastställas att EU-lagstiftningen entydigt har företräde framför avtalets bestämmelser,
– alla åtgärder för att genomföra avtalet ska vidtas i enlighet med relevanta förfaranden i EU:s fördrag,
– avtalet måste vara förenligt med EU:s lagstiftning, särskilt med siffrorna i stabilitets- och tillväxtpakten, samt att avtalsparter, i de fall då de vill fastställa mål som inte överensstämmer med EU:s lagstiftning, måste följa tillämpliga rättsliga EU‑förfaranden, och att detta inte får leda till dubbla måttstockar,
– demokratisk ansvarighet måste respekteras genom ett ökat deltagande från Europaparlamentets sida i alla aspekter av EU:s ekonomiska samordning och styrning,
– samarbetet mellan nationella parlament och Europaparlamentet måste ske inom ramen för EU:s fördrag, i enlighet med artikel 9 i protokoll nr 1 till fördraget,
– det nya avtalet måste innehålla ett juridiskt bindande åtagande från avtalsparterna om att de kommer att vidta alla sådana åtgärder som krävs för att avtalet i allt väsentligt införlivas i fördraget inom fem år.
om möjligheten att införa stabilitetsobligationer ( 2011/2959(RSP) )
Sharon Bowles
,
Sylvie Goulard
för utskottet för ekonomi och valutafrågor
PE479.453v01-00 B7‑0016/2012 Europaparlamentets resolution om möjligheten att införa stabilitetsobligationer ( 2011/2959(RSP) )
Europaparlamentet utfärdar denna resolution
– med beaktande av Europaparlamentets och rådets förordning (EU) nr 1173/2011 av den 16 november 2011 om effektiv övervakning av de offentliga finanserna i euroområdet, som är en del av det så kallade ”sexpacket”,
– med beaktande av kommissionens grönbok av den 23 november 2011 om möjligheten att införa stabilitetsobligationer,
– med beaktande av presentationen av den 23 november 2011 av kommissionens vice ordförande Olli Rehn i utskottet för ekonomi och valutafrågor och av diskussionerna av den 29 november 2011 med det tyska rådet av ekonomiska experter om en europeisk skuldinlösenfond,
– med beaktande av Europeiska rådets ordförande Herman Van Rompuys interimsrapport av den 6 december 2011: Mot en starkare ekonomisk union,
1.
Europaparlamentet är mycket oroat över de fortsatta spänningarna på euroområdets statsobligationsmarknader, vilket återspeglats i större spreadar, hög volatilitet och sårbarhet för spekulativa attacker under de två senaste åren.
2.
Europaparlamentet understryker att det ligger i euroområdets och medlemsstaternas långsiktiga intresse att utnyttja alla fördelar med att ge ut euron, som har förutsättning att bli en internationell reservvaluta.
Parlamentet påpekar att det kunde vara i euroområdets intresse att utveckla en gemensam likvid och diversifierad obligationsmarknad.
Europaparlamentet anser också att euroområdet och medlemsstaterna bär ansvaret för att en valuta som används av mer än 330 miljoner människor och många företag och investerare är stabil på lång sikt, något som indirekt påverkar resten av världen.
Parlamentet är öppet och angeläget att aktivt diskutera alla frågor – både styrkor och svagheter – rörande möjligheten att införa stabilitetsobligationer i olika former.
Europaparlamentet tar del av kommissionens bedömning, som utgör en del av kommissionens grönbok om möjligheten att införa stabilitetsobligationer, att stabilitetsobligationer skulle underlätta penningpolitiken i euroområdet och även effektivisera statsobligationsmarknaden och det finansiella systemet i hela euroområdet.
Europaparlamentet anser att de mål som ligger till grund för besluten i Europeiska rådet av den 8–9 december 2011 om att ytterligare stärka de offentliga finansernas hållbarhet också bidrar till att skapa nödvändiga villkor för ett eventuellt införande av stabilitetsobligationer.
– Effektiva marknadsincitament för att minska skulderna.
– Kriterier för inträde och utträde, överenskommelser om villkor och löptid, omfördelning av finansieringsfördelar för de nuvarande AAA-länderna.
– Ett system för differentiering av räntesatser mellan medlemsstater med olika kreditbetyg.
– Budgetdisciplin och ökad konkurrenskraft.
– Procykliska effekter och effekter av skulddeflation.
– Tillräcklig attraktionskraft för marknadsinvesterare, samtidigt som man är försiktig med eller undviker alltför högt ställda säkerheter eller en omfördelning av riskerna mellan länderna.
– Förmånsrätt för stabilitetsobligationer i förhållande till nationella obligationer om medlemsstaten inte kan betala sin skuld.
– Kriterier för tilldelning av lån till medlemsstater och kapaciteten att hantera skulden.
– Mätbara och genomförbara skuldprogram.
– Formaliteterna för en bindande färdplan, i likhet med Maastrichtkriterierna för införandet av den gemensamma valutan.
– Samverkan mellan EFSF och ESM för medlemsstater som har likviditetsproblem.
– Lämpliga rättsliga krav, inklusive ändringar av fördrag och konstitutioner.
om den gemensamma fiskeripolitikens bidrag till produktionen av kollektiva nyttigheter ( 2011/2899(RSP) )
Pat the Cope Gallagher
,
Giommaria Uggias
,
Filiz Hakaeva Hyusmenova
för ALDE-gruppen
PE483.126v01-00 B7‑0067/2012 Europaparlamentets resolution om den gemensamma fiskeripolitikens bidrag till produktionen av kollektiva nyttigheter ( 2011/2899(RSP) )
Europaparlamentet utfärdar denna resolution
– med beaktande av rådets förordning (EG) nr 2371/2002 av den 20 december 2002 om bevarande och hållbart utnyttjande av fiskeresurserna inom ramen för den gemensamma fiskeripolitiken EGT L 358, 31.12.2002. s.
59.
,
– med beaktande av FN:s havsrättskonvention av den 10 december 1982,
– med beaktande av FN:s livsmedels- och jordbruksorganisations (FAO) uppförandekod för ansvarsfullt fiske, som antogs den 31 oktober 1995,
– med beaktande av kommissionens meddelande till Europaparlamentet, rådet, Europeiska ekonomiska och sociala kommittén och Regionkommittén med titeln ”Rio+20: mot en grön ekonomi och bättre styrning” ( COM(2011)0363 ),
– med beaktande av kommissionens meddelande om Europa 2020 ( COM(2010)2020 ),
A. Fiskerisektorn bidrar till EU:s ekonomiska tillväxt genom produktion, förädling och marknadsföring av fisk.
B. EU:s fiskerisektor är en mångfunktionell sektor som vid sidan av den huvudsakliga verksamheten även inbegriper fritidsfiske och vattenbruk.
D. Fiskets mångfunktionella karaktär bör erkännas och stödjas inom ramen för reformen av den gemensamma fiskeripolitiken.
E. Även i kustsamhällen är fritidsfiske ett centralt inslag i fiskeverksamheten.
F. Kustsamhällen har drabbats hårt av nedgången inom fiskerisektorn som helhet, vilket i hög grad har påverkat små fiskehamnar runtom i EU.
Europaparlamentet uppmanar kommissionen att bekräfta att fritidsfiske är förenligt med Europa 2020-strategin och tjänar målen i meddelandet ”Rio+20: mot en grön ekonomi och bättre styrning”.
om den senaste politiska utvecklingen i Ungern ( 2012/2511(RSP) )
Hannes Swoboda
,
Sylvie Guillaume
,
Juan Fernando López Aguilar
,
Claude Moraes
,
Csaba Sándor Tabajdi
,
Kinga Göncz
för S&D-gruppen
Guy Verhofstadt
,
Renate Weber
,
Louis Michel
,
Alexander Alvaro
,
Sonia Alfano
,
Ramon Tremosa i Balcells
,
Kristiina Ojuland
, Sophia in ’t Veld
för ALDE-gruppen
Daniel Cohn-Bendit
,
Rebecca Harms
,
Judith Sargentini
,
Rui Tavares
,
Ulrike Lunacek
för Verts/ALE-gruppen
Cornelia Ernst
,
Marie-Christine Vergiat
för GUE/NGL-gruppen
PE483.154v01-00 B7‑0095/2012 Europaparlamentets resolution om den senaste politiska utvecklingen i Ungern ( 2012/2511(RSP) )
Europaparlamentet utfärdar denna resolution
– med beaktande av artiklarna 2, 3, 4, 6 och 7 i fördraget om Europeiska unionen (EU‑fördraget), artiklarna 49, 56, 114, 167 och 258 i fördraget om Europeiska unionens funktionssätt (EUF-fördraget), Europeiska unionens stadga om de grundläggande rättigheterna samt den europeiska konventionen om skydd för de mänskliga rättigheterna (Europakonventionen), vilka rör respekten för och främjande och skydd av de grundläggande rättigheterna,
– med beaktande av Ungerns grundlag som antogs av republiken Ungerns nationalförsamling den 18 april 2011 (nedan kallad ”den nya författningen”) samt de övergångsbestämmelser till denna som antogs av nationalförsamlingen den 30 december 2011 (nedan kallade ”övergångsbestämmelserna”),
– med beaktande av yttrandena CDL(2011)016 och CDL(2011)001 från Europeiska kommissionen för demokrati genom lag (Venedigkommissionen) över den nya ungerska författningen och de tre rättsliga frågor som utarbetandet av den nya ungerska författningen väcker,
– med beaktande av sin resolution av den 10 mars 2011 om den ungerska medielagen samt sin resolution av den 5 juli 2011 om Ungerns reviderade författning,
– med beaktande av kommissionens meddelande ”Artikel 7 i Fördraget om Europeiska unionen – Att respektera och främja unionens värden” ( COM(2003)0606 ),
– med beaktande av den högnivågrupp för mediefrihet och mediepluralism som kommissionens vice ordförande Neelie Kroes inrättade i oktober 2011,
– med beaktande av rådets och kommissionens uttalanden inför kammaren vid parlamentets plenardebatt den 18 januari 2012 om den senaste politiska utvecklingen i Ungern samt med beaktande av den utfrågning som utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor anordnade den 9 februari 2012,
– med beaktande av kommissionens beslut av den 17 januari 2012 att inleda påskyndade överträdelseförfaranden mot Ungern med anledning av frågor beträffande den ungerska nationalbankens och de ungerska dataskyddsmyndigheternas oberoende samt beträffande landets rättsväsende,
A. Europeiska unionen är grundad på värdena demokrati och rättsstatliga principer, vilket fastställs i artikel 2 i EU-fördraget, på en entydig respekt för de grundläggande fri- och rättigheterna, vilket fastställs i Europeiska unionens stadga om de grundläggande rättigheterna och i Europakonventionen, samt på ett erkännande av dessa rättigheters, friheters och principers rättsliga värde, vilket EU:s förestående anslutning till Europakonventionen är ytterligare ett bevis på.
B. Såväl nuvarande som blivande medlemsstater liksom EU har en skyldighet att se till att innehållet och processerna i medlemsstaternas författningar överensstämmer med EU:s rättsordning och värderingar, i första hand som de kommer till uttryck i Köpenhamnskriterierna, Europeiska unionens stadga om de mänskliga rättigheterna och Europakonventionen, samt att bokstaven och andan i antagna författningar inte strider mot dessa värden och instrument.
Det gäller i första hand rättsväsendets, centralbankens och dataskyddsmyndighetens oberoende, förutsättningarna för rättvis politisk konkurrens och maktskifte liksom de s.k. stabilitetslagarna, enligt vilka beslut om systemet för inkomstbeskattning kan fattas med två tredjedels majoritet i nationalförsamlingen, samt kardinallagar som ger den rådande majoriteten i församlingen ensamrätt att tillsätta offentliga befattningar under ovanligt lång tid, med konsekvenser för framtida regeringars maktutövning.
E. Tilldelningen av mål till domstol kommer att ankomma på det nya överhuvudet för den nationella rättsliga myndigheten och högste allmänne åklagaren, en ordning som undergräver principerna om rätten att vända sig till domstol, rätten till rättvis rättegång och rättsväsendets oberoende.
F. Genom den nya författningen och dess genomförandebestämmelser döps landets högsta domstol om till ”kúria” och domstolens – nu före detta – ordförandes sexåriga tjänsteperiod avbröts i förtid efter två år.
G. Enligt den nya författningen ska den obligatoriska pensionsåldern för domare och åklagare – med undantag för kúrians ordförande och högste allmänne åklagaren – sänkas från 70 till 62 år.
I. Den ungerska nationalförsamlingen har antagit ett antal lagar med retroaktiv verkan och har därmed agerat i strid med en av de grundläggande principerna för EU:s rättsordning, nämligen att retroaktivt verkande lagstiftning inte ska antas.
J. I den nyligen antagna lagen om kyrkor och religiösa samfund ingår ovanligt stränga bestämmelser om registrering av kyrkosamfund, bl.a. ska sådan registrering vara föremål för nationalförsamlingens godkännande med två tredjedels majoritet.
K. Enligt bestämmelser i den nya författningen har den ungerska författningsdomstolens befogenheter när det gäller att granska budgetrelaterad lagstiftning reducerats avsevärt.
L. Den påfallande stora mängden lagstiftningsområden som enligt den nya författningen ska regleras genom kardinallagar, med två tredjedels majoritet i nationalförsamlingen, härunder även ärenden som bör vara föremål för ordinarie politiska förfaranden och som vanligtvis regleras genom enkel majoritet, reser ett antal farhågor, vilket bl.a. kommer till uttryck i Venedigkommissionens rapport.
P. I sitt betänkande ”Situationen för de grundläggande rättigheterna i Europeiska unionen (2009) – institutionella aspekter efter Lissabonfördragets ikraftträdande” ( 2009/2161(INI) efterlyste Europaparlamentet ”en uppföljning av kommissionens meddelande om artikel 7 i Fördraget om Europeiska unionen från 2003 för att fastställa ett transparent och enhetligt sätt att bemöta eventuella brott mot de mänskliga rättigheterna och använda artikel 7 i FEU på grundval av den nya strukturen för de mänskliga rättigheterna”.
Q. I en skrivelse till kommissionen och i ett anförande inför Europaparlamentet har Ungerns premiärminister signalerat att hans regering är beredd att åtgärda de problem som föranledde överträdelseförfarandena, ändra lagstiftningen i fråga och i övrigt samarbeta med EU:s institutioner utöver vad de rättsliga förfarandena kräver.
Europaparlamentet uttrycker allvarlig oro över situationen i Ungern för demokratin, rättsstaten, respekten för och skyddet av mänskliga och sociala rättigheter, kontrollsystemet för maktdelning, jämlikhet och icke-diskriminering.
Europaparlamentet noterar kommissionens, Europarådets och Venedigkommissionens åtagande att noga granska huruvida den ungerska lagstiftningen överensstämmer inte bara med andan utan även med bokstaven i EU:s regelverk.
a. rättsväsendets fullständiga oberoende garanteras, och i första hand att förvaltningen av den nationella rättsliga myndigheten, det allmänna åklagarämbetet och landets domstolar sker helt utan politiskt inflytande och att tjänsteperioden för domare som utsetts genom oberoende förfaranden inte kan reduceras på ett godtyckligt sätt,
b. den ungerska nationalbanken regleras i enlighet med EU:s lagstiftning,
c. det institutionella oberoendet för skyddet av personuppgifter och informationsfrihet återupprättas och garanteras i den relevanta lagens bokstav och genomförande,
d. författningsdomstolens rätt att granska all lagstiftning återupprättas helt och fullt, härmed även rätten att granska budget- och skattelagstiftning,
e. mediernas frihet och pluralism garanteras i såväl genomförandet som ordalydelsen av den ungerska medielagen, särskilt vad gäller medverkan av företrädare för det civila samhället och den politiska oppositionen i landets medieråd,
f. den nya vallagen uppfyller europeiska demokratiska normer och respekterar principen om maktskifte,
g. rätten att med demokratiska medel utöva politisk opposition såväl i som utanför institutioner garanteras,
h. lagen om kyrkor och religiösa samfund ändras så att den respekterar principerna om samvetsfrihet och inte längre kräver att nationalförsamlingen måste godkänna kyrkor med två tredjedels majoritet för att de ska kunna registreras.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, Europarådet, medlemsstaternas regeringar och parlament, byrån för grundläggande rättigheter, OSSE och FN:s generalsekreterare.
om finansiering av vetenskaplig forskning om flytande tvål med tillsatt järn
Sergio Paolo Francesco Silvestris
PE483.173v01-00 B7‑0128/2012 Förslag till Europaparlamentets resolution om finansiering av vetenskaplig forskning om flytande tvål med tillsatt järn
Europaparlamentet utfärdar denna resolution
– med beaktande av artikel 120 i arbetsordningen, och av följande skäl:
A. En av medlemsstaternas prioriteringar är att skydda det marina ekosystemet.
B. Utsläpp av tvål i havet kan ofta vara starkt förorenande och inte mindre farliga än oljeutsläpp.
Europaparlamentet uppmanar kommissionen att finansiera ytterligare forskning och försök på detta område för att undersöka egenskaperna hos flytande tvål med tillsatt järn.
SKRIFTLIG FRÅGA E-2814/05
från Hynek Fajmon (PPE-DE)
till kommissionen
(27 juli 2005)
Angående: Inrättande av Europeiska försvarsbyrån
Även om ratificeringsprocessen för fördraget om upprättande av en konstitution för Europa inte är avslutad ännu, beslutade försvarsministrarna att redan inrätta en sådan byrå, vilken formellt inledde sin verksamhet i juli 2004.
Mot denna bakgrund ber jag kommissionen besvara följande frågor: 1.
Hur är det möjligt att Europeiska försvarsbyrån kunde inrättas, utan att Fördraget om upprättande av en konstitution för Europa har trätt i kraft? 2.
Kommer Europeiska försvarsbyrån att avvecklas om Fördraget om upprättande av en konstitution för Europa inte ratificeras? 3.
Vilka finansiella medel går till Europeiska försvarsbyråns verksamhet, och varifrån kommer dessa medel?
SKRIFTLIG FRÅGA E-0576/07
från Libor Rouček (PSE) , Jan Marinus Wiersma (PSE) och Marek Siwiec (PSE)
till rådet
(13 februari 2007)
Angående: Amerikanskt missilförsvarssystem i Tjeckien och Polen
Den 20 januari 2007 rapporterade medierna att USA hade framfört en förfrågan till två EU-medlemsstater (Tjeckien och Polen) om tillstånd att placera (en del av) ett missilförsvarssystem på deras territorier.
Detta missilförsvarssystem skulle bli det första i sitt slag utanför amerikanskt territorium.
Har detta eventuella bilaterala samarbete mellan USA och de två EU-medlemsstaterna diskuterats i rådet?
Hur ställer sig rådet till den här typen av bilaterala överenskommelser?
Och hur skulle det inverka på den europeiska säkerhetsstrategin?
Den amerikanska regeringen ansåg uppenbarligen att missilförsvarssystemet även kunde bidra till att skydda europeiska länder mot eventuella anfall från Nordkorea eller Iran.
Har någon diskussion förts mellan USA och EU om ett eventuellt samarbete på detta område?
Har några transatlantiska överenskommelser ingåtts på detta område?
Tänker rådet föra upp frågan om missilförsvarssystemet på föredragningslistan för diskussionerna mellan EU och USA respektive EU och Nato?
SKRIFTLIG FRÅGA E-3431/10
från Cornelis de Jong (GUE/NGL) , Jaromír Kohlíček (GUE/NGL) , Sabine Wils (GUE/NGL) och Jacky Hénin (GUE/NGL)
till kommissionen
(14 maj 2010)
Angående: Nationella hinder för den gränsöverskridande småskaliga inlandssjöfarten
1.
Känner kommissionen till att franska fartyg för inlandssjöfart har stoppats ett antal gånger på Rhen vid Wageningen, Nederländerna, av Nationella vattenstyrelsen i Nederländerna, för att man på dessa fartyg inte behärskat det nederländska språket tillräckligt bra för kommunikationen fartyg till kust?
2.
Är den situation som avses i punkt 1 sällsynt, eller hindrar sådan språkförbistring också den gränsöverskridande inlandssjöfarten inom andra små språkområden, som Ungern och Tjeckien?
3.
Hur förklarar kommissionen att det blir allt svårare för fartyg från andra medlemsstater att få tillgång till de inre vattenvägarna i EU-medlemsstaterna?
Innebär detta att man föredrar att gränsöverskridande godstransport i allt högre grad ska ske genom vägtrafik?
Hur passar denna utveckling ihop med den politik som förordas på området för transport och miljö?
4.
Hur kan EU-medlemsstaternas agerande i fråga om inlandssjöfarten anpassas bättre inbördes, så att de små företagen inom denna sektor kan fortsätta att existera på ett drägligt sätt?
Vad gör kommissionen för att bidra till detta?
Frågor för skriftligt besvarande E-005448/2011
till kommissionen
Artikel 117 i arbetsordningen
Olga Sehnalová (S&D)
(14 juni 2011)
Angående: Märkning av batterier med tillverkningsdatum eller bäst före‑datum
Enligt min åsikt är den nuvarande EU‑lagstiftningen som avser (icke‑)märkning av ackumulatorer med tillverkningsdatum eller bäst före‑datum otillräcklig.
För närvarande är denna uppgift dold i streckkoden eller saknas helt, vilket gör det möjligt att sälja mycket gamla batterier.
Normalkonsumenten har inte möjlighet att kontrollera detta vid köpet.
Enligt tillgängliga uppgifter förlorar blyackumulatorer sin kapacitet när de ligger på lager, även om de är i så kallat torrt tillstånd.
De flesta av dem är när de säljs åtminstone delvis fyllda med elektrolyt, men ändå köper kunden en produkt med kortare livslängd än normalt.
Detta gäller även batterier med en cell, och liknande problem kan även uppträda hos fotoceller, vätedrivna bränsleceller och andra elkällor.
En meningsfull lösning skulle vara att ändra lagstiftningen så att batterierna måste vara märkta med tillverkningsdatum, varigenom batteriets kapacitet kan fastställas och livslängden garanteras.
Uppgiften om batteriets kapacitet är nämligen endast användbar om tillverkningsdatum samtidigt anges.
Hur ser kommissionen på detta problem?
Planerar kommissionen att ändra EU‑lagstiftningen så att tillverkare av ackumulatorer av alla typer blir skyldiga att märka produkterna med tillverkningsdatum eller bäst före‑datum?
Vilka andra eventuella åtgärder tänker kommissionen vidta i detta avseende?
SKRIFTLIG FRÅGA P-6294/07
från Tomáš Zatloukal (PPE-DE)
till kommissionen
(11 december 2007)
Angående: Utomhusmarknader i Tjeckien
Det finns över 50 utomhusmarknader i Tjeckien som säljer varor som vanligtvis är piratkopierade, varumärkesförfalskade eller insmugglade.
Marknaderna ligger längs gränserna mot Tyskland och Österrike och utövar en magnetisk dragningskraft på både lokalbefolkningen och utlänningar som kommer för att köpa varumärkesförfalskade och piratkopierade varor.
Dessa marknader undergräver EU:s trovärdighet då man tar upp frågor om varumärkesförfalskning och piratkopiering med tredjeländer, t.ex. med Ryssland, Kina och Ukraina.
Det är helt uppenbart en EU-fråga eftersom flera medlemsstater berörs.
Vilka åtgärder avser kommissionen att vidta för att komma åt denna varumärkesförfalskning och piratkopiering inom sina gränser?
Kommer kommissionen i sin översyn av tullförordningen eventuellt täppa till det kryphål (rådets förordning (EG) nr 1383/2003 EUT L 298, 17.11.2003, s.
– Nirj Deva och Tokia Saïfi, för PPE-DE-gruppen
– Miguel Angel Martínez Martínez, för PSE-gruppen
– Fiona Hall och Thierry Cornillet, för ALDE-gruppen
– Caroline Lucas, Frithjof Schmidt och Margrete Auken, för Verts/ALE-gruppen
– Luisa Morgantini, Gabriele Zimmer, Feleknas Uca och Vittorio Agnoletto, för GUE/NGL-gruppen
– Eoin Ryan, Roberta Angelilli och Ģirts Valdis Kristovskis, för UEN-gruppen
som ersätter resolutionsförslagen från följande grupper:
– PPE-DE (B6‑0119/2006)
– GUE/NGL (B6‑0121/2006)
– ALDE (B6‑0124/2006)
– PSE (B6‑0142/2006)
– Verts/ALE (B6‑0143/2006)
om nya ekonomiska instrument för utveckling i samband med millennieutvecklingsmålen
Europaparlamentets resolution om nya ekonomiska instrument för utveckling i samband med millennieutvecklingsmålen
Europaparlamentet utfärdar denna resolution
–
med beaktande av den internationella konferensen om innovativa källor till biståndsfinansiering, avsedd att hållas den 28 februari–1 mars 2006 i Paris,
–
med beaktande av millennieutvecklingsmålen och FN:s sammankomst på hög nivå i september 2005 för översyn av framstegen på väg mot millennieutvecklingsmålen,
–
med beaktande av Landaurapporten om nya internationella ekonomiska bidrag till utveckling, en rapport som givits i uppdrag i november 2003 av president Chirac,
–
med beaktande av New York-deklarationen om åtgärder mot hunger och fattigdom, vilken undertecknats av över 120 länder vid FN:s generalförsamling 2004,
–
med beaktande av Förenade kungarikets finansminister Gordon Browns förslag om en internationell finansieringsmekanism, något som kunde leda till en fördubbling av utvecklingsbiståndet,
–
med beaktande av solidaritetsavgiften på franska flygbiljetter, vilken kommer att träda i kraft den 1 juli 2006,
–
med beaktande av kommissionens dokument med en undersökning av hur en eventuell avgift på flygbiljetter kunde fungera som ny källa till biståndsfinansiering,
–
med beaktande av den ”förklaring om innovativa källor till biståndsfinansiering”, som undertecknats av 79 regeringar före FN:s sammankomst på hög nivå i september 2005 för översyn av millennieutvecklingsmålen,
–
A.
För att man skall kunna bryta spiralen av fattigdom och ge utvecklingsländerna medel att förverkliga sina inneboende ekonomiska möjligheter och gå med i globaliseringen behövs det ofrånkomligen en sund utvecklingspolitik som stöds av ett massivt och verkningsfullt utvecklingsbistånd.
B.
Hur mycket man än ger i utvecklingsbistånd kommer man på det sättet aldrig att få bukt med fattigdomen i utvecklingsländerna, förrän dessa har tillräcklig kapacitet för att ta emot biståndet, genomföra en sund förvaltning och bekämpa korruptionen.
C.
I rapporten om framsteg på väg mot millennieutvecklingsmålen 2005 finns det klara belägg för att man inte kommer att kunna hjälpa de fattiga länderna att nå dessa mål fram till den fastställda tidsgränsen 2015, om man inte tar på sig ytterligare politiska och ekonomiska åtaganden, i fråga såväl om biståndets kvantitet som dess kvalitet.
D.
I New York-deklarationen om åtgärder mot hunger och fattigdom uppmanas regeringarna i de utvecklade länderna att ingå konkreta åtaganden för finansiering av millennieutvecklingsmålen.
E.
F.
Enligt Världsbankens uppskattningar kommer det att behövas minst 50 miljarder USD mer per år i offentligt utvecklingsbistånd för att millennieutvecklingsmålen skall kunna nås.
G.
Bidragen till världsfonden för kampen mot aids, tuberkulos och malaria uppgick till mindre än 15 procent av vad som hade behövts.
H.
I.
1.
Europaparlamentet välkomnar den konferens som skall hållas i Paris den 28 februari–1 mars, med avsikt att det skall göras framsteg i riktning mot en överenskommelse om internationella avgifter och särskild inriktning på en eventuell avgift på flygbiljetter.
2.
Europaparlamentet vidhåller att eventuella alternativa metoder för biståndsfinansiering måste leda till att det frigörs ytterligare nya medel för biståndet och inte ersätta det offentliga utvecklingsbiståndet.
3.
Europaparlamentet välkomnar varmt rådets överenskommelse från i juni 2005 om att fördubbla EU:s bistånd till utvecklingsländerna samt om att medlemsstaterna skall öka sitt officiella utvecklingsbistånd till 0,56 procent av BNI senast 2010 och 0,7 procent av BNI senast 2015.
4.
5.
Europaparlamentet uppmanar de utvecklade länderna att fullgöra sina åligganden och uppfylla sina åtaganden om att i statsbudgetarna höja anslagen till utvecklingsbistånd till 0,7 procent av BNI.
6.
7.
8.
9.
10.
11.
Europaparlamentet uppmanar EU:s institutioner och regeringarna inom EU att grundligt utreda om åtgärderna mot hunger skulle kunna finansieras med hjälp av ett världslotteri, såsom det förslagits av FN:s världslivsmedelsprogram i form av ett livsmedelsprojekt.
12.
Europaparlamentet understryker att man i dagens ytterst ansträngda budgetläge behöver unionsmedborgarnas fulla stöd, för att eventuella nya initiativ skall kunna handhas med omsorg så att det inte uppstår risker för att allmänna opinionen i Europa inte längre skall acceptera utvecklingspolitikens mål.
13.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, EU:s alla statsöverhuvuden, FN:s generalsekreterare, FN:s särskilda sändebud för millennieutvecklingsmålen, Världsbanken och OECD:s sekretariat.
– Astrid Lulling och Bernd Posselt, för PPE-DE-gruppen
– Pasqualina Napoletano och Martine Roure, för PSE-gruppen
– Graham Watson, Alexander Lambsdorff och Cecilia Malmström, för ALDE‑gruppen
– Raül Romeva i Rueda och Eva Lichtenberger, för Verts/ALE-gruppen
– Bastiaan Belder, för IND/DEM-gruppen
– Cristiana Muscardini, Konrad Szymański och Roberts Zīle, för UEN-gruppen
som ersätter resolutionsförslagen från följande grupper:
– ALDE (B6‑0284/2006)
– Verts/ALE (B6‑0285/2006)
om Taiwan
Europaparlamentets resolution om Taiwan
Europaparlamentet utfärdar denna resolution
–
med beaktande av sin resolution av den 14 mars 2002 om Taiwans observatörsstatus vid Världshälsoförsamlingens årliga möte i maj 2002 i Genève,
–
med beaktande av sin resolution av den 15 maj 2003 om observatörsstatus för Taiwan vid WHO:s 56:e möte,
–
med beaktande av sitt betänkande av den 5 september 2002 om kommissionens meddelande ”Europa och Asien: en strategisk ram för förbättrade partnerskap”, där det konstaterades att det behövs ett nära samarbete med Asien inom multilaterala organisationer, exempelvis för att inom ramen för WHO bekämpa aids/hiv i regionen, och att alla demokratier i Asien, även Taiwan, därför bör kunna delta i WHO,
–
med beaktande av sin resolution av den 7 juli 2005 om förbindelserna mellan EU, Kina och Taiwan samt säkerheten i Fjärran Östern,
–
A.
Det är nödvändigt att alla delar av världen har möjlighet att direkt och obehindrat delta i internationella samarbetsnätverk, forum och program på hälso- och sjukvårdsområdet, i synnerhet med tanke på att det i dag är lättare för olika infektionssjukdomar (som fågelinfluensa och sars) att sprida sig över gränserna.
B.
WHO har gjort det möjligt för observatörer att delta i dess verksamhet.
C.
Kommissionen har också redan ställt sig positiv till att förbättra kontakterna mellan Taiwan och WHO, i den mån WHO:s bestämmelser medger detta, och är intresserad av att finna en ”praktisk lösning” tillsammans med medlemsstaterna.
D.
Den största risken för en influensapandemi kommer från asiatiska länder, där ett mycket patogent fågelinfluensavirus har spridits i två år trots behöriga myndigheters oavbrutna insatser för att hejda sjukdomen.
E.
Infektionssjukdomar som hiv/aids, tuberkulos, malaria och sars når allt större utbredning över hela världen.
F.
En pandemi utanför EU skulle även utgöra ett allvarligt hot mot EU-medborgarnas hälsa.
G.
H.
Taiwans hälso- och sjukvård är en av de bästa och mest avancerade i regionen, och de taiwanesiska myndigheterna vill låta sina specialister delta i WHO:s förberedande expertmöten om situationen när det gäller fågelinfluensan.
1.
Europaparlamentet kräver att Taiwan skall bli bättre representerat i internationella organisationer och anser det orättvist att fortsätta att utesluta mer än 20 miljoner människor från världssamfundet.
2.
Europaparlamentet uppmanar WHO:s generaldirektör att omedelbart låta Taiwans centrum för sjukdomskontroll (Taiwan CDC) ingå i WHO:s globala nätverk för varningar och motåtgärder (GOARN), så att snabbt utbyte av relevant information kan möjliggöras på regional och global nivå.
3.
Europaparlamentet uppmanar WHO:s generaldirektör och alla dess medlemsstater att se till att Taiwan får direkt tillträde till och kan närvara vid alla WHO:s tekniska möten som är av betydelse för att den offentliga hälso- och sjukvården skall kunna upprätthållas och förbättras både i Taiwan och i resten av världen samt att låta Taiwan delta på meningsfullt vis i den tekniska verksamhet och de arrangemang som WHO:s berörda regionkontor anordnar.
4.
Europaparlamentet uppmanar Folkrepubliken Kina att undersöka alla möjligheter att ge Taiwan observatörsstatus i Världshälsoorganisationen eller åtminstone i Världshälsoförsamlingen, dess viktigaste beslutsfattande organ, för att skydda hälsan hos det taiwanesiska folket, hos internationella representanter och utländska arbetstagare på ön liksom hos hela världens befolkning.
5.
Europaparlamentet upprepar sin uppmaning till kommissionen och medlemsstaterna att stödja Taiwans ansökan om observatörsstatus i WHO.
6.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, medlemsstaternas och anslutningsländernas regeringar och parlament, Folkrepubliken Kinas regering och parlament, Taiwans myndigheter, FN:s generalsekreterare samt WHO:s generaldirektör.
– Hubert Pirker, Georg Jarzembowski, Bernd Posselt, Charles Tannock och Albert Jan Maat för PPE-DE-gruppen
– Pasqualina Napoletano för PSE-gruppen
– István Szent-Iványi, Marios Matsakis och Frédérique Ries för ALDE-gruppen
– Gérard Onesta och Gisela Kallenbach för Verts/ALE-gruppen
– Giusto Catania och Jonas Sjöstedt för GUE/NGL-gruppen
– Bastiaan Belder för IND/DEM-gruppen
som ersätter resolutionsförslagen från följande grupper:
– ALDE ( B6‑0341/2006 )
– GUE/NGL ( B6‑0361/2006 )
– PSE ( B6‑0363/2006 )
– PPE-DE ( B6‑0366/2006 )
– IND/DEM ( B6‑0368/2006 )
– Verts/ALE ( B6‑0369/2006 )
om Nordkorea
Europaparlamentets resolution om Nordkorea
Europaparlamentet utfärdar denna resolution
–
med beaktande av sina tidigare resolutioner om Nordkorea,
–
med beaktande av EU:s riktlinjer om dödsstraff gentemot tredje land (1998), om tortyr och annan omänsklig eller förnedrande behandling (2001), om människorättsdialog med tredjeländer (2001) och om människorättsförsvarare (2004),
–
med beaktande av resolutionen av den 16 april 2003 från FN:s människorättskommission,
–
med beaktande av uttalandet av den 31 maj 2006 från FN:s särskilde rapportör för utomrättsliga, summariska eller godtyckliga avrättningar, ordföranden och rapportören i FN:s arbetsgrupp för godtyckligt frihetsberövande, FN:s särskilde rapportör för tortyrfrågor och FN:s särskilde rapportör för människorättsläget i Nordkorea,
–
A.
FN:s människorättskommission uttrycker i sin resolution djup oro över Nordkoreas tillämpning av tortyr och annan grym, omänsklig eller förnedrande behandling eller bestraffning samt offentliga avrättningar liksom över landets omfattande och allvarliga inskränkningar av tankefriheten, samvetsfriheten, religionsfriheten, åsiktsfriheten och yttrandefriheten.
B.
C.
Ingen form av opposition tillåts och alla personer som uttrycker en åsikt som strider mot det regerande nordkoreanska arbetarpartiets riskerar stränga straff, vilket i många fall även deras familjemedlemmar gör.
D.
Son Jong Nam, som bott i Kina och gått i kyrkan och blivit kristen i landet, skall enligt rapporter ha torterats av den nationella säkerhetstjänsten och sedan dömts till döden för påstått högförräderi, utan rättegång och utan tillgång de rättsliga garantier som krävs i internationell humanitär rätt.
E.
Fyra FN-experter på människorättsområdet, däribland den särskilde rapportören för människorättsläget i Nordkorea, som uppmanat Nordkoreas regering att skjuta upp avrättningen och ompröva domen, har med bestörtning tagit emot regeringens svar, i vilket deras skrivelse betecknas som ett led i en konspiration med det illasinnade syftet att sprida falska uppgifter och bistå de fientliga krafter som vill förtala, sönderdela och störta den nordkoreanska staten och dess sociala system med mänskliga rättigheter som förevändning.
F.
Nordkorea har ratificerat den internationella konventionen om medborgerliga och politiska rättigheter.
G.
Nordkoreas regering har sedan 2001 minskat antalet brott som föranleder dödsstraff från 33 till fem, men fyra av dessa brott är huvudsakligen av politisk natur.
H.
I.
J.
Vittnen uppskattar antalet människor som befinner sig i ”omskolningsläger” (arbetsläger), fångläger och fängelser till upp till 200 000, och rapporter från bland annat personer som nyligen frigivits från läger som Kang Chol Hwan vittnar om omfattande tortyr och misshandel och om mycket svåra förhållanden.
K.
Många människor i Nordkorea lider brist på mat och är beroende av det humanitära bistånd som landet får från givare som EU, som beslutade att anslå 13 715 000 euro till Nordkorea under 2005, och FN:s världslivsmedelsprogram, som den 10 maj 2006 nådde en överenskommelse med regeringen om att förse 1,9 miljoner nordkoreaner med 150 000 ton förnödenheter under två års tid.
L.
Tiotusentals nordkoreaner har flytt till Kina och lämnat sitt land på grund av förtryck och omfattande hungersnöd.
1.
Europaparlamentet beklagar att Nordkorea inte samarbetar med internationella institutioner på människorättsområdet och framför allt att landet vägrar att följa de förfaranden som FN:s människorättskommission föreskriver.
2.
Europaparlamentet uppmanar Nordkoreas regering att
∙ efterleva principerna i de fördrag inom ramen för internationell humanitär rätt som landet ratificerat (exempelvis den internationella konventionen om medborgerliga och politiska rättigheter) och att införliva dessa principer i sin nationella lagstiftning,
∙ avskaffa dödsstraffet,
∙ frige alla människor som frihetsberövats eller fängslats sedan de fredligt utövat sina grundläggande mänskliga rättigheter,
∙ garantera yttrande- och rörelsefriheten för alla nordkoreaner,
∙ se över befintlig lagstiftning så att den görs förenlig med normerna i internationell humanitär rätt och införa säkerhetsmekanismer för att ge medborgarna skydd och rättsmedel mot människorättsbrott.
3.
Europaparlamentet uppmanar Nordkoreas regering att lämna information om fallet med Son Jong Nam och att stoppa hans avrättning.
4.
Europaparlamentet uppmanar kommissionen och rådet att kräva att Nordkoreas regering upphör med sina brott mot de mänskliga rättigheterna, lämnar information om fallet med Son Jong Nam och stoppar hans avrättning.
5.
Europaparlamentet uppmanar Nordkoreas regering att noga se över situationen för alla dem som dömts till döden och att bevilja uppskov med avrättningen och kräver att FN:s särskilde rapportör för människorättsläget i Nordkorea, Vitit Muntarbhorn, skall tillåtas besöka dem.
6.
Europaparlamentet uppmanar med eftertryck Nordkoreas regering att upphöra med de svåra brott mot de mänskliga rättigheterna – bland annat fängslingarna och avrättningarna på grund av religion eller tro – som drabbar medborgare som inte tillhör de statligt understödda religiösa sammanslutningarna, och att låta troende personer mötas för att utöva sin tro, inrätta och underhålla platser för religiös verksamhet och fritt ge ut religiös litteratur.
7.
8.
Europaparlamentet uppmanar Nordkoreas regering att fullgöra sina skyldigheter enligt de akter på människorättsområdet som den anslutit sig till och att se till att humanitära organisationer, oberoende människorättsinspektörer, FN:s särskilde rapportör för människorättsläget i Nordkorea och FN:s särskilde rapportör för religions- och trosfrihet har fritt tillträde till landet.
9.
10.
Europaparlamentet uppmanar Nordkoreas regering att slutgiltigt och utan inskränkningar lämna över all information om de medborgare i Sydkorea och Japan som bortförts under de senaste årtiondena och att omedelbart frige de bortförda personer som fortfarande kvarhålls i landet.
11.
12.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, Nordkoreas regering, Sydkoreas regering, Kinas regering, FN:s särskilde rapportör för utomrättsliga, summariska eller godtyckliga avrättningar, ordföranden och rapportören för FN:s arbetsgrupp för godtyckligt frihetsberövande, FN:s särskilde rapportör för tortyrfrågor och FN:s särskilde rapportör för människorättsläget i Nordkorea.
GEMENSAMT FÖRSLAG TILL RESOLUTION
– Godelieve Quisthoudt-Rowohl, Ria Oomen-Ruijten och Maria Martens, för PPE-DE-gruppen
– Antolín Sánchez Presedo, Jan Andersson, Erika Mann och Stephen Hughes, för PSE-gruppen
– Jean-Louis Bourlanges och Bernard Lehideux, för ALDE-gruppen
– Caroline Lucas och Jean Lambert, för Verts/ALE-gruppen
– Helmuth Markov, för GUE/NGL-gruppen
– Mieczysław Edmund Janowski, Eugenijus Maldeikis och Roberta Angelilli, för UEN-gruppen
som ersätter resolutionsförslagen från följande grupper:
– GUE/NGL ( B6‑0578/2006 )
– PPE-DE ( B6‑0579/2006 )
– UEN ( B6‑0580/2006 )
– Verts/ALE ( B6‑0581/2006 )
– PSE ( B6‑0582/2006 )
– ALDE ( B6‑0583/2006 )
om Europeiska unionens allmänna preferenssystem
Europaparlamentets resolution om Europeiska unionens allmänna preferenssystem
Europaparlamentet utfärdar denna resolution
–
–
med beaktande av kommissionens beslut 2005/924/EG EUT L 337, 22.12.2005, s.
–
A.
Den särskilda stimulansordningen för hållbar utveckling och gott styre (GSP+) ger varor från utvecklingsländer, som tillämpar vissa internationella standarder för mänskliga rättigheter, arbetstagares rättigheter, miljöskydd, narkotikabekämpning och gott styre, förmånstillträde till europeiska marknader.
B.
Bland kriterierna för att erhålla tullförmåner enligt GSP+ ingår ratificering och effektivt genomförande av centrala FN- och ILO-konventioner samt miljöavtal, enligt förteckningen i del A i förordningens bilaga III.
C.
Kommissionen beviljade i sitt beslut av den 21 december 2005 förmåner enligt den särskilda stimulansordningen till Bolivia, Colombia, Costa Rica, Ecuador, Georgien, Guatemala, Honduras, Sri Lanka, Moldavien, Mongoliet, Nicaragua, Panama, Peru, El Salvador och Venezuela.
D.
Det nya GSP+-systemet bör fungera som incitament för förmånsländerna att uppnå utvecklingsmål, inklusive inrättandet av lämpliga institutioner för att fullt ut respektera de rättigheter som följer av FN:s och ILO:s konventioner.
E.
Effektiviteten i genomförandet av de aktuella FN- och ILO-konventionerna bör utvärderas regelbundet genom de slutsatser som dras av behöriga övervakningsorgan, bland annat i den årliga rapporten från ILO:s expertkommitté för tillämpning av konventioner och rekommendationer, och vederbörlig hänsyn bör tas till Europaparlamentets ståndpunkt.
F.
Enligt artikel 16 i förordningen om Allmänna preferenssystemet (GSP) kan skyddsklausuler och tillfälliga upphävanden tillämpas för länder som allvarligt och systematiskt kränker bestämmelserna i de internationella konventioner som finns uppräknade i bilaga III i rådets förordning (EG) nr 980/2005.
1.
Europaparlamentet noterar kommissionens beslut att bevilja förmåner enligt GSP+ till de länder som är uppräknade i kommissionens beslut 2005/924/EG.
2.
Europaparlamentet konstaterar att den ekonomiska utvecklingen i de länder som omfattas av GSP+ och deras integration i det globala handelssystemet är avgörande för att uppnå målsättningarna om en hållbar utveckling, inklusive stabilitet och god samhällsstyrning.
3.
4.
Europaparlamentet konstaterar att uppgifter förekommit om upprepade fall av överträdelser av arbetstagarnas rättigheter i flera av de länder som ratificerat de aktuella ILO‑konventionerna, och att dessa överträdelser, om de visar sig utgöra allvarliga och systematiska kränkningar av ILO:s grundläggande arbetstagarrättigheter, i enlighet med artikel 16 i förordningen skulle kunna motivera ett tillfälligt upphävande av GSP+‑förmånerna.
5.
Europaparlamentet uppmanar kommissionen att skärpa sin övervakning av genomförandet av ILO:s konventioner samt konventioner om miljö och god samhällsstyrning i GSP+-länderna, och att i synnerhet fullgöra sina skyldigheter enligt artikel 18 i förordningen, nämligen informera kommittén för allmänna tullförmåner om de brott mot arbetstagarnas rättigheter och miljökonventionerna som rapporterats och samråda om huruvida en undersökning bör genomföras av om det förekommit allvarliga och systematiska kränkningar av ILO:s konventioner om grundläggande arbetstagarrättigheter, särskilt när det gäller barnarbete och tvångsarbete.
6.
7.
Europaparlamentet uppmanar kommissionen att regelbundet informera parlamentet om vad den har kommit fram till under sin övervakning av tillämpningen av FN- och ILO‑konventionerna och efterlevnadsnivån i GSP+-länderna, särskilt på områdena föreningsfrihet, kollektiva förhandlingar, icke-diskriminering i arbetslivet och avskaffande av barn- och tvångsarbete, och framför allt uppge om det i något av de nuvarande GSP+‑länderna förekommer allvarliga och systematiska kränkningar av de principer som fastlagts i internationella konventioner om de mänskliga rättigheterna och arbetstagarnas rättigheter samt miljöavtal.
8.
9.
10.
Europaparlamentet uppmanar kommissionen att varje år utarbeta en heltäckande rapport där varje enskilt land behandlas och inte bara situationen i förmånsländerna beskrivs utan även kommissionens åtgärder.
11.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet och kommissionen.
GEMENSAMT FÖRSLAG TILL RESOLUTION
– Michael Gahler, Mario Mauro och Bernd Posselt, för PPE-DE-gruppen
– Pasqualina Napoletano och Ana Maria Gomes, för PSE-gruppen
– Marios Matsakis, för ALDE-gruppen
– Marie-Hélène Aubert, Margrete Auken och Raül Romeva i Rueda, för Verts/ALE-gruppen
– Luisa Morgantini, för GUE/NGL-gruppen
– Eoin Ryan, Roberts Zīle, Michał Tomasz Kamiński, Adam Jerzy Bielan och Romano Maria La Russa, för UEN-gruppen
som ersätter resolutionsförslagen från följande grupper:
– GUE/NGL ( B6‑0596/2006 )
– UEN ( B6‑0598/2006 )
– ALDE ( B6‑0600/2006 )
– PSE ( B6‑0603/2006 )
– PPE-DE ( B6‑0606/2006 )
– Verts/ALE ( B6‑0613/2006 )
om Etiopien
Europaparlamentets resolution om Etiopien
Europaparlamentet utfärdar denna resolution
–
med beaktande av sina tidigare resolutioner om den kris som uppstått efter valet och de allvarliga kränkningarna av de mänskliga rättigheterna i Etiopien, och särskilt resolutionerna av den 7 juli 2005 om mänskliga rättigheter i Etiopien, av den 13 oktober 2005 om situationen i Etiopien, och av den 15 december 2005 om situationen i Etiopien och den nya gränskonflikten,
–
A.
Två tjänstemän från Europeiska kommissionen har arresterats och utvisats från Etiopien under förevändningen att ha försökt att hjälpa Yalemzewd Bekele, advokat och kvinnorättsaktivist, som arbetar för Europeiska kommissionen i Addis Abeba, att ta sig ut ur landet.
B.
Enligt rapporter förekommer det fortfarande arresteringar, trakasseringar, godtyckliga frihetsberövanden, förnedring av och hot mot oppositionspolitiker samt mot personer verksamma inom det civila samhället, studenter och andra vanliga medborgare.
C.
Efter att EU intervenerat på hög nivå för att få Yalemzewd Bekele frisläppt, frigavs hon den 27 oktober 2006, efter att ha kvarhållits utan kontakt med yttervärlden under ett par dagar.
D.
Det etiopiska parlamentet inrättade en regeringsstödd utredningskommission i slutet av november 2005 som fått i uppdrag att utreda morden i juni och november 2005.
E.
Medlemmar av utredningskommissionen utsattes för påtryckningar av den etiopiska regeringen att göra ändringar i utredningens slutsatser och tre av dem, inkluderande ordföranden och vice ordföranden, har lämnat landet efter att ha motsatt sig regeringens order att ändra slutsatserna i den slutgiltiga rapporten.
F.
Dessa tjänstemän har lyckats lämna landet med den slutgiltiga rapporten, som i kraftfulla ordalag fördömer regeringens handläggning av krisen som krävt 193 människoliv i samband med demonstrationerna i juni och november 2005.
G.
Till följd av massarresteringarna av regeringsmotståndare, människorättsaktivister och journalister i samband med demonstrationerna i juni och november 2005, hålls fortfarande 111 oppositionsledare, journalister och människorättsaktivister fängslade, anklagade bl.a. för ”grov kränkning av konstitutionen”, ”uppvigling, organisering eller ledning av väpnat uppror” och ”försök till folkmord”.
H.
I.
Senaste tidens arresteringar av Wassihun Melese och Anteneh Getne, medlemmar av Etiopiska lärarförbundet, och dessa nya arresteringar förefaller att utgöra en reaktion på lärarförbundets beskyllningar mot regeringen om inblandning i dess verksamhet och hot mot dess ledare.
J.
Premiärminister Meles Zenawi är en av Europeiska kommissionens gäster vid de Europeiska utvecklingsdagar som anordnas 13-17 november 2006 i Bryssel.
K.
Etiopien har undertecknat partnerskapsavtalet mellan AVS-länderna, å enda sidan, och Europeiska kommissionen och dess medlemsstater, å andra sidan, vars artikel 96 (Cotonouavtalet) föreskriver att respekten för de mänskliga rättigheterna och de grundläggande friheterna utgör ett viktigt element i AVS-EU samarbetet.
1.
Europaparlamentet välkomnar EU:s ansträngningar att försöka få Yalemzewd Bekele frigiven och beklagar djupt att Bjorn Jonsson och Enrico Sborgi, två EU-tjänstemän som arbetat i Etiopien, utvisats.
2.
Europaparlamentet uppmanar Etiopiens regering att omedelbart och utan ändringar offentliggöra utredningskommissionens slutgiltiga rapport i dess helhet.
Europaparlamentet uppmanar berörda domstolar att införskaffa rapporten och ta vederbörlig hänsyn till denna så att en rättvis rättegång kan hållas.
3.
Europaparlamentet uppmanar de etiopiska myndigheterna att avhålla sig från hot och trakasserier mot nationella ledare, inkluderande domare vid domstol och medlemmar av lärarförbundet, i samband med utövandet av de skyldigheter som åligger dem genom yrket.
4.
5.
6.
Europarlamentet uppmanar den etiopiska regeringen att respektera den allmänna förklaringen om mänskliga rättigheter och den Afrikanska unionens stadga om mänskliga rättigheter och folkens rättigheter, inkluderande rätten till fredliga sammankomster, yttrandefrihet, samt garantera rättsväsendets oberoende.
Europaparlamentet uppmanar kommissionen och rådet att ingående följa situationen i Etiopien och anser att utarbetandet av samarbetsprogram inom ramen för Cotonouavtalet skall vara beroende av huruvida mänskliga rättigheter och principen om god förvaltning respekteras, vilket klart framgår av klausulen om att respekt för dessa faktorer utgör en ”väsentlig beståndsdel” av avtalet.
9.
Europaparlamentet uppmanar kommissionen och rådet att utreda på vilket sätt det går att få igång en övergripande dialog mellan olika parter i Etiopien under medverkan av politiska partier, det civila samhällets organisationer och alla intressenter för att kunna få till stånd en hållbar lösning på den nuvarande politiska krisen.
10.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, Etiopiens regering, FN:s generalsekreterare och Afrikanska unionen.
– Françoise Grossetête och Hans-Gert Poettering, för PPE-DE-gruppen
– Martin Schulz och Hannes Swoboda, för PSE-gruppen
– Silvana Koch-Mehrin och Graham Watson, för ALDE-gruppen
– Pierre Jonckheer, Monica Frassoni och Daniel Cohn-Bendit, för Verts/ALE‑gruppen
– Brian Crowley, Roberta Angelilli, Zdzisław Zbigniew Podkański, Roberts Zīle och Gintaras Didžiokas, för UEN-gruppen
som ersätter resolutionsförslagen från följande grupper:
– Verts/ALE ( B6‑0630/2006 )
– ALDE ( B6‑0634/2006 )
– UEN ( B6‑0635/2006 )
– PPE-DE ( B6‑0640/2006 )
– PSE ( B6‑0642/2006 )
om kommissionens lagstiftnings- och arbetsprogram för 2007 (KOM(2006)0629)
Europaparlamentets resolution om kommissionens lagstiftnings- och arbetsprogram för 2007 (KOM(2006)0629)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens meddelande av den 24 oktober 2006 om sitt lagstiftnings- och arbetsprogram för 2007, som lades fram av kommissionen och diskuterades under parlamentets sammanträdesperiod i november,
–
med beaktande av kommissionens strategiska politiska riktlinjer för 2004–2009, kommissionens årliga politiska strategi för 2007 och de bidrag från parlamentsutskotten som överlämnats till kommissionen av talmanskonferensen, i överensstämmelse med ramavtalet mellan parlamentet och kommissionen,
–
A.
B.
Det är oerhört viktigt att kommissionen förmår uppnå ambitiösa politiska, ekonomiska och sociala mål för medborgarna och att man tillvaratar de europeiska gemensamma intressena genom att göra unionen till en ledande global aktör som verkar för gemensamma lösningar såsom fred, säkerhet, globalt välstånd och en hållbar ekonomisk och social utveckling.
C.
Det är angeläget att anpassa utgifterna efter de politiska prioriteringarna, eftersom de medel som tillhandahålls i den nya budgetplanen är otillräckliga för att möta alla utmaningar framöver.
D.
Det är nödvändigt att EU vidtar åtgärder för att infria medborgarnas ökade förväntningar och för att förstärka sin roll som ledande aktör på världsnivå.
1.
2.
3.
Europaparlamentet gläds åt att kommissionen har ställt sig bakom flera av de förslag som parlamentsutskotten har lagt fram i samband med den nya ”strukturerade dialogen” och som beskrivs i utskottsordförandekonferensens kortfattade rapport.
4.
Europaparlamentet ber dock kommissionen att informera parlamentet om varför man i arbetsprogrammet för 2007 inte inkluderade följande lagstiftningsinitiativ som föreslogs av parlamentets utskott: ömsesidigt erkännande inom varuhandeln, förslag om förbättring av EU-märkningen, revidering av stadgan för Europabolag, utveckling av mikrolån, möjligheter att kombinera yrkes- och familjeliv, skydd för arbetstagare med atypiska anställningsformer, ett nytt förslag till europeiska ömsesidiga bolag, gränser för utsäde innehållande genmodifierade organismer och ett förslag avseende initiativet om insyn.
5.
Europaparlamentet anser att tillämpningen av ramavtalet om förbindelserna mellan parlamentet och kommissionen kan och bör förbättras genom att man engagerar de politiska grupperna på ett mer konsekvent sätt och i ett tidigt stadium av förfarandet.
6.
Parlamentet efterlyser, i överensstämmelse med ramavtalet mellan Europaparlamentet och kommissionen, en bättre samordning mellan de båda förfarandena, och ser fram emot en diskussion om hur detta kan uppnås.
7.
Europaparlamentet uppmanar kommissionen att i ett tidigt skede inleda en dialog med parlamentet om den mycket viktiga översynen av EU:s budgetram och av budgetplanen, halvtidsöversynen av den gemensamma jordbrukspolitiken och diskussionen om nya mekanismer för de egna resurserna.
8.
9.
10.
11.
Prioriteringar för 2007
Modernisera EU:s ekonomi
12.
13.
Europaparlamentet uppmanar kommissionen att förbättra samordningen av den ekonomiska politiken, särskilt när det gäller att främja nationella och europeiska initiativ som syftar till att stödja forskning, kompetens och ny teknik och när det gäller att utbyta bästa praxis om hur man kan förbättra effektiviteten och kvaliteten i de offentliga utgifterna och att förbättra statistikens kvalitet.
Forskning och utveckling
14.
Europaparlamentet påpekar att det är hög tid att stödja samordnad forskningsverksamhet för att förbättra den europeiska ekonomins konkurrenskraft, inte minst på området för avancerad teknik, och efterlyser fler samordnade insatser för att främja telekommunikations- och IT‑sektorerna.
15.
16.
17.
Europaparlamentet understryker den strategiska betydelsen av en mycket expansiv rymdsektor och stöder därmed helhjärtat kommissionens initiativ att utarbeta en sammanhängande och övergripande europeisk rymdpolitik.
Inre marknad
18.
19.
Europaparlamentet begär återigen att kommissionen skall utforska alla tänkbara möjligheter att förbättra patentsystemet och systemet för att lösa patenttvister.
20.
Bemöta de samhälleliga utmaningarna i EU
21.
22.
Europaparlamentet efterlyser en lämplig uppföljning av kommissionens meddelande om aktiv integration av de personer som befinner sig längst ifrån arbetsmarknaden.
23.
Europaparlamentet uppmanar kommissionen att utarbeta en tydlig rättslig grund för kampen mot alla former av våld, särskilt mot kvinnor och barn.
24.
Parlamentet välkomnar i detta sammanhang kommissionens avsikt att undersöka olika vägar att förstärka flexicurityn och hjälpa medlemsstaterna att uppnå både en hög produktivitet och ett gott socialt skydd.
Konsumentskydd
25.
26.
Europaparlamentet välkomnar därför handlingsplanen för hållbar produktion och konsumtion, eftersom den innehåller både den sociala och ekonomiska dimensionen.
Medborgarnas säkerhet, rättvisa och migration
27.
Europaparlamentet efterlyser ett åtagande från EU:s medlemsstater och från kommissionen att ta itu med de strukturella orsakerna till de stora migrationsströmmarna genom att anpassa och uppdatera sin nuvarande politik för att göra det möjligt för utvecklingsländerna att skydda och bygga upp sina ekonomier och garantera rimliga inkomster för sina befolkningar, vilket är det enda alternativet om man vill minska den illegala invandringen.
28.
29.
30.
31.
32.
Europaparlamentet påpekar att det är angeläget att bekämpa IT-brottslighet och förbättra gränskontrollerna och handläggningen av visumansökningarna, och betonar vikten av ett snabbt ikraftträdande av både SIS II och VIS.
33.
Europaparlamentet uppmanar kommissionen att 2007 lägga fram ett förslag till rapport om hur säsongarbetares rättigheter i EU kan skyddas, för att undvika missbruk och överträdelser av grundläggande arbetsmarknadsnormer, vilket förekommer i dagsläget.
34.
Trygg, konkurrenskraftig och hållbar energi
35.
Europaparlamentet välkomnar kommissionens förslag om att göra utvecklingen av den europeiska energipolitiken till ett strategiskt mål för 2007 med utgångspunkt i principerna om en tryggad och diversifierad försörjning, hållbarhet, effektivitet och större energiberoende.
36.
37.
38.
Europaparlamentet uppmanar medlemsstaterna att skapa en inre energimarknad i EU genom att skapa jämvikt mellan inre och yttre försörjningskällor och säkra driftskompatibiliteten mellan nationella kraftledningsnät.
39.
Europaparlamentet uppmanar kommissionen att utveckla en bättre samverkan mellan å ena sidan ekonomisk utveckling och å ena sidan utveckling och användning av ren och energisnål teknik, eftersom det finns stark komplementaritet och detta utgör en potentiell källa till ökad konkurrenskraft.
Göra Europa till en bättre plats att leva i
Miljö och hållbar utveckling
40.
41.
Europaparlamentet uppmanar kommissionen att stödja en stark roll för EU vid utformningen av politiska strategier och nya mål efter Kyoto.
42.
43.
Europaparlamentet uppmanar kommissionen att bättre samordna transport- och miljöpolitiken i syfte att uppnå en hållbar utveckling, och att föreslå konkreta mål för minskningen av koldioxidutsläppen för hela fordonsparken samt att inkludera flygtransporterna i de bindande åtagandena i Kyotoprotokollet.
44.
45.
Hälsa
46.
Europaparlamentet välkomnar kommissionens bidrag när det gäller att mejsla ut EU:s hälsopolitik, och är fast beslutet om att skyddet och främjandet av hälsan bör vara ett centralt inslag i EU-politiken.
47.
Europaparlamentet betonar att en effektiv europeisk hälsostrategi kräver ett bättre samarbete mellan hälsotjänsterna, särskilt när det gäller patientrörlighet och patientsäkerhet (t.ex. läkemedelsförfalskning), information till patienter om läkemedel och livsstilsförändringar, och när det gäller att möta utmaningarna med ett hälsosamt åldrande.
Jordbruk och fiske
48.
49.
50.
EU:s ställning som partner i världen
Grannskapspolitik
51.
52.
Europaparlamentet uppmanar kommissionen att utarbeta en årlig rapport om efterlevnaden av de klausuler i avtalen som behandlar mänskliga rättigheter och demokrati, tillsammans med en detaljerad utvärdering och rekommendationer rörande de vidtagna åtgärdernas effektivitet och samstämmighet.
Stabilitet och demokrati i sydöstra Europa
53.
Europaparlamentet konstaterar att länderna i sydöstra Europa kommer allt närmare anslutningen, vilket förutspåddes i Thessalonikiförklaringen, och förväntar sig att unionen skall gå i bräschen för att befästa stabiliteten och öka välståndet i västra Balkan och på så sätt hjälpa länderna i regionen att komma närmare ett EU-medlemskap.
Ryssland
54.
Utvecklingspolitik
55.
Europaparlamentet uppmanar medlemsstaterna och kommissionen att i större utsträckning respektera sina åtaganden i samband med millennieutvecklingsmålen, och uppmanar kommissionen att lägga fram konkreta förslag till alternativ finansiering av utvecklingsprogram.
56.
För att göra det möjligt för AVS-länderna att uppnå utvecklingsmålen anser Europaparlamentet att den regionala utvecklingsaspekten bör respekteras i samband med förhandlingarna om avtalen om ekonomiskt partnerskap.
Handelspolitik och WTO-förhandlingar
57.
ESFP
58.
Europaparlamentet betonar behovet av att stärka mekanismerna för parlamentarisk tillsyn över utvecklingen av den europeiska säkerhets- och försvarspolitiken (ESFP) i allmänhet och ESFP-uppdragen i synnerhet, och understryker behovet av att tillhandahålla proaktiv information och av att föra diskussioner innan det fattas beslut om gemensamma åtgärder inom området för ESFP så att parlamenten kan uttrycka sina åsikter och ta upp eventuella problem.
Bättre lagstiftning
59.
60.
Europaparlamentet vidhåller att alla förenklingsinitiativ skall vara helt förenliga med alla de principer och villkor som lades fast i parlamentets resolution av den 16 maj 2006 om strategin för enklare lagstiftning.
Konsekvensutredningar
61.
Icke-bindande regler
62.
Europaparlamentet beklagar att kommissionen alltmer använder icke-bindande regler, såsom rekommendationer och tolkningsmeddelanden, vilket medför att den lagstiftande myndighetens privilegier kringgås.
Övervakning av genomförandet och efterlevnaden av gemenskapens regelverk
63.
Europaparlamentet beklagar att kommissionen har varit tämligen ointresserat av att stödja parlamentets krav när det gäller genomförandet av EU-lagstiftningen i medlemsstaterna.
64.
Europaparlamentet uppmanar kommissionen att göra hela processen för införlivande och genomförande mera öppen för insyn och att förmå medlemsstaterna att utarbeta de så kallade jämförelsetabellerna som visar exakt vilka delar av lagen som härstammar från EU och vilka delar som härstammar från medlemsstaterna.
Budgetansvar
65.
Europaparlamentet förväntar sig att alla nya reformer som fastställs i det interinstitutionella avtalet av den 17 maj 2006 om budgetdisciplin och sund ekonomisk förvaltning skall genomföras fullt ut under 2007, så att det blir möjligt att uppnå snabba resultat när det gäller att förbättra kvaliteten i budgetgenomförandet.
66.
67.
68.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen och medlemsstaternas parlament.
9.7.2008
GEMENSAMT FÖRSLAG TILL RESOLUTION
– Laima Liucija Andrikienė, Bernd Posselt, Eija-Riitta Korhola och Tadeusz Zwiefka, för PPE-DE-gruppen
– Pasqualina Napoletano, Ana Maria Gomes, Józef Pinior och Marianne Mikko, för PSE-gruppen
– Marco Pannella, Marco Cappato, Frédérique Ries och Marios Matsakis, för ALDE-gruppen
– Roberta Angelilli, för UEN-gruppen
– Hélène Flautre, Monica Frassoni, Raül Romeva i Rueda, Milan Horáček, Kathalijne Maria Buitenweg, Pierre Jonckheer, Caroline Lucas och Claude Turmes, för Verts/ALE-gruppen
– Vittorio Agnoletto, för GUE/NGL-gruppen
som ersätter resolutionsförslagen från följande grupper:
– ALDE ( B6‑0350/2008 )
– UEN ( B6‑0357/2008 )
– Verts/ALE ( B6‑0358/2008 )
– GUE/NGL ( B6‑0363/2008 )
– PPE-DE ( B6‑0369/2008 )
– PSE ( B6‑0370/2008 )
om dödsstraff, särskilt Troy Davis fall
Europaparlamentets resolution om dödsstraff, särskilt Troy Davis fall
Europaparlamentet utfärdar denna resolution
–
med beaktande av sina tidigare resolutioner om avskaffande av dödsstraff och behovet av ett omedelbart moratorium för avrättningar i de länder där dödsstraffet fortfarande tillämpas,
–
med beaktande av FN:s generalförsamlings resolution 62/149 av den 18 december 2007 om dödsstraffets användning i världen,
–
med beaktande av den uppdaterade versionen av EU:s riktlinjer av den 5 juni 2008 avseende dödsstraff, och av följande skäl:
A.
Troy Davis dömdes till döden 1991 av Georgias högsta domstol för mord på en polisman och planeras avrättas i slutet av juli 2008.
B.
C.
Georgias högsta domstol gick den 4 augusti 2007 med på att granska de nya faktorer som gör att Davis skuld kan ifrågasättas.
D.
Den 17 mars 2008 beslöt Georgias högsta domstol att neka Troy Davis en ny rättegång, trots att domstolens ordförande var av avvikande mening
E.
Sedan 1975 har i USA mer än 120 personer befunnits oskyldiga och släppts fria från cellerna där de väntat på sin avrättning.
F.
I USA finns för dödsdomar en befogenhet att bevilja nåd som en säkerhetsåtgärd för att avvärja oåterkalleliga misstag som domstolar inte kunnat eller inte velat avhjälpa.
G.
New Jersey är den första delstaten som i sin lagstiftning avskaffar dödsstraffet sedan detta återinfördes i USA 1972, och man refererar till den oundvikliga risken att felaktigt dömda personer avrättas.
1.
Europaparlamentet uppmanar de länder där dödsstraffet tillämpas att vidta nödvändiga åtgärder för att avskaffa det.
2.
Mot bakgrund av de många bevis som kan ändra Troy Davis dom, anser Europaparlamentet att de berörda domstolarna bör erbjuda honom en ny rättegång och att hans dödsstraff därför bör ändras.
3.
Europaparlamentet vädjar till Georgiadomstolens nådeansökningsnämnd (Board of Pardons and Paroles) att ändra dödsstraffet.
4.
Europaparlamentet uppmanar rådets ordförandeskap och Europeiska kommissionens delegation i Förenta staterna att snabbt ta upp ärendet med de amerikanska myndigheterna.
5.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, Förenta staternas regering och Georgias Board of Pardons and Paroles samt till Georgias statsåklagare.
22.10.2008
GEMENSAMT FÖRSLAG TILL RESOLUTION
– Joseph Daul, Charles Tannock, Jacek Saryusz-Wolski, José Ignacio Salafranca Sánchez-Neyra, Tunne Kelam, Urszula Gacek och Zita Pleštinská, för PPE‑DE-gruppen
– Hannes Swoboda, Jan Marinus Wiersma och Adrian Severin, för PSE-gruppen
– Annemie Neyts-Uyttebroeck, Grażyna Staniszewska, Janusz Onyszkiewicz, István Szent-Iványi och Šarūnas Birutis, för ALDE-gruppen
– Rebecca Harms och Milan Horáček, för Verts/ALE-gruppen
– Adam Bielan, Wojciech Roszkowski, Konrad Szymański och Mieczysław Edmund Janowski, för UEN-gruppen
som ersätter resolutionsförslagen från följande grupper:
– Verts/ALE ( B6‑0571/2008 )
– ALDE ( B6‑0572/2008 )
– UEN ( B6‑0573/2008 )
– PPE-DE ( B6‑0574/2008 )
om minnesdagen för holodomor – den framtvingade hungersnöden i Ukraina 1932–1933
Europaparlamentets resolution om minnesdagen för holodomor – den framtvingade hungersnöden i Ukraina 1932–1933
Europaparlamentet utfärdar denna resolution
–
med beaktande av EU-fördraget,
–
med beaktande av Europeiska konventionen om skydd för de mänskliga rättigheterna och de grundläggande friheterna,
–
med beaktande av FN:s konvention om förebyggande och bestraffning av brottet folkmord,
–
med beaktande av det gemensamma uttalandet om 70-årsdagen av holodomor i Ukraina som gjordes vid FN:s generalförsamlings 58:e session och som understöddes av 63 stater, däribland alla EU:s (då) 25 medlemsstater,
–
med beaktande av den ukrainska lagen om holodomor i Ukraina 1932–1933 som antogs den 28 november 2006,
–
med beaktande av uttalandet av Europaparlamentets talman den 21 november 2007 som markerade inledningen av firandet av 75-årsdagen av holodomor i Ukraina,
–
med beaktande av slutdeklarationen och rekommendationerna från det tionde mötet i den parlamentariska samarbetskommittén EU–Ukraina som antogs den 27 februari 2008,
–
med beaktande av artikel 103.4 i arbetsordningen, och av följande skäl:
A.
Svälten (holodomor) 1932–1933, som kostade miljontals ukrainare livet, hade på ett cyniskt och grymt sätt planerats av den stalinistiska regimen för att genomdriva Sovjetunionens politik för en kollektivisering av jordbruket mot landsbygdsbefolkningens vilja i Ukraina.
D.
Att komma ihåg brott mot mänskligheten i Europas historia bör hjälpa oss att förebygga liknande brott i framtiden.
E.
1.
Europaparlamentet gör följande uttalande till folket i Ukraina och särskilt till dem som överlevde holodomor och fortfarande lever och deras familjer och släktingar:
a) Europaparlamentet erkänner holodomor (den framtvingade hungersnöden 1932–1933 i Ukraina) som ett avskyvärt brott mot det ukrainska folket och mot mänskligheten.
b) Europaparlamentet fördömer kraftfullt dessa gärningar mot de ukrainska bönderna, i form av massförintelse, brott mot de mänskliga rättigheterna och friheterna.
c) Europaparlamentet uttrycker sin medkänsla med det ukrainska folket, som drabbades av denna tragedi, och visar sin aktning för dem som dog till följd av den framtvingade hungersnöden 1932–1933.
d) Europaparlamentet uppmanar de före detta länderna i Sovjetunionen att ge full tillgång till arkiven om holodomor i Ukraina 1932–1933 för en omfattande undersökning för att avslöja och grundligt undersöka alla orsaker och följder.
2.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet och kommissionen och till Ukrainas regering och parlament, FN:s generalsekreterare, OSSE:s generalsekreterare och Europarådets generalsekreterare.
GEMENSAMT FÖRSLAG TILL RESOLUTION
– Michael Gahler, Mario Mauro, Laima Liucija Andrikienė, Bernd Posselt och Eija‑Riitta Korhola, för PPE-DE-gruppen
– Pasqualina Napoletano och Alain Hutchinson, för PSE-gruppen
– Marios Matsakis, Marco Cappato och Marco Pannella, för ALDE-gruppen
– Eoin Ryan, Mieczysław Edmund Janowski och Ryszard Czarnecki, för UEN‑gruppen
– Marie-Hélène Aubert och Margrete Auken, för Verts/ALE-gruppen
– Vittorio Agnoletto, för GUE/NGL-gruppen
som ersätter resolutionsförslagen från följande grupper:
– ALDE ( B6‑0602/2008 )
– Verts/ALE ( B6‑0603/2008 )
– PSE ( B6‑0604/2008 )
– UEN ( B6‑0605/2008 )
– GUE/NGL ( B6‑0606/2008 )
– PPE-DE ( B6‑0607/2008 )
om dödsstraffet i Nigeria
Europaparlamentets resolution om dödsstraffet i Nigeria
Europaparlamentet utfärdar denna resolution
–
med beaktande av sina tidigare resolutioner om brott mot de mänskliga rättigheterna i Nigeria,
–
med beaktande av att Nigerias förbundsregering utfärdat ett moratorium för tillämpningen av dödsstraffet,
–
med beaktande av den allmänna förklaringen om de mänskliga rättigheterna,
–
med beaktande av den internationella konventionen om medborgerliga och politiska rättigheter, som ratificerats den 29 oktober 1993,
–
med beaktande av den afrikanska stadgan om mänskliga rättigheter och folkens rättigheter, som ratificerats den 22 juni 1983,
–
med beaktande av den afrikanska stadgan om barnets rättigheter och välfärd, som ratificerats den 23 juli 2001,
–
med beaktande av konventionen mot tortyr och annan grym, omänsklig eller förnedrande behandling eller bestraffning, som ratificerats den 28 juli 2001,
–
med beaktande av konventionen om avskaffande av all slags diskriminering av kvinnor, som ratificerats den 13 juni 1985, och dess fakultativa tilläggsprotokoll, som ratificerades den 22 november 2004,
–
med beaktande av konventionen om barnets rättigheter, som ratificerats den 19 april 1991,
–
A.
I dag uppgår antalet dödsdömda i Nigerias fängelser till över 720 män och 11 kvinnor.
B.
Nigerias nationella arbetsgrupp för utredning av dödsstraffet och presidentens kommission för reform av rättsväsendet har kommit fram till att dödsfångarna nästan undantagslöst är fattiga som inte har någon som driver deras sak inför rätta.
C.
Folkrätten förbjuder visserligen att dödsstraffet tillämpas mot underåriga förbrytare, men minst 40 av dödsfångarna var mellan 13 och 17 år gamla då de föregivna brotten begåtts.
D.
E.
F.
Nigerias system för rättskipning i brottmål utmärks av florerande rättsröta, slarv och kännbar brist på resurser.
G.
H.
Många som i fängelse väntar på rättegång eller på att avrättas utsätts för utpressning från polisers sida, som vill att de ska betala poliserna för att försättas på fri fot.
I
Över hälften av landets 40 000 fängelseinterner har inte rannsakats eller dömts.
J.
Kroniska sjukdomar, som dock går att förebygga, såsom hiv, malaria, tuberkulos, influensa och lunginflammation förekommer också i fängelserna.
K.
Nigerias nationella arbetsgrupp 2004 för utredning av dödsstraffet och presidentens kommission för reform av rättsväsendet 2007 betvivlade att dödsstraffet bidrog till att minska brottsfrekvensen och den grasserande brottsligheten i landet, men varken förbundsregeringen eller delstatsregeringarna har gjort något åt de brännande problem som påtalats vid de båda undersökningarna.
L.
Nigeria har officiellt inte rapporterat några avrättningar sedan 2002.
M.
Endast sju av Afrikanska unionens 53 medlemsstater har, såvitt veterligt, verkställt några avrättningar under 2007, medan 13 afrikanska länder avskaffat dödsstraffet i sin lagstiftning och ytterligare 22 i praktiken inte verkställer några dödsdomar.
N.
Medan bara 16 länder avskaffat dödsstraffet för alla brott 1977 har i dag 137 av FN:s 192 medlemsstater avskaffat detta straff i sin lagstiftning eller i praktiken.
1.
Europaparlamentet uppmanar Nigerias förbundsregering och delstatsregeringar att avskaffa dödsstraffet.
2.
Europaparlamentet uppmanar Nigerias förbundsregering och delstatsregeringar att, i avvaktan på att dödsstraffet avskaffas, utfärda ett omedelbart moratorium för alla avrättningar, såsom det föreskrivs i FN:s generalförsamlings resolution nr 62/149 och utan dröjsmål omvandla alla dödsstraff till fängelsestraff.
3.
Europaparlamentet uppmanar Nigerias förbundsregering och delstatsregeringar att utveckla en helhetssyn på brottsligheten och förklara hur situationen i fråga om brottslighet kommer att åtgärdas.
4.
Europaparlamentet uppmanar med kraft Nigerias förbundsregering och delstatsregeringar att ta bort alla stadganden både i förbundsstatens lagstiftning och i delstaternas lagstiftning enligt vilka dödsdomar kan avkunnas mot personer som ej fyllt 18 år vid tidpunkten för det föregivna brottets begående.
5.
Europaparlamentet uppmanar Nigerias förbundsregering och delstatsregeringar att se till att de mest rigorösa internationellt erkända och i statsförfattningen förankrade normerna för opartisk rättegång respekteras i sådana mål där den åtalade riskerar dödsstraff, framför allt i fråga om att mindre bemedlade interner inte kan få sin talan adekvat förd inför rätta samt i fråga om att bekännelser eller bevis utverkats genom våld, tvång eller tortyr, att rättegångarna och överklagandena drar orimligt ut på tiden och att underåriga döms.
6.
Europaparlamentet uppmanar Nigerias förbundsregering att ratificera det andra fakultativa tilläggsprotokollet till Internationella konventionen om medborgerliga och politiska rättigheter samt det fakultativa tilläggsprotokollet till FN:s konvention mot tortyr.
7.
Europaparlamentet uppmanar med kraft Nigerias delstatsregeringar att avskaffa alla stadganden om att dödsstraff alltid ska utdömas.
8.
Europaparlamentet uppmanar Nigerias förbundsregering och delstatsregeringar att genomföra rekommendationerna från den nationella arbetsgruppen 2004 för utredning av dödsstraffet och presidentens kommission för reform av rättsväsendet (2007), framför allt att införa ett moratorium för alla avrättningar och omvandla alla dödsstraff.
9.
Europaparlamentet uppmanar rådet, kommissionen och medlemsstaterna att ge Nigerias myndigheter tekniskt stöd för att de ska kunna se över lagstiftning med stadganden om dödsstraff för att avskaffa dödsstraffet, samt kunna förbättra den nigerianska polisens utredningsarbete.
10.
Europaparlamentet uppmanar till att Afrikanska kommissionens arbetsgrupp för dödsstraffet ska få hjälp med att utarbeta ett protokoll till den afrikanska stadgan om förbud mot dödsstraffet, så att detta straff inte heller kan återinföras.
11.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till kommissionen, rådet, medlemsstaterna, Ecowas, Nigerias förbundsregering och parlament, Afrikanska unionen och Panafrikanska parlamentet.
P6_TA(2004)0078
Protokoll till avtalet EU/San Marino *
A6-0062/2004
Europaparlamentets lagstiftningsresolution om förslaget till rådets beslut om ingående på Europeiska gemenskapens och dess medlemsstaters vägnar av ett protokoll till avtalet om samarbete och tullunion mellan Europeiska ekonomiska gemenskapen och Republiken San Marino, rörande Republiken Tjeckiens, Republiken Estlands, Republiken Cyperns, Republiken Lettlands, Republiken Litauens, Republiken Ungerns, Republiken Maltas, Republiken Polens, Republiken Sloveniens och Republiken Slovakiens deltagande som avtalsslutande parter till följd av deras anslutning till Europeiska unionen ( KOM(2004)0258 – C6-0048/2004 – 2004/0083(CNS))
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till rådets beslut ( KOM(2004)0258 ) Ännu ej offentliggjort i EUT.
,
–
–
–
–
med beaktande av betänkandet från utskottet för internationell handel ( A6-0062/2004 ).
1.
Europaparlamentet godkänner ingåendet av protokollet till avtalet.
2.
Europaparlamentet uppdrar åt talmannen att delge rådet, kommissionen samt medlemsstaternas och Republiken San Marinos regeringar och parlament parlamentets ståndpunkt.
P6_TA(2004)0103
Förslag till allmän budget 2005, ändrad av rådet
A6-0068/2004
Europaparlamenttes resolution om rådets ändrade förslag till Europeiska unionens allmänna budget för budgetåret 2005 (alla avsnitt) (15178/2004 – C6-0225/2004 – 2004/2001(BUD) – 2004/2002(BUD)) och om ändringsskrivelserna nr 1/2005 (15180/2004 – C6-0216/2004 ), 2/2005 (15181/2004 – C6-0217/2004 ) och 3/2005 (15182/2004 – C6-0218/2004 ) till förslaget till Europeiska unionens allmänna budget för budgetåret 2005
Europaparlamentet utfärdar denna resolution
–
–
med beaktande av Fördraget om upprättandet av Europeiska atomenergigemenskapen, särskilt artikel 177,
–
med beaktande av rådets beslut 2000/597/EG, Euratom av den 29 september 2000 om systemet för gemenskapernas egna medel EGT L 253, 7.10.2000, s.
42.
,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
, särskilt artikel 40,
–
med beaktande av det interinstitutionella avtalet av den 6 maj 1999 mellan Europaparlamentet, rådet, och kommissionen om budgetdisciplin och förbättring av budgetförfarandet EGT C 172, 18.6.1999, s.
1.
Avtal ändrat genom Europaparlamentets och rådets beslut 2003/429/EG (EUT L 147, 14.6.2003, s.
25).
samt justeringen och översynen den 19 maj 2003 av budgetplanen inför utvidgningen,
–
det preliminära budgetförslag till Europeiska unionens allmänna budget för budgetåret 2005 som kommissionen lagt fram,
–
med beaktande av det förslag till Europeiska unionens allmänna budget för budgetåret 2005 som rådet fastställde den 16 juli 2004 ( C6-0123/2004 ),
–
med beaktande av parlamentets resolution av den 28 oktober 2004 om förslaget till Europeiska unionens allmänna budget för budgetåret 2005, avsnitt III – kommissionen Antagna texter, P6_TA(2004)0038.
,
–
med beaktande av parlamentets resolution av den 28 oktober 2004 om förslaget till Europeiska unionens allmänna budget för budgetåret 2005, avsnitt I – Europaparlamentet, avsnitt II – rådet, avsnitt IV – domstolen, avsnitt V – revisionsrätten, avsnitt VI – Europeiska ekonomiska och sociala kommittén, avsnitt VII – Regionkommittén, avsnitt VIII (A) – Europeiska ombudsmannen, avsnitt VIII (B) – Europeiska datatillsynsmannen Antagna texter, P6_TA(2004)0039.
,
–
med beaktande av de ändringar i och ändringsförslag till förslaget till allmän budget som parlamentet antog den 28 oktober 2004,
–
med beaktande av rådets modifieringar av parlamentets ändringar i och ändringsförslag till förslaget till allmän budget (15178/2004 – C6-0225/2004 ),
–
med beaktande av resultaten av medlingen den 25 november 2004,
–
med beaktande av Europaparlamentets och rådets beslut av den 16 december 2004 om användning av mekanismen för flexibilitet enligt punkt 24 i det ovannämnda interinstitutionella avtalet av den 6 maj 1999 för utökning av Peace II-programmet, bidrag till decentraliserade organ och återanpassning och återuppbyggnad i Irak,
–
med beaktande av ändringsskrivelserna nr 1/2005 (15180/2004 - C6-0216/2004 ), 2/2005 (15181/2004 - C6-0217/2004 ) och 3/2005 (15182/2004 - C6-0218/2004 ) till förslaget till Europeiska unionens allmänna budget för budgetåret 2005,
–
med beaktande av artikel 69 och bilaga IV i arbetsordningen,
–
med beaktande av budgetutskottets betänkande ( A6-0068/2004 ), och av följande skäl:
A.
B.
Kommissionens skrivelse angående genomförbarheten av de ändringar som antagits till budgetförslaget för 2005 har beaktats.
1.
Europaparlamentet beslutar att bekräfta sina prioriteringar och ändringar från första behandlingen såsom ändrade till följd av den överenskommelse som nåddes med rådet vid medlingssammanträdet den 25 november 2004.
Rubrik 1: Jordbruk
2.
3.
Europaparlamentet stöder den överenskommelse som nåddes av parlamentets delegation vid medlingssammanträdet den 25 november 2004 om att finansiera pilotprojektet om kvalitetsförbättring och pilotprojektet om en riskfinansieringsmodell för boskapsepidemier som en fortsättning på initiativ som genomfördes under 2004.
Rubrik 2: Strukturåtgärder
4.
5.
Europaparlamentet bekräftar sitt beslut att garantera ett effektivt genomförande av strukturåtgärder och godkänner det gemensamma uttalandet (se bilaga) som kommer att säkerställa att ytterligare betalningsbemyndiganden vid behov kan tillgängliggöras genom en ändringsbudget under 2005.
6.
Europaparlamentet ställer sig bakom rådet när det gäller att garantera att Peace II-programmet till stöd för fredsprocessen på Nordirland kan fortsätta under 2005 och 2006 samt när det gäller att tillgängliggöra 50 miljoner euro för 2005.
Rubrik 3: Inre politik
7.
Europaparlamentet välkomnar den överenskommelse som nåddes vid medlingssammanträdet den 25 november 2004 som innebär att ett belopp på ytterligare 40 miljoner euro kommer att göras tillgängligt för 2005 för att finansiera decentraliserade organ, samtidigt som parlamentets prioriteringar skyddas och stärks, särskilt när det gäller Lissabonstrategin för att främja ekonomisk tillväxt, hållbar utveckling och sysselsättning, rättsliga och inrikes frågor (inbegripet bekämpande av terrorism) samt informationspolitiken (inbegripet information till medborgarna och debatten om den framtida unionen).
8.
Europaparlamentet beklagar emellertid att rådet knappt har godkänt någon av parlamentets enskilda ändringar och är särskilt bekymrat över att rådet är ovilligt att till fullo erkänna konsekvenserna av att en allt större del av utgiftskategori 3 används för decentraliserade organ.
9.
Europaparlamentet har beslutat att för de decentraliserade organen föra in anslag motsvarande nivån i det preliminära budgetförslaget.
10.
11.
12.
13.
Europaparlamentet bekräftar den vikt det lägger vid åtgärder för att förhindra föroreningar till havs, och har tagit upp 17,8 miljoner euro i såväl åtagandebemyndiganden som betalningsbemyndiganden för det program som förvaltas av Europeiska sjösäkerhetsbyrån.
14.
Europaparlamentet godkänner förslagen för de budgetposter som är knutna till inrättandet av genomförandeorganen, i enlighet med ändringsskrivelse nr 2/2005.
Rubrik 4: Externa åtgärder
15.
16.
17.
Europaparlamentet uppmanar kommissionen att noggrant följa utvecklingen i Ukraina och garantera att tillräckliga anslag ställs till förfogande för att stödja ytterligare demokratiseringssträvanden i landet.
18.
19.
20.
Europaparlamentet uppmanar kommissionen att, i enlighet med den information om finansiering av icke-statliga aktörer som tillhandahölls efter parlamentets första behandling, senast i april 2005 lägga fram en rapport som utreder möjliga ändringar i tillämpningen av gemenskapens regler och bestämmelser, med särskild hänvisning till följande:
a)
Färre direktöverenskommelser med icke-statliga aktörer ifråga om externt bistånd, bl.a. genom en översyn av bidraget till internationella organisationer, vilket också kan minska EU-biståndets synlighet,
b)
Sänkning av EU:s maximala bidrag till projekt som genomförs av icke-statliga aktörer i förhållande till den maximinivå på 85 procent som för närvarande tillämpas samt garantier för att återstoden finansieras med icke offentliga medel,
c)
Förbättring av den ekonomiska styrningen av icke-statliga aktörer och samordning mellan internationella givare för att bemöta den allvarliga oro som kommer till uttryck i EU:s bedrägeribekämpningsbyrås femte verksamhetsrapport.
Rubrik 5: Administrativa utgifter
21.
22.
23.
Som ett resultat av lönejusteringen, besparingar och tidigareläggande av vissa investeringar, uppskattar Europaparlamentet att en betydande marginal kan skapas under taket i utgiftskategori 5, dels i budgeten för 2005 dels genom en ändringsbudget som justerar löner och pensioner under 2005.
24.
25.
Europaparlamentet uppmanar institutionernas generalsekreterare att senast den 1 april 2005 lägga fram den fjärde rapporten om tendenserna i utgiftskategori 5 tillsammans med en uppdatering av rekryteringsläget.
Övriga avsnitt
26.
Europaparlamentet har återinfört sina ändringsförslag från första behandlingen med några ändringar för att beakta att några av de andra institutionerna har tidigarelagt utgifter från 2005 till 2004.
27.
Rubrik 7: Föranslutningsstrategi
28.
Europaparlamentet stödjer den överenskommelse som nåddes av parlamentets delegation vid medlingssammanträdet den 25 november 2004 om att föra in 120 miljoner euro för att stimulera den ekonomiska utvecklingen inom den turkcypriotiska befolkningsgruppen.
Parlamentet beslutar även att öka anslagen till Kroatien till 105 miljoner euro, i överensstämmelse med strategin inför anslutningen av detta land, och att föra över befintliga anslag från utgiftskategori 4 till utgiftskategori 7.
°
29.
Europaparlamentet uppdrar åt talmannen att förklara att budgeten slutgiltigt har antagits och se till att den offentliggörs i Europeiska unionens officiella tidning.
30.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, domstolen, revisionsrätten, Europeiska ekonomiska och sociala kommittén, Regionkommittén, Europeiska ombudsmannen och Europeiska datatillsynsmannen samt till övriga berörda institutioner och organ.
BILAGA
Gemensamt uttalande
1.
Budgetmyndigheten uppmanar kommissionen att varje år tillsammans med sitt preliminära budgetförslag lägga fram en uppdaterad lägesbeskrivning avseende de tjänster som inte kan tillsättas eller som har omvandlats till följd av inrättandet av genomförandeorgan.
Ändringsbudget för 2005 om anslagen för institutionernas administration
2.
Budgetmyndigheten uppmanar kommissionen att senast i mars 2005 lägga fram en ändringsbudget som endast får omfatta minskningen av anslagen för institutionernas administration till följd av den årliga justeringen av löner och pensioner.
Betalningsbemyndiganden för utgiftskategori 2
3.
Om genomförandet av betalningsbemyndigandena för strukturfonderna överskrider 40 % i slutet av juli 2005, eller om kommissionen på annat sätt blir övertygad om att en brist på betalningsbemyndiganden kommer att uppstå, bör den efter att ha undersökt möjligheterna till omfördelning av betalningsbemyndiganden inom den totala budgeten inklusive utgiftskategori 2, och efter att ha utvärderat möjliga källor till andra inkomster, så snart som möjligt lägga fram ett preliminärt förslag till ändringsbudget för budgetmyndigheten.
Rådet och Europaparlamentet kommer att fatta beslut vid en enda behandling om det preliminär förslaget till ändringsbudget så att ytterligare nödvändiga anslag finns tillgängliga senast i början av november 2005.
Detta preliminära förslag till ändringsbudget som läggs fram och fastställs vid en enda behandling avser uteslutande de anslag som krävs under utgiftskategori 2.
P6_TA(2005)0216
Utbyte av uppgifter i fråga om grova brott, inbegripet terroristdåd *
A6-0162/2005
Europaparlamentets lagstiftningresolution om Konungariket Sveriges initiativ till rådets antagande av ett rambeslut om förenklat uppgifts- och underrättelseutbyte mellan de brottsbekämpande myndigheterna i Europeiska unionens medlemsstater, särskilt i fråga om grova brott, inbegripet terroristdåd (10215/2004 – C6-0153/2004 – 2004/0812(CNS) )
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
–
med beaktande av Konungariket Sveriges initiativ (10215/2004) EUT C 281, 18.11.2004, s.
5.
,
–
–
–
med beaktande av artiklarna 93 och 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor ( A6-0162/2005 ).
1.
Europaparlamentet godkänner Konungariket Sveriges initiativ såsom ändrat av parlamentet.
2.
Rådet uppmanas att ändra texten i överensstämmelse härmed.
3.
Rådet uppmanas att underrätta Europaparlamentet om rådet har för avsikt att avvika från den text som parlamentet har godkänt.
4.
Rådet uppmanas att på nytt höra Europaparlamentet om rådet har för avsikt att väsentligt ändra Konungariket Sveriges initiativ.
5.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen och Konungariket Sveriges regering parlamentets ståndpunkt.
Konungariket Sveriges initiativ Parlamentets ändringar Ändring 24 Skäl 1 (1)
Ett av unionens centrala mål är att inom ett område med frihet, säkerhet och rättvisa ge medborgarna en hög skyddsnivå.
(1)
Ett av unionens centrala mål är att inom ett område med frihet, säkerhet och rättvisa ge medborgarna en hög skyddsnivå
med samtidig respekt för deras integritet
.
Ändring 1 Skäl 6 (6)
För närvarande hindras ett effektivt och snabbt uppgifts- och underrättelseutbyte mellan de brottsbekämpande myndigheterna allvarligt av formella förfaranden, administrativa strukturer och juridiska hinder i medlemsstaternas lagstiftning.
Detta förhållande
är oacceptabelt för medborgarna i Europeiska unionen, som begär
större säkerhet och effektivare brottsbekämpning samtidigt som de mänskliga rättigheterna värnas.
(6)
För närvarande hindras ett effektivt och snabbt uppgifts- och underrättelseutbyte mellan de brottsbekämpande myndigheterna allvarligt av formella förfaranden, administrativa strukturer och juridiska hinder i medlemsstaternas lagstiftning.
Detta förhållande
måste vägas mot behoven av
större säkerhet och effektivare brottsbekämpning samtidigt som de mänskliga rättigheterna värnas
, i synnerhet artikel 8 i Europakonventionen om mänskliga rättigheter samt artiklarna 7 och 8 i stadgan om de grundläggande rättigheterna
(8a) En hög nivå av förtroende måste skapas mellan medlemsstaternas brottsbekämpande myndigheter och med Europol och Eurojust, eftersom en brist på sådant förtroende hittills har hindrat ett effektivt uppgifts- och underrättelseutbyte.
Dessa åtgärder bör inbegripa:
– inrättande av gemensamma normer när det gäller skydd av personuppgifter inom den tredje pelaren under överinseende av en oberoende gemensam tillsynsmyndighet,
– införande av en handbok för goda metoder avsedd för polistjänstemän, i vilken deras ansvar och skyldigheter när det gäller uppgiftsskydd fastställs på ett lättfattligt och mycket konkret sätt,
– fastställande av minimistandarder inom straff- och processrätten,
– fastställande av allmän behörighet för EG-domstolen inom tredje pelaren,
– garanti för fullständig parlamentarisk kontroll.
Ändring 3 Skäl 9a (nytt)
(9a) Genom detta rambeslut, i vilket den uppgiftsskyddsnivå som genom Europaparlamentets och rådets direktiv 95/46/EG av den 24 oktober 1995 om skydd för enskilda personer med avseende på behandling av personuppgifter och om det fria flödet av sådana uppgifter
1
_________________
1
EUT L 281, 23.11.1995, s.
31.
Ändring 4 Skäl 12 (12)
De personuppgifter som behandlas i samband med genomförandet av rambeslutet kommer att skyddas i enlighet med
(12)
De personuppgifter som behandlas i samband med genomförandet av rambeslutet kommer att skyddas i enlighet med
EU:s gemensamma normer när det gäller skydd av personuppgifter under överinseende av den gemensamma tillsynsmyndigheten för skydd
av personuppgifter
.
Ändring 5 Artikel 1, punkt 1 1.
Detta rambeslut syftar till att fastställa bestämmelser enligt vilka medlemsstaternas brottsbekämpande myndigheter effektivt och snabbt kan utbyta befintliga uppgifter och underrättelser för genomförandet av brottsutredningar eller kriminalunderrättelseåtgärder, särskilt i fråga om grova brott, inbegripet terroristdåd.
Det påverkar inte mer fördelaktiga bestämmelser i nationell lagstiftning, bilaterala eller multilaterala avtal eller överenskommelser mellan medlemsstaterna eller mellan medlemsstaterna och tredjeländer och påverkar inte heller tillämpningen av Europeiska unionens rättsakter om ömsesidig rättslig hjälp eller ömsesidigt erkännande av domar i brottmål.
1.
Detta rambeslut syftar till att fastställa bestämmelser enligt vilka medlemsstaternas brottsbekämpande myndigheter effektivt och snabbt kan utbyta befintliga uppgifter och underrättelser för genomförandet av brottsutredningar eller kriminalunderrättelseåtgärder, särskilt i fråga om grova brott, inbegripet terroristdåd.
och inte heller de bestämmelser och instrument som rör tillhandahållandet av uppgifter och underrättelser till Europol och Eurojust
Uppgifts- och underrättelseutbyte i enlighet med detta rambeslut får ske i fråga om brott som enligt lagstiftningen i den ansökande medlemsstaten är belagda med frihetsstraff eller är föremål för ett beslut om frihetsberövande som avser minst 12 månader.
Medlemsstaterna får bilateralt komma överens om en utvidgad tillämpning av förfarandena enligt detta rambeslut.
Uppgifts- och underrättelseutbyte i enlighet med detta rambeslut får ske i fråga om brott som enligt lagstiftningen i den ansökande medlemsstaten är belagda med frihetsstraff eller är föremål för ett beslut om frihetsberövande som avser minst 12 månader
och i fråga om alla de brott som anges i artiklarna 1−3 i rådets rambeslut 2002/475/RIF
1
.
Medlemsstaterna får bilateralt komma överens om en utvidgad tillämpning av förfarandena enligt detta rambeslut.
__________
1
EGT L 164, 22.6.2002, s.
3.
Ändring 7 Artikel 4, punkt 2 2.
Medlemsstaterna skall se till att villkoren för att tillhandahålla övriga medlemsstaters behöriga brottsbekämpande myndigheter uppgifter och underrättelser
, inte är strängare än de
som tillämpas på nationell nivå för tillhandahållande av eller begäran om uppgifter eller underrättelser.
2.
Medlemsstaterna skall se till att villkoren för att tillhandahålla övriga medlemsstaters behöriga brottsbekämpande myndigheter uppgifter och underrättelser
motsvarar de villkor
3a.
1.
1a.
Om uppgifter eller underrättelser inte kan lämnas omgående skall den behöriga brottsbekämpande myndighet som mottagit en begäran om uppgifter eller underrättelser omgående ange den tidsfrist inom vilken dessa kan lämnas.
Medlemsstaterna skall se till att de förfogar över förfaranden för att inom högst tolv timmar kunna besvara en begäran om uppgifter och underrättelser när den ansökande staten anger att den genomför en brottsutredning eller en kriminalunderrättelseåtgärd som rör följande brott enligt definitionen i den ansökande statens lagstiftning:
2.
Medlemsstaterna skall se till att de förfogar över förfaranden för att inom högst tolv timmar
eller, vid uppgifter eller underrättelser som förutsätter att formella förfaranden tillämpas eller att förhandskontakter tas med andra myndigheter, inom högst 48 timmar i brådskande fall och tio arbetsdagar i andra fall,
kunna besvara en begäran om uppgifter och underrättelser när den ansökande staten anger att den genomför en brottsutredning eller en kriminalunderrättelseåtgärd som rör följande brott enligt definitionen i den ansökande statens lagstiftning:
2a.
1.
.
Ändring 14 Artikel 5, punkt 3a (ny)
3a.
1.
Varje medlemsstat skall
, i överensstämmelse med de principer som anges i artiklarna 9a och 9b,
2.
utgår
3.
Uppgifter och underrättelser, inklusive personuppgifter, som lämnats enligt detta rambeslut får användas av de behöriga brottsbekämpande myndigheterna i den medlemsstat till vilken de har lämnats för
a) förfaranden på vilka rambeslutet är tillämpligt,
b) andra brottsbekämpningsförfaranden som direkt rör de som anges i a,
c) förebyggande av ett omedelbart och allvarligt hot mot den allmänna säkerheten,
d) varje annat ändamål, inklusive lagföring eller administrativa förfaranden, endast med uttryckligt förhandsmedgivande av den behöriga brottsbekämpande myndighet som har lämnat uppgifterna eller underrättelserna.
4.
När uppgifter eller underrättelser lämnas i enlighet med detta rambeslut får den lämnande behöriga brottsbekämpande myndigheten, i enlighet med sin nationella lagstiftning, ställa villkor för den mottagande behöriga brottsbekämpande myndighetens användning av uppgifterna eller underrättelserna.
Villkor får även ställas när det gäller rapportering av resultatet av den brottsutredning eller kriminalunderrättelseåtgärd inom vilken uppgifts- eller underrättelseutbytet har ägt rum.
2a.
Uppgifter och underrättelser som lämnats enligt detta rambeslut får ej användas för att lagföra andra brott än det som informationen erhållits för.
Överskottsinformation får överhuvudtaget inte användas för lagföring.
Ändring 18 Artikel 9a (ny)
Artikel 9a
Principer gällande insamling och behandling av uppgifter
1.
Uppgifter och underrättelser, inbegripet personuppgifter, som utbyts eller tillhandahålls i enlighet med detta rambeslut skall
a) vara korrekta, adekvata och relevanta med hänsyn till det syfte för vilka de insamlas och därefter behandlas,
b) insamlas och behandlas enbart i syfte att fullgöra de åligganden som föreskrivs i lag.
Uppgifter som hänför sig till privatlivet samt uppgifter som rör icke misstänkta enskilda personer får endast insamlas i absolut nödvändiga fall och under beaktande av strikta villkor.
2.
Uppgifter som tillhandahålls i enlighet med detta beslut skall på alla nivåer av utbytet och behandlingen garanteras rättrådig och konfidentiell hantering.
Källorna skall skyddas.
Ändring 19 Artikel 9b (ny)
Artikel 9b
Den person vars uppgifter har insamlats skall
a) informeras om att uppgifter om honom/henne insamlats, utom när det föreligger betydande hinder,
b) beredas rätt till kostnadsfri tillgång till de uppgifter som berör honom/henne och ges rätt att rätta felaktiga uppgifter, utom när sådan tillgång kan tänkas påverka allmän säkerhet och ordning eller tredje mans rättigheter och friheter eller hindra pågående utredningar,
c) få rätt, i samband med felaktig användning av uppgifter enligt denna artikel, att kostnadsfritt överklaga för att se till att lagen efterlevs och i förekommande fall erhålla skadestånd om de principer som föreskrivs i denna artikel inte följs.
Ändring 20 Artikel 9c (ny)
Artikel 9c
Gemensam tillsynsmyndighet för skydd för personuppgifter
1.
En gemensam tillsynsmyndighet för skydd av personuppgifter, nedan kallad tillsynsmyndigheten, skall inrättas.
Tillsynsmyndigheten skall vara ett fristående rådgivande organ.
2.
Tillsynsmyndigheten skall vara sammansatt av en företrädare för den tillsynsmyndighet eller de tillsynsmyndigheter som varje enskild medlemsstat utser, en företrädare för den myndighet eller de myndigheter som institutionerna inrättar, den europeiska datatillsynsmannen och gemenskapsorganen samt en företrädare för kommissionen.
Varje medlem i tillsynsmyndigheten skall utses av den institution, den myndighet eller de myndigheter som han/hon företräder.
Om en medlemsstat utsett flera tillsynsmyndigheter skall de välja en gemensam företrädare.
Detta gäller även de myndigheter som inrättats för institutionerna eller gemenskapsorgan.
3.
Tillsynsmyndigheten skall fatta beslut med enkel majoritet av företrädarna för tillsynsmyndigheterna.
4.
Tillsynsmyndigheten skall välja en ordförande.
Mandatperioden är två år.
Mandatet kan förnyas.
5
1
.
Sekretariatet skall överföras till kommissionen så snart som möjligt.
____________
1
EGT L 271, 24.10.2000, s.
1.
Ändring 21 Artikel 9d (ny)
Artikel 9d
Ansvarsområdet för den gemensamma tillsynsmyndigheten för skydd av personuppgifter
1.
Tillsynsmyndigheten skall ha till uppgift att
a) utreda varje fråga som avser tillämpningen av de nationella bestämmelser som antas för genomförandet av detta rambeslut,
b) avge yttranden till kommissionen om skyddsnivån inom EU,
c) ge råd om alla förslag till ändring av detta rambeslut, om alla förslag till ytterligare eller särskilda åtgärder som skall vidtas för att tillvarata fysiska personers rättigheter och friheter i samband med behandling av personuppgifter och om alla andra förslag till gemenskapslagstiftning som påverkar dessa rättigheter och friheter,
d) avge yttranden om de uppförandekoder som tagits fram på EU-nivå,
2.
Om tillsynsmyndigheten fastställer att det förekommer olikheter mellan medlemsstaternas lagstiftning och praxis som kan leda till skillnader när det gäller skydd för enskilda med avseende på behandling av personuppgifter inom EU, skall tillsynsmyndigheten informera kommissionen om detta.
3.
Tillsynsmyndigheten kan på eget initiativ utfärda rekommendationer i alla frågor om skydd för enskilda med avseende på behandling av personuppgifter inom ramen för tredje pelaren.
4.
De yttranden och rekommendationer som avges av tillsynsmyndigheten skall vidarebefordras till kommissionen.
De begärda uppgifterna eller underrättelserna
helt klart
inte står i proportion till eller är irrelevanta för de syften som ledde till begäran.
En behörig brottsbekämpande myndighet kan även vägra lämna uppgifter om den har skäl att misstänka att den uppgiftsbegärande staten ämnar använda dessa uppgifter för lagföring av andra brott än det som angivits vid ansökan.
Ändring 23 Artikel 11a (ny)
Artikel 11a
EG-domstolens behörighet
P6_TA(2005)0338
Hungersnöd i Niger
B6-0460 , 0464 , 0470 , 0473 , 0476 och 0479/2005
Europaparlamentets resolution om hungersnöden i Niger
Europaparlamentet utfärdar denna resolution
–
med beaktande av FN:s vädjan till givarländer om pengar till livsmedelshjälp till Niger, där beloppet ligger på 80,9 miljoner US-D,
–
A.
Niger var det näst fattigaste landet i världen även innan de uteblivna regnen och invasionen av gräshoppor förstörde förra årets skördar, vilket lett till att uppskattningsvis en tredjedel av landets nära tolv miljoner invånare lider allvarlig brist på mat, av vilka 800 000 är akut undernärda barn.
B.
Sedan 1900 har Niger nio gånger drabbats av svår torka och allvarlig hungersnöd och åtta gånger av gräshoppsinvasioner.
C.
Det är också känt att områden som drabbats av torka i sin tur kan medföra utbrott av ett antal smittsamma sjukdomar såsom malaria, gulsot, kolera, tyfoidfeber och diarré.
D.
Nigers livsmedelskris är sammansatt av många faktorer som alla spelar in: väderförhållanden, livsmedelsproduktion, marknader, teknik, hygien, hälsovård, utbildning, barnalstring, landets stora utlandsskuld och den utbredda fattigdomen.
E.
Ända till juni månad 2005 vägrade Nigers regering att dela ut gratis matransoner.
F.
Motivet för denna vägran var att man inte ville destabilisera marknaden och att man förnekade hur allvarlig krisen var.
G.
Livsmedel till rimliga priser, subventionerade av regeringen, har varit sällsynta och oåtkomliga för de fattigaste.
H.
När dödstalet stiger dramatiskt kan det inte vara fråga om att utdelning av katastrofhjälp i form av gratis livsmedel skall stå åt sidan för att den framtida livsmedelsförsörjningen skall tryggas.
I.
FN:s upprepade vädjanden som inleddes i november 2004 förblev i stort sett ohörda ända tills situationen blev helt krisartad.
J.
Behoven av humanitär hjälp är enorma och gäller allt från mat, dricksvatten och medicin till vaccin för barn för att förhindra epidemier.
K.
L.
Ökenspridningen och utarmningen av jordarna i Sahel är ett resultat av ohållbart utnyttjande av naturresurserna, med förstörelse av skogarna och bushen, och även av effekterna av klimatförändringarna.
M.
1.
2.
Europaparlamentet begär att undernäringen i Niger skall erkännas vara av extremt endemisk karaktär, så att man kan inrätta ett övergripande ansvarssystem med möjlighet till vård för barn under fem år och ställa terapeutiska livsmedel som visat sig effektiva till förfogande.
3.
Europaparlamentet begär att man skall prioritera förebyggande insatser, så att man minskar beroendet av de oregelbundet förekommande regnen, genom att utveckla bevattningssystemet (mikrodammar), förbättra livsmedelsproduktiviteten, använda gödsel, konstgödsel samt verktyg och öka kapaciteten i de lokala spannmålsreserverna.
4.
Europaparlamentet välkomnar att kommissionen öronmärkt 4,6 miljoner EUR till humanitärt bistånd till Niger, och även det löfte som gavs den 1 juli 2005 att ge ytterligare humanitär hjälp om situationen skulle förvärras ännu mer.
5.
Europaparlamentet beklagar Nigers regerings otillräckliga och långsamma reaktion på den annalkande krisen och myndigheternas försummelse att dela ut gratis mat i ett tidigt skede av krisen.
6.
Europaparlamentet beklagar att staten inte ingripit tillräckligt för att förhindra spekulation och kris och önskar att Nigers regering inrättar mekanismer som gör det möjligt att undvika att liknande situationer upprepar sig.
7.
Europaparlamentet ifrågasätter det välgrundade i den totala avreglering av jordbruksmarknaderna som inleddes inom ramen för den "strukturanpassningspolitik" som förespråkats av Internationella valutafonden.
8.
Europaparlamentet varnar samtidigt för risken att ge missriktad livsmedelshjälp och uppmanar det internationella samfundet att avsluta matbiståndet så snart de anser att situationen har förbättrats.
9.
10.
Europaparlamentet begär att de reserver som finns i FN:s hjälpfonder skall ökas markant, för att tillräckligt mycket pengar skall finnas tillgängliga i förväg och därmed möjliggöra för FN:s stödorganisationer att snabbt sätta igång sina hjälpinsatser.
11.
Europaparlamentet beklagar djupt att afrikanska katastrofer medför en sådan påtvingad mobilisering, medan tsunamin och dess offer, varav många var västerlänningar, fick oerhörd uppmärksamhet i medierna.
12.
Europaparlamentet välkomnar samordningen av ECHO:s katastrofhjälp med mer långsiktiga insatser för tryggad livsmedelsförsörjning som handläggs av kommissionen, liksom ett klart åtagande att se landsbygdsutveckling och tryggad livsmedelsförsörjning som en prioritet i landstrategidokumentet för Niger.
13.
Europaparlamentet uppmanar de internationella givarna att även fokusera på hälsorelaterat stöd, till exempel att underlätta tillgången till rent vatten, dela ut vattenreningstabletter och stödja och utvidga befintlig hälsovård för att förhindra utbrott av smittsamma sjukdomar.
14.
15.
Europaparlamentet är oroat över tillgången till mat i grannstaterna Mali och Burkina Faso och önskar att man noggrant skall övervaka situationen i detta större område.
16.
Europaparlamentet uppmanar kommissionen och rådet att förbättra systemet för tidig varning så att man övervakar känsliga regioner där svält kan uppstå för att göra det möjligt att vidta tidiga åtgärder och förhindra katastrofer.
17.
Europaparlamentet betonar att huvudproblemet i Niger är den kroniska utbredda fattigdomen och att landet inte har några marginaler att bygga upp beredskapslager för att möta detta slags krisbehov.
18.
Europaparlamentet uppmanar kommissionen och rådet att erkänna effekterna av den globala uppvärmningen i Afrika söder om Sahara och att agera i Europa för att mildra effekterna genom att anta strängare EU-strategier för att minska koldioxidutsläppen.
19.
Europaparlamentet anser att frågan om exploatering av naturresurserna är en faktor som måste beaktas i handelsförhandlingarna med de afrikanska länderna.
20.
Europaparlamentet begär att åtgärder vidtas för att se till att den avskrivning av Nigers utlandsskulder som annonserades vid G8-toppmötet verkligen kommer att genomföras.
21.
Europaparlamentet uppmanar kommissionen att när nödsituationen är över börja tillämpa en övergripande politik för att angripa krisens grundorsaker, ta itu med bakomliggande strukturella orsaker och förbättra jordbrukets produktivitet i regionen.
22.
Europaparlamentet uppmanar regeringarna i regionen att börja tillämpa en politik för hållbar utveckling inom jordbruket.
23.
Europaparlamentet begär att FN:s generalförsamling i september 2005 skall fastställa villkor och verktyg för det internationella stödet i syfte att utrota fattigdomen och svälten i världen, i enlighet med millenniemålen.
24.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, Afrikanska unionen, FN:s generalsekreterare, medordförandena i AVS-EG:s gemensamma parlamentariska församling samt regeringarna i Niger, Mali, Burkina Faso och Mauretanien.
P6_TA(2005)0416
Fallet Tenzin Delek Rinpoche
B6-0562 , 0565 , 0567 , 0570 , 0575 och 0581/2005
Europaparlamentets resolution om fallet Tenzin Delek Rinpoche
Europaparlamentet utfärdar denna resolution
–
med beaktande av sina tidigare resolutioner om Tibet och situationen i fråga om de mänskliga rättigheterna i Kina,
–
med beaktande av sina resolutioner av den 18 november 2004 om Tibet och fallet Tenzin Delek Rinpoche EUT C 201 E, 18.8.2005, s.
122.
och den 13 januari 2005 om Tibet EUT C 247 E, 6.10.2005, s.
158.
,
–
med beaktande av sin resolution av den 28 april 2005 om årsrapporten om de mänskliga rättigheterna i världen 2004 och EU:s politik på detta område Antagna texter, P6_TA(2005)0150 .
,
–
med beaktande av dialogen om mänskliga rättigheter mellan EU och Kina,
–
med beaktande av rapporten och rekommendationerna från seminariet om EU:s och Kinas dialog om mänskliga rättigheter den 20–21 juni 2005,
–
med beaktande av det gemensamma uttalandet från det åttonde toppmötet mellan EU och Kina den 5 september 2005,
–
A.
Den 2 december 2002 dömde folkdomstolen i den tibetanska självständiga prefekturen Kardze i provinsen Sichuan den inflytelserika och respekterade buddhistiska laman Tenzin Delek Rinpoche till döden med två års uppskov, och hans assistent Lobsang Dhondup till döden utan uppskov.
B.
Det har inte kunnat bevisas att vare sig Tenzin Delek Rinpoche eller Lobsang Dhondup varit inblandade i bombattentat eller i uppmaningar till separatism.
C.
Lobsang Dhondup avrättades den 26 januari 2003.
D.
E.
F.
Informationen om Tenzin Deleks Rinpoches hälsotillstånd kan inte kontrolleras av oberoende observatörer eftersom den kinesiska regeringen nekar tillträde.
G.
H.
Det embargo som man 1989 beslutade om och började tillämpa mot försäljning av vapen till Kina, på grund av massakern på Himmelska fridens torg och de fortsatta kränkningarna av de mänskliga rättigheterna och religionsfriheten, är fortfarande i kraft.
1.
Europaparlamentet är mycket oroat över Tenzin Delek Rinpoches hälsotillstånd.
2.
Europaparlamentet uppmanar de ansvariga myndigheterna att göra allt för att förbättra Tenzin Deleks Rinpoches levnadsvillkor och hälsotillstånd.
3.
Europaparlamentet begär att den kinesiska regeringen låter Manfred Nowak, FN:s särskilde rapportör om tortyr, besöka Tenzin Delek Rinpoche under sin inspektionsresa till Kina den 21 november till 2 december 2005 och rapportera om hans hälsotillstånd.
4.
Europaparlamentet upprepar sitt stöd för rättssäkerheten och uppskattar att Tenzin Delek Rinpoches dödsstraff har omvandlats.
5.
Icke desto mindre uppmanar Europaparlamentet den kinesiska regeringen att upphäva alla domar mot Tenzin Delek Rinpoche och omedelbart släppa honom fri.
6.
Europaparlamentet upprepar sitt krav på att dödsstraffet skall avskaffas och vill omedelbart se ett moratorium för dödsstraff i Kina.
7.
Europaparlamentet beklagar bristen på konkreta resultat i EU:s och Kinas dialog om mänskliga rättigheter och uppmanar på nytt Kinas regering att förbättra de omänskliga villkoren i fängelserna, att upphöra med och avskaffa tortyren av fångarna och att stoppa de fortsatta kränkningarna av det tibetanska folkets och andra minoriteters mänskliga rättigheter, samt att följa internationella bestämmelser om mänskliga rättigheter och människorättslagstiftning.
8.
Europaparlamentet uppmanar rådet och medlemsstaterna att bibehålla EU:s vapenembargo mot Kina och att inte lätta på de befintliga nationella begränsningarna av sådan vapenförsäljning.
9.
Europaparlamentet uppmanar Kinas regering att intensifiera den pågående dialogen med Dalai Lamas företrädare i syfte att utan ytterligare dröjsmål uppnå en ömsesidigt acceptabel lösning på Tibetfrågan.
10.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, FN:s generalsekreterare, den kinesiska regeringen, guvernören för provinsen Sichuan och chefsåklagaren i folkets rättsliga övervakningsmyndighet i provinsen Sichuan.
P6_TA(2005)0441
Nyligen gjorda uttalanden av Irans president Mahmoud Ahmadinejad
B6-0585 , 0608 , 0609 , 0610 , 0611 och 0612/2005
Europaparlamentets resolution om Iran
Europaparlamentet utfärdar denna resolution
-
med beaktande av sina tidigare resolutioner om Iran, särskilt sin resolution av den 13 oktober 2005 Antagna texter, P6_TA(2005)0382 .
,
-
med beaktande av slutsatserna från rådets (allmänna frågor) möte den 7 november 2005,
-
med beaktande av sina tidigare resolutioner om Mellanöstern, i synnerhet de av den 23 oktober 2003 EUT C 82 E, 1.4.2004, s.
610.
och den 27 januari 2005 EUT C 253 E, 13.10.2005, s.
35.
,
-
A.
Vid en konferens i Teheran kallad "En värld utan sionism" onsdagen den 26 oktober 2005 citerade Irans president Mahmoud Ahmadinejad Irans före detta revolutionsledare ayatolla Ruhollah Khomeini och fastslog att Israel måste strykas från världskartan.
B.
Det internationella samfundet har omedelbart och med kraft tillbakavisat denna typ av uppmuntran till våld och förstörelse av en stat.
C.
Även i Iran har kritiska röster höjts mot president Ahmadinejads uttalande, bland annat från ingen mindre än Irans förre president Mohammad Khatami.
D.
Iran håller på att förhandla med EU om en föreslagen omfattande dialog som rör känsliga ämnen som kärnprogrammet, bekämpningen av den internationella terrorismen, ekonomiskt samarbete samt mänskliga rättigheter.
1.
2.
Europaparlamentet uppmanar Irans regering att uppfylla sina internationella förpliktelser enligt artikel 2 i FN:s stadga, och att i sina internationella förbindelser avhålla sig från hot om eller bruk av våld, vare sig riktat mot någon annan stats territoriella integritet eller politiska oberoende, eller på annat sätt agera oförenligt med Förenta Nationernas ändamål.
3.
Europaparlamentet uttrycker sin oro over de möjliga följder som denna typ av kommentarer kan få i en region som fortfarande är utsatt för våld, terroristattacker och extremistiska och fundamentalistiska uppmaningar till våld.
4.
Europaparlamentet bekräftar på nytt sin oföränderliga utfästelse när det gäller Israels existensberättigande inom internationellt erkända gränser och i säkerhet vid sidan av en palestinsk självständig och livskraftig stat.
5.
Europaparlamentet uppmanar Iran att erkänna staten Israel och dess rätt att leva i fred och säkerhet och att använda sitt inflytande i Mellanöstern till att övertyga de rörelser som den har kontakt med att avstå från våldshandlingar.
6.
7.
Europaparlamentet välkomnar det internationella samfundets mycket kritiska reaktioner och stöder till fullo FN:s säkerhetsråds förklaring i vilket man fördömer den iranske presidenten för hans uttalande och stöder FN:s generalsekreterare, som påmint Iran om dess skyldigheter i enlighet med FN:s stadga.
8.
9.
Europaparlamentet välkomnar den ståndpunkt som ett flertal äldre palestinska tjänstemän och företrädare intog då de fördömde president Ahmedinejads attityd och uttalade sig för en fredlig samexistens mellan en palestinsk och israelisk stat.
10.
11.
12.
Europaparlamentet uppmanar rådet och kommissionen att handla enligt slutsatserna från rådet (allmänna frågor) den 7 november 2005 och Europaparlamentets resolution av den 13 oktober 2005 för att komma fram till en diplomatisk lösning på problemen med Irans kärnprogram och att behålla denna position i den fortsatta utvecklingen av den omfattande dialogen.
13.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till kommissionen, rådet, medlemsstaternas regeringar och parlament, Irans och Israels regeringar och parlament samt till generaldirektören för IAEA och FN:s generalsekreterare.
P6_TA(2005)0459
Återbetalning av mervärdesskatt till personer etablerade i en annan medlemsstat *
A6-0324/2005
Europaparlamentets lagstiftningsresolution om förslaget till rådets direktiv om fastställande av närmare regler för återbetalning enligt direktiv 77/388/EEG av mervärdesskatt till beskattningsbara personer som inte är etablerade inom landets territorium men etablerade i en annan medlemsstat ( KOM(2004)0728 – C6-0251/2005 – 2005/0807(CNS) )
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till rådet ( KOM(2004)0728 ) Ännu ej offentliggjort i EUT.
,
–
med beaktande av artikel 93 i EG-fördraget, i enlighet med vilken rådet har hört parlamentet (C6–0251/2005),
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för ekonomi och valutafrågor ( A6-0324/2005 ).
1.
Europaparlamentet godkänner kommissionens förslag såsom ändrat av parlamentet.
2.
3.
Rådet uppmanas att underrätta Europaparlamentet om rådet har för avsikt att avvika från den text som parlamentet har godkänt.
4.
Rådet uppmanas att på nytt höra Europaparlamentet om rådet har för avsikt att väsentligt ändra kommissionens förslag.
5.
Den medlemsstat där mervärdesskatten betalades skall meddela den sökande sitt beslut beträffande ansökan om återbetalning inom tre månader från den dag då ansökan lämnades in.
1.
Den medlemsstat där mervärdesskatten betalades skall meddela den sökande sitt beslut beträffande ansökan om återbetalning inom tre månader från den dag då ansökan lämnades in.
Överföringen av det återbetalade beloppet skall genomföras inom en vecka efter att tremånadsperioden för beslut löpt ut.
ytterligare
uppgifter inom tre månader från
den dag då ansökan
lämnades in.
4.
den dag då ansökan
P6_TA(2006)0086
Tvångsprostitution
B6-0160/2006
Europaparlamentets resolution om tvångsprostitution i samband med internationella idrottsevenemang
Europaparlamentet utfärdar denna resolution
–
med beaktande av den Internationella kvinnodagen den 8 mars 2006,
–
med beaktande av Europeiska unionens stadga om de grundläggande rättigheterna EGT C 364, 18.12.2000, s.
1.
–
med beaktande av Internationella konventionen om avskaffande av all slags rasdiskriminering som trädde i kraft den 4 januari 1969,
–
med beaktande av FN-konventionen om avskaffande av all slags diskriminering av kvinnor av den 18 december 1979,
–
med beaktande av det meddelande som kommissionen nyligen lagt fram om kampen mot människohandel – en integrerad strategi och förslag till handlingsplan ( KOM(2005)0514 ),
–
med beaktande av den handlingsplan som rådet nyligen offentliggjort om bästa metoder, standarder och förfaranden för att bekämpa och förhindra människohandel EUT C 311, 9.12.2005, s.
1.
,
–
,
–
med beaktande av Europarådets konvention om åtgärder mot människohandel,
–
med beaktande av FN:s konvention om barnets rättigheter och ILO:s konvention om de värsta formerna av barnarbete,
–
A.
B.
Tvångsprostitution som en form av utnyttjande av kvinnor och barn är ett betydande problem som inte bara drabbar enskilda kvinnor och barn utan också skadar samhället i stort.
C.
Erfarenheten visar att efterfrågan på sexuella tjänster tillfälligt ökar dramatiskt under varje större idrottsevenemang som drar till sig många besökare.
D.
E.
Om alla medlemsstater följde samma praxis och på ett effektivt sätt använde de medel för kommunikation som finns samt genomförde samordnade kampanjer, med deltagande av massmedia och idrottsstjärnor, i syfte att höja medvetandenivån, så skulle detta på ett positivt sätt kunna påverka allmänheten att ändra mentalitet och beteende.
1.
2.
Europaparlamentet uppmanar Tyskland och de andra medlemsstaterna att inrätta en flerspråkig hotline och genomföra en väl synlig informationskampanj i syfte att erbjuda den information, den rådgivning, det trygga boende och den rättshjälp som krävs för de kvinnor, barn och andra offer som tvingats in i prostitution, samt för att informera andra offer som ofta sitter isolerade i bostads- eller industriområden, inte kan tala transit- eller destinationslandets språk och inte har tillgång till de mest grundläggande upplysningarna, som vem man skall kontakta och vilka åtgärder som kan vidtas.
3.
Europaparlamentet uppmanar Internationella olympiska kommittén, förbund som FIFA, UEFA, det tyska fotbollsförbundet m.fl. och idrottsmännen själva att stödja Rött kort-kampanjen och att fördöma människohandel och tvångsprostitution.
4.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att genomföra kampanjer över hela Europa i samband med alla internationella idrottsevenemang i syfte att informera allmänheten, i synnerhet idrottsutövare, idrottsentusiaster och supportrar, och därigenom öka kunskaperna om problematiken och omfattningen av tvångsprostitution och människohandel, men framför allt för att minska efterfrågan genom att höja de potentiella kundernas medvetande.
5.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att inleda en förebyggande kampanj som riktar sig till potentiella offer, där man informerar dem om riskerna och farorna med att låta sig snärjas av människohandelsnätverk och därigenom falla offer för tvångsprostitution och sexuellt utnyttjande, samt att tillhandahålla information om deras rättigheter och var i destinationsländerna de kan få hjälp och stöd.
6.
7.
Europaparlamentet uppmanar samtliga medlemsstater att ratificera Europarådets konvention om åtgärder mot människohandel, i vilken det fastställs miniminormer för skydd av offren för människohandel som syftar till sexuellt utnyttjande, samt att genomföra rådets direktiv 2004/81/EG om uppehållstillstånd till offer för människohandel EUT L 261, 6.8.2004, s.
19.
.
8.
Europaparlamentet uppmanar de medlemsstater som inte respekterat tidsfristen den 1 augusti 2004 för genomförande av rådets rambeslut 2002/629/RIF om bekämpande av människohandel EUT L 203, 1.8.2002, s.
1.
9.
P6_TA(2006)0089
Socialt skydd och social integration
A6-0028/2006
Europaparlamentets resolution om socialt skydd och social integration ( 2005/2097(INI) )
–
med beaktande av kommissionens meddelande med titeln "Utkast till gemensam rapport om socialt skydd och social integration" ( KOM(2005)0014 ),
–
med beaktande av kommissionens arbetsdokument med titeln "Bilaga till utkastet till gemensam rapport om socialt skydd och social integration" ( SEK(2005)0069 ),
–
med beaktande av kommissionens arbetsdokument om social integration i de nya medlemsstaterna: Sammanfattning av de gemensamma meddelandena om social integration ( SEK(2004)0848 ),
–
med beaktande av ordförandeskapets slutsatser från Europeiska rådets möte i Bryssel den 22–23 mars 2005,
–
med beaktande av sin resolution av den 9 mars 2005 om halvtidsöversynen av Lissabonstrategin EUT C 320 E, 15.12.2005, s.
164.
,
–
med beaktande av ordförandeskapets slutsatser från Europeiska rådets möte i Santa Maria da Feira den 19–20 juni 2000 och särskilt överenskommelsen om att man bör definiera indikatorer som gemensamma referenser i kampen mot social utslagning och utrotandet av fattigdom,
–
med beaktande av kommissionens meddelande om den socialpolitiska agendan ( KOM(2005)0033 ),
–
med beaktande av rådets beslut 2005/600/EG av den 12 juli 2005 om riktlinjer för medlemsstaternas sysselsättningspolitik EUT L 205, 6.8.2005, s.
21.
,
–
med beaktande av Europaparlamentet och rådets beslut nr 50/2002/EG av den 7 december 2001 om inrättande av ett program för gemenskapsåtgärder som skall uppmuntra medlemsstaterna att samarbeta för att motverka social utslagning EGT L 10, 12.1.2002, s.
1.
,
–
–
–
med beaktande av kommissionens meddelande "Stärka Lissabonstrategins sociala dimension – Rationalisera den öppna samordningen inom socialt skydd" ( KOM(2003)0261 ),
–
med beaktande av kommissionens meddelande om att modernisera de sociala trygghetssystemen för att utveckla högkvalitativ, tillgänglig och hållbar vård och omsorg: stöd till de nationella strategierna genom den öppna samordningsmetoden ( KOM(2004)0304 ),
–
–
med beaktande av sin resolution av den 11 juni 2002 om kommissionens meddelande till rådet, Europaparlamentet, Ekonomiska och sociala kommittén och Regionkommittén om förslag till gemensam rapport om social integration EUT C 261 E, 30.10.2003, s.
136.
,
–
med beaktande av sin resolution av den 5 juni 2003 om tillämpningen av den öppna samordningsmetoden EUT C 68 E, 18.3.2004, s.
604.
,
–
med beaktande av sin resolution av den 24 september 2003 om den gemensamma rapporten från kommissionen och rådet om adekvata och hållbara pensioner EUT C 77 E, 26.3.2004, s.
251.
,
–
med beaktande av sin resolution av den 28 april 2005 om modernisering av det sociala skyddet och utvecklingen av en högkvalitativ hälsovård EUT C 45 E, 23.2.2006, s.
134.
,
–
P6_TA(2005)0210 .
,
–
P6_TA(2005)0244 .
,
–
med beaktande av artikel 45 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för sysselsättning och sociala frågor samt yttrandet från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män ( A6-0028/2006 ), och av följande skäl:
A.
B.
Medlemsstaterna åtog sig vid Europeiska rådets möte i Nice 2000 att till 2010 uppvisa en betydande och mätbar minskning av fattigdom och social utestängning.
C.
Social integration handlar om mänsklig värdighet, vilket är en grundläggande rättighet.
D.
Social integration kan i vissa fall bidra direkt och effektivt till den ekonomiska utvecklingen.
E.
F.
Enligt statistik från OECD åldras befolkningen i de länder som ingår i denna organisation, och även om det för närvarande går 38 pensionstagare på 100 arbetstagare kan denna siffra komma att stiga till hela 70 pensionstagare på 100 arbetstagare om sysselsättningspolitiken inte förändras.
G.
Moderniseringen av de sociala skyddssystemen borde inte enbart handla om att garantera ekonomisk hållbarhet, utan även om att dela på riskerna som enskilda individer har svårt att hantera på egen hand, och om att främja ekonomisk tillväxt och sysselsättning så att systemen blir hållbara.
H.
Därför bekräftas det på nytt att sociala skyddssystem som bygger på allmängiltighet, rättvisa och solidaritet är en viktig del av den europeiska sociala modellen.
Allmänna synpunkter
1.
2.
3.
4.
5.
Europaparlamentet understryker att sysselsättning måste betraktas som det effektivaste skyddet mot fattigdom och att man därför även i fortsättningen, genom åtgärder för att få in fler kvinnor på arbetsmarknaden och genom att ställa upp mål för kvaliteten på de arbetstillfällen som erbjuds, måste se till att det lönar sig att arbeta.
Social integration
6.
Europaparlamentet anser att åtgärderna mot fattigdom och social utestängning måste fullföljas och utökas för att förbättra situationen för de människor som i första hand riskerar fattigdom och utestängning, till exempel tillfälligt anställda, arbetslösa, ensamstående hushåll (som oftast förestås av kvinnor), ensamstående äldre personer, kvinnor, familjer med stor försörjningsbörda, missgynnade barn samt etniska minoriteter, sjuka eller funktionshindrade individer, bostadslösa samt personer som är offer för människohandel och för droger och alkoholberoende.
7.
8.
9.
Europaparlamentet betonar i detta sammanhang att det för romerna vore önskvärt om medlemmar ur denna minoritet motiverades på alla sätt att intressera sig för sina barns vidareutbildning, för barnens utveckling av sina positiva egenskaper och färdigheter.
10.
11.
Europaparlamentet rekommenderar medlemsstaterna att motverka riskerna med avbrott i yrkeslivet och utöka möjligheterna till livslångt lärande, för att på det sättet minska den social utestängningen av personer som är äldre än 50 år och göra det lättare för dem att stanna kvar på arbetsmarknaden.
12.
Europaparlamentet anser det därför självklart att arbetsgivarna borde vara mer engagerade i livslångt lärande, med tanke på de fördelar som det innebär för dem att ha kvalificerad arbetskraft.
13.
14.
Europaparlamentet understryker att i 14 av de 17 medlemsstater för vilka uppgifter finns att tillgå Unicef:s rapport nr 6: Barnfattigdom i rika länder 2005.
15.
16.
17.
Europaparlamentet uppmanar kommissionen att lägga fram en grönbok om barnfattigdom med tydliga mål och lämpliga åtgärder för att eliminera barnfattigdomen och verka för den sociala integrationen av fattiga barn.
18.
Europaparlamentet uppmanar kommissionen att göra mera för att införa en stadga för barnens rättigheter i syfte att nå framsteg när det gäller att försvara barnens rättigheter som en del av Europeiska unionens in- och utrikespolitik.
19.
20.
Europaparlamentet uppmanar medlemsstaterna att utveckla integrerade strategier för att ekonomiskt, socialt, kulturellt och miljömässigt försöka främja utvecklingen av geografiskt avlägsna och underutvecklade städer, öar och landsbygdsområden i syfte att ta itu med problemen med utestängning och fattigdom så att inte problemen kvarstår från en generation till nästa.
21.
Europaparlamentet understryker behovet av att få fler kvinnor i arbete genom att avlägsna sådant som hindrar dem från att komma in på arbetsmarknaden, framför allt genom att uppmuntra äldre kvinnor att stanna längre på arbetsmarknaden.
22.
Europaparlamentet rekommenderar medlemsstaterna att stödja en politik som gynnar tillväxt och kvinnors sysselsättning och underlättar kvinnors tillgång till kvalificerade arbeten samt lika lön för kvinnor.
23.
Europaparlamentet understryker att ökningen av andelen yrkesverksamma kvinnor inte enbart skall ses som ett nödvändigt skydd mot risken för fattigdom, som i huvudsak drabbar kvinnor, utan även som ett sätt att bevara balansen mellan andelen yrkesverksamma och inte yrkesverksamma, en balans som hotas av den åldrande befolkningen.
24.
25.
Europaparlamentet uppmanar vidare medlemsstaterna att vidta åtgärder för att se till att inte kvinnor får sämre pensionsrättigheter till följd av avbrott i anställningen på grund av mamma- eller föräldraledighet.
26.
Europaparlamentet uppmanar medlemsstaterna att utveckla och genomföra åtgärder, inklusive medvetandehöjande åtgärder, som ett led i deras kamp mot den omfattande utestängning som drabbar etniska minoriteter och invandrare, för att integrera dessa målgrupper på den formella arbetsmarknaden, genomdriva lagstiftning mot människohandel och diskriminering och underlätta dessa gruppers sociala integration genom särskilda bestämmelser om och omfattande program för speciella utbildningsprogram och anständiga levnads- och bostadsförhållanden som en förutsättning för social integration.
27.
Europaparlamentet uppmanar med kraft kommissionen att lägga fram förslag som syftar till att skapa en lämplig rättslig ram för att utrota diskrimineringen av funktionshindrade personer och främja dessa personers lika möjligheter och fulla deltagande på arbetsmarknaden, i samhället och i politiken, särskilt med hjälp av ett förslag till direktiv som bygger på artikel 13 i EG-fördraget för att täcka de områden som ännu inte har behandlats.
28.
29.
Europaparlamentet anser därför dessutom att undervisning i sådana grundläggande färdigheter inte bara skulle syfta till att öva upp folks förmåga att klara sig själva utan också skulle skapa solidaritet med dem som är mer sårbara, och att sådan undervisning fortgående bör ges åt hela det europeiska samhället, ända från grundskolan.
30.
31.
Europaparlamentet välkomnar erkännandet att det vanligtvis är just de människor som är socialt sett mest illa däran som har det svårast i samhällsmiljön och att man borde ta ordentlig hänsyn till detta när man bekämpar social utestängning.
32.
Europaparlamentet uppmanar kommissionen att vidta rättsliga åtgärder mot de medlemsstater som inom den obligatoriska tidsfristen inte tillämpar eller underlåtit att införliva anti-diskrimineringsdirektivet som bygger på artikel 13 i EU-fördraget.
33.
Europaparlamentet upprepar behovet av en effektivare insamling av harmoniserade uppgifter och en utveckling av gemensamma indikatorer som tar hänsyn till ålders- och könsskillnader eftersom den här sortens indikatorer spelar en viktig roll i övervakningen och utvärderingen av politiska åtgärder mot fattigdom och social utestängning.
34.
35.
Europaparlamentet påpekar att den sociala integrationsprocessen verkligen måste omfatta nyckelaktörer på lokal och regional nivå, till exempel lokala myndigheter som är ansvariga för den sociala integrationspolitiken, arbetsmarknadens parter, icke-statliga organisationer samt personer som är drabbade av fattigdom och social utestängning.
36.
Europaparlamentet stöder kommissionens avsikter att ägna särskild uppmärksamhet åt arbetet med att bekämpa fattigdom genom att arrangera Europeiska året för bekämpning av utestängning och fattigdom.
Socialt skydd
37.
Europaparlamentet anser att den snabba förändringen till följd av globaliseringen och den vidsträckta användningen av informations- och kommunikationsteknik ökar sårbarheten för sociala risker och skapar ett behov av effektivare åtgärder för socialt skydd för att garantera allas rätt till socialt skydd.
38.
39.
Europaparlamentet anser att de nuvarande demografiska trenderna – en åldrande arbetskraft och en krympande arbetsför andel av befolkningen – innebär en utmaning för de sociala trygghetssystemens ekonomiska hållbarhet på medellång och lång sikt.
40.
Europaparlamentet pekar i detta avseende på behovet av att främja utveckling och tillämpning av heltäckande åldrandestrategier för att de anställda skall kunna förbli aktiva längre och uppmuntra arbetsgivarna att anställa eller ha kvar äldre personer.
41.
Europaparlamentet uppmanar med kraft kommissionen att lägga fram förslag till lämpliga rättsliga ramar för att utrota åldersdiskriminering.
42.
Europaparlamentet anser i detta avseende att Europeiska socialfonden kan spela en viktig roll för att integrera och återinslussa äldre människor på arbetsmarknaden, och mer allmänt, när det gäller den sociala integrationen av sårbara och/eller socialt utestängda grupper.
43.
Europaparlamentet anser att det behövs ekonomisk tillväxt och tillräcklig produktivitet, liksom höga sysselsättningsnivåer och ett aktivt främjande av livslångt lärande, arbetskvalitet samt en trygg och hälsosam arbetsmiljö för att pensionssystemen skall bli ekonomiskt hållbara.
44.
Europaparlamentet rekommenderar att pensionssystemen inte enbart skall bestå av ett stort antal olika former av socialförsäkringar och tilläggsförsäkringar (antingen lagstadgade eller privata), utan även garantera maximal social rättvisa i dessa system.
45.
Europaparlamentet är av den åsikten att reformerna av de offentliga pensionssystemen inte bör öka den totala beskattningen av arbete, utan skapa en lämplig balans mellan skatten på arbete och beskattningen av andra resurser för att kunna förhindra negativa effekter på sysselsättningen.
46.
Europaparlamentet uppmanar medlemsstaterna att bygga ut sin administrativa och institutionella kapacitet, bland annat genom en mer jämlik tillgång till högkvalitativa tjänster, framför allt inom områdena för hälso- och långtidsvård, social trygghet, sociala tjänster, bland dem även rådgivning om sociala rättigheter, barnrelaterade tjänster, transport och rörlighet, tjänster för återintegrering koncentrerade på integration på arbetsmarknaden samt yrkesutbildning.
47.
Europaparlamentet ser fram emot kommissionens dokument om minimiinkomst som ett möjligt användbart bidrag till debatten om social integration och socialt skydd.
48.
49.
50.
Europaparlamentet förespråkar vidare en utbyggnad av alla de samhällstjänster som behövs för omsorg av vårdberoende, dvs. sådana som inte kan klara sina grundläggande vardagsgöromål själva.
51.
Europaparlamentet konstaterar att även om offentliga pensionssystem bör förbli en viktig inkomstkälla för pensionärerna, så kan privata bidrag via arbetsanknutna eller privata försäkringssystem spela en kompletterande roll som källa till högre pension.
52.
Europaparlamentet påpekar i detta sammanhang behovet av samordnade heltäckande informations- och övervakningssystem som betonar följderna för enskilda individers inkomst- och levnadsstandard.
53.
Europaparlamentet understryker betydelsen av en kontinuerlig effektivitetsutvärdering av pensionssystemen, med hänsyn till deras ekonomiska hållbarhet och förmåga att uppnå de sociala målen.
54.
Europaparlamentet uppmanar Europeiska rådet att vid sitt vårmöte 2006 anta ett integrerat ramverk inom området socialt skydd och social integration och enas om en enhetlig förteckning över gemensamma mål inom området social integration, pensioner och hälso- och långtidsvård, i syfte att rationalisera och förenkla den öppna samordningsmetoden.
55.
Europaparlamentet anser att upprättandet av ett integrerat ramverk och rationaliseringen av samordningen inom områdena socialt skydd och social integration innebär en möjlighet att, inom ramarna för Lissabonprocessen, ge socialskyddet en ökad social dimension så att det får en egen självständig samhällsekonomisk betydelse, i motsats till samordningen av den sociala politiken och sysselsättningspolitiken.
56.
Europaparlamentet uppmanar medlemsstaterna och kommissionen att i framtiden fästa större uppmärksamhet vid frågor som rör möjligheterna att förena arbete och familjeliv när de tillämpar den öppna samordningsmetoden för socialt skydd och social integration, med särskild betoning på tillgången till barnomsorg, familjers inkomstsituationer och mödrarnas sysselsättningsgrad.
57.
Europaparlamentet uppmanar medlemsstaterna att på bästa sätt utnyttja de möjligheter som erbjuds genom den öppna samordningsmetoden, som ett verktyg för politiskt beslutsfattande inom områdena sysselsättning, socialt skydd, social integration, pensioner och hälsa.
58.
Europaparlamentet uppmanar medlemsstaterna – i synnerhet de nya medlemsstaterna – att se över sina pensionssystem och att i samband med detta ta hänsyn till männens betydligt kortare medellivslängd och till de stora löneskillnaderna mellan män och kvinnor som återspeglas av storleken på kvinnors efterlevandepensioner och som ofta leder till att de hamnar under gränsen för fattigdom.
59.
Europaparlamentet framhåller att utvecklingen och upprätthållandet av de sociala trygghetssystemen hänger nära samman med Lissabonmålen och att de kan bidra starkt till ökad sysselsättning och tillväxt, mer solidaritet och bättre social integration.
60.
Europaparlamentet upprepar sin övertygelse om att parlamentets roll i tillämpningen av den öppna samordningsmetoden – i egenskap av det organ som direkt representerar Europas medborgare – måste förtydligas och stärkas för att processen skall kunna bli demokratiskt berättigad.
61.
Europaparlamentet uppmanar rådet och kommissionen att inleda förhandlingar med Europaparlamentet om ett interinstitutionellt avtal som fastställer reglerna för hur man skall välja ut de politiska områden som den öppna samordningsmetoden skall tillämpas på och som gör det möjligt att tillämpa metoden konsekvent, med oinskränkt och jämlikt deltagande från Europaparlamentets sida.
62.
Europaparlamentet betonar att ett sådant interinstitutionellt avtal måste innehålla regler för Europaparlamentets deltagande vid fastställandet av mål och indikatorer och för parlamentets tillgång till handlingar, deltagande i sammanträden, tillsyn och övervakning av utvecklingen, information om rapporter och bästa metoder och ett förfarande som gör att den öppna samordningsmetoden kan utvecklas till en gemenskapsmetod.
°
° °
63.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, Kommittén för socialt skydd, regeringarna och parlamenten i medlemsstaterna, anslutningsländerna och kandidatländerna.
P6_TA(2006)0117
A6-0084/2006
Europaparlamentets beslut om begäran om fastställelse av Witold Tomczaks immunitet och privilegier ( 2005/2129(IMM) )
Europaparlamentet fattar detta beslut
–
med beaktande av Witold Tomczaks begäran om fastställelse av hans immunitet, med anledning av att åtal har väckts mot honom vid distriktsrätten i Ostrów Wielkopolski i Polen, daterad den 29 april 2005 och tillkännagiven i kammaren den 12 maj 2005,
–
–
med beaktande av den skrivelse från Witold Tomczak, undertecknad den 20 mars 2006, i vilken han uttryckte sitt önskemål att dra tillbaka begäran om fastställelse av hans immunitet,
–
–
med beaktande av EG-domstolens domar av den 12 maj 1964 och 10 juli 1986 Mål 101/63, Wagner mot Fohrmann och Krier, svensk specialutgåva I, s.
203 och mål 149/85, Wybot mot Faure m.fl., svensk specialutgåva VIII, s.
703.
,
–
–
med beaktande av betänkandet från utskottet för rättsliga frågor ( A6-0084/2006 ).
A.
B.
Witold Tomczak anklagas för att ha förolämpat två polismän i tjänst i Ostrów Wielkopolski den 26 juni 1999, vilket innebär ett brott mot artikel 226.1 i den polska strafflagen.
Witold Tomczak gick den 4 oktober 2000 med på att ställas till svars i ärendet, i enlighet med artikel 105.4 i Polens konstitution.
C.
D.
Witold Tomczak hävdar att allmänna åklagaren borde ha ingett en begäran om upphävande av hans immunitet till Polens parlament innan åtal väcktes, och eftersom han valts till ledamot av Europaparlamentet var det till detta parlament och inte till det polska parlamentet Sejm som han ställt sin begäran om fastställelse av hans immunitet.
E.
Witold Tomczak uppger att det straffrättsliga förfarandet mot honom inte är opartiskt, att det utövas politiska påtryckningar på de rättsvårdande myndigheterna, att förfalskade bevis inges och att opålitliga vittnen framträder i rättegången.
F.
Mot bakgrund av den information som inkommit skyddas Witold Tomczak inte av parlamentarisk immunitet med avseende på något av de krav som kommit till Europaparlamentets talmans kännedom.
G.
H.
Utan att det påverkar Witold Tomczaks skrivelse om att han önskar dra tillbaka begäran om fastställelse av hans immunitet, betonas att ärendet icke desto mindre måste prövas uttömmande för att garantera att parlamentets privilegier har respekterats på ett korrekt sätt.
1.
Europaparlamentet beslutar att inte fastställa Witold Tomczaks immunitet och privilegier.
P6_TA(2006)0151
Unescos konvention om främjande av och skydd för mångfalden av kulturella uttryck *
A6-0079/2006
Europaparlamentets lagstiftningsresolution om förslaget till rådets beslut om ingående av Unescos konvention om främjande av och skydd för mångfalden av kulturella uttryck (5067/2006 - KOM(2005)0678 – C6-0025/2006 – 2005/0268(CNS) )
(Samrådsförfarandet)
–
med beaktande av förslaget till rådets beslut ( KOM(2005)0678 ) Ännu ej offentliggjort i EUT.
,
–
med beaktande av Unescos konvention om främjande av och skydd för mångfalden av kulturella uttryck, som antogs av Unescos generalkonferens den 20 oktober 2005,
–
–
–
–
med beaktande av betänkandet från utskottet för kultur och utbildning ( A6-0079/2006 ).
1.
Europaparlamentet godkänner ingåendet av Unescos konvention om främjande av och skydd för mångfalden av kulturella uttryck.
2.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen samt regeringarna och parlamenten i medlemsstaterna och Unesco parlamentets ståndpunkt.
P6_TA(2006)0221
Budgeten för 2007: Kommissionens rapport om den årliga politiska strategin
A6-0154/2006
Europaparlamentets resolution om budgeten för 2007: Kommissionens rapport om den årliga politiska strategin ( 2006/2020(BUD) )
–
med beaktande av kommissionens meddelande till Europaparlamentet, rådet, Europeiska ekonomiska och sociala kommittén och regionkommittén - Årlig politisk strategi för 2007: Öka förtroendet genom handling ( KOM(2006)0122 ),
–
med beaktande av det interinstitutionella avtalet av den 6 maj 1999 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och förbättring av budgetförfarandet EGT C 172, 18.6.1999, s.
1.
Avtalet senast ändrat genom Europaparlamentets och Rådets beslut 2005/708/EG (EUT L 269, 14.10.2005, s.
24).
,
–
med beaktande av det reviderade förslaget till ett förnyat interinstitutionellt avtal om budgetdisciplin och förbättring av budgetförfarandet ( KOM(2006)0036 ),
–
,
–
med beaktande av artikel 272 i EG-fördraget och artikel 177 i Euratomfördraget,
–
–
med beaktande av budgetutskottets betänkande och yttrandena från utskottet för utveckling och utskottet för internationell handel ( A6-0154/2006 ).
A.
Institutionerna har kommit fram till en kompromiss om ett nytt interinstitutionellt avtal och en ny flerårig budgetram precis innan budgetförfarandet för 2007 skall inledas.
B.
I avsaknad av ett gällande interinstitutionellt avtal finns bestämmelser för det årliga budgetförfarandet fastlagt i EG-fördraget, särskilt artikel 272.
C.
Mycket av gemenskapslagstiftningen kommer att förnyas 2007, vilket gör det möjligt att i budgeten för 2007 införa nya prioriteringar för den kommande finansiella perioden.
D.
Utvidgningen med Bulgarien och Rumänien torde äga rum 2007.
E.
Valet av prioriteringar för 2007 års budget, den första inom den kommande fleråriga budgetramen, kommer inte bara att lägga fast EU:s politik under det kommande året, utan kommer otvivelaktigt också att få en strategisk roll för kommande år.
F.
G.
Sammanhang
1.
Europaparlamentet uttrycker oro avseende den tydliga diskrepansen mellan de globala utmaningar som Europeiska unionen står inför och de anslag som kan bli tillgängliga under de tillämpliga rubrikerna i en flerårig budgetram 2007–2013 utan ambitioner för att effektivt möta dessa utmaningar, särskilt vad gäller konkurrenskraft, forskning och innovationer som rådet och kommissionen själva har angett som prioriteringar.
2.
3.
Europaparlamentet anser att om man utgår från att 2007 kommer att bli den första budgeten i en ny budgetram bör denna budget vara strategisk till sin karaktär och inriktas mot de interna och externa politikområden där finansiering kan vara av avgörande betydelse och som kan ge verklig valuta för pengarna.
4.
5.
6.
Europaparlamentet anse att när det gäller att slå fast de politiska prioriteringarna bör budgeten för 2007 under de reducerade taken, jämfört med de ursprungliga förväntningarna, koncentreras på ett begränsat antal prioriteringar, särskilt
–
Yttre förbindelser – EU:s roll i en globaliserad värld
-
Partnerskap/Samarbetsavtal
-
Gemenskapens grannskapspolitik och föranslutningsinstrumenten
-
Utvecklingspolitik, demokratisering och mänskliga rättigheter, millennieutvecklingsmålen
-
Den gemensamma utrikes- och säkerhetspolitiken (GUSP)
–
Säkerhets-, frihets- och solidaritetsdimensionen (både extern och intern)
-
Extern, t.ex. energisäkerhet, förebyggande av, förberedelser för och hantering av konsekvenserna av terroristhot
-
Intern, t.ex. invandringspolitik för integration av medborgare i tredjeländer, solidarisk gränsbevakning, säkerhet och försvar för friheter
-
Sammanhållning
–
EU-intern politik
-
Lissabonmålen (tillväxt, sysselsättning, utbildning, transporter, forskning och innovationer)
-
Miljö och landsbygdens utveckling
-
Medborgare (bland annat kultur och ungdom) och kommunikation
-
Anpassning av mål och resurser för den europeiska offentliga förvaltningen inklusive Europeiska gemenskapens organ
7.
8.
9.
Beslut om politiska prioriteringar
A.
Yttre förbindelser – Europa som en global partner
10.
11.
12.
Europaparlamentet välkomnar att kommissionen prioriterar större politisk sammanhållning och effektivare bistånd när det gäller de externa åtgärderna.
13.
Europaparlamentet framhåller sin oro för fågelinfluensans fortsatta utveckling i och utanför Europeiska unionen och understryker att det krävs ett nära samarbete med FAO, WHO, Världsorganisationen för djurens hälsa (OIE) och länderna i de drabbade regionerna.
14.
15.
16.
Europaparlamentet påminner kommissionen och rådet om deras åtaganden att förse de länder som omfattas av sockerprotokollet med adekvat och lämplig finansiering för kompletterande åtgärder som skall hjälpa dem att möta de utmaningar som uppstår under en övergångsperiod till följd av EU:s interna reformering av sockerordningen och de tillämpliga WTO-bestämmelserna.
17.
18.
B.
Säkerhetsdimensionen – Säkerhet, frihet och medborgarskap
19.
20.
21.
22.
23.
Europaparlamentet betonar att målet att integrera invandrarna samt hanteringen av gränserna är viktigt under de kommande åren.
24.
25.
C.
Intern politik – välstånd och solidaritet
26.
27.
28.
29.
30.
31.
D.
Sammanhållning
32.
Kvalitativ valuta för pengarna
33.
34.
35.
36.
Europaparlamentet avser att begära kostnads-nyttoanalyser inom specifika budgetområden genom att använda delar av de resurser som anslagits till parlamentets utskott, för att utvärdera den genomförda politikens efterlevnad (efterlevnad av budgetförordningen, ekonomiska rapportsystem) och resultat (effektivitet i samband med resursanvändning och projekt, administrationskostnader) och att dra de politiska slutsatserna av en sådan utvärdering.
37.
Förberedelse för översynen 2008/2009
38.
39.
Europaparlamentet anser att budgeten för 2007, som den första budgeten under kommande period, innebär ett tillfälle att starta de nya programmen inom ramen för justeringarna till de behov som kan tänkas uppkomma under periodens första del.
40.
EU:s styrning: personella och finansiella resurser för 2007
41.
42.
Europaparlamentet betonar att efter resultaten av förhandlingarna om den nya fleråriga budgetramen bör budgetutskottet se till att de nya bestämmelserna och de kvalitativa reformerna i det nya interinstitutionella avtalet tillämpas i budgeten för 2007.
43.
44.
45.
46.
47.
48.
o
o o
49.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen och revisionsrätten.
P6_TA(2006)0245
Kvinnor i väpnade konflikter och deras roll i återuppbyggnaden efter konflikter
A6-0159/2006
Europaparlamentets resolution om kvinnornarnas situation i väpnade konflikter och deras roll i återuppbyggnaden och den demokratiska processen i länder som just genomgått en konflikt ( 2005/2215(INI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av resolution 1325 (2000) som antogs av FN:s säkerhetsråd den 31 oktober 2000 om kvinnor i fred och säkerhet (nedan kallad UNSCR 1325 (2000)), i vilken betonas vikten av att kvinnor jämställs med män i arbetet med att bevara och främja fred och säkerhet och att de är fullt delaktiga i detta arbete,
–
med beaktande av sin resolution av den 30 november 2000 om kvinnors deltagande i fredlig lösning av konflikter EGT C 228, 13.8.2001, s.
186.
,
–
med beaktande av FN:s allmänna förklaring av den 10 december 1948 om de mänskliga rättigheterna och den förklaring och det handlingsprogram som följde efter världskonferensen om mänskliga rättigheter i Wien den 14–25 juni 1993,
–
med beaktande av FN:s generalsekreterares bulletin om särskilda åtgärder för skydd mot sexuellt utnyttjande och sexuella övergrepp (ST/SGB/2003/13),
–
med beaktande av FN:s förklaring av den 20 december 1993 FN:s generalförsamlings resolution 48/104.
och FN:s konvention av den 20 november 1989 om barnets rättigheter,
–
med beaktande av FN:s konvention om avskaffande av all slags diskriminering av kvinnor (CEDAW) av den 18 december 1979 samt tillhörande fakultativt protokoll,
–
med beaktande av FN:s konvention av den 10 december 1984 mot tortyr och annan grym, omänsklig eller förnedrande behandling eller bestraffning och FN:s förklaring av den 14 december 1974 om skydd av kvinnor och barn i nöd eller väpnade konflikter FN:s generalförsamlings resolution 3318 (XXIX).
, särskilt artikel 4 som innehåller en uppmaning till effektiva åtgärder för att förbjuda förföljelse, tortyr, våld och förnedrande behandling av kvinnor,
–
med beaktande av FN:s säkerhetsråds resolution 1265 (1999) av den 17 september 1999 om skydd av civila vid väpnade konflikter, särskilt artikel 14 i vilken föreskrivs att FN-personal som deltar i fredsbevarande och fredsskapande verksamhet skall ha en lämplig utbildning i människorätt inbegripet könsrollsrelaterade bestämmelser,
–
med beaktande av FN:s resolution av den 15 december 1975 om kvinnors delaktighet i stärkandet av internationell fred och säkerhet FN:s generalförsamlings resolution 3519 (XXX).
, FN:s förklaring av den 3 december 1982 om kvinnors delaktighet i främjandet av internationell fred och internationellt samarbete FN:s generalförsamlings resolution 37/63.
, särskilt artikel 12 om praktiska åtgärder för att öka kvinnors representation i samband med fredsinsatser,
–
med beaktande av den förklaring och det handlingsprogram som följde efter FN:s fjärde världskvinnokonferens i Beijing den 4–15 september 1995, särskilt det kritiska problemområdet E om kvinnor och väpnade konflikter, och resultatdokumentet från FN:s specialsession Beijing + 5 och Beijing + 10 den 5–9 juni 2000 om ytterligare åtgärder och initiativ för att genomföra förklaringen och handlingsprogrammet från Beijing, särskilt artikel 13 om hinder för kvinnors lika deltagande i fredsskapande insatser och artikel 124 om en 50/50-fördelning mellan könen i fredsbevarande uppdrag och vid fredsförhandlingar,
–
med beaktande av Romstadgan som antagits den 17 juli 1998 genom vilken Internationella brottmålsdomstolen inrättades, särskilt artiklarna 7 och 8, i vilka slås fast att våldtäkt, sexuellt slaveri, påtvingat havandeskap eller påtvingad sterilisering och alla andra former av sexuellt våld utgör brott mot mänskligheten och krigsförbrytelser och även skall anses som en särskild form av tortyr och allvarliga krigsförbrytelser, oavsett om de begås på ett systematiskt eller icke-metodiskt sätt, och oavsett om dessa handlingar begås i internationella eller inbördes konflikter,
–
med beaktande av Genèvekonventionerna från 1949 och tilläggsprotokollen från 1977 i vilka anges att kvinnor skall skyddas mot våldtäkt och alla andra former av sexuella övergrepp,
–
med beaktande av resolution 1385 (2004) och rekommendation 1665 (2004) från Europarådets parlamentariska församling om förebyggande och lösning av konflikter: kvinnornas roll, vilken antogs den 23 juni 2004,
–
med beaktande av den resolution som antogs vid den femte europeiska ministerkonferensen om jämställdhet mellan kvinnor och män den 22–23 januari 2003 i Skopje om kvinnors och mäns roll i arbetet med att förebygga konflikter, säkra freden och demokratiseringsprocessen efter konflikter – ur ett jämställdhetsperspektiv,
–
med beaktande av förklaringen om jämställdhet mellan könen: en viktig fråga i samhällen under omvandling, och handlingsprogrammet i samma ämne, vilket antogs vid den ovannämnda femte europeiska ministerkonferensen,
–
med beaktande av beslut nr 14/04 som antogs av OSSE:s ministerråd den 7 december 2004 i Sofia om OSSE:s handlingsplan 2004 för att främja jämställdhet,
–
med beaktande av beslut nr 14/05 som antogs av OSSE:s ministerråd den 6 december 2005 i Ljubljana om kvinnor i konfliktförebyggande arbete, krishantering och återuppbyggnadsarbetet efter konflikter,
–
med beaktande av Europarådets rekommendation nr 5/2002 från ministerkommittén till medlemsstaterna om skydd av kvinnor mot våld under och efter konflikter,
–
med beaktande av rådets "operativa dokument" om genomförandet av UNSCR 1325 (2000) inom ramen för den europeiska säkerhets- och försvarspolitiken (ESFP), såsom det antogs i november 2005,
–
med beaktande av artikel 45 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män och yttrandena från utskottet för utrikesfrågor och utskottet för utveckling ( A6-0159/2006 ), och av följande skäl:
A.
Under konflikter utsätts civila kvinnor, i likhet med barn och äldre, för många övergrepp, däribland sexuella.
B.
Våld mot kvinnor under väpnade konflikter innebär inte bara fysisk och/eller sexuell misshandel, utan kränker också kvinnors ekonomiska, sociala och kulturella rättigheter.
C.
D.
Våldtäkter och sexuella övergrepp används som ett vapen i krig för att förödmjuka och försvaga motståndaren psykologiskt, men offren för dessa metoder blir ofta stämplade, utstötta, misshandlade eller till och med dödade av sina egna, för att det samhälle de lever i skall återvinna sin heder.
E.
Historien har visat att krigföring tycks vara starkt mansdominerad och att det därför finns anledning att tro att kvinnors särskilda förmåga till dialog och icke-våld på ett mycket positivt sätt kan bidra till förebyggande och hantering av konflikter på ett fredligt sätt.
F.
I konflikttider är det svårt för kvinnor att få tillgång till den reproduktiva vård de behöver, till exempel preventivmedel, behandling av sexuellt överförbara sjukdomar, mödravård, abort om kvinnan så önskar, förlossning, eftervård och behandling för klimakteriebesvär.
G.
Frivilligt eller påtvingat sex när kvinnan inte har tillgång till skydd kan främja spridningen av sexuellt överförbara sjukdomar, till exempel hiv, vilket särskilt är fallet vid konflikter och i flyktingläger.
H.
Kvinnor som drabbats av sexuell misshandel i konflikttider får sällan skydd, psykologiskt stöd, läkarvård eller rättshjälp, för att de skall kunna övervinna sina lidanden och för att gärningsmännen skall kunna straffas.
I.
Våld inom äktenskapet, som förekommer under alla konflikter, minskar inte efter en konflikt när de stridande återvänder hem.
J.
Kvinnor som arbetar för fred har i hela världen använt sig av ett föreningsnätverk för att bygga en bro mellan de krigförande och för att kräva rättvisa för sina försvunna anhöriga.
K.
Kvinnliga fredsrörelser arbetar inte alltid medvetet för att förändra de regler och sociala band som definierar maktförhållandena mellan kvinnor och män.
L.
Att kvinnor deltar vid förhandlingsbordet och har aktiva roller under en fredlig övergång är ett nödvändigt men otillräckligt steg på vägen mot demokrati, och dessa kvinnor behöver därför stöd och hjälp med sitt politiska arbete.
M.
I ett fåtal undantagsfall har kvinnor gått från ställningen som politiska motståndare till höga offentliga ämbeten, som Ellen Johnson-Sirleaf i Liberia och Micheline Bachelet i Chile, men dessa fall är fortfarande alltför sällsynta.
N.
Sannings- och försoningskommissioner understödjer försoningsprocessen i samhällen som varit med om en konflikt, men kvinnor deltar alltför sällan i dessa sammanhang.
O.
Vissa länders eller internationella organisationers initiativ till att få med detta könsperspektiv bör välkomnas och fungera som exempel på god praxis.
P.
Det har alltid funnits kvinnor som har varit soldater och tillhört motståndsrörelsen, men i dag ingår de officiellt i många länders väpnade styrkor av jämställdhetsskäl.
Q.
Företeelsen självmordsbombare är relativt ny, begränsad och lokaliserad till länder med islamisk tradition, och antalet kvinnliga självmordsbombare är mycket litet.
R.
Att dessa kvinnor ofta befinner sig i en hopplös situation på det politiska, personliga och sociala planet är en avgörande faktor för deras agerande.
S.
Dagens fundamentalism försöker rättfärdiga martyrdöden, vilket motståndskvinnor och militanta kvinnor som strävar efter social rättvisa är mottagliga för.
T.
Mediernas extrema uppmärksammande av företeelsen gör att självmordsattacker lockar mottagliga ungdomar alltmer, med tanke på den ära som familjen kommer att få efter deras död.
1.
Europaparlamentet understryker att man måste föra in ett genusperspektiv i fredsforskning, i konfliktförebyggande, konfliktlösande och fredsbevarande arbete samt i återanpassning och återuppbyggnad efter konflikter och att man även bör se till att genusaspekten beaktas i fältprogram.
Kvinnor som krigsoffer
2.
3.
4.
5.
Europaparlamentet prioriterar att barnsoldater inte skall användas i konflikter, bland dem flickor som i realiteten fungerar som veritabla sexslavar i dessa sammanhang.
6.
7.
8.
Europaparlamentet understryker att det stora antalet kvinnor och barn bland flyktingar och internt fördrivna som registrerats av internationella organ som resultat av väpnade konflikter och inbördeskrig är mycket oroväckande.
9.
Kvinnor som fredsfaktorer
10.
Europaparlamentet understryker den positiva roll som kvinnor spelar i samband med konfliktlösning, och uppmanar kommissionen och medlemsstaterna att garantera tillräckliga tekniska och ekonomiska bidrag till program som gör det möjligt för kvinnor att delta fullt ut i fredsförhandlingar och att ge kvinnor större ansvar i det civila samhället som helhet.
11.
12.
12 Parlamentet uttrycker sitt starka stöd för den uppmaning som framfördes av en kraftfull koalition av kvinnoorganisationer från Kosovo den 8 mars 2006, i fråga om att inkludera kvinnor i den internationella grupp på sju personer från Kosovo som skall förhandla om regionens framtida status.
13.
Parlamentet välkomnar olika internationella initiativ som verkar i denna riktning, till exempel de australiska organisationerna i Papua Nya Guinea och de norska organisationerna i Sri Lanka.
14.
Europaparlamentet välkomnar olika initiativ för att ta fram könsrelaterade indikatorer för snabba insatser vid och övervakning av konflikter, i likhet med FN:s utvecklingsfond för kvinnor (UNIFEM), Europarådet, Swisspeace, International Alert och Forum on Early Warning and Early Response.
15.
16.
Europaparlamentet upprepar sina tidigare uppmaningar om en effektiv parlamentarisk kontroll av ESFP.
17.
Europaparlamentet betonar att en allmän uppförandekodex för insatser som genomförs inom ramen för ESFP måste tillämpas och utvecklas, varvid man bör se till att kodexen överensstämmer med de bestämmelser som reglerar andra typer av EU-insatser i tredjeländer, liksom med riktlinjerna om skydd för civilbefolkningen i samband med EU-ledda krishanteringsinsatser.
18.
Europaparlamentet välkomnar varmt rådets "operativa rapport" som antogs i november 2005 om genomförandet av UNSCR 1325 (2000) i samband med ESFP.
19.
Europaparlamentet uppmanar EU att stödja åtgärder för att kraftigt öka antalet kvinnor på alla nivåer i ESFP-uppdragen, framför allt att uppmuntra kvinnor att söka sådana befattningar genom att skicka in sina namn för att kandidera till militära, polisiära och politiska tjänster i samband med ESFP-uppdrag, och att göra detta i ett så tidigt skede som möjligt av planeringen av sådana uppdrag.
20.
Europaparlamentet är övertygat om att lokala kvinnoorganisationers delaktighet i en fredsprocess bör vägas in i uppdragsplaneringen inom ESFP i syfte att bygga vidare på det särskilda bidrag som dessa organisationer kan ge och erkänna att kvinnor drabbas på särskilda sätt av en konflikt.
21.
Europaparlamentet uppmanar EU att ägna större uppmärksamhet åt närvaro, förberedelse, utbildning och utrustning för polisstyrkor i militära uppdrag, eftersom polisenheter är det bästa sättet att garantera säkerheten för den civila befolkningen, framför allt kvinnor och barn.
22.
Europaparlamentet välkomnar att det i de nya fredsstyrkorna inom FN:s fredsuppdrag sedan år 2000 finns rådgivare i jämställdhetsfrågor och att en sådan tjänst inrättades 2003 inom avdelningen för fredsbevarande operationer.
23.
Europaparlamentet begär att man inte glömmer bort de modiga kvinnor som valt fredliga former för motstånd och som har betalat, eller fortfarande betalar för detta, genom att fängslas, hållas inspärrade i sina bostäder eller kidnappas.
24.
25.
Europaparlamentet anser det nödvändigt att främja ett ökat deltagande och en ökad närvaro av kvinnor i medierna och i opinionsplattformar genom vilka kvinnor kan föra fram sin åsikt.
26.
27.
Kvinnor som krigsfaktorer
28.
29.
30.
31.
Europaparlamentet uppmanar till en närmare granskning av självmordsattacker som begås av hämnd och av politiska skäl och uppmanar ihärdigt det internationella samfundet att följa internationell rätt och sträva efter fred i framför allt Palestina och Tjetjenien där kvinnor rekryterats eller löper risk att rekryteras för självmordsattacker.
Rekommendationer
32.
Europaparlamentet stöder alla rekommendationer som efter UNSCR 1325 (2000) har syftat till att förbättra kvinnornas öde i konflikter och uppmanar rådet och kommissionen att utan ytterligare dröjsmål infoga och genomföra dessa rekommendationer, framför allt rekommendationerna i dess ovannämnda resolution av den 30 november 2000, i samtliga politikområden.
33.
34.
Europaparlamentet betonar vikten av att kvinnor deltar i diplomatiska insatser och uppmanar medlemsstaterna att rekrytera fler kvinnor som diplomater och utbilda kvinnor inom diplomatin i förhandlings- och medlingsteknik och på så sätt skapa förteckningar över kvinnor som är kvalificerade för freds- och säkerhetsrelaterade befattningar.
35.
Europaparlamentet kräver att begreppen för "övergångsrättvisa" tillämpas på freds- och övergångsprocesser på väg mot en demokrati och en rättsstat, med respekt för offren och kvinnliga vittnens värdighet, och att de innebär att kvinnor deltar i de undersökningskommissioner för försoning som nu håller på att bildas, och att målet om jämställdhet mellan kvinnor och män ingår i de åtgärder som vidtas av dessa kommissioner.
36.
Europaparlamentet föreslår att rekommendationerna begränsas till det absolut viktigaste, nämligen att uppmana institutionerna att söka samverkansvinster genom att vidta konkreta åtgärder tillsammans med andra internationella institutioner som strävar mot samma mål samt att i största möjliga utsträckning utnyttja de nya finansiella instrumenten i budgetramen 2007–2013 som incitament och hävstänger.
37.
Parlamentet föreslår att man i detta projekt anlitar lokala kvinnoorganisationer, sammanslutningar av mödrar, ledare vid ungdomsläger och lärare.
38.
Europaparlamentet uppmanar kommissionen att rapportera till parlamentet om genomförandet av 2003 års riktlinjer om barn och väpnade konflikter.
39.
40.
41.
Europaparlamentet uppmanar kommissionen och andra bidragsgivare att kanalisera resurserna så att de stöder organisationer i det civila samhället att bygga upp kapacitet, och i synnerhet när det gäller lokala kvinnogrupper som arbetar för att lösa konflikter utan våld, samt att erbjuda tekniskt bistånd och yrkesutbildning.
42.
43.
Europaparlamentet begär att integreringen av ett jämställdhetsperspektiv sprids på ett synligt och verifierbart sätt inom samtliga finansiella instrument, särskilt i föranslutningsinstrumentet, den europeiska grannskapspolitiken, instrumentet för utvecklingssamarbete och ekonomiskt samarbete (DCECI) och stabilitetsinstrumentet och att den integreras i villkoren för associeringsavtal.
44.
45.
Europaparlamentet begär att rätten till reproduktiv hälsa skyddas och prioriteras av kommissionen i dess samarbetsinsatser och i stabilitetsinstrumentet, i konfliktdrabbade områden, vilket bör avspeglas i kommissionens budgetposter.
46.
Europaparlamentet betonar att det är nödvändigt att bättre kontrollera fördelningen av livsmedel, kläder och hälsovårdsartiklar såsom sanitetsbindor under krisinsatser, och ber de internationella hjälporganisationerna att verka för säkerhetsinsatser i flyktingläger och att bidra till att förbättra sådana åtgärder i syfte att minska riskerna för våld och sexuella övergrepp mot kvinnor och flickor och att inrätta program för reproduktiv hälsa i flyktingläger och se till att alla kvinnor och flickor som har blivit våldtagna får omedelbar tillgång till bromsmediciner mot HIV (post-exposure prophylaxis).
47.
Europaparlamentet rekommenderar att ett samarbete inleds mellan Europaparlamentet, Europarådet, Nato, alla behöriga FN-organ inklusive UNIFEM, OSSE och eventuellt andra organisationer för införandet av könsspecifika indikatorer som kan övervakas vid konflikter och kunde inlemmas i utrikes- och utvecklingspolitikens nya instrument eller fungera som tidig varning.
48.
Parlamentet uppmanar därför kommissionen att främja en ökning av andelen kvinnor som deltar vid genomförandet av UNSCR 1325 (2000) i sina handlingsplaner och att övervaka utvecklingen mot jämställdhet och lägga fram resultaten för Europaparlamentet.
49.
Europaparlamentet stöder att man i avtal med tredjeländer i tillbörlig utsträckning tillämpar människorättsklausuler och principerna i den internationella människorättslagstiftningen samt tillhörande internationella avtal, och att man därvid ägnar särskild uppmärksamhet åt kvinnornas rättigheter och behov.
50.
Europaparlamentet anser att Europeiska unionens uppförandekod för vapenexport bör göras rättsligt bindande eftersom detta kommer att minska antalet väpnade konflikter runtom i världen och på så sätt avsevärt bidra till att minska kvinnornas lidande.
51.
Europaparlamentet rekommenderar att Europaparlamentet tar upp problemet med självmordsattacker bland kvinnor, inleder en undersökning i ämnet som skall avslutas med en konferens med forskare och andra personer med genuskompetens från berörda länder och från islamska religiösa myndigheter.
o
o o
52.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen och till regeringarna i medlemsstaterna, de anslutande länderna och kandidatländerna.
P6_TA(2006)0257
Europeiska centrumet för kontroll av narkotika och narkotikamissbruk ***I
A6-0124/2006
Europaparlamentets lagstiftningsresolution om förslaget till Europaparlamentets och rådets förordning om Europeiska centrumet för kontroll av narkotika och narkotikamissbruk ( KOM(2005)0399 – C6-0256/2005 – 2005/0166(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2005)0399 ) Ännu ej offentliggjort i EUT.
,
–
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor och yttrandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A6-0124/2006 ).
1.
Europaparlamentet godkänner kommissionens förslag såsom ändrat av parlamentet.
2.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om kommissionen har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
3.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
P6_TC1-COD(2005)0166
Europaparlamentets ståndpunkt fastställd vid första behandlingen den 14 juni 2006 inför antagandet av Europaparlamentets och rådets förordning (EG) nr .../2006 om Europeiska centrumet för kontroll av narkotika och narkotikamissbruk (omarbetning)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 152,
med beaktande av kommissionens förslag,
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande EUT C 69, 21.3.2006, s.
22.
,
med beaktande av Regionkommitténs yttrande,
i enlighet med förfarandet i artikel 251 i fördraget Europaparlamentets ståndpunkt av den 14 juni 2006.
, och
av följande skäl: (1)
Vid mötet i Luxemburg den 28 och 29 juni 1991 godkände Europeiska rådet planen på inrättande av ett europeiskt centrum för kontroll av narkotika.
Ett sådant organ, kallat Europeiska centrumet för kontroll av narkotika och narkotikamissbruk ("centrumet"), inrättades genom rådets förordning (EEG) nr 302/93, av den 8 februari 1993 EGT L 36, 12.2.1993, s.
1.
Förordningen senast ändrad genom förordning (EG) nr 1651/2003 (EGT L 245, 29.9.2003, s.
30).
som har ändrats väsentligt flera gånger Se bilaga II.
.
Med anledning av kommande ändringar bör den av tydlighetsskäl omarbetas.
(2)
På gemenskapsnivå krävs saklig, objektiv, tillförlitlig och jämförbar information om narkotika, narkotikamissbruk och konsekvenser av detta för att ge gemenskapen och medlemsstaterna en heltäckande bild, och därmed förbättra effekten av de åtgärder som de vidtar eller beslutar om inom respektive behörighetsområde för att bekämpa narkotika.
(3)
Narkotikabruket som företeelse innefattar många komplexa och inbördes sammanvävda faktorer som inte utan vidare kan avskiljas.
Centrumet bör därför få i uppgift att sprida allmänna upplysningar till gemenskapen och dess medlemsstater om alla aspekter av problemen med narkotika och narkotikamissbruk.
Denna uppgift bör inte påverka ansvarsfördelningen mellan gemenskapen och dess medlemsstater vad gäller lagstiftning som rör utbudet av och efterfrågan på narkotika.
(4)
Genom beslut nr 2367/2002/EG av den 16 december 2002 EGT L 358, 31.12.2002, s.
1.
Beslutet ändrat genom beslut nr 787/2004/EG (EUT L 138, 30.4.2004, s.
12).
fastställde Europaparlamentet och rådet gemenskapens statistiska program för perioden 2003−2007, som också omfattar gemenskapens statistikinsatser på området hälsa och säkerhet.
(5)
I rådets beslut 2005/387/RIF av den 10 maj 2005 om informationsutbyte, riskbedömning och kontroll avseende nya psykoaktiva ämnen EUT L 127, 20.5.2005, s.
32.
fastställs vilka uppgifter centrumet och dess vetenskapliga kommitté skall ha i systemet för tidig varning och vid utvärderingen av riskerna med nya ämnen.
(6)
Hänsyn bör tas till nya konsumtionsmönster, särskilt blandmissbruk av olaglig narkotika och laglig narkotika eller läkemedel.
(7)
En av centrumets uppgifter bör vara att tillhandahålla information om bästa praxis och riktlinjer i medlemsstaterna och underlätta ömsesidigt utbyte av sådan praxis.
(8)
I rådets resolution av den 10 december 2001 om genomförande av de fem viktigaste epidemiologiska indikatorerna för narkotika uppmanas medlemsstaterna att, särskilt med stöd av nationella kontaktpunkter, se till att det finns jämförbar informationen om dessa indikatorer.
Att medlemsstaterna genomför dessa indikatorer är en förutsättning för att centrumet skall kunna utföra sina uppgifter enligt denna förordning.
(9)
Det är önskvärt att kommissionen till centrumet direkt kan överföra ansvaret för att genomföra gemenskapsprojekt för strukturstöd på området för informationssystem om narkotika i tredje länder, såsom kandidatländerna eller de länder i västra Balkan som efter godkännande av Europeiska rådet får delta i gemenskapens program och organ.
(10)
Centrumets organisation och arbetssätt bör vara inrättade för att uppnå objektiva resultat, dvs. källor och metoder när det gäller information om narkotika måste vara jämförbara och kompatibla.
(11)
Den information som sammanställs av centrumet bör innehålla uppgifter om prioriterade områden, vars innehåll, omfattning och tillämpningsbestämmelser bör definieras.
(12)
Det finns nationella, europeiska och internationella organisationer och organ som redan tillhandahåller sådan information, och centrumet måste kunna utföra sina uppgifter i intimt samarbete med dessa.
(13)
Europaparlamentets och rådets förordning (EG) nr 45/2001 av den 18 december 2000 om skydd för enskilda då gemenskapsinstitutionerna och gemenskapsorganen behandlar personuppgifter och om den fria rörligheten för sådana uppgifter EGT L 8, 12.1.2001, s.
1.
bör tillämpas på centrumets behandling av personuppgifter.
(14)
Centrumet bör även tillämpa de allmänna principer och gränser för rätten till tillgång till handlingar som avses i artikel 255 i fördraget och som har fastställts genom Europaparlamentets och rådets förordning (EG) nr 1049/2001 av den 30 maj 2001 om allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar EGT L 145, 31.5.2001, s.
43.
.
(15)
Centrumet bör vara en juridisk person.
(16)
Med hänsyn till dess storlek bör centrumets styrelse bistås av en verkställande kommitté.
(17)
För att Europaparlamentet skall hållas välinformerat om situationen på narkotikaområdet inom Europeiska unionen, bör parlamentet ha rätt att höra centrumets direktör.
(18)
Centrumets arbete bör vara öppet för insyn och dess ledning bör omfattas av alla gällande bestämmelser om sund förvaltning och bedrägeribekämpning, särskilt Europaparlamentets och rådets förordning (EG) nr 1073/1999 av den 25 maj 1999 om utredningar som utförs av Europeiska byrån för bedrägeribekämpning (OLAF) EGT L 136, 31.5.1999, s.
1.
och det interinstitutionella avtalet av den 25 maj 1999 mellan Europaparlamentet, Europeiska unionens råd och europeiska gemenskapernas kommission om interna utredningar som utförs av Europeiska byrån för bedrägeribekämpning (OLAF) EGT L 136, 31.5.1999, s.
15.
, till vilket centrumet har anslutit sig och för vilket centrumet har utfärdat de nödvändiga genomförandebestämmelserna.
(19)
Centrumets arbete bör regelbundet utvärderas externt, och på grundval av denna utvärdering bör denna förordning i förekommande fall ändras.
(20)
Eftersom målen för denna förordning inte i tillräcklig utsträckning kan uppnås av medlemsstaterna och de därför, på grund av förordningens omfattning och verkningar, bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget.
I enlighet med proportionalitetsprincipen i samma artikel går denna förordning inte utöver vad som är nödvändigt för att uppnå dessa mål.
(21)
Denna förordning står i överensstämmelse med de grundläggande rättigheter och principer som erkänns särskilt i Europeiska unionens stadga om de grundläggande rättigheterna.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Mål
1.
I denna förordning föreskrivs ett Europeiskt centrum för kontroll av narkotika och narkotikamissbruk (nedan kallat centrumet).
2.
Målet med centrumet är att inom de områden som avses i artikel 3 förse gemenskapen och dess medlemsstater med saklig, objektiv, tillförlitlig och jämförbar information på europeisk nivå om narkotika och narkotikamissbruk och konsekvenser av detta.
3.
Syftet med den statistiska, dokumentariska och tekniska information som behandlas eller tas fram är att hjälpa gemenskapen och medlemsstaterna att få en god översikt över situationen vad gäller narkotika och narkotikamissbruk när de vidtar åtgärder eller fattar beslut inom respektive behörighetsområden.
Den statistiska delen av denna information skall utformas i samarbete med de relevanta statistiska myndigheterna, vid behov med hjälp av gemenskapens statistikprogram, så att synergieffekter främjas och dubbelarbete undviks.
Hänsyn skall tas till ytterligare, globalt tillgängliga uppgifter från Världshälsoorganisationen och Förenta nationerna (FN).
4.
5.
Centrumet skall inte samla in några data som gör det möjligt att identifiera enskilda personer eller mindre grupper av personer.
Centrumet skall inte överföra information som hänför sig till specifikt namngivna fall.
Artikel 2
Uppgifter
För att uppfylla målet enligt artikel 1 skall centrumet utföra följande typer av uppgifter inom sitt verksamhetsområde:
a)
Insamling och analys av befintliga data
i)
ii)
iii)
Tillhandahålla ett organisatoriskt och tekniskt system som är i stånd att sprida information om liknande eller kompletterande program eller åtgärder i medlemsstaterna.
iv)
Upprätta och samordna det nätverk som anges i artikel 5 i samarbete med behöriga myndigheter och organisationer i medlemsstaterna.
v)
Underlätta utbyte av information mellan beslutsfattare, forskare, specialister och de personer som arbetar med narkotikarelaterade frågor inom statliga och icke-statliga organ
b)
Förbättring av metoderna för jämförelse av data
i)
ii)
Underlätta och strukturera informationsutbyte, både ur kvalitativ och kvantitativ synvinkel (databaser).
c)
Förmedling av data
i)
Göra den information som tas fram tillgänglig för gemenskapen, medlemsstaterna och behöriga organisationer.
ii)
Se till att arbete som utförts av medlemsstaterna, gemenskapen eller, i förekommande fall, av tredjeländer eller internationella organisationer får stor spridning.
iii)
Se till att de tillförlitliga och icke-konfidentiella uppgifter som samlas in får stor spridning samt på grundval av de uppgifter som centrumet samlar in publicera en årsrapport över situationen på narkotikaområdet, bland annat med uppgifter om nya trender.
d)
Samarbete med europeiska och internationella organ och organisationer och med tredjeländer
i)
Bidra till en bättre samordning av medlemsstaternas och gemenskapens åtgärder på området.
ii)
Arbeta för en integrering av de data om narkotika och narkotikamissbruk som samlas in i medlemsstaterna eller av gemenskapen i internationella program för kontroll av narkotika, i synnerhet de som fastställts av FN och dess särskilda byråer, utan att det påverkar medlemsstaternas skyldigheter när det gäller att lämna uppgifter enligt bestämmelserna i FN:s konventioner om narkotika.
iii)
Bedriva ett aktivt samarbete med Europol för att övervaka narkotikaproblemet så effektivt som möjligt.
iv)
Bedriva ett aktivt samarbete med de organisationer och organ som anges i artikel 20.
v)
På begäran av kommissionen, och med godkännande av den styrelse som avses i artikel 9, överföra sin kunskap till vissa tredjeländer, såsom kandidatländerna eller länderna i västra Balkan, samt bidra till skapande och förstärkande av strukturella kopplingar till det nätverk som avses i artikel 5 samt inrättande och stärkande av de nationella kontaktpunkter som avses i den artikeln.
e)
Informationsskyldighet
Centrumet skall i princip ha skyldighet att informera de behöriga myndigheterna i medlemsstaterna om det får kännedom om ny utveckling och trendförändringar.
Artikel 3
Prioriterade verksamhetsområden
Centrumets mål och uppgifter såsom de definieras i artiklarna 1 och 2 skall genomföras enligt den prioritering som anges i bilaga I.
Artikel 4
Arbetsmetod
1.
2.
För att undvika dubbelarbete skall centrumet, i sin verksamhet, ta hänsyn till det arbete som genomförts av befintliga organisationer eller skall genomföras av framtida organisationer, särskilt Europol, och sträva efter att tillföra något till detta arbete.
Artikel 5
Europeiskt nätverk för information om narkotika och narkotikamissbruk (Reitox)
1.
Till centrumets förfogande skall stå Europeiska nätverket för information om narkotika och narkotikamissbruk (Reitox).
Nätverket skall bestå av en kontaktpunkt för varje medlemsstat och för varje land som har ingått ett avtal enligt artikel 21 samt en kontaktpunkt för kommissionen.
Ansvaret för att utse de nationella kontaktpunkterna skall helt och hållet ligga hos de berörda länderna.
2.
De nationella kontaktpunkterna skall utgöra en länk mellan de deltagande länderna och centrumet.
De skall bidra till utarbetandet av nyckelindikatorer och data, samt av riktlinjer för genomförandet av dessa, i syfte att erhålla tillförlitlig och jämförbar information på unionsnivå.
Kontaktpunkterna skall, på ett objektivt sätt och på nationell nivå, samla in och analysera all relevant information om narkotika och narkotikamissbruk och om den politik och de lösningar som valts, varvid erfarenheter från olika sektorer, såsom hälsovård, rättsväsende och brottsbekämpning, skall samlas i samarbete med experter och nationella organisationer inom det narkotikapolitiska området.
De nationella kontaktpunkterna får till centrumet också lämna information om nya trender när det gäller missbruk av befintliga psykoaktiva ämnen och/eller nya former av kombinationer av psykoaktiva ämnen, som utgör en potentiell folkhälsorisk, samt information om eventuella åtgärder på folkhälsoområdet.
3.
De nationella myndigheterna skall säkerställa att deras kontaktpunkt samlar in och analyserar informationen på nationell nivå på grundval av de riktlinjer som centrumet har antagit.
4.
5.
Samtidigt som centrumet fullt ut skall respektera de nationella kontaktpunkternas företräde, får centrumet, i nära samarbete med kontaktpunkterna, använda sig av kompletterande expertis och informationskällor på området för narkotika och narkotikamissbruk.
Artikel 6
Konfidentialitet och skydd av data
1.
Data om narkotika och narkotikamissbruk som tillhandahålls till eller av centrumet får publiceras under förutsättning att gemenskapsregler och nationella regler om spridning av information och om konfidentialitet är uppfyllda.
Personuppgifter får inte publiceras eller göras tillgängliga för allmänheten.
Medlemsstaterna och de nationella kontaktpunkterna skall inte ha någon skyldighet att tillhandahålla uppgifter som är konfidentiella enligt nationell lagstiftning
2.
Förordning (EG) nr 45/2001 skall tillämpas på centrumet.
Artikel 7
Tillgång till handlingar
1.
Förordning (EG) nr 1049/2001 skall tillämpas på de handlingar som finns hos centrumet.
2.
3.
De beslut som fattas av centrumet i enlighet med artikel 8 i förordning (EG) nr 1049/2001 kan överklagas hos ombudsmannen eller genom att väcka talan inför Europeiska gemenskapernas domstol i enlighet med villkoren i artiklarna 195 och 230 i EG-fördraget.
Artikel 8
Rättskapacitet och lokalisering
1.
Centrumet skall vara en juridisk person.
Det skall i varje medlemsstat ha den mest vittgående rättskapacitet som tillerkänns juridiska personer enligt den nationella lagstiftningen.
Det skall särskilt kunna förvärva och avyttra fast och lös egendom samt föra talan inför domstolar och andra myndigheter.
2.
Centrumet skall ha sitt säte i Lissabon.
Artikel 9
Styrelse
1.
Centrumet skall ha en styrelse som består av en företrädare för varje medlemsstat, två företrädare för kommissionen, två oberoende experter med särskild kompetens inom narkotikaområdet, vilka skall utses av Europaparlamentet, samt en företrädare för varje land som har ingått ett avtal enligt artikel 21.
Varje ledamot av styrelsen skall ha en röst, med undantag för företrädarna för de länder som har ingått avtal enligt artikel 21 som inte skall ha någon rösträtt.
Styrelsen skall fatta beslut med två tredjedels majoritet av dess ledamöter med rösträtt, utom i de fall som avses i punkt 6 i denna artikel och i artikel 20.
Varje ledamot av styrelsen får biträdas eller företrädas av en suppleant.
Suppleanten skall ha rätt att rösta för den ordinarie ledamoten med rösträtt i ledamotens frånvaro.
Styrelsen får bjuda in företrädare för internationella organisationer med vilka man samarbetar i enlighet med artikel 20; dessa deltar då i egenskap av observatörer och har inte rösträtt.
2.
Styrelsens ordförande och vice ordförande skall väljas bland och av ledamöterna för en period av tre år.
De skall kunna omväljas en gång.
Ordföranden och vice ordföranden har rösträtt.
Styrelsen skall själv anta sin arbetsordning.
3.
Styrelsens möten skall sammankallas av ordföranden.
Den skall hålla ett ordinarie möte minst en gång om året.
4.
Styrelsen skall anta ett treårigt arbetsprogram med utgångspunkt från ett utkast som lagts fram av direktören, efter samråd med den vetenskapliga kommitté som avses i artikel 13 och yttrande från kommissionen, och skall översända programmet till Europaparlamentet, rådet och kommissionen.
5.
Medan det treåriga arbetsprogrammet löper skall styrelsen varje år anta centrumets årliga arbetsprogram med utgångspunkt från ett utkast som lagts fram av direktören, efter samråd med den vetenskapliga kommittén och yttrande från kommissionen.
Arbetsprogrammet skall översändas till Europaparlamentet, rådet och kommissionen.
Det får justeras under årets gång enligt samma förfarande.
6.
Om kommissionen reserverar sig mot det treåriga eller årliga arbetsprogrammet, skall styrelsen anta programmen med tre fjärdedels majoritet av ledamöterna med rösträtt.
7.
Styrelsen skall anta årsrapporten om centrumets verksamhet och senast den 15 juni översända den till Europaparlamentet, rådet, kommissionen, revisionsrätten och medlemsstaterna.
8.
Centrumet skall varje år till budgetmyndigheten översända alla uppgifter som rör utvärderingsresultaten.
Artikel 10
Verkställande kommitté
1.
Styrelsen skall biträdas av en verkställande kommitté.
Den skall bestå av styrelsens ordförande och vice ordförande, två andra styrelseledamöter som företräder medlemsstaterna och som har utsetts av styrelsen samt två företrädare för kommissionen.
Direktören skall delta i den verkställande kommitténs möten.
2.
Den verkställande kommittén skall sammanträda minst två gånger om året, och därutöver vid behov, för att förbereda styrelsens beslut och för att bistå och ge direktören råd.
Beslut skall fattas med enhällighet.
Artikel 11
Direktör
1.
Centrumet skall ledas av en direktör som skall utses av styrelsen på förslag av kommissionen för en period på fem år som kan förlängas.
2.
Före sin utnämning till den första av högst två mandatperioder skall styrelsens kandidat till direktörstjänsten omgående uppmanas att göra ett uttalande inför Europaparlamentet och besvara frågor från parlamentets ledamöter.
3.
Direktören skall ansvara för
a)
förberedelse och genomförande av de beslut och program som antas av styrelsen,
b)
den löpande administrationen,
c)
förberedelse av centrumets arbetsprogram,
d)
upprättande av utkastet till beräkning av centrumets intäkter och utgifter samt budgetens genomförande,
e)
förberedelse och publicering av de rapporter som föreskrivs i denna förordning,
f)
hantering av alla personalfrågor, särskilt utövandet av de befogenheter som gäller för en tillsättningsmyndighet,
g)
fastställande av centrumets organisationsstruktur och framläggande av denna inför styrelsen för godkännande,
h)
utförande av de uppgifter som anges i artiklarna 1 och 2,
i)
regelbunden utvärdering av centrumets arbete.
4.
Direktören skall för sin verksamhet vara ansvarig inför styrelsen.
5.
Direktören skall vara centrumets juridiska företrädare.
Artikel 12
Europaparlamentets utfrågning av direktören och styrelsens ordförande
Direktören skall varje år lägga fram den allmänna rapporten över centrumets verksamhet för Europaparlamentet.
Europaparlamentet får dessutom begära att höra direktören och styrelsens ordförande om en fråga som har samband med centrumets verksamhet.
Artikel 13
Vetenskaplig kommitté
1.
Styrelsen och direktören skall biträdas av en vetenskaplig kommitté som i enlighet med denna förordning och på begäran av styrelsen eller direktören skall avge yttrande i vetenskapliga frågor som rör centrumets verksamhet.
Den vetenskapliga kommitténs yttranden skall offentliggöras.
2.
Den vetenskapliga kommittén skall bestå av högst 15 välkända forskare som utsetts av styrelsen på grundval av sin vetenskapliga expertis och oavhängighet, efter det att en uppmaning till intresseanmälan offentliggjorts i Europeiska unionens officiella tidning.
Urvalsförfarandet skall säkerställa att de specialområden som den vetenskapliga kommitténs medlemmar representerar täcker de mest relevanta vetenskapliga områden som har anknytning till narkotika och narkotikamissbruk.
Medlemmarna i den vetenskapliga kommittén skall utses personligen och skall avge sina yttranden helt oavhängigt av medlemsstaterna och gemenskapens institutioner.
Den vetenskapliga kommittén skall ta hänsyn till de olika ståndpunkter som framförs i nationella expertyttranden, då sådana finns, innan den lämnar något yttrande.
3.
Medlemmarna skall utses för en period på tre år, som skall kunna förnyas.
4.
Vetenskapliga kommittén skall välja sin ordförande för en period på tre år.
Kommittén skall sammankallas av ordföranden minst en gång om året.
Artikel 14
Upprättande av budgeten
1.
För varje budgetår, vilket skall motsvara kalenderåret, skall det upprättas en beräkning av centrumets intäkter och utgifter, vilka skall tas upp i centrumets budget.
2.
Det skall råda balans mellan intäkter och utgifter i centrumets budget.
3.
Centrumets intäkter skall, utan att detta påverkar övriga resurser, bestå av bidrag från gemenskapen som tas upp i Europeiska unionens allmänna budget (kommissionens avsnitt), betalningar för utförda tjänster och finansiella bidrag från sådana organisationer, organ och tredje länder som anges i artikel 20 respektive artikel 21.
4.
Centrumets utgifter skall bland annat omfatta
a)
löner till personal och utgifter för administration och infrastruktur samt driftskostnader,
b)
utgifter för stöd till kontaktpunkterna inom Reitox.
5.
Varje år skall styrelsen, på grundval av ett utkast utarbetat av direktören, upprätta en beräkning av centrumets intäkter och utgifter för nästkommande budgetår.
Senast den 31 mars skall styrelsen till kommissionen översända denna beräkning, inklusive ett förslag till tjänsteförteckning, tillsammans med centrumets arbetsprogram.
Kommissionen skall, tillsammans med det preliminära förslaget till Europeiska unionens allmänna budget, översända denna beräkning till Europaparlamentet och rådet (nedan kallade "budgetmyndigheten").
6.
På grundval av den upprättade beräkningen skall kommissionen i det preliminära förslaget till Europeiska unionens allmänna budget ta upp de medel som den betraktar som nödvändiga med avseende på tjänsteförteckningen och storleken på det bidrag som skall belasta den allmänna budgeten, och som den skall förelägga budgetmyndigheten enligt artikel 272 i fördraget.
7.
Budgetmyndigheten skall bevilja de anslag som utgör bidrag till centrumet och anta centrumets tjänsteförteckning.
8.
Styrelsen skall fastställa budgeten.
Den blir definitiv när Europeiska unionens allmänna budget slutligen fastställs.
Den skall i tillämpliga fall anpassas i enlighet därmed.
9.
Styrelsen skall så snart som möjligt underrätta budgetmyndigheten om sin avsikt att genomföra projekt som kan ha betydande ekonomiska konsekvenser för finansieringen av budgeten, särskilt projekt som rör fast egendom, t.ex. hyra eller förvärv av fastigheter.
Den skall informera kommissionen om detta.
Om en enhet inom budgetmyndigheten har meddelat att den har för avsikt att avge ett yttrande, skall den översända detta yttrande till styrelsen inom sex veckor från och med dagen för underrättelse om projektet.
Artikel 15
Genomförande av budgeten
1.
Direktören skall genomföra centrumets budget.
2.
Senast den 1 mars efter utgången av det berörda budgetåret skall centrumets räkenskapsförare till kommissionens räkenskapsförare översända de preliminära räkenskaperna, tillsammans med en rapport om budgetförvaltningen och den finansiella förvaltningen under budgetåret.
Kommissionens räkenskapsförare skall konsolidera institutionernas och de decentraliserade organens preliminära räkenskaper i enlighet med artikel 128 i rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
(nedan kallad den allmänna budgetförordningen).
3.
Senast den 31 mars efter utgången av det berörda budgetåret skall kommissionens räkenskapsförare till revisionsrätten översända de preliminära räkenskaperna, tillsammans med en rapport om budgetförvaltningen och den finansiella förvaltningen under budgetåret.
Rapporten om budgetförvaltningen och den finansiella förvaltningen skall också översändas till Europaparlamentet och rådet.
4.
Efter det att revisionsrättens synpunkter på centrumets preliminära räkenskaper enligt bestämmelserna i artikel 129 i den allmänna budgetförordningen inkommit, skall direktören ansvara för upprättandet av de slutliga räkenskaperna och översända dem till styrelsen för ett yttrande.
5.
Styrelsen skall lämna ett yttrande om centrumets slutliga räkenskaper.
6.
Senast den 1 juli efter utgången av det berörda budgetåret skall direktören översända de slutliga räkenskaperna tillsammans med styrelsens yttrande till Europaparlamentet, rådet, kommissionen och revisionsrätten.
De slutliga räkenskaperna skall offentliggöras.
7.
Senast den 30 september skall direktören till revisionsrätten översända ett svar på dess synpunkter.
Han skall även översända detta svar till styrelsen.
8.
9.
Europaparlamentet skall före den 30 april år n+ 2, på rekommendation av rådet som skall fatta sitt beslut med kvalificerad majoritet, bevilja direktören ansvarsfrihet för budgetens genomförande budgetår n.
10.
Styrelsen skall anta centrumets finansiella regler efter samråd med kommissionen.
Vid utformningen av dessa regler får styrelsen avvika från kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002 EGT L 357, 31.12.2002, s.
72.
, endast om centrumets särskilda förvaltningsbehov kräver detta och efter det att kommissionen gett sitt godkännande.
Artikel 16
Bedrägeribekämpning
1.
När det gäller kampen mot bedrägeri, korruption och annan olaglig verksamhet som påverkar gemenskapens finansiella intressen skall förordning (EG) nr 1073/1999 tillämpas på centrumet utan inskränkning.
2.
I finansieringsbeslut och i avtal och bestämmelser om tillämpning av dessa beslut skall det uttryckligen föreskrivas att revisionsrätten och OLAF vid behov får utföra kontroller på plats hos dem som tar emot medel från centrumet.
Artikel 17
Privilegier och immunitet
Protokollet om Europeiska gemenskapernas immunitet och privilegier skall tillämpas på centrumet.
Artikel 18
Tjänsteföreskrifter
Tjänsteföreskrifterna för tjänstemän i Europeiska gemenskaperna och anställningsvillkoren för övriga anställda i Europeiska gemenskaperna samt de regler som har antagits gemensamt av gemenskapens institutioner för tillämpningen av tjänsteföreskrifterna och anställningsvillkoren skall tillämpas på centrumets personal.
Om centrumet anställer personal från tredjeländer efter ingående av avtal enligt artikel 21, skall det under alla omständigheter rätta sig efter de tjänsteföreskrifter och anställningsvillkor som avses i punkt 1 i den här artikeln.
Centrumet skall gentemot sin personal utöva de befogenheter som gäller för en tillsättningsmyndighet.
Styrelsen skall anta lämpliga tillämpningsbestämmelser i samråd med kommissionen i enlighet med de tjänsteföreskrifter, artikel 110, och anställningsvillkor som avses i punkt 1.
Styrelsen får anta bestämmelser som gör det möjligt att anställa nationella experter från andra medlemsstater genom utstationering vid centrumet.
Artikel 19
Ansvar
1.
Centrumets avtalsrättsliga ansvar skall regleras av den lagstiftning som är tillämplig på avtalet i fråga.
Domstolen skall vara behörig att träffa avgöranden i enlighet med en skiljedomsklausul som ingår i ett avtal som centrumet ingått.
2.
Vad beträffar utomobligatoriskt ansvar skall centrumet ersätta skada som orsakats av centrumet eller av dess anställda under tjänsteutövning, i enlighet med de allmänna principer som är gemensamma för medlemsstaternas rättsordningar.
Domstolen skall ha behörighet att pröva tvister som rör ersättning för sådan skada.
3.
Personalens personliga ansvar gentemot centrumet regleras av de bestämmelser som gäller för centrumets personal.
Artikel 20
Samarbete med andra organisationer och organ
Centrumet skall aktivt söka samarbete med internationella organisationer och andra, särskilt europeiska statliga eller icke-statliga organ med uppgifter på narkotikaområdet, utan att det påverkar de förbindelser som kommissionen får ha i enlighet med artikel 302 i fördraget.
Samarbetet skall bygga på samarbetsarrangemang med de organisationer och organ som avses i första stycket.
Styrelsen skall anta arrangemangen på grundval av ett utkast från direktören efter att ha inhämtat ett yttrande från kommissionen.
Om kommissionen reserverar sig mot arrangemangen, skall styrelsen anta dem med tre fjärdedels majoritet av ledamöterna med rösträtt.
Artikel 21
Tredjeländers deltagande
Tredjeländer som delar gemenskapens och medlemsstaternas intressen och målsättningar med uppgifterna och arbetet inom centrumet skall få möjlighet att delta i centrumets arbete på grundval av avtal som ingåtts mellan sådana tredjeländer och gemenskapen på grundval av artikel 300 i fördraget.
Artikel 22
Domstolens behörighet
Domstolen skall i enlighet med artikel 230 i fördraget vara behörig då talan förs mot centrumet.
Artikel 23
Utvärderingsrapport
Kommissionen skall vart sjätte år ta initiativ till en extern utvärdering av centrumets verksamhet samtidigt med att centrumets treåriga arbetsprogram avslutas.
Utvärderingen skall också omfatta Reitox-systemet.
Kommissionen skall överlämna utvärderingsrapporten till Europaparlamentet, rådet och styrelsen.
Vid behov skall kommissionen i samband med detta lägga fram ett förslag till ändring av bestämmelserna i denna förordning för att ta hänsyn till utvecklingen i fråga om tillsynsmyndigheter, i enlighet med förfarandet i artikel 251 i fördraget.
Artikel 24
Upphävande
Förordning (EEG) nr 302/93 skall upphöra att gälla.
Hänvisningar till den upphävda förordningen skall anses som hänvisningar till denna förordning och skall läsas i enlighet med jämförelsetabellen i bilaga III.
Artikel 25
Ikraftträdande
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Utfärdad i ... den ...
På Europaparlamentets vägnar På rådets vägnar
Ordförande Ordförande
BILAGA I
A.
Centrumets arbete skall utföras med vederbörlig hänsyn till gemenskapens och medlemsstaternas befogenheter på området narkotika, såsom dessa befogenheter definieras i fördraget.
Det skall omfatta de olika aspekterna av problemet med narkotika och narkotikamissbruk och de åtgärder som vidtas för att avhjälpa problemet.
Därvid skall centrumet vägledas av Europeiska unionens narkotikastrategier och handlingsplaner.
Följande områden skall vara prioriterade för centrumet.
1.
Uppföljning av narkotikaproblemet, särskilt genom epidemiologiska indikatorer eller andra indikatorer och uppföljning av nya trender, i synnerhet när det gäller blandmissbruk.
2.
Uppföljning av åtgärder som har vidtagits för att avhjälpa narkotikarelaterade problem; tillhandahållande av information om bästa praxis i medlemsstaterna och underlättande av ömsesidigt utbyte av sådan praxis.
3.
Utvärdering av riskerna med nya psykoaktiva ämnen och bibehållande av ett system för tidig varning avseende användning av sådana ämnen och avseende nya former av missbruk av befintliga psykoaktiva ämnen.
4.
Framtagande av verktyg och instrument som hjälper medlemsstaterna att övervaka och utvärdera respektive lands nationella politik samt kommissionen att övervaka och utvärdera Europeiska unionens politik.
B.
Kommissionen skall till centrumet för vidare spridning överlämna den information och de statistiska data som den till följd av sin behörighet förfogar över.
BILAGA II
Upphävda förordningar med senare ändringar
Rådets förordning (EEG) nr 302/93
EGT L 36, 12.2.1993, s.
1.
Rådets förordning (EG) nr 3294/94
EGT L 341, 30.12.1994, s.
7.
Rådets förordning (EG) nr 2220/2000
EGT L 253, 7.10.2000, s.
1.
Rådets förordning (EG) nr 1651/2003
EUT L 245, 29.9.2003, s.
30.
BILAGA III
JÄMFÖRELSETABELL
Rådets förordning (EEG) nr 302/93
Denna förordning
Artikel 1
Artikel 1
–
Artikel 2 A.1
–
Artikel 2 a i, andra och tredje meningen
Artikel 2 a ii–v
–
Artikel 2 B.7
Artikel 2 b ii
Artikel 2 C.8–10
Artikel 2 c i–iii
Artikel 2 D.11–13
–
Artikel 2 d iii och v
–
Artikel 2 e
Artikel 3
Artikel 4
Artikel 4
Artikel 3
–
–
Artikel 6a
Artikel 7
Artikel 7
Artikel 8
–
–
–
–
–
–
Artikel 10
–
–
–
–
–
Artikel 12
–
Artikel 11a.6 och 11a.7
Artikel 15.6
–
Artikel 16
Artikel 12
Artikel 20
–
Artikel 21
–
Artikel 14
Artikel 17
Artikel 15
–
Artikel 16
Artikel 19
Artikel 17
Artikel 22
Artikel 18
–
–
–
Artikel 24
Artikel 19
Artikel 25
Bilaga, punkt A första stycket
Bilaga I, punkt A, första stycket, första meningen
–
Bilaga I, punkt A, första stycket, andra och tredje meningen
–
Annex I, punkt A, andra stycket, led 1–4
Bilaga, punkt A, andra stycket, led 1–5
–
Bilaga, punkt B
Bilaga I, punkt B
Bilaga, punkt C
–
–
Bilaga II
–
Bilaga III
P6_TA(2006)0304
Ett partnerskap för tillväxt, stabilitet och utveckling mellan EU och Västindien
A6-0211/2006
Europaparlamentets resolution om partnerskapet för tillväxt, stabilitet och utveckling mellan EU och Västindien ( 2006/2123(INI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens meddelande av den 2 mars 2006 till rådet, Europaparlamentet och Europeiska ekonomiska och sociala kommittén "Ett partnerskap för tillväxt, stabilitet och utveckling mellan EU och Västindien", KOM(2006)0086 (nedan kallat "kommissionens meddelande"),
–
med beaktande av kommissionens utvärderingsrapport om en regional strategi för Västindien, volymerna 1 och 2 från april 2005,
–
med beaktande av rådets slutsatser (allmänna frågor och yttre förbindelser) av den 10 april 2006 och dess bekräftande av den gemensamma ståndpunkten om Kuba av den 2 december 1996,
–
med beaktande av den gemensamma förklaringen från rådet och företrädarna för medlemsstaternas regeringar, församlade i rådet, Europaparlamentet och kommissionen om Europeiska unionens utvecklingspolitik "Europeiskt samförstånd" EUT C 46, 24.2.2006, s.
1.
,
–
med beaktande av förklaringen från det tredje forumet för det civila samhället mellan EU och Latinamerika/Västindien i Wien den 1 april 2006,
–
med beaktande av sin resolution av den 23 mars 2006 om utvecklingspåverkan av avtalen om ekonomiskt partnerskap Antagna texter, P6_TA(2006)0113 .
,
–
med beaktande av artikel 45 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för utveckling ( A6-0211/2006 ), och av följande skäl:
A.
Fram till 2020 kommer många västindiska stater att kunna ansluta sig till skaran av industriländer, medan andra riskerar att gå från att ha tillhört gruppen medelinkomstländer till att klassas som låginkomstländer.
B.
Dessa små östater är på grund av sina särdrag sårbara för naturkatastrofer och annan extern påverkan.
C.
D.
Caricoms gemensamma marknad och ekonomi (CSME), som de västindiska staterna själva beslutat att upprätta, utgör ett viktigt instrument för den regionala integrationen.
E.
Cariforum-staterna vill införa en tydlig utvecklingspolitisk dimension i förhandlingarna om ett ekonomiskt partnerskap med EU för att kunna bekämpa den ökande fattigdomen och ojämlikheten, främja den sociala sammanhållningen och genomföra millennieutvecklingsmålen.
F.
Över 60 procent av befolkningen i regionen är under 30 år, och bortsett från Kuba har staterna i Västindien inte löst problemet med utbildning för alla.
G.
Den belgiska regeringen har positiva erfarenheter av den kritiska dialogen och av utvecklingssamarbetet med den kubanska regeringen.
H.
1.
Europaparlamentet uppskattar att Cariforum-gruppen togs med i diskussionen om förslaget till kommissionens meddelande och välkomnar att de flesta av de angelägenheter som regionens stater framfört beaktats i meddelandet.
2.
Europaparlamentet välkomnar att kommissionen i sin strategi lyfter fram den etiska grundsynen om jämlikhet, partnerskap och ägarskap.
3.
Europaparlamentet anser att den faktiska marginaliseringen av parlamentet, genom en tidsplan som omöjliggjorde dess medverkan i formuleringen av samarbetsstrategin för Västindien, på ett högst beklagligt sätt strider mot det förfaringssätt som de tre EU-institutionerna kommit överens om, och som bekräftats i såväl formuleringen av Afrikastrategin som i det europeiska samförståndet om Europeiska unionens utvecklingspolitik.
4.
Europaparlamentet beklagar att kommissionen inte tagit tillräcklig hög grad beaktat rekommendationerna i sin utvärderingsrapport.
5.
Europaparlamentet instämmer i kommissionens analys om att samarbetet mellan de båda regionerna hittills inte har åtföljts av en tillräcklig politisk dialog och anser att nuvarande praxis att en gång vartannat år hålla ett timslångt möte mellan EU-trojkan och regeringscheferna i Cariforum är otillräcklig och välkomnar avsikten att i framtiden avsätta den tid som krävs åt en sådan dialog på alla nivåer.
6.
3)
7.
Europaparlamentet delar uppfattningen hos staterna i Afrika, Västindien och Stillahavsområdet (AVS) att EU:s utformande av olika politiska program för de tre AVS-regionerna ingalunda får leda till en underminering av de övergripande förbindelserna mellan Europeiska unionen och AVS-länderna och välkomnar det extra forum för politisk dialog som skapas genom toppmöten mellan Europeiska unionen och Latinamerikas stater och Västindien, men yrkar dock på de prioriteringar som man enats om inom ramen för Cotonouavtalet.
8.
Europaparlamentet gläder sig över att kommissionen i sitt meddelande gav uttryck för sin avsikt att främja tillförlitliga institutioner och goda styrelseformer samt transparens i de västindiska staterna inom finans- och skatteområdet och det rättsliga området.
9.
Europaparlamentet stöder kommissionens avsikt att prioritera Caricoms nybildade gemensamma marknad och ekonomi, och bekräftar återigen sin åsikt att förhandlingarna om ett ekonomiskt partnerskapsavtal med EU måste föras i enlighet med centralt bestämda utvecklingsmål, att den unga västindiska inhemska marknaden är i behov av handelsrelaterat stöd och kapacitetsuppbyggnad och att liberaliseringen av handeln måste planeras ordentligt.
10.
11.
12.
13.
Europaparlamentet anser att åtgärder för handelsrelaterad kapacitetsuppbyggnad måste beakta begränsningarna på utbudssidan, bland annat genom att stödja bearbetningen av basprodukter och diversifieringen av produktionen, genom att främja samråd med och stöd till små och medelstora företag och genom att avskaffa byråkratiska hinder för investeringar och därmed främja utvecklingen av företagslivet i regionen.
14.
Europaparlamentet uppmanar kommissionen eftertryckligen att genomföra rekommendation 7 i kommissionens utvärderingsrapport, att beakta principerna i Förenta nationernas nätverk av små östater under utveckling och uppmanar kommissionen att offentliggöra den studie som utförts om vilka effekter handelsliberalisering och globalisering har för dessa staters långsiktiga utveckling.
15.
Europaparlamentet ser att det avsatts för små medel till de kompensations- och anpassningsprogram som skall mildra följderna av marknadsförändringarna för socker och bananer och befarar med tanke på den senaste tidens demonstrationer i regionen att den sociala sammanhållningen, som utgör ett mål för utvecklingssamarbetet, allvarligt kan äventyras.
16.
Europaparlamentet uppmanar kommissionen att utveckla program för att främja en omställning av jordbruket, som ur ett socialpolitiskt, energipolitiskt och miljöpolitiskt perspektiv samt ur ett livsmedelsförsörjningsperspektiv gör det möjligt att bibehålla och skapa människovärdiga arbetsplatser på jordbruksföretag som för närvarande drivs med konventionella metoder som inte är konkurrenskraftiga.
17.
Europaparlamentet kräver att sociala, kulturella och miljömässiga konsekvenser ges större tyngd i samarbetsstrategin och att det skapas en systematisk konsekvensanalys och utvärdering baserad på kriterierna i millennieutvecklingsmålen.
18.
Europaparlamentet välkomnar att viktiga miljöskyddsuppgifter tas upp i utvecklingssamarbetet med den västindiska regionen och kräver att utbyggnaden av användningen av förnybara energikällor och energieffektivitet intensivt främjas för att förhindra negativa konsekvenser av prishöjningarna på råolja och för att fördröja klimatförändringen.
19.
20.
Europaparlamentet ställer sig kritisk till att strategin för Västindien inte tillräckligt handlar om att bekämpa problemen med ungdomsarbetslösheten och med den växande frustrationen bland ungdomar och är bekymrad över att situationen ytterligare kommer att förvärras av den förestående krisen i det västindiska jordbruket.
21.
22.
Europaparlamentet välkomnar kommissionens erbjudande om att hålla dörren öppen för en politisk dialog med Kuba, men ställer sig kritisk till att denna begränsas till att hållas inom ramen för den gemensamma ståndpunkten från 1996.
23.
Europaparlamentet påpekar att om Europeiska unionen skulle lyckas påverka Förenta staterna att upphöra med sin embargopolitik skulle detta kunna innebära betydande ekonomiska möjligheter för hela regionen, och rekommenderar i enlighet med en politik som är inriktad på politiska, sociala, individuella och ekonomiska mänskliga rättigheter att det inleds en kritisk dialog med den kubanska regeringen.
24.
Europaparlamentet betonar hur viktigt det är att även samordna utvecklingsåtgärderna med utomeuropeiska aktörer i regionen, särskilt med Kanada, Kina, Brasilien och Venezuela, och beklagar i detta sammanhang att kommissionens beskrivning av andra aktörers engagemang snarast präglas av misstro.
25.
26.
27.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet och kommissionen och till medlemsstaternas regeringar och parlament samt till de västindiska staternas regeringar och parlament.
P6_TA(2006)0350
Uppskjutna förhandlingar i Doharundan för utveckling
B6-0465 , 0468 , 0470 , 0480 och 0484/2006
Europaparlamentets resolution om beslutet att tills vidare skjuta upp förhandlingarna om utvecklingsagendan från Doha
Europaparlamentet utfärdar denna resolution
–
med beaktande av Världshandelsorganisationens (WTO) ministerdeklaration från Doha av den 14 november 2001,
–
,
–
med beaktande av ministerdeklarationen från WTO:s sjätte ministerkonferens som antogs den 18 december 2005 Dokumentnummer 05-6248, dokumentsymbol WT/MIN(05)/DEC).
,
–
A.
Doharundan inleddes 2001 med målet att rätta till den befintliga obalansen i det multilaterala handelssystemet, med utgångspunkt i den allmänna övertygelsen att endast ett multilateralt system som bygger på rättvis handel och rättvisa och rimliga regler kan driva på en verklig utveckling, och placera utvecklingsländernas behov och intressen i centrum för Dohaarbetsporgrammet.
B.
Ett misslyckande med att slutföra Doharundan skulle äventyra det multilaterala handelssystemets trovärdighet och leda till en övergång till bilaterala och regionala handelsavtal, som ofta framhäver obalanserna mellan industriländerna och utvecklingsländerna.
C.
Utvecklingsländerna och de minst utvecklade länderna skulle förlora mest på att rundan skjuts upp, eftersom det länge emotsedda återupprättandet av balansen i handelsbestämmelserna, främjandet av en hållbar utveckling genom handel och beaktandet av det mer omfattande globala styrsystemet inte kan uppnås utanför den multilaterala ramen.
D.
En förlängning av den nuvarande osäkra situationen om framtiden för multilateralismen och själva WTO skulle öka den globala ekonomiska och politiska osäkerheten och få ekonomiska, finansiella och sociala konsekvenser.
E.
WTO:s nuvarande struktur måste reformeras för att underlätta förhandlingarna och öka ansvarsskyldigheten och insynen.
1.
2.
3.
Europaparlamentet betonar att konsekvenserna av uppskjutandet på kort och medellång sikt i första hand kommer att drabba utvecklingsländerna och de minst utvecklade länderna, särskilt om de utvecklingsinriktade åtaganden som gjordes i Hongkong inte längre iakttas.
4.
Parlamentet är bekymrat över att uppskjutandet av de multilaterala förhandlingarna skulle kunna leda till att handelsdispyterna ökar och att WTO:s medlemmar då genom rättsliga processer försöker uppnå det som inte kunde uppnås förhandlingsvägen.
5.
6.
7.
8.
Parlamentet är övertygat om att vi måste utnyttja det nuvarande avbrottet i förhandlingarna till att fundera över vad som krävs för att förbättra de framtida handelsförhandlingarna.
9.
Europaparlamentet uppmanar kommissionen och rådet att ingå ett avtal så att ett fullt deltagande för Europaparlamentet i Europeiska unionens internationella handelsförhandlingar garanteras.
10.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, medlemsstaternas regeringar och parlament samt WTO:s generalsekreterare.
P6_TA(2006)0432
Stödprogram för den europeiska audiovisuella sektorn (Media 2007) ***II
A6-0337/2006
Europaparlamentets lagstiftningsresolution om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets beslut om genomförandet av ett stödprogram för den europeiska audiovisuella sektorn (Media 2007) (6233/2/2006 – C6-0271/2006 – 2004/0151(COD) )
(Medbeslutandeförfarandet: andra behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av rådets gemensamma ståndpunkt (6233/2/2006 – C6-0271/2006 ),
–
med beaktande av parlamentets ståndpunkt vid första behandlingen av ärendet Antagna texter, 25.10.2005, P6_TA(2005)0398 .
, en behandling som avsåg kommissionens förslag till Europaparlamentet och rådet ( KOM(2004)0470 ) Ännu ej offentliggjort i EUT.
,
–
–
med beaktande av artikel 67 i arbetsordningen,
–
med beaktande av andrabehandlingsrekommendationen från utskottet för kultur och utbildning ( A6-0337/2006 ).
1.
Europaparlamentet godkänner den gemensamma ståndpunkten.
2.
Europaparlamentet konstaterar att rättsakten är antagen i enlighet med den gemensamma ståndpunkten.
3.
4.
5.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
P6_TA(2006)0443
Programmet "Ett Europa för medborgarna" (2007-2013) ***II
A6-0342/2006
Europaparlamentets lagstiftningsresolution om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets beslut om inrättande av programmet "Ett Europa för medborgarna" för åren 2007−2013 i syfte att främja ett aktivt europeiskt medborgarskap (9575/1/2006 – C6-0316/2006 – 2005/0041(COD) )
(Medbeslutandeförfarandet: andra behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av rådets gemensamma ståndpunkt (9575/1/2006 – C6-0316/2006 ),
–
med beaktande av parlamentets ståndpunkt vid första behandlingen av ärendet
Antagna texter
, 5.4.2006, P6_TA(2006)0127 .
, en behandling som avsåg kommissionens förslag till Europaparlamentet och rådet ( KOM(2005)0116 ) Ännu ej offentliggjort i EUT.
,
–
–
med beaktande av artikel 62 i arbetsordningen,
–
med beaktande av andrabehandlingsrekommendationen från utskottet för kultur och utbildning ( A6-0342/2006 ).
1.
Europaparlamentet godkänner den gemensamma ståndpunkten såsom ändrad av parlamentet.
2.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
P6_TC2-COD(2005)0041
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artiklarna 151 och 308,
med beaktande av kommissionens förslag,
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande EUT C 28.
,
med beaktande av Regionkommitténs yttrande EUT C 115, 16.5.2006, s.
81.
,
i enlighet med förfarandet i artikel 251 i fördraget Europaparlamentets
ståndpunkt
av den 5 april 2006 (ännu ej offentliggjord i EUT), rådets gemensamma ståndpunkt av den
25 september 2006
(ännu ej offentliggjord i EUT) och Europaparlamentets ståndpunkt av den
25 oktober 2006
(ännu ej offentliggjord i EUT).
, och
av följande skäl: (1)
Genom fördraget inrättas ett medborgarskap i unionen som kompletterar det nationella medborgarskapet.
Det är ett viktigt redskap för att stärka och garantera den europeiska integrationsprocessen.
(2)
Gemenskapen bör göra medborgarna fullt medvetna om deras europeiska medborgarskap, dess fördelar och de rättigheter och skyldigheter som det medför och som bör främjas med vederbörlig hänsyn till subsidiariteten och i sammanhållningens intresse.
(3)
Det är särskilt viktigt att göra unionens medborgare fullt medvetna om deras medborgarskap i Europeiska unionen mot bakgrund av den omfattande reflektion över Europas framtid som inleddes av Europeiska rådet i Bryssel den 16–17 juni 2005.
Programmet "Ett Europa för medborgarna" bör därför vara ett komplement till, men inte överlappa, andra initiativ i detta sammanhang.
(4)
För att medborgarna till fullo skall stödja den europeiska integrationen bör därför större vikt läggas vid deras gemensamma värderingar, historia och kultur såsom centrala inslag i deras tillhörighet till ett samhälle som grundas på principerna om frihet, demokrati och respekt för mänskliga rättigheter, kulturell mångfald, tolerans och solidaritet, i enlighet med Europeiska unionens stadga om de grundläggande rättigheterna EGT C 364, 18.12.2000, s.
1.
(5)
Främjandet av ett aktivt medborgarskap är en avgörande faktor inte bara för att intensifiera kampen mot rasism, främlingsfientlighet och intolerans, utan även för att stärka sammanhållningen och utvecklingen av demokratin.
(6)
Det bör säkerställas att den verksamhet som programmet stöder får bred spridning och stor genomslagskraft inom ramen för EU:s informations- och kommunikationsstrategi.
(7)
För att föra Europa närmare medborgarna och göra det möjligt för dem att full ut delta i uppbyggnaden av ett allt närmare Europa måste man vända sig till alla medborgare och lagligt bosatta i de deltagande länderna och engagera dem i gränsöverskridande utbyten och samarbete och på så sätt bidra till att skapa en känsla av tillhörighet till gemensamma europeiska ideal.
(8)
Europaparlamentet anser i resolutionen som antogs 1988 att betydande ansträngningar bör göras för att intensifiera kontakterna mellan medborgarna i olika medlemsstater och att det både är motiverat och önskvärt att Europeiska unionen särskilt stöder utvecklingen av vänortsverksamhet i medlemsstaterna.
(9)
Europeiska rådet har vid flera tillfällen betonat behovet av att föra Europeiska unionen och dess institutioner närmare medlemsstaternas medborgare.
Rådet har uppmuntrat unionens institutioner att föra och utveckla en öppen, tydlig och regelbunden dialog med det organiserade civila samhället och därigenom främja medborgarnas deltagande i det offentliga livet och i beslutsfattandet, alltmedan man betonar de väsentliga värderingar som är gemensamma för Europas medborgare.
(10)
Rådet upprättade genom sitt beslut 2004/100/EG av den 26 januari 2004 om upprättande av gemenskapens åtgärdsprogram för att främja ett aktivt europeiskt medborgarskap (medborgardeltagande) EUT L 30, 4.2.2004, s.
6.
ett åtgärdsprogram vilket har bekräftat behovet av att främja en kontinuerlig dialog med det civila samhällets organisationer och med lokalsamhällen och att stödja medborgarnas aktiva engagemang.
(11)
Gränsöverskridande och sektorsövergripande medborgarprojekt är viktiga redskap för att nå medborgarna och för att främja den europeiska medvetenheten, den politiska integrationen i Europa samt social integration och ömsesidig förståelse.
(12)
De är också länkar mellan Europa och dess medborgare.
Deras gränsöverskridande samarbete bör därför främjas och uppmuntras.
(13)
Organisationer som bedriver forskning om europeisk offentlig politik kan tillhandahålla idéer och funderingar för att näring åt debatten på europeisk nivå.
De utgör en länk mellan EU-institutionerna och medborgarna och man bör därför stödja sådan verksamhet som speglar deras engagemang i skapandet av en europeisk identitet och ett europeiskt medborgarskap genom att inrätta förfaranden med tydliga kriterier för att främja nätverk för information och utbyte.
(14)
Det är också värdefullt att fortsätta den verksamhet som Europeiska unionen påbörjade inom ramen för Europaparlamentets och rådets beslut nr 792/2004/EG av den 21 april 2004 om upprättande av ett handlingsprogram för gemenskapen för att främja organisationer verksamma på europeisk nivå inom kulturområdet EUT L 138, 30.4.2004, s.
40.
för att bevara och upprätthålla minnet av de viktigaste platserna och arkiven med anknytning till deportationer.
Medvetenheten om andra världskrigets fulla omfattning och tragiska följder kan på så sätt vidmakthållas och den allmänna hågkomsten främjas som ett medel att gå vidare och bygga framtiden.
(15)
I det uttalande om idrott som antogs av Europeiska rådet i Nice den 7–9 december 2000 noterades att "även om gemenskapen inte har direkta befogenheter på detta område bör den i åtgärder i enlighet med fördragets olika bestämmelser beakta idrottens sociala, fostrande och kulturella funktion."
(16)
Särskild uppmärksamhet bör ägnas åt en balanserad integrering av medborgare och det civila samhällets organisationer från alla medlemsstater i gränsöverskridande projekt och insatser.
(17)
Kandidatländerna och de Eftaländer som är parter i EES-avtalet erkänns som potentiella deltagare i gemenskapens program i enlighet med de avtal som ingåtts med dessa länder.
(18)
(19)
Kommissionen och medlemsstaterna bör samarbeta om regelbunden övervakning och oberoende utvärdering av detta program för att möjliggöra de anpassningar som krävs för att åtgärderna skall kunna genomföras på rätt sätt.
(20)
I förfarandena för att följa upp och utvärdera programmet bör det ingå specifika, mätbara, uppnåeliga och tidsbestämda mål och indikatorer för olika tidpunkter.
(21)
Rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 om budgetförordningen för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
(nedan kallad "budgetförordningen") och kommissionens förordning (EG, Euratom) nr 2342/2002 av den 23 december 2002 om genomförandebestämmelser för rådets förordning (EG, Euratom) nr 1605/2002 EGT L 357, 31.12.2002, s.
1.
Förordningen ändrad genom förordning (EG, Euratom) nr 1261/2005 (EUT L 201, 2.8.2005, s.
3).
, vilka slår vakt om gemenskapens finansiella intressen, måste tillämpas med beaktande av principerna om enkelhet och konsekvens i valet av budgetinstrument, en begränsning av antalet fall där kommissionen behåller direkt ansvar för genomförande och administration och den nödvändiga proportionaliteten mellan mängden resurser och den administrativa bördan i samband med användningen av dessa.
(22)
Lämpliga åtgärder bör också vidtas för att förebygga oegentligheter och bedrägeri och för återkrav av medel som försvunnit, betalats ut felaktigt eller använts otillbörligt.
(23)
I enlighet med principen om sund ekonomisk förvaltning kan genomförandet av programmet förenklas genom att man väljer finansiering med ett standardbelopp, antingen för stöd till deltagare i programmet eller stöd från gemenskapen till de organisationer som inrättas på nationell nivå för att förvalta programmet.
(24)
I detta direktiv fastställs en finansieringsram för hela den tid programmet pågår, vilken utgör den särskilda referensen för budgetmyndigheten under det årliga budgetförfarandet enligt punkt 37 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning EUT C 139, 14.6.2006, s.
1.
.
(25)
Eftersom målen för detta beslut inte i tillräcklig utsträckning kan uppnås av medlemsstaterna och de därför, på grund av den gränsöverskridande och mångsidiga arten hos programmets insatser och åtgärder, bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget.
I enlighet med proportionalitetsprincipen i samma artikel går detta beslut inte utöver vad som är nödvändigt för att uppnå dessa mål.
(26)
De åtgärder som är nödvändiga för att genomföra detta beslut bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter EGT L 184, 17.7.1999, s.
23.
Beslutet ändrat genom beslut 2006/512/EG (EUT L 200, 22.7.2006, s.
11).
.
(27)
Övergångsbestämmelser för övervakning av sådana insatser som påbörjas före den 31 december 2006 bör antas i enlighet med beslut 2004/100/EG,
1.
Genom detta beslut inrättas programmet "Ett Europa för medborgarna" (nedan kallat "programmet") för perioden från och med den 1 januari 2007 till och med den 31 december 2013.
2.
Programmet skall bidra till följande allmänna mål:
a)
Att ge medborgarna möjlighet att samarbeta och delta i uppbyggandet av ett allt närmare Europa, som är demokratiskt och öppet mot omvärlden och som enas och berikas genom sin kulturella mångfald, och därigenom utveckla unionsmedborgarskapet.
b)
Att utveckla en känsla av europeisk identitet, grundad på gemensamma värderingar och gemensam historia och kultur.
c)
Att främja medborgarnas känsla av delaktighet i Europeiska unionen.
d)
Att öka
toleransen och
den ömsesidiga förståelsen mellan Europas medborgare och respektera och främja den kulturella och språkliga mångfalden och samtidigt bidra till den interkulturella dialogen.
Programmet skall, i linje med de grundläggande målen i fördraget, ha följande specifika mål, vilka skall genomföras via gränsöverskridande samarbete:
a)
Att föra samman människor från lokalsamhällen i hela Europa, så att de kan dela och utbyta erfarenhet, åsikter och värderingar, lära av historien och bygga för framtiden.
b)
Att genom samarbete inom det civila samhällets organisationer på europeisk nivå främja verksamhet, debatt och reflektion med koppling till EU-medborgarskap, demokrati, gemensamma värderingar och en gemensam historia och kultur.
c)
Att föra Europa närmare medborgarna genom främjande av Europas värderingar och landvinningar, samtidigt som minnet av det förflutna värnas.
d)
Att uppmuntra samverkan mellan medborgare och det civila samhällets organisationer från alla deltagande länder, bidra till interkulturell dialog och framhäva såväl Europas mångfald som dess enighet, med särskild uppmärksamhet på verksamhet vars syfte är att utveckla närmare band mellan medborgare från de medlemsstater som ingick i Europeiska unionen den 30 april 2004 och medborgare från medlemsstater som har anslutit sig efter detta datum.
1.
Programmets mål skall uppnås via stöd till följande insatser, vilka beskrivs utförligare i del I i bilagan:
a)
"Aktiva medborgare för Europa", bestående av
–
vänortssamarbete,
–
medborgarprojekt och stödåtgärder.
b)
"Aktivt civilt samhälle i Europa", bestående av
–
strukturellt stöd till organisationer som bedriver forskning om europeisk offentlig politik (tankesmedjor),
–
strukturellt stöd till det civila samhällets organisationer på europeisk nivå,
–
stöd till projekt till vilka det civila samhällets organisationer tar initiativet.
c)
"Tillsammans för Europa", bestående av
–
mycket synliga evenemang, exempelvis minneshögtider, prisutdelningar, konstnärliga evenemang, Europaomfattande konferenser,
–
studier, undersökningar och opinionsmätningar,
–
verktyg för information och informationsspridning.
d)
"Aktivt europeiskt ihågkommande", bestående av
–
2.
1.
Gemenskapens åtgärder kan genomföras i form av bidrag eller avtal om offentlig upphandling.
2.
Gemenskapens bidrag kan tillhandahållas i specifika former, exempelvis driftsbidrag, bidrag till insatser, stipendier eller priser.
3.
Avtal om offentlig upphandling kommer att täcka inköp av tjänster, exempelvis anordnande av evenemang, studier och undersökningar, verktyg för information och informationsspridning, övervakning och utvärdering.
4.
För att komma i fråga för bidrag måste de sökande uppfylla kraven i del II i bilagan.
Programmet skall vara öppet för deltagare från följande länder, nedan kallade "de deltagande länderna":
a)
Medlemsstaterna.
b)
De Eftaländer som är parter i EES-avtalet, i enlighet med bestämmelserna i avtalet.
c)
De kandidatländer som omfattas av en föranslutningsstrategi, i enlighet med de allmänna principerna och allmänna villkoren i de ramavtal som ingåtts med dessa länder för deras deltagande i gemenskapens program.
d)
Länderna på västra Balkan, i enlighet med de arrangemang som skall fastställas tillsammans med dessa länder enligt ramavtalen om de allmänna principerna för deras deltagande i gemenskapens program.
Programmet skall vara öppet för alla berörda parter som främjar ett aktivt europeiskt medborgarskap, särskilt lokala myndigheter och organisationer, organisationer för forskning om europeisk offentlig politik (tankesmedjor), medborgargrupper och det civila samhällets övriga organisationer.
Programmet får omfatta gemensam och innovativ verksamhet inom aktivt europeiskt medborgarskap tillsammans med berörda internationella organisationer, till exempel Europarådet och Unesco, vilken genomförs på grundval av gemensamma bidrag och enligt budgetförordningen samt varje institutions eller organisations bestämmelser.
1.
Kommissionen skall anta de bestämmelser som är nödvändiga för genomförandet av programmet på det sätt som anges i bilagan.
2.
a)
Bestämmelserna för genomförandet av programmet, inbegripet den årliga arbetsplanen, urvalskriterierna och urvalsförfarandena.
b)
En allmän avvägning mellan programmets olika insatser.
c)
Förfaranden för övervakning och utvärdering av programmet.
d)
Ekonomiskt stöd (belopp, varaktighet, fördelning och bidragsmottagare) från gemenskapen vad gäller alla driftsbidrag, fleråriga vänortsavtal enligt insats 1 och mycket synliga evenemang enligt insats 3.
3.
4.
Som del i det förfarande som avses i punkt 2 får kommissionen fastställa riktlinjer för var och en av insatserna i bilagan för att anpassa programmet till eventuella ändringar i prioriteringarna när det gäller aktivt europeiskt medborgarskap.
Artikel 9
1.
Kommissionen skall biträdas av en kommitté.
2.
3.
När det hänvisas till denna punkt skall artiklarna 3 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
4.
Kommittén skall själv anta sin arbetsordning.
1.
Kommissionen skall se till att detta program stämmer överens med och kompletterar instrument på andra områden som omfattas av gemenskapens insatser, särskilt allmän och yrkesinriktad utbildning, kultur, ungdom, idrott, miljö, audiovisuell sektor och medier, grundläggande fri- och rättigheter, social integrering, jämställdhet, bekämpning av alla former av diskriminering, rasism och främlingsfientlighet, vetenskaplig forskning, informationssamhället samt gemenskapens yttre insatser, särskilt inom den europeiska grannskapspolitiken.
2.
Programmet får dela medel med gemenskapens eller Europeiska unionens övriga instrument för att genomföra insatser som motsvarar målen såväl i detta program som i dessa övriga instrument.
1.
.
2.
De årliga anslagen skall godkännas av budgetmyndigheten inom budgetramen.
1.
Det ekonomiska stödet skall utges i form av bidrag till juridiska personer.
Allt efter insatsens art och mål får bidrag även beviljas fysiska personer.
2.
Kommissionen får dela ut priser till fysiska eller juridiska personer för insatser eller projekt som genomförs inom ramen för programmet.
3.
I enlighet med artikel 181 i förordning (EG, Euratom) nr 2342/2002 får schablonfinansiering eller tillämpning av enhetskostnadstariffer tillåtas, allt efter insatsens art.
4.
Samfinansiering in natura får tillåtas.
5.
Allt efter bidragsmottagarnas egenskaper och insatsernas art får kommissionen besluta att undanta bidragsmottagarna från kontroll av att de förfogar över den yrkeskompetens och de yrkeskvalifikationer som krävs för att genomföra den föreslagna insatsen eller arbetsprogrammet.
6.
Den mängd information som skall lämnas av bidragsmottagaren får begränsas när det rör sig om små bidrag.
7.
I särskilda fall, t.ex. vid beviljandet av små bidrag, behöver bidragsmottagaren inte avkrävas bevis på ekonomisk förmåga att utföra det planerade projektet eller arbetsprogrammet.
8.
Driftsbidrag som beviljas inom programmet till organisationer som arbetar för mål av allmänt europeiskt intresse enligt definitionen i artikel 162 i förordning (EG, Euratom) nr 2342/2002 skall inte minskas automatiskt vid förlängning.
1.
Kommissionen skall när åtgärder enligt detta beslut genomförs se till att gemenskapens ekonomiska intressen skyddas, genom förebyggande åtgärder mot bedrägeri, korruption och annan olaglig verksamhet, genom verkningsfulla kontroller och återkrävande av orättmätigt utbetalda belopp och, om oegentligheter påvisas, verkningsfulla, proportionella och avskräckande påföljder i enlighet med rådets förordning (EG, Euratom) nr 2988/95 av den 18 december 1995 om skydd av Europeiska gemenskapernas finansiella intressen EGT L 312, 23.12.1995, s.
1.
, rådets förordning (Euratom, EG) nr 2185/96 av den 11 november 1996 om de kontroller och inspektioner på platsen som kommissionen utför för att skydda Europeiska gemenskapernas finansiella intressen mot bedrägerier och andra oegentligheter EGT L 292, 15.11.1996, s.
2.
och Europaparlamentets och rådets förordning (EG) nr 1073/1999 av den 25 maj 1999 om utredningar som utförs av Europeiska byrån för bedrägeribekämpning (OLAF) EGT L 136, 31.5.1999, s.
1.
.
2.
unionens
allmänna budget eller budgetar som
gemenskaperna
förvaltar, genom en otillbörlig utgift.
3.
Kommission skall sänka, hålla inne eller återkräva ekonomiskt stöd som har beviljats för en insats, om det visar sig att oegentligheter har förekommit, exempelvis att bestämmelserna i detta beslut, ett enskilt beslut eller avtalet om stöd inte har följts eller om det framkommer att insatsen har ändrats på ett sätt som står i strid med projektets art eller genomförandevillkor, utan att kommissionens godkännande har sökts.
4.
Om tidsfristerna inte har iakttagits eller om verksamheten utvecklas så att endast en del av det tilldelade ekonomiska stödet är berättigat, skall kommissionen begära att bidragsmottagaren yttrar sig inom en viss tid.
Om bidragsmottagaren inte ger en tillfredsställande förklaring, kan kommissionen annullera det resterande ekonomiska stödet och kräva återbetalning av tidigare utbetalda belopp.
5.
Alla felaktigt utbetalda belopp skall återbetalas till kommissionen.
Ränta skall läggas till belopp som inte återbetalas i tid enligt villkoren i budgetförordningen.
1.
Kommissionen skall se till att programmet regelbundet följs upp.
Resultaten av uppföljningen och utvärderingen skall tas tillvara då programmet genomförs.
De specifika målen får ses över i enlighet med artikel 251 i fördraget.
2.
Kommissionen skall se till att det görs regelbundna, externa och oberoende utvärderingar av programmet och regelbundet lämna rapporter till Europaparlamentet.
3.
Kommissionen skall till Europaparlamentet, rådet, Europeiska ekonomiska och sociala kommittén samt Regionkommittén överlämna följande:
a)
En utvärderingsrapport efter halva tiden om resultaten och om de kvalitativa och kvantitativa aspekterna av genomförandet av programmet, senast den 31 december 2010.
b)
Ett meddelande om fortsättningen av programmet, senast den 31 december 2011.
c)
En utvärderingsrapport efter programmets avslutning, senast den 31 december 2015.
För insatser som påbörjas före den 31 december 2006 i enlighet med beslut 2004/100/EG skall det beslutet fortsätta att tillämpas tills de avslutas.
I enlighet med artikel 18 i budgetförordningen kan anslag som motsvarar inkomster som avsatts för ett särskilt ändamål och kommer från återbetalning av belopp som betalats ut på felaktiga grunder enligt beslut 2004/100/EG göras tillgängliga för programmet.
Detta beslut träder i kraft
dagen
Ordförande Ordförande
BILAGA
I.
BESKRIVNING AV INSATSERNA
Kompletterande information om tillträde till programmet
De civila samhällets organisationer som avses i artikel 6 kan bland annat innefatta fackföreningar, utbildningsinstitutioner och organisationer för frivilligt arbete samt amatöridrott.
INSATS 1: Aktiva medborgare för Europa
Denna insats utgör den del av programmet som är särskilt inriktad på verksamhet i vilken medborgarna medverkar.
Denna verksamhet delas in i följande två slags åtgärder:
Vänortssamarbete
Denna åtgärd avser verksamhet som inbegriper eller främjar direkt utbyte mellan Europas medborgare genom deltagande i vänortssamarbete.
Det kan röra sig om enstaka insatser eller pilotverksamhet eller strukturerade, fleråriga arrangemang med flera partner vilka följer ett mer planerat tillvägagångssätt och inbegriper en rad aktiviteter, från möten mellan medborgare till specifika konferenser eller seminarier, anordnade inom ramen för vänortssamarbete, kring ämnen av gemensamt intresse tillsammans med därtill kopplade publikationer.
Denna åtgärd kommer att aktivt bidra till att öka kunskaperna och förståelsen mellan medborgare och kulturer.
Medborgarprojekt och stödåtgärder
Denna åtgärd omfattar stöd till en rad olika transnationella och sektorsövergripande projekt i vilka medborgare medverkar direkt.
Projekt vilkas syfte är att främja deltagande på lokal nivå kommer att prioriteras.
Projektens omfattning och räckvidd kommer att bero på utvecklingen i samhället och de kommer att inriktas på att via innovativa tillvägagångssätt söka möjliga lösningar på kartlagda behov.
Man kommer att uppmuntra användningen av ny teknik, särskilt informationssamhällets teknik (IST).
Projekten kommer att samla medborgare med olika bakgrund, vilka tillsammans kommer att arbeta med eller diskutera gemensamma europeiska frågor och på så sätt utveckla ömsesidig förståelse och göra människor mer uppmärksamma på den europeiska integrationsprocessen.
För att förbättra vänortssamarbete och medborgarprojekten är det också nödvändigt att utarbeta stödåtgärder för utbyte av bästa praxis, dela erfarenheter mellan berörda partner på lokal och regional nivå, inbegripet offentliga myndigheter, samt utveckla nya färdigheter, till exempel genom utbildning.
45 %
INSATS 2: Aktivt civilt samhälle i Europa
Strukturellt stöd till organisationer för forskning om europeisk offentlig politik (tankesmedjor)
Organisationer med nya idéer och funderingar kring europeiska frågor är viktiga institutionella samtalspartner, vilka kan lämna oberoende strategiska och sektorsövergripande rekommendationer till EU-institutionerna.
De kan företa insatser som ger näring till debatten, särskilt om EU-medborgarskap och om europeiska värderingar och kulturer.
Denna åtgärd syftar till att stärka den institutionella kapaciteten hos de organisationer som är representativa, tillhandahåller ett verkligt europeiskt mervärde, kan få till stånd betydande multiplikatoreffekter och kan samarbeta med övriga bidragsmottagare inom programmet.
Förstärkningen av Europaomfattande nätverk är ett viktigt inslag på detta område.
Bidrag får beviljas på grundval av fleråriga arbetsprogram där en rad teman eller aktiviteter ingår.
Strukturellt stöd till det civila samhällets organisationer på europeisk nivå
Det civila samhällets organisationer är en viktig del av medborgerlig, kulturell och politisk verksamhet och utbildning för delaktighet i samhället.
De behöver finnas och ha möjlighet att fungera och samarbeta på europeisk nivå.
De bör även kunna delta i det politiska beslutsfattandet i egenskap av rådgivande organ.
Denna åtgärd kommer att ge dem kapacitet och stabilitet att på ett sektorsöverskridande och övergripande sätt fungera som katalysatorer över gränserna för sina medlemmar och för det civila samhället på europeisk nivå och därigenom bidra till programmets mål.
Förstärkningen av Europaomfattande nätverk och europeiska föreningar är ett viktigt inslag på detta verksamhetsområde.
Bidrag får beviljas på grundval av fleråriga arbetsprogram där en rad teman eller aktiviteter ingår.
Det civila samhällets organisationer på lokal, regional, nationell eller europeisk nivå engagerar medborgarna eller företräder deras intressen genom debatt, publikationer, opinionsbildning och andra konkreta gränsöverskridande projekt.
Att införa eller bygga vidare på en europeisk dimension i verksamheten hos det civila samhällets organisationer kommer att göra det möjligt för dem att öka sin kapacitet och nå en större publik.
Direkt samarbete mellan det civila samhällets organisationer från olika medlemsstater kommer att bidra till ömsesidig förståelse för olika kulturer och ståndpunkter och till fastställandet av gemensamma angelägenheter och värderingar.
Även om detta kan ske i form av enskilda projekt, kommer ett mer långsiktigt tillvägagångssätt att säkerställa en mer hållbar effekt och utveckling av nätverk och synergieffekter.
Som vägledning kan nämnas att cirka
31 %
av programmets sammanlagda budget kommer att användas till denna insats.
INSATS 3: Tillsammans för Europa
Mycket synliga evenemang
Inom denna åtgärd stöds evenemang som anordnas av kommissionen, om lämpligt i samarbete med medlemsstaterna eller andra relevanta partner, vilka är av betydande skala och räckvidd, berör Europas folk, bidrar till att öka deras känsla av att tillhöra samma gemenskap, gör dem medvetna om Europeiska unionens historia, resultat och värderingar, engagerar dem i den i interkulturella dialogen och bidrar till utvecklingen av deras europeiska identitet.
Dessa evenemang kan exempelvis vara minneshögtider kring historiska händelser, uppmärksammande av europeiska framgångar, konstnärliga evenemang, medvetandegörande kring bestämda frågor, Europaomfattande konferenser samt prisutdelningar för att uppmärksamma betydande resultat.
Användning av ny teknik, särskilt IST, skall uppmuntras.
Studier
För att få en bättre insikt i aktivt medborgarskap på europeisk nivå kommer kommissionen att utföra studier, undersökningar och opinionsmätningar.
Verktyg för information och informationsspridning
Med tanke på programmets inriktning på medborgare och de olika initiativen inom aktivt medborgarskap måste övergripande information om verksamheten inom programmet, övriga insatser i Europa i samband med medborgarskap och andra relevanta initiativ tillhandahållas via en Internetportal och andra verktyg.
Som vägledning kan nämnas att cirka 10 % av programmets sammanlagda budget kommer att användas till denna insats.
INSATS 4: Aktivt Europeiskt ihågkommande
Inom denna åtgärd kan projekt av följande slag få stöd:
–
Projekt för att bevara de viktigaste platserna och minnesmärkena med anknytning till massdeportationerna, de tidigare koncentrationslägren och andra platser för martyrskap och massutrotning under nazismen och de arkiv som dokumenterar dessa händelser samt för att bevara minnet av offren och av dem som under extrema förhållanden räddade människor undan förintelsen.
–
Projekt för att bevara minnet av offren för massutrotningar och massdeportationer med anknytning till stalinismen samt bevarande av de minnesmärken och arkiv som dokumenterar dessa händelser.
Cirka 4 % av programmets sammanlagda budget kommer att användas till denna insats.
II.
PROGRAMMETS FÖRVALTNING
Programmet kommer att genomföras enligt principerna om öppenhet och tydlighet och omfatta en bred skala av organisationer och projekt.
Undantag blir möjliga bara under mycket speciella omständigheter och helt i enlighet med artikel 168.1 c och 168.1 d i förordning (EG, Euratom) nr 2342/2002.
Programmet kommer att tillämpa principen med fleråriga partnerskap som baseras på överenskomna mål och bygger på analyser av resultat, så att både det civila samhället och Europeiska unionen får nytta av det.
Finansiering som tilldelas genom ett avtal om engångsbidrag inom detta program får ha varaktighet på högst tre år.
För vissa insatser kan det bli nödvändigt med indirekt centraliserad förvaltning, genom ett verkställande organ eller, särskilt för insats 1, genom nationella organ.
Alla insatser kommer att genomföras via samarbete över gränserna.
De kommer att främja rörlighet för medborgare och idéer inom Europeiska unionen.
Arbete i nätverk och inriktning på multiplikatoreffekterna, inbegripet användning av informations- och kommunikationsteknik (IKT), blir viktigt och kommer att återspeglas både i typen av verksamhet och raden av medverkande organisationer.
Man kommer att uppmuntra till samverkan och synergi mellan de olika berörda parterna i programmet.
Ur programmets budget får man även täcka de utgifter i samband med förberedelser, uppföljning, övervakning, revision och utvärdering som är direkt nödvändiga för förvaltningen av programmet och förverkligandet av dess mål, särskilt studier, möten, informations- och publikationsverksamhet, utgifter i samband med IKT-nätverken för utbyte av information och alla övriga utgifter för administrativt och tekniskt stöd som kommissionen kan besluta om för programmets förvaltning.
De totala administrativa kostnaderna för programmet bör stå i proportion till de uppgifter som fastställs i det berörda programmet och bör, som vägledning, utgöra cirka 10 % av den totala budgeten för programmet.
Kommissionen kan även bedriva sådan verksamhet som avser information, publikation och spridning och därigenom säkerställa en bred kunskap om och stor genomslagskraft för de verksamheter som stöds genom programmet.
III.
GRANSKNINGAR OCH REVISIONER
För projekt som väljs ut i enlighet med detta beslut kommer man att fastställa ett revisionssystem baserat på stickprov.
Bidragsmottagarna måste för kommissionen lägga fram alla verifikationer i samband med utgifter under fem år efter den sista utbetalningen.
Mottagaren skall i förekommande fall se till att styrkande handlingar som innehas av dennes partner eller medlemmar görs tillgängliga för kommissionen.
Kommissionen får genomföra en granskning av hur bidraget har använts, antingen direkt av kommissionens egen personal eller av någon kvalificerad extern organisation som den väljer.
En sådan granskning får utföras under hela avtalets löptid samt under fem år efter den dag då slutbetalning sker.
Resultaten av dessa revisioner kan eventuellt leda till att kommissionen fattar beslut om återkrav.
Kommissionens personal och extern personal som bemyndigas av kommissionen måste få tillträde till bidragsmottagarens lokaler och tillgång till all information som behövs för att genomföra sådana revisioner, inbegripet information i elektronisk form.
Revisionsrätten och Europeiska byrån för bedrägeribekämpning (Olaf) bör ha samma rättigheter som kommissionen, särskilt vad gäller tillträde.
P6_TA(2006)0452
Förslag till allmän budget 2007 (avsnitt I, II, IV, V, VI, VII, VIII)
A6-0356/2006
Europaparlamentets resolution om förslaget till Europeiska unionens allmänna budget för budgetåret 2007, Avsnitt I - Europaparlamentet, Avsnitt II - Rådet, Avsnitt IV - Domstolen, Avsnitt V - Revisionsrätten, Avsnitt VI - Europeiska ekonomiska och sociala kommittén, Avsnitt VII - Regionkommittén, Avsnitt VIII (A) - Europeiska ombudsmannen - Avsnitt VIII (B) -Europeiska datatillsynsmannen ( C6-0300/2006 - 2006/2018(BUD) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av artikel 272 i EG-fördraget,
–
med beaktande av rådets beslut 2000/597/EG, Euratom av den 29 september 2000 om systemet för Europeiska gemenskapernas egna medel EGT L 253, 7.10.2000, s.
42.
,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
,
–
med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning EUT C 139, 14.6.2006, s.
1.
,
–
med beaktande av det interinstitutionella avtalet av den 6 maj 1999 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och förbättring av budgetförfarandet EGT C 172, 18.6.1999, s.
1.
Avtalet senast ändrat genom Europaparlamentets och rådets beslut 2005/708/EG (EUT L 269, 14.10.2005, s.
24).
, särskilt punkt 26,
–
med beaktande av parlamentets resolution av den 15 mars 2006 om riktlinjerna för 2007 års budgetförfarande – avsnitt II, IV, V, VI, VII, VIII (A) och VIII (B) och om det preliminära förslaget till Europaparlamentets budgetberäkning (avsnitt I) för budgetförfarandet för budgetåret 2007 Antagna texter, P6_TA(2006)0090 .
,
–
med beaktande av parlamentets resolution av den 1 juni 2006 om Europaparlamentets beräknade inkomster och utgifter för budgetåret 2007 Antagna texter, P6_TA(2006)0241 .
,
–
med beaktande av det preliminära förslag till Europeiska unionens allmänna budget för budgetåret 2007 som kommissionen lade fram den 3 maj 2006 ( SEK(2006)0531 ),
–
med beaktande av det förslag till Europeiska unionens allmänna budget för budgetåret 2007 som rådet fastställde den 14 juli 2006 ( C6-0300/2006 ),
–
med beaktande artikel 69 och bilaga IV i arbetsordningen,
–
med beaktande av betänkandet från budgetutskottet och yttrandena från utskottet för internationell handel, utskottet för utveckling, utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor och utskottet för framställningar ( A6-0356/2006 ), och av följande skäl:
A.
År 2007 är det första året under den nya budgetramen 2007–2013 för vilket taket för rubrik 5 (administrativa utgifter) har fastställts till 7 115 000 000 EUR i löpande priser.
B.
I det preliminära budgetförslaget för samtliga institutioner lämnades en marginal på 160 750 000 EUR under taket för budgetramens rubrik 5 för budgetåret 2007.
C.
Efter rådets beslut har budgetförslaget en marginal på 285 190 000 EUR under taket för rubrik 5 för 2007.
Allmän ram
1.
2.
3.
4.
5.
Parlamentet rekommenderar att 30 389 840 EUR återinförs utav den minskning på 47 812 781 EUR som rådet gjorde i budgeten för övriga institutioner (med undantag av kommissionen).
6.
7.
Europaparlamentet välkomnar att institutionerna antagit en ny kontoplan som gör presentationen av budgetdokument mer begriplig och tydlig för medborgarna men anser att den kan förbättras ytterligare.
8.
9.
10.
Dessa rapporter kunde användas för att bättre motivera äskanden om extraanslag och samtidigt göra det möjligt för budgetmyndigheten att fatta mer rationella beslut när det gäller tilldelning av sådana anslag.
11.
12.
13.
Europaparlamentet hävdar att anslag så långt som möjligt skall knytas till specifika verksamheter så att annulleringar av anslag och uppsamlingsöverföringar i slutet av året kan undvikas.
14.
Europaparlamentet stöder inte rådets beslut att öka "schablonminskningen" till en relativt hög nivå och basera den på det befintliga antalet lediga tjänster eftersom detta potentiellt skulle kunna skapa en del onödiga problem, särskilt om godkända sökande inte kan anställas på grund av brist på anslag.
15.
Europaparlamentet rekommenderar former av samarbete mellan institutioner vilka nödvändigtvis måste skapa synergieffekter och bidra till ekonomiska besparingar och större effektivitet, samtidigt som det hjälper medborgarna att bättre förstå EU:s roll i deras vardagsliv.
16.
Europaparlamentet uppmanar institutionerna att använda sig av ett mer harmoniserat och standardiserat tillvägagångssätt när de utarbetar sina budgetberäkningar, med tydliga och exakta motiveringar, eftersom detta skulle underlätta deras analys.
Avsnitt I — Europaparlamentet
Budgeteringsnivå
17.
Europaparlamentet uppmanar presidiet att åter diskutera det självpåtagna taket på 20 procent av rubrik 5 under de kommande åren, där man beaktar utvecklingen och de åtföljande behoven för parlamentet för 2009 och därefter.
18.
19.
20.
Informations- och kommunikationspolitiken
21.
22.
Europaparlamentet beslutar att ändra kontoplanen och inrätta två nya budgetposter för besökscentrumet och webb-TV i syfte att förbättra insynen i ekonomin samt ansvars- och redovisningsskyldigheten.
23.
24.
25.
26.
27.
28.
Europaparlamentet har beslutat att följa presidiets förslag angående följande anslag:
-
Att anslå ett extra belopp på 2 700 000 EUR för besöksprogrammet.
-
-
Att i kapitel 10 4 ("Reserv för informations- och kommunikationspolitiken") bibehålla ett belopp på 15 700 000 EUR för audiovisuell utrustning i D5-byggnaden.
29.
Utvidgningen
30.
Europaparlamentet bekräftar sitt beslut att införa ett anslag på 48 000 000 EUR för utvidgningsrelaterade utgifter (Rumänien och Bulgarien) när det gäller följande:
1.
Utgifter knutna till nya ledamöter (35 rumäner och 18 bulgarer).
2.
Ytterligare personal (de återstående 113 utav 226 fasta tjänster och 22 tillfälliga tjänster för de politiska grupperna).
3.
Tolkning och konferenstekniker.
4.
Utrustning och möbler.
5.
Verksamhetsutgifter.
6.
Information och stadgeenlig finansiering av politiska grupper och partier.
31.
Tjänsteförteckningen
32.
33.
-
Iriska: 3 AD5 (granskningsjurister), 3 AD5 (översättare) och 3 AST3.
-
-
Kommittéförfarande: 5 AD5 och 2 AST3.
-
Bättre lagstiftning: 1 AD5.
-
Budgetkontroll: 1 AD5 och direktorat D: 1 AST3.
-
Utbyggnad av KAD-fastigheten: 1 AD5 och 2 AST3, av vilka en förs till reserven.
-
Webb-TV: 1 AD9, 2 AD5 och 2 AST3 i reserven.
-
EMAS: 1 AST3.
34.
Europaparlamentet har beslutat att frigöra följande från reserven:
-
-
Underhåll av fastigheter: 3 AST3, av vilka en förblir i reserven.
-
Besökscentrumet: 1 AD5 och 1 AST3.
-
Övriga: 1 AST3 (audiovisuella sektorn) och 1 AST3 (läkarmottagningen)
-
De 47 återstående tjänsterna i reserven utgår.
35.
36.
37.
Europaparlamentet har också beslutat att bekräfta följande uppgraderingar som begärts av de politiska grupperna: 8 AD12 till AD13, 9 AD11 till AD12, 6 AD10 till AD11, 1 AD9 till AD10, 4 AD6 till AD7, 9 AD5 till AD6, 10 AST10 till AST11, 1 AST9 till AST10, 5 AST8 till AST9, 5 AST7 till AST8, 14 AST6 till AST7, 14 AST5 till AST6, 1 AST4 till AST5, 9 AST3 till AST4, 7 AST2 till AST3, 2 AST1 till AST2.
38.
Europaparlamentet har beslutat att bekräfta följande omvandlingar och att frigöra motsvarande anslag:
-
4 AST3 till AD5.
-
2 AST och 2 AD5 tidsbegränsade tillfälliga tjänster till tillfälliga tjänster utan tidsbegränsning.
39.
40.
Europaparlamentet påpekar att anslagen för den ändrade tjänsteförteckningen därför har minskat från 2 760 616 EUR till 1 608 096 EUR, vilket motsvarar besparingar som uppgår till 1 152 520 EUR.
41.
Europaparlamentet välkomnar att de utbildnings och introduktionskurser, bland annat i samband med arbetsrotation (rörlighet) och omfördelning av personal, som Europeiska förvaltningsskolan givit personalen, har utvecklats på ett framgångsrikt sätt under de senaste åren.
42.
43.
Europaparlamentet välkomnar det faktum att praktikprogram för personer med funktionshinder, såsom omnämndes i riktlinjerna för 2007, har utformats och utvecklas relativt väl.
Fastighetspolitiken
44.
45.
Europaparlamentet uppmanar administrationen, i synnerhet efter "Strasbourg-erfarenheterna", att tillämpa mer stringenta, vattentäta och tydliga förfaranden när man förvärvar fastigheter.
46.
47.
48.
Europaparlamentet gör det mycket klart att det till fullo kommer att ge sitt stöd till att outnyttjade medel inom 20 procent av rubrik 5 – genom ändringsbudgetar – används i den händelse att parlamentet behöver extra kapitalutlägg för oförutsedda utgifter, särskilt i samband med köp och förvärv av väsentliga nya byggnader.
49.
om att en rapport skall utarbetas om huruvida det skulle vara möjligt att inrätta ett fastighetsorgan för EU med ansvar för byggnad och underhåll av EU-institutionernas och EU-organens fastigheter och begär att denna rapport skall läggas fram inför budgetutskottet.
50.
Europaparlamentet noterar presidiets begäran om tilldelning av ett specifikt belopp för att köpa följande fastigheter och har beslutat att godkänna följande:
-
Ytterligare 4 000 000 EUR för utbyggnaden av KAD-byggnaden i Luxemburg.
-
7 832 000 EUR för inredning och iordningställande av D4-byggnaden till följd av en tidig överlåtelse.
-
350 000 EUR för ombyggnader i plenisalen i Bryssel till följd av anslutningen av Rumänien och Bulgarien.
51.
Säkerhet
52.
Preliminärt anslag
Flerspråkigheten
53.
54.
55.
Europaparlamentet har, när det gäller iriskan, beslutat att följande anslag skall godkännas:
-
100 000 EUR under budgetpost 1 4 2 0 "Externa tjänster".
-
150 000 EUR under budgetpost 3 2 4 0 "Europeiska unionens officiella tidning".
-
112 000 EUR under budgetpost 2 1 0 0 "Inköp, installation, service och underhåll av utrustning och programvara"
-
50 000 EUR under budgetpost 3 2 2 2 "Utgifter för arkivsamlingar".
Stöd och tjänster till ledamöterna
56.
57.
Europaparlamentet anser fortfarande att en bättre användning kan ske både av parlamentets resurser och av intern specialiserad personal, i synnerhet då viktigare parlamentsbetänkanden skall utarbetas.
58.
59.
60.
61.
Europaparlamentet uppmanar generalsekreteraren att göra regelbundet återkommande granskningar av de tjänster som tillhandahålls ledamöterna, särskilt när det gäller datorer, resebyrån, telefoner, biltjänster och rättstjänsten.
62.
Parlamentet beslutar att till reserven föra 2 000 000 EUR från budgetpunkt 2 1 0 2 ("
Övrigt
63.
64.
65.
Avsnitt IV — Domstolen
66.
Andra extra utgifter (översättning/tolkning)
"), som vanligtvis täcker extra behov inom korrekturläsningen.
67.
68.
Europaparlamentet har fattat beslut om följande tjänsteförteckningsåtgärder:
-
-
Inrättande av 115 fasta tjänster för Rumänien och Bulgarien.
69.
70.
Avsnitt V — Revisionsrätten
71.
Europaparlamentet har beslutat att inrätta två tjänster för personalenheten för att underlätta moderniseringen av personalförvaltningen och förpliktar sig att inrätta ytterligare två tjänster som kommer att behövas under budgetåret 2008.
72.
Europaparlamentet har beslutat om att inrätta en tjänst inom vidareutbildningsenheten för att tillhandahålla adekvata utbildningsprogram för unga revisorer.
73.
Europaparlamentet har därför fattat beslut om följande tjänsteförteckningsåtgärder:
-
Inrättandet av 3 nya fasta tjänster (1 AST3 och 2 AST1) vid sidan av de 3 nya tjänster som rådet redan godkänt i sitt budgetförslag.
-
Inrättande av 41 fasta tjänster för Rumänien och Bulgarien.
74.
75.
Europaparlamentet har ökat de anslag som rådet avsatt i budgetförslaget med 3 579 729 EUR vilket motsvarar en ökning med 3,12 procent, exklusive kostnaderna i samband med utvidgningen.
Europeiska ekonomiska och sociala kommittén och Regionkommittén
76.
77.
78.
Europaparlamentet konstaterar att Regionkommittén beställde två oberoende externa utvärderingar av den gemensamma tjänsten, från Joan Colom i Naval och Robert Reynders, och uppmanar Regionkommitténs generalsekreterare att vidarebefordra dessa rapporter till Europaparlamentets budgetutskott.
Avsnitt VI — Europeiska ekonomiska och sociala kommittén
79.
Europaparlamentet begär att Europeiska ekonomiska och sociala kommittén skall lägga fram en årlig rapport före den 1 september varje år om effekterna av det rådgivande arbete som denna institution utför för Europaparlamentet, rådet och kommissionen.
80.
Europaparlamentet har beslutat att godkänna en tidigareläggning av utgifter på 1 995 120 EUR från budgeten för 2006 för att täcka en del av kommitténs behov för 2007 och minska dess äskanden för 2007 i motsvarande grad.
81.
Europaparlamentet anser att om Europeiska ekonomiska och sociala kommittén skall kunna klara av sin ökande arbetsbörda, måste kommittén begränsa längden på sina yttranden och andra publikationer, såsom de andra institutionerna gjort.
82.
Europaparlamentet har fattat beslut om följande tjänsteförteckningsåtgärder:
-
Inrättande av 5 nya fasta tjänster (1 AD5 och 4 AST3) vid sidan av de 13 nya tjänster som rådet redan godkänt i sitt budgetförslag.
-
Inrättande av 6 fasta tjänster för Rumänien och Bulgarien.
83.
Europaparlamentet har ökat de anslag som rådet avsatt i budgetförslaget med 1 529 115 EUR vilket motsvarar en ökning med 1,12 procent, exklusive kostnaderna i samband med utvidgningen.
Avsnitt VII — Regionkommittén
84.
Europaparlamentet är överens med rådet om den begäran om uppgraderingar som är knuten till tjänsteföreskrifterna och också om en begäran att uppgradera en enhetschefstjänst vid Regionkommittén till en direktörstjänst för den gemensamma tjänsten, under förutsättning att detta inte kommer att leda till behov av ytterligare personal och att inget förslag om att splittra upp den gemensamma tjänsten kommer att läggas fram till följd av denna uppgradering innan en djupgående och noggrann analys och bedömning av den gemensamma tjänsten genomförts.
85.
Europaparlamentet noterar att ingen begäran om nya tjänster i samband med utvidgningen till Bulgarien och Rumänien har inlämnats.
86.
Europaparlamentet har fattat beslut om följande tjänsteförteckningsåtgärder:
-
Inrättande av 3 nya fasta tjänster (2 AD5 och 1 AST3) och en tillfällig tjänst (AD5) vid sidan av de 3 nya tjänster som rådet redan godkänt i sitt budgetförslag.
87.
Europaparlamentet har ökat de anslag som rådet avsatt i budgetförslaget med 581 684 EUR vilket motsvarar en ökning med 2,53 procent, exklusive kostnaderna i samband med utvidgningen.
Avsnitt VIII (A) — Ombudsmannen
88.
Europaparlamentet noterar att bara 10 uppgraderingar har begärts av ombudsmannen och att dessa uppgraderingar fått rådets godkännande.
89.
Europaparlamentet har beslutat att begränsa anslaget till seminariet för de nationella ombudsmännen, som äger rum vartannat år och för vars organisation ombudsmannen ansvarar i år, till 45 000 EUR.
90.
Europaparlamentet har ökat anslagen som rådet avsatt i budgetförslaget med 150 000 EUR i syfte att fylla på anslaget till översättning.
Avsnitt VIII (B) — Europeiska datatillsynsmannen
91.
92.
Europaparlamentet har fattat beslut om följande tjänsteförteckningsåtgärder:
-
Inrättande av 2 nya fasta tjänster (1 AD9 och 1 AST5) vid sidan av de 3 nya tjänster (1AD9, 1 AD8 och 1 AD7) som rådet redan godkänt i sitt budgetförslag.
93.
o o
94.
Europaparlamentet uppdrar åt talmannen att översända denna resolution, tillsammans med ändringarna i avsnitt I, II, IV, V, VI, VII, VIII (A) och VIII (B) i förslaget till allmän budget, till rådet, kommissionen samt övriga berörda institutioner och organ.
P6_TA(2006)0512
Rumäniens anslutning
A6-0421/2006
Europaparlamentets resolution om Rumäniens anslutning till Europeiska unionen ( 2006/2115(INI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av fördraget om Republiken Bulgariens och Rumäniens anslutning till Europeiska unionen som undertecknades den 25 april 2005 EUT L 157, 21.6.2005, s.
11.
,
–
,
–
med beaktande av ordförandeskapets slutsatser från Europeiska rådets möte i Bryssel den 15-16 juni 2006,
–
med beaktande av slutsatserna från rådsmötet (allmänna frågor och yttre förbindelser) om utvidgningen den 17 oktober 2006,
–
med beaktande av kommissionens uppföljningsrapport om Rumänien av den 26 september 2006 ( KOM(2006)0549 ) och tidigare uppföljningsrapporter,
–
med beaktande av skriftväxlingen mellan Europaparlamentets talman och kommissionens ordförande om parlamentets fulla medverkan i övervägandena om att eventuellt tillämpa en av skyddsklausulerna i anslutningsfördraget,
–
med beaktande av artikel 45 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för utrikesfrågor och yttrandena från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor och utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män ( A6-0421/2006 ), och av följande skäl:
A.
B.
Rumäniens integration i Europeiska unionen kommer att bidra till stabiliteten och välståndet i sydöstra Europa.
C.
Rumäniens införlivande i Europeiska unionen kommer att stärka den politiska och kulturella dimensionen av den europeiska integrationsprocessen.
D.
Den första etappen av den femte utvidgningen 2004 har haft positiva återverkningar för både gamla och nya medlemsstater, vilket tveklöst även kommer att vara fallet för den aktuella utvidgningen som avslutar den femte utvidgningsomgången.
E.
Sedan kommissionens rapport från maj 2006 kan man återigen konstatera betydande förbättringar, vilket fastställs i kommissionens senaste uppföljningsrapport av den 26 september 2006.
F.
1.
Europaparlamentet uppskattar den noggrannhet och stringens som präglat hela kommissionens uppföljning av reformerna i Rumänien.
2.
Europaparlamentet lyckönskar Rumänien, välkomnar dess anslutning den 1 januari 2007 och ser fram emot den förestående ankomsten av landets trettiofem ledamöter av Europaparlamentet, dess kommissionsledamot och EU-tjänstemän i EU:s institutioner, samt värdesätter de rumänska medlemmarnas utmärkta insatser i egenskap av observatörer i Europaparlamentet sedan september 2005.
3.
Europaparlamentet betonar att denna utvidgning av Europeiska unionen, i likhet med tidigare utvidgningar, förverkligar den europeiska enhets- och solidaritetstanken som är till gagn för samtliga parter och främjar värden som demokrati, jämlikhet, mångfald och icke-diskriminering.
4.
Europaparlamentet välkomnar att kommissionen i sin rapport av den 26 september 2006 förordat att Bulgarien och Rumänien skall anslutas samtidigt.
5.
Europaparlamentet välkomnar de avsevärda framsteg som landet gjort sedan den senaste rapporten från maj 2006 och godkänner således den 1 januari 2007 som anslutningsdatum för Rumänien, men erinrar de rumänska myndigheterna om nödvändigheten av att fortsätta reformarbetet i samma takt efter anslutningen.
6.
Europaparlamentet välkomnar de ansträngningar som Rumänien gjort för att genomföra ett stort antal reformer inför anslutningen och uttalar sin uppskattning till de rumänska myndigheterna för de stora framsteg som gjorts på kort tid.
7.
Europaparlamentet betonar att reformprocessen är till stor fördel för Rumänien i samband med anslutningen till EU och även bidrar till den ekonomiska tillväxten och säkerheten i landet.
8.
Europaparlamentet konstaterar att det gjorts stora framsteg på de områden som kommissionen, i sin rapport från maj 2006, bedömt vara i behov av omedelbara åtgärder, nämligen: reform av rättsväsendet, korruptionsbekämpning, inrättande av utbetalningsorgan samt integrerat system för administration och kontroll, TSE, och sammankoppling av skatteuppbördssystemen.
9.
Europaparlamentet konstaterar med tillfredsställelse att Rumänien har en fungerande marknadsekonomi med en BNP-tillväxt på nära 7 procent och en arbetslöshet på cirka 5,5 procent.
10.
Europaparlamentet uppmuntrar medlemsstaterna att öppna sina arbetsmarknader för rumänsk arbetskraft från den 1 januari 2007 i enlighet med principen om arbetskraftens fria rörlighet, som garateras i gemenskapslagstiftningen.
11.
Europaparlamentet betonar nödvändigheten av att, med hänvisning till de finansiella transaktionerna från EU och Rumäniens nödvändiga medfinansiering i samband med de förväntade budgetomfördelningarna, detta inte enbart får ske på bekostnad av de sociala utgifterna och leda till nedskärningar av de sociala utgifterna.
12.
13.
14.
Om den romska minoriteten: Europaparlamentet uppmanar med kraft de rumänska myndigheterna att konsolidera de påbörjade reformerna för skydd mot institutionaliserat våld, förbättring av levnadsstandard och boende och tillgång till sysselsättning och hälso- och sjukvårdssystem, genom att tillräckliga medel ställs till förfogande.
15.
Om den ungerska minoriteten: Europaparlamentet uppmanar de rumänska myndigheterna att beakta den ungerska minoritetens förväntningar, i enlighet med subsidiaritetsprincipen och principen om kulturellt självstyre, särskilt genom att tillräckliga medel ställs till förfogande för förbättring av utbildningsstandarden.
16.
Europaparlamentet föreslår att utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor från den 1 januari 2007 gör en uppföljning av reformerna i fråga om adoption och skydd för barn i Rumänien.
17.
18.
19.
15.
20.
Europaparlamentet konstaterar att kommissionen fastställt tre områden där väsentliga framsteg gjorts sedan rapporten från maj 2006, men som fortfarande kräver ytterligare åtgärder:
–
reformen av rättsväsendet och kampen mot korruption,
–
utnyttjandegraden och hanteringen av gemenskapsstödet inom jordbrukssektorn och strukturfonderna,
–
21.
Europaparlamentet understryker att av dessa tre områden är det slutliga genomförandet av reformen av rättsväsendet och kampen mot korruption av avgörande betydelse och måste därför bli föremål för särskilda insatser från de rumänska myndigheternas sida.
22.
Europaparlamentet stöder att kommissionen inrättar kontroll- och uppföljningsmekanismer för dessa områden som särskilt baserar sig på fastställandet av vissa bestämda kriterier, och uppmanar mycket kraftfullt den rumänska regeringen att vidta alla erforderliga åtgärder för att uppfylla de uppställda förväntningarna och därmed undvika att skyddsklausuler tillämpas.
23.
24.
25.
Europaparlamentet kräver att kommissionen systematiskt håller parlamentet underrättat om de framsteg som Rumänien gör under de kommande månaderna och att parlamentet involveras på nära håll i den övervakningsmekanism som kommissionen föreslår för tiden efter anslutningen.
26.
Europaparlamentet betonar att Rumäniens regering bör vara medveten om att den återstående tiden måste utnyttjas till fullo för fortsatta insatser för att konsolidera de uppnådda resultaten.
27.
Europaparlamentet kräver att anslutningsfördraget snarast ratificeras av de två medlemsstater som ännu inte gjort detta.
28.
Europaparlamentet uppmanar kommissionen att avsätta lämpliga medel för informationskampanjer för att förbättra allmänhetens medvetenhet i samband med Rumäniens (och Bulgariens) anslutning.
29.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen och regeringarna och parlamenten i medlemsstaterna och Rumänien.
P6_TA(2006)0569
De institutionella aspekterna av Europeiska unionens kapacitet att integrera nya medlemsstater
A6-0393/2006
Europaparlamentets resolution om institutionella aspekter på Europeiska unionens förmåga att integrera nya medlemsstater ( 2006/2226(INI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av artikel 49 i EG-fördraget,
–
med beaktande av ordförandeskapets slutsatser från Europeiska rådets möte i Köpenhamn i juni 1993, i Madrid i december 1995, i Luxemburg i december 1997, i Thessaloniki i juni 2003, och i Bryssel i december 2004, i juni 2005 och juni 2006,
–
med beaktande av Europeiska unionens stadga om de grundläggande rättigheterna,
–
med beaktande av 2005 års strategidokument för utvidgningen från kommissionen ( KOM(2005)0561 ),
–
med beaktande av sin resolution av den 12 januari 2005 om fördraget om upprättande av en konstitution för Europa EUT C 247 E, 6.10.2005, s.
88.
,
–
med beaktande av sin resolution av den 28 september 2005 om inledandet av förhandlingar med Turkiet EUT C 227 E, 21.9.2006, s.
163.
,
–
med beaktande av förhandlingsramarna för Turkiet och Kroatien som rådet antog den 3 oktober 2005,
–
med beaktande av sin resolution av den 19 januari 2006 om perioden av eftertanke: struktur, teman och ramar för en utvärdering av debatten om Europeiska unionen EUT C 287 E, 24.11.2006, s.
306.
,
–
,
–
,
–
,
–
med beaktande av artikel 45 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för konstitutionella frågor ( A6-0393/2006 ), och av följande skäl:
A.
Vid sitt möte i Thessaloniki den 19-20 juni 2003 gav Europeiska rådet tydligt uttryck för ett europeiskt perspektiv för länderna på västra Balkan, med EU-medlemskap för dessa länder som slutmål (Tessalonikiagendan).
B.
Europeiska rådet bekräftade vid sitt möte den 16-17 juni 2005 sitt åtagande att fullt ut genomföra Thessalonikiagendan, och bekräftade vid sitt möte den 15-16 juni 2006 sin avsikt att respektera de åtaganden som gjorts gentemot länderna i sydöstra Europa (Turkiet och Kroatien såsom länder med vilka förhandlingar har inletts, f.d. jugoslaviska republiken Makedonien/FYROM såsom kandidatland samt övriga länder i västra Balkan såsom möjliga kandidatländer) i fråga om utvidgningen samtidigt som det underströk behovet att se till att unionen fungerar politiskt, ekonomiskt och institutionellt medan utvidgningen pågår.
C.
Den 3 oktober 2005 inledde rådet formellt anslutningsförhandlingar med Turkiet och Kroatien.
D.
Vid sitt möte den 15-16 december 2005 gav rådet f.d. jugoslaviska republiken Makedonien (FYROM) status som kandidatland.
E.
Iakttagandet av samtliga Köpenhamnskriterier har varit utgångspunkten för medlemskap i EU sedan 1993 och bör även vara det vid framtida utvidgningar.
F.
I Köpenhamnskriterierna betonas även betydelsen av unionens förmåga att ta emot nya medlemmar utan att den europeiska integrationen förlorar i kraft.
G.
EU:s institutionella förmåga att integrera nya medlemsstater har i stigande grad blivit föremål för diskussion i samband med utvidgningar efter Bulgariens och Rumäniens tillträde.
H.
I sin ovannämnda resolution om kommissionens strategidokument inför utvidgningen (2005) inbjöd parlamentet kommissionen att senast vid utgången av 2006 lägga fram en rapport i vilken den redogör för de principer som EU:s absorptionsförmåga baseras på.
I.
J.
Enligt Europeiska rådet bör denna rapport även innehålla en redogörelse för medborgarnas uppfattning om utvidgningen nu och i framtiden samt beakta nödvändigheten att förklara utvidgningsprocessen på ett lämpligt sätt till allmänheten inom EU.
K.
Enligt ordförandeskapets slutsatser från Europeiska rådet möte i Bryssel den 16-17 december 2004 "kan anslutningsförhandlingar som ännu inte har inletts med kandidatstater vilkas anslutning kan få betydande finansiella konsekvenser inte slutföras förrän finansieringsramen från och med 2014 har fastställts, tillsammans med eventuella finansiella följdreformer".
L.
M.
Det pågår en diskussion om EU:s så kallade "absorptionsförmåga" när det gäller framtida utvidgningar.
N.
Kommissionens ordförande har inför parlamentet förklarat att han anser att de institutionella frågorna bör lösas innan någon ytterligare utvidgning tar vid, och har uttryckt sin förhoppning om att denna lösning, såsom den fastställdes vid Europeiska rådets möte den 15-16 juni 2006, kan uppnås före utgången av 2008 och därmed tillåta EU att respektera sina åtaganden gentemot de länder som inlett förhandlingar liksom de för vilka det förespeglat möjligheten till anslutning.
O.
En institutionell lösning av detta slag behövs framför allt för att bibehålla takten i den europeiska integrationen, såsom medlemsstaternas stats- och regeringschefer noterade vid Europeiska rådets möte i Köpenhamn 1993.
1.
Europaparlamentet påpekar att utvidgningen har tenderat att stärka unionen, främja dess ekonomiska tillväxt, stärka dess roll i internationellt hänseende och påskynda utvecklingen av EU:s politik inom nya områden.
2.
Europaparlamentet erinrar om att begreppet "absorptionsförmåga" användes för första gången 1993 då Europeiska rådet vid sitt möte i Köpenhamn erkände att vid sidan om de politiska och ekonomiska kriterier som kandidatländerna måste uppfylla för att kunna tillträda unionen utgör även "unionens förmåga att ta emot nya medlemmar, utan att takten i den europeiska integrationen blir lidande en viktig faktor som ligger i både EU:s och kandidatländernas allmänna intresse".
3.
Europaparlamentet erinrar om att även om varje utvidgning av unionen har medfört ändringar av dess institutionella, politiska och ekonomiska ramar har dessa ändringar inte varit tillräckliga för att säkra effektiviteten i unionens beslutsfattande.
4.
Europaparlamentet anser att termen "absorptionsförmåga" är missvisande eftersom EU på intet sätt "absorberar" sina medlemmar, och föreslår därför att den ersätts med termen "integrationsförmåga" som på ett bättre sätt ger uttryck för innebörden av EU-medlemskap.
5.
6.
Europaparlamentet anser att "integrationskapacitet" efter utvidgningen innebär att
–
EU:s institutioner kan fungera som de skall och fatta beslut på ett effektivt och demokratiskt sätt och i enlighet med de specifika förfaranden de har att följa,
–
EU:s ekonomiska resurser räcker till för att finansiera dess verksamhet,
–
unionen kan fortsätta att utveckla sin politik på ett framgångsrikt sätt och att uppnå sina målsättningar och därmed förverkliga sitt politiska syfte.
7.
8.
Europaparlamentet erkänner att EU idag står inför svårigheter att uppfylla sina åtaganden gentemot länderna i sydöstra Europa på grund av att dess institutionella, ekonomiska och politiska struktur är otillräcklig för ytterligare utvidgningar och måste förbättras.
Integrationskapacitetens institutionella aspekter
9.
a)
Ett nytt system för kvalificerad majoritetsröstning bör antas som ger rådet bättre möjlighet att fatta beslut.
b)
En rejäl utökning bör ske av de politikområden som är föremål för kvalificerad majoritetsomröstning.
c)
Europaparlamentet bör ges betydligt större möjlighet att delta i budget- och lagstiftningsarbetet på lika villkor med rådet.
d)
Rotationssystemet för Europeiska rådets ordförandeskap bör ändras.
e)
En befattning som utrikesminister bör inrättas.
f)
Kommissionens sammansättning bör ändras utöver vad som föreskrivs i Nicefördraget.
g)
Kommissionens ordförandes roll och demokratiska legitimitet bör stärkas genom att han/hon väljs av Europaparlamentet.
h)
EG-domstolens domsrätt bör utvidgas till att omfatta unionens samtliga verksamhetsområden, inklusive övervakningen av respekten för de grundläggande rättigheterna.
i)
Mekanismer bör skapas för att involvera medlemsstaternas parlament i granskningen av EU:s åtgärder.
j)
Mer flexibla arrangemang bör införas som svar på den växande möjligheten att inte alla medlemsstater kan eller vill föra politiken på vissa områden vidare på samma gång.
k)
Förfarandet för att göra ändringar i fördragen bör ändras i syfte att göra det enklare och mer effektivt och för att stärka det demokratiska tillvägagångssättet liksom insynen och öppenheten.
l)
"Pelarstrukturen" bör avskaffas och ersättas med ett verksamhetsfält med enhetlig struktur och rättslig status.
m)
En klausul bör införas som ger medlemsstaterna möjlighet att lämna EU.
n)
De värderingar som ligger till grund för EU, liksom dess målsättningar, bör definieras klart och tydligt.
o)
EU:s befogenheter och de principer som ligger till grund för såväl unionens åtgärder som dess förbindelser med medlemsstaterna bör definieras klart och tydligt.
p)
Insynen i EU:s förfaranden för beslutfattande bör stärkas, i första hand genom offentlig granskning av rådets verksamhet i egenskap av lagstiftande myndighet.
q)
De instrument med vilka EU utövar sina befogenheter bör definieras klart och tydligt och därtill förenklas.
Parlamentet påpekar att alla dessa reformer redan ingår i konstitutionsfördraget och att om de genomförs skulle det göra det möjligt för ett utvidgat EU att fungera som det skall och fatta beslut på ett effektivt och demokratiskt sätt.
Andra relevanta aspekter av integrationskapaciteten
10.
a)
Europeiska unionens stadga om de grundläggande rättigheterna om de grundläggande rättigheterna bör antas och solidaritetspolitiken bör stärkas mellan medlemsstaterna.
b)
373.
samt med bestämmelserna enligt det interinstitutionella avtalet av den 17 maj 2006 om budgetdisciplin och sund ekonomisk förvaltning EUT C 139, 14.6.2006, s.
1.
.
c)
Ett flertal av unionens politikområden, varav somliga fastställdes för över 50 år sedan, bör omdefinieras så att unionen får möjlighet att genomföra Lissabonstrategin, stärka sin handlingsförmåga i internationella sammanhang och anpassa sig efter de nya utmaningar som en mycket större och mer heterogen union står inför i en globaliserad värld.
d)
Europeiska grannskapspolitiken bör stärkas i syfte att skapa ett lämpligt instrument för att upprätta ömsesidigt fördelaktiga förbindelser med de europeiska länder som inte har omedelbara utsikter till EU-medlemskap på grund av att de inte uppfyller villkoren för medlemskap eller väljer att inte ansluta sig.
11.
12.
Europaparlamentet upprepar dock att varje beslut av EU om att godkänna en ny medlemsstat fattas genom ett förfarande som säkerställer en rad garantier, det vill säga enhälligt beslut av samtliga medlemsstater att inleda och avsluta anslutningsförhandlingar, Europaparlamentets godkännande och ratificering av varje anslutningsavtal av samtliga medlemsstater.
13.
Europaparlamentet betonar under alla omständigheter att det faktum att medlemsstaternas regeringar undertecknar ett anslutningsfördrag innebär att dessa regeringar fullt ut åtar sig att agera i enlighet med det aktuella fördraget för att se till att man på ett framgångsrikt sätt lyckas genomföra ratificeringsprocessen enligt de förfaranden som tillämpas i respektive land.
14.
Europaparlamentet anser att Europaparlamentets samtycke, som krävs för att rådet skall kunna agera enligt artikel 49 i fördraget om Europeiska unionen i frågan om anslutningen av nya medlemsstater, bör gälla såväl beslutet att inleda förhandlingar som förhandlingarnas slutförande.
Slutsatser
15.
16.
Europaparlamentet understryker att EU måste kunna anpassa sin institutionella, ekonomiska och politiska struktur i god tid för att undvika att anslutningen av kandidatländer försenas efter det att det har slagits fast att de uppfyllt samtliga kriterier för medlemskap.
17.
Europaparlamentet bekräftar åter att Nicefördraget inte utgör tillräcklig grund för ytterligare utvidgningar.
18.
Europaparlamentet bekräftar åter sitt stöd för konstitutionsfördraget, som redan erbjuder lösningar på flertalet av de reformer som EU måste genomföra för att kunna uppfylla sina åtaganden vad gäller den nu aktuella utvidgningen och som utgör ett konkret uttryck för sambandet mellan fördjupning och utvidgning, och varnar för att varje försök att bit för bit genomföra delar av det åtgärdspaket som konstitutionsfördraget avser riskerar att undergräva den kompromiss om helheten som fördraget vilar på.
19.
Europaparlamentet noterar den tidsplan som Europeiska rådet fastslog vid sitt möte den 15-16 juni 2006 för att senast under hösten 2008 finna en lösning på den konstitutionella krisen.
20.
Europaparlamentet bekräftar åter sitt åtagande att snarast möjligt finna en konstitutionell lösning för EU och under alla omständigheter innan Europas medborgare kallas att avge sin röst vid Europavalen 2009, för att unionen skall kunna uppfylla sina åtaganden gentemot kandidatländerna och vara redo att ta emot dem.
o
o o
21.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, parlamenten och regeringarna i medlemsstaterna, parlamenten och regeringarna i Turkiet, Kroatien, före detta jugoslaviska republiken Makedonien, Albanien, Bosnien och Hercegovina, Serbien, Montenegro, Kosovos provisoriska institutioner för självstyre samt FN:s interimadministration i Kosovo (UNMIK).
P6_TA(2006)0599
Kärnsäkerhetsstöd *
A6-0397/2006
Europaparlamentets lagstiftningsresolution om förslaget till rådets förordning om inrättande av ett instrument för kärnsäkerhetsstöd (9037/2006 – C6-0153/2006 – 2006/0802(CNS) )
(Samrådsförfarandet)
–
med beaktande av rådets text (9037/2006),
–
med beaktande av kommissionens förslag till rådet ( KOM(2004)0630 ) Ännu ej offentliggjort i EUT.
,
–
med beaktande av artiklarna 177 och 203 i fördraget om upprättandet av Europeiska atomenergigemenskapen, i enlighet med vilken rådet har hört parlamentet ( C6-0153/2006 ),
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för industrifrågor, forskning och energi och yttrandena från utskottet för utrikesfrågor, utskottet för miljö, folkhälsa och livsmedelssäkerhet och budgetutskottet ( A6-0397/2006 ).
1.
Europaparlamentet godkänner rådets text såsom ändrad av parlamentet.
2.
Europaparlamentet anser att det vägledande referensbelopp som anges i lagstiftningstexten måste stämma överens med taket i utgiftskategori 4 i den nya fleråriga budgetramen och påpekar att beslut om det årliga beloppet kommer att fattas inom ramen för det årliga budgetförfarandet i enlighet med bestämmelserna i punkt 38 i det interinstitutionella avtalet mellan Europaparlamentet, rådet och kommissionen av den 17 maj 2006 om budgetdisciplin och sund ekonomisk förvaltning EUT C 139, 14.6.2006, s.
1.
.
3.
4.
Rådet uppmanas att underrätta Europaparlamentet om rådet har för avsikt att avvika från den text som parlamentet har godkänt.
5.
Rådet uppmanas att på nytt höra Europaparlamentet om rådet har för avsikt att väsentligt ändra den text som är föremål för samråd.
6.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
Rådets förslag Parlamentets ändringar Ändring 1 Skäl 1 (1)
Europeiska gemenskapen är en av de främsta givarna av ekonomiskt, finansiellt, tekniskt, humanitärt och makroekonomiskt bistånd till tredjeländer.
I syfte att effektivisera Europeiska gemenskapens bistånd till tredjeländer har det utarbetats en ny ram med bestämmelser om hur stödinsatser skall planeras och tillhandahållas.
Genom rådets förordning (EG) nr … av den … upprättas ett föraranslutningsinstrument, vilket skall täcka gemenskapens stöd till kandidatländer och potentiella kandidatländer.
Genom Europaparlamentets och rådets förordning (EG) nr … av den … upprättas ett europeiskt grannskaps- och partnerskapsinstrument.
Europaparlamentets och rådets förordning (EG) nr … av den … är inriktad på utvecklingssamarbete
och
ekonomiskt samarbete med övriga tredjeländer.
Genom Europaparlamentets och rådets förordning (EG) nr ... av den ... inrättas ett stabilitetsinstrument.
Europeiska gemenskapen är en av de främsta givarna av ekonomiskt, finansiellt, tekniskt, humanitärt och makroekonomiskt bistånd till tredjeländer.
I syfte att effektivisera Europeiska gemenskapens bistånd till tredjeländer har det utarbetats en ny ram med bestämmelser om hur stödinsatser skall planeras och tillhandahållas.
Genom rådets förordning (EG) nr … av den … upprättas ett föraranslutningsinstrument, vilket skall täcka gemenskapens stöd till kandidatländer och potentiella kandidatländer.
Genom Europaparlamentets och rådets förordning (EG) nr … av den … upprättas ett europeiskt grannskaps- och partnerskapsinstrument.
Europaparlamentets och rådets förordning (EG) nr … av den … är inriktad på utvecklingssamarbete
med tredjeländer
1
.
Genom rådets förordning (EG) nr … av den … främjas
ekonomiskt samarbete med övriga tredjeländer.
Genom Europaparlamentets och rådets förordning (EG) nr ... av den ... inrättas ett stabilitetsinstrument.
Genom Europaparlamentets och rådets förordning (EG) nr … av den … inrättas ett finansieringsinstrument för främjande av demokrati och mänskliga rättigheter i hela världen (Europeiska instrumentet för demokrati och mänskliga rättigheter)
2
_______________
1
EUT L …, …, s. … .
2
EUT L …, …, s. … .
Ändring 3 Skäl 2a (nytt)
(2a) Kärnmaterial blir allt tillgängligare, vilket ökar risken för spridning av kärnvapen och därför får tydliga följder för kärnsäkerheten, något som bör tas upp i detta instrument.
Ändring 4 Skäl 3a (nytt)
(3a) Det är mycket viktigt att sekretessen för uppgifter om kärn- och strålsäkerhet, som måste vara exakta och bekräftade, garanteras, särskilt uppgifter som kan vara av stort intresse för terrorister.
Ändring 5 Skäl 4 (4)
I enlighet med
kapitel X
i fördraget bedriver gemenskapen ett nära samarbete med Internationella atomenergiorganet (IAEA), både vad avser kärnämneskontroller (för främjande av syftena i fördragets
del två kapitel VII
) och vad avser kärnsäkerhet.
(4)
I enlighet med
avdelning II kapitel 10
i fördraget bedriver gemenskapen ett nära samarbete med Internationella atomenergiorganet (IAEA), både vad avser kärnämneskontroller (för främjande av syftena i fördragets
avdelning II kapitel 7
) och vad avser kärnsäkerhet.
Gemenskapen stöder därför aktivt ett utarbetande av en uppförandekod för ett internationellt övervakningssystem avseende kärnkraftsolyckor under IAEA:s överinseende.
Ändring 6 Skäl 7 (7)
Utöver internationella konventioner och fördrag har några medlemsstater ingått bilaterala överenskommelser om tillhandahållande av tekniskt stöd.
(7)
Utöver internationella konventioner och fördrag har några medlemsstater ingått bilaterala överenskommelser om tillhandahållande av tekniskt stöd.
En samordning mellan åtgärder som vidtas med stöd av sådana överenskommelser och gemenskapsåtgärderna är önskvärd.
Ändring 7 Skäl 9 (9)
skall ha
maximal effekt, dock utan att ge avkall på principen att ansvaret för anläggningens säkerhet bör vila på den driftsansvarige och den stat som har behörighet över anläggningen.
(9)
Det är underförstått att när stöd lämnas till den berörda kärnenergianläggningen är det i syfte att det
skulle kunna få
maximal effekt, dock utan att ge avkall på principen att
"förorenaren betalar" och att
ansvaret för anläggningens säkerhet
, avvecklingen av den och för det avfall den genererat
bör vila på den driftsansvarige och den stat som har behörighet över anläggningen.
Dessutom bör företräde ges åt stöd till sådana kärnenergianläggningar och sådan verksamhet på kärnenergins område som sannolikt kan få betydande konsekvenser för medlemsstaterna.
Ändring 8 Skäl 13 (13)
Denna förordning som föreskriver ekonomiskt bistånd till stöd för syftena i fördraget påverkar inte gemenskapens och medlemsstaternas respektive behörighet på de berörda områdena, särskilt vad avser kärnämneskontroller.
(13)
Denna förordning som föreskriver ekonomiskt bistånd till stöd för syftena i fördraget påverkar inte
medlemsstaternas exklusiva behörighet att själva välja energiformer och
gemenskapens och medlemsstaternas respektive behörighet på de berörda områdena, särskilt vad avser kärnämneskontroller.
Ändring 9 Skäl 13a (nytt)
(13a) Ett ekonomiskt referensbelopp av det slag som avses i artikel 38 i det interinstitutionella avtalet av den 17 maj 2006 om budgetdisciplin och sund ekonomisk förvaltning
1
EUT C 139, 14.6.2006, s.
1.
hög
kärnsäkerhetsnivå, strålskydd och tillämpning av effektiva och verkningsfulla säkerhetskontroller av kärnmaterial i tredjeländer.
Gemenskapen
finansiera åtgärder som främjar
, strålskydd och tillämpning av effektiva och verkningsfulla säkerhetskontroller av kärnmaterial i tredjeländer.
Främjande av
på alla nivåer, särskilt genom
effektiva kärnsäkerhetsåtgärder
på alla nivåer, särskilt genom
Ändring 13 Artikel 2, led a, strecksats 3
utformning,
drift och underhåll av befintliga
kärnkraftsverk
eller andra befintliga kärnenergianläggningar så att
höga
säkerhetsnivåer kan uppnås,
– bättre säkerhetsaspekter vid drift
, modernisering
som är i drift, med hänsyn tagen till de erfarenheter som vunnits vid driften av dem,
så att
högsta möjliga
– stöd till säker transport, behandling och bortskaffande av kärnbränsle och radioaktivt avfall,
– stöd till
utveckling av korrekta metoder och korrekt teknik för
säker transport, behandling och bortskaffande av
använt
kärnbränsle och radioaktivt avfall
och
– utveckling och genomförande av strategier för avveckling av befintliga anläggningar och sanering av f.d. kärnenergianläggningar
, för att uppnå en hög säkerhetsnivå till ett rimligt pris under en överskådlig tid
.
Ändring 16 Artikel 2, led b (b)
Främjande av effektiva regelverk, förfaranden och system för att säkerställa ett tillräckligt skydd mot joniserande strålning från radioaktivt material, särskilt från radioaktiva strålkällor med hög aktivitet, och bortskaffande
Ändring 17 Artikel 2, led d d)
d)
Upprättande av effektiva arrangemang för
katastrofberedskap, beredskaps- och insatsplanering, räddningstjänst
, skadebegränsning
och saneringsåtgärder.
Ändring 18 Artikel 2, led e e)
och
Åtgärder för att främja internationellt samarbete (bland annat inom berörda internationella organisationer, särskilt IAEA) på ovannämnda områden, bl.a. genom genomförande och övervakning av internationella konventioner och fördrag, informationsutbyte,
utbildning
forskning.
Mål, åtgärdsområden, planerade åtgärder, förväntade resultat, förvaltningsformer samt beräknat totalt finansieringsbelopp skall anges i dessa handlingsprogram.
Vid behov kan
de innehålla resultaten av erfarenheter från tidigare stöd.
2.
Mål, åtgärdsområden, planerade åtgärder, förväntade resultat, förvaltningsformer samt beräknat totalt finansieringsbelopp skall anges i dessa handlingsprogram.
De skall också innehålla en kortfattad beskrivning av de insatser som skall finansieras samt uppgifter om finansieringsbelopp för dem och en vägledande tidsplan för deras genomförande.
de innehålla resultaten av erfarenheter från tidigare stöd.
3.
och med hänsyn tagen till artikel 18
, i förekommande fall efter samråd med det eller de partnerländer i regionen som berörs.
Europeiska unionens organ.
–
Gemenskapens gemensamma forskningscenter och
Europeiska unionens organ.
Skuldlättnadsprogram.
, som skall komma i fråga i undantagsfall och genomföras i enlighet med ett internationellt överenskommet skuldlättnadsprogram
.
2a.
Gemenskapsfinansieringen skall i princip inte användas för betalning av skatter, tullavgifter eller andra avgifter av skatterättslig natur i mottagarländerna.
Ändring 24 Artikel 18
I syfte att kontrollera om målen har nåtts och för att utarbeta rekommendationer om hur verksamheten kan förbättras i framtiden skall kommissionen regelbundet utvärdera resultaten av strategier och program samt effektiviteten i programplaneringen.
Kommissionen skall för kännedom överlämna mer betydelsefulla utvärderingsrapporter till den kommitté som inrättas i enlighet med artikel 20.
I syfte att kontrollera om målen har nåtts och för att utarbeta rekommendationer om hur verksamheten kan förbättras i framtiden skall kommissionen
med biträde av oberoende sakkunniga
regelbundet
, utgående från de enskilda projekten tagna vart för sig,
utvärdera resultaten av strategier och program samt effektiviteten i programplaneringen.
Kommissionen skall för kännedom överlämna mer betydelsefulla utvärderingsrapporter till
Europaparlamentet, rådet och
den kommitté som inrättas i enlighet med artikel 20.
Ändring 25 Artikel 20a (ny)
Artikel 20a
Ekonomiskt referensbelopp
Det ekonomiska referensbeloppet för genomförandet av denna förordning under perioden 2007–2013 skall uppgå till 524 miljoner EUR.
De årliga anslagen skall godkännas av den budgetansvariga myndigheten, inom de gränser som uppställs av budgetramen.
Ändring 26 Artikel 21
Kommissionen skall senast den 31 december 2010 till Europaparlamentet och rådet lägga fram en rapport med en utvärdering av genomförandet av förordningen under de första tre åren, vid behov tillsammans med ett lagstiftningsförslag om införande av nödvändiga ändringar i instrumentet.
Kommissionen skall senast den 31 december 2010 till Europaparlamentet och rådet lägga fram en rapport med en utvärdering av genomförandet av förordningen under de första tre åren
och därefter rapportera vartannat år
, vid behov tillsammans med ett lagstiftningsförslag om införande av nödvändiga ändringar i instrumentet.
P6_TA(2007)0018
Moratorium för dödsstraff
B6-0032 , 0033 , 0034 , 0035 och 0036/2007
Europaparlamentets resolution angående initiativet till ett allmänt moratorium för dödsstraff
Europaparlamentet utfärdar denna resolution
-
med beaktande av sina tidigare resolutioner om ett allmänt moratorium för dödsstraff, särskilt resolutionerna av den 23 oktober 2003 EUT C 82 E, 1.4.2004, s.
609.
, 6 maj 1999 EGT C 279, 1.10.1999, s.
421.
och 18 juni 1998 EGT C 210, 6.7.1998, s.
207.
,
-
med beaktande av de resolutioner om ett moratorium för dödsstraff som antagits av flera FN-organ, bland annat FN:s kommission för mänskliga rättigheter,
-
med beaktande av EU:s uttalanden till stöd för ett allmänt moratorium för dödsstraffet, och det uttalande om avskaffande av dödsstraffet som gjordes den 19 december 2006 vid FN:s generalförsamling och som undertecknades av 85 länder från samtliga geografiska grupper,´
-
med beaktande av riktlinjerna för EU:s politik gentemot tredjeländer avseende dödsstraffet som antogs av rådet (allmänna frågor) den 29 juni 1998,
–
A.
Dödsstraff är en grym och omänsklig bestraffning och ett brott mot rätten till liv.
B.
Dödsstraffets avskaffande är en grundläggande värdering för Europeiska unionen och är ett krav för länder som söker medlemskap i EU.
C.
Det är mycket oroväckande att dussintals länder i världen än i dag har, eller har återinfört, lagar som föreskriver dödsstraff och att tusentals människor således avrättas varje år enligt dessa lagar.
D.
E.
EU beslutade i sina riktlinjer om EU:s politik gentemot tredje länder beträffande dödsstraff, som antagits av Europeiska rådet, att inom internationella organisationer verka för att dödsstraffet avskaffas.
F.
Den 9 januari 2007 beslutade den italienska regeringen och Europarådet att gemensamt försöka samla så mycket stöd som möjligt för ett initiativ i FN:s pågående generalförsamling för ett världsomspännande moratorium för avrättningar i syfte att helt avskaffa dödsstraffet.
G.
H.
Avrättningen av Saddam Hussein och mediernas exploatering av hängningen kan inte annat än fördömas, och det sätt på vilket den genomfördes är beklagansvärt.
1.
Europaparlamentet erinrar om sin orubbliga inställning till dödsstraff i alla lägen och under alla omständigheter, och uttrycker ännu en gång sin övertygelse att om dödsstraffet avskaffas kommer detta att bidra till att människovärdet stärks och de mänskliga rättigheterna fortsätter att utvecklas.
2.
3.
4.
Europaparlamentet uppmanar alla EU:s institutioner och medlemsstater att politiskt och diplomatiskt göra allt för att denna resolution skall få tillräckligt stöd i FN:s pågående generalförsamling.
5.
Europaparlamentet stöder aktivt den italienska deputeradekammarens och den italienska regeringens initiativ som även har Europeiska rådets, kommissionens och Europarådets stöd.
6.
Europaparlamentet uppmanar alla EU:s medlemsstater att utan dröjsmål ratificera det andra frivilliga protokollet till Internationella konventionen om medborgerliga och politiska rättigheter som syftar till att dödsstraffet skall avskaffas helt.
7.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, FN:s generalsekreterare, ordföranden i FN:s generalförsamling och alla FN:s medlemsstater.
P6_TA(2007)0068
Saluföring av kött från nötkretaur som är högst tolv månader *
A6-0006/2007
Europaparlamentets lagstiftningsresolution av den 14 mars 2007 om förslaget till rådets förordning om saluföring av nötkött från djur på högst tolv månader ( KOM(2006)0487 – C6-0330/2006 – 2006/0162(CNS) )
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till rådet ( KOM(2006)0487 ) Ännu ej offentliggjort i EUT.
,
–
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för jordbruk och landsbygdens utveckling ( A6-0006/2007 ).
1.
Europaparlamentet godkänner kommissionens förslag såsom ändrat av parlamentet.
2.
3.
Rådet uppmanas att underrätta Europaparlamentet om rådet har för avsikt att avvika från den text som parlamentet har godkänt.
4.
Rådet uppmanas att på nytt höra Europaparlamentet om rådet har för avsikt att väsentligt ändra kommissionens förslag.
5.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
Kommissionens förslag Parlamentets ändringar Ändring 1 Skäl 5 (5)
För att förbättra den inre marknadens funktion bör saluföringen av nötkött från djur på högst tolv månader organiseras på ett så genomsynligt sätt som möjligt.
Det blir därigenom också möjligt att organisera produktionen på ett bättre sätt.
Det måste definieras vilka handelsbeteckningar som skall användas i var och en av medlemsstaterna för saluföringen av nötkött från djur på högst tolv månader.
Kvaliteten på konsumentupplysningarna förbättras också genom detta.
(5)
För att förbättra den inre marknadens funktion bör saluföringen av nötkött från djur på högst tolv månader organiseras på ett så genomsynligt sätt som möjligt.
Det blir därigenom också möjligt att organisera produktionen på ett bättre sätt.
Det måste definieras vilka handelsbeteckningar som skall användas i var och en av medlemsstaterna för saluföringen av nötkött
eller beredningar därav avsedda för mänsklig konsumtion
från djur på högst tolv månader.
Kvaliteten på konsumentupplysningarna förbättras också genom detta.
Ändring 2 Skäl 12 (12)
Det bör också föreskrivas att nötkött från djur på högst tolv månader bör märkas med en bokstavsbeteckning som anger vilken underkategori köttet tillhör
,
samt att märkningen av köttet skall innehålla uppgift om slaktåldern.
(12)
Det bör också föreskrivas att nötkött från djur på högst tolv månader bör märkas med en bokstavsbeteckning som anger vilken underkategori köttet tillhör
Dessa uppgifter bör också anges i samtliga handelsdokument.
Ändring 3 Skäl 13 (13)
Aktörer som önskar komplettera de handelsbeteckningar som föreskrivs i denna förordning med frivilliga uppgifter bör kunna göra detta i enlighet med förfarandet i artikel 16 och 17 i Europaparlamentets och rådets förordning (EG) nr 1760/2000 av den 17 juli 2000 om upprättande av ett system för identifiering och registrering av nötkreatur samt märkning av nötkött och nötköttsprodukter och om upphävande av rådets förordning (EG) nr 820/97.
(13)
Aktörer som önskar komplettera de handelsbeteckningar som föreskrivs i denna förordning med frivilliga uppgifter
, såsom typ av foder,
bör kunna göra detta i enlighet med förfarandet i artikel 16 och 17 i Europaparlamentets och rådets förordning (EG) nr 1760/2000 av den 17 juli 2000 om upprättande av ett system för identifiering och registrering av nötkreatur samt märkning av nötkött och nötköttsprodukter och om upphävande av rådets förordning (EG) nr 820/97.
Ändring 4 Skäl 14 (14)
För att säkra att uppgifterna i märkningen används på det sätt som avses i denna förordning bör det föreskrivas att de uppgifter lagras som behövs för att det i varje etapp av produktionen och saluföringen skall vara möjligt att kontrollera att uppgifterna i märkningen stämmer.
(14)
För att säkra att uppgifterna i märkningen används på det sätt som avses i denna förordning bör det föreskrivas att de uppgifter lagras som behövs för att det i varje etapp av produktionen och saluföringen skall vara möjligt att kontrollera att uppgifterna i märkningen stämmer.
Vissa av dessa uppgifter behöver dock inte lämnas vid den etapp då produkten saluförs till slutkonsumenten.
Ändring 5 Skäl 15a (nytt)
(15a) Medlemsstaterna bör fastställa vilka sanktioner som skall tillämpas vid överträdelser av bestämmelserna i denna förordning och se till att påföljderna verkställs.
Sanktionerna bör vara proportionerliga men tillräckligt avskräckande.
Förordningen skall tillämpas på kött från nötdjur
produceras i gemenskapen eller importeras från tredjeland.
____________
* Datum för ikraftträdandet av denna förordning.
rådets förordning (EEG) nr 1208/81
10
.
2.
Denna förordning skall tillämpas utan att det påverkar tillämpningen av
rådets förordning (EG) nr 1183/2006 av den 24 juli 2006 om fastställande av en gemenskapsskala för klassificering av slaktkroppar av vuxna nötkreatur
1
.
_____________________
10
EUT L 123, 7.5.1981, s.
3.
EUT L 214, 4.8.2006, s.
1.
3.
Ändring 9 Artikel 2
I denna förordning avses med kött oförpackade eller förpackade färska, kylda och frysta slaktkroppar, oförpackat eller förpackat färskt, kylt och fryst kött med ben och urbenat kött och oförpackade eller förpackade färska, kylda och frysta styckade och hela slaktbiprodukter från nötdjur på högst tolv månader.
I denna förordning avses med kött oförpackade eller förpackade färska, kylda och frysta slaktkroppar, oförpackat eller förpackat färskt, kylt och fryst kött med ben och urbenat kött och oförpackade eller förpackade färska, kylda och frysta styckade och hela slaktbiprodukter
som är avsedda för mänsklig konsumtion
från nötdjur på högst tolv månader.
Bestämmelserna i denna förordning gäller också för förädlade, bearbetade eller tillagade produkter som innehåller kött.
Ändring 10 Artikel 3
Kött från nötdjur på högst tolv månader får endast saluföras i medlemsstaterna under de för varje medlemsstat fastställda handelsbeteckningar som anges i bilaga II.
1.
Kött från nötdjur på högst tolv månader får endast saluföras i medlemsstaterna under de för varje medlemsstat fastställda handelsbeteckningar som anges i bilaga II.
Dessa beteckningar skall anges i samtliga handelsdokument.
2a.
Denna förordning skall tillämpas på kött från nötkreatur på mer än åtta månader endast när det saluförs under en annan beteckning än "nötkött" (eller motsvarande term för kött från vuxna nötkreatur på andra gemenskapsspråk).
1.
a)
Bokstavsbeteckning för aktuell kategori enligt bilaga I till denna förordning
, vid varje etapp av produktionen och saluföringen, utom vid saluföringen till slutkonsumenten
.
Ändring 15 Artikel 5, punkt 1, led b b)
Handelsbeteckning enligt artikel 4 i denna förordning
.
Ändring 16 Artikel 5, punkt 1a (ny)
1a.
utgår
Djurens identifieringsnummer och födelsedata
, som endast skall uppges vid slakterierna
.
Medlemsstaterna skall före den
[1 juli 2007]
1.
Medlemsstaterna skall före den
…*
utse den eller de myndigheter som skall ansvara för
de officiella kontrollerna
av tillämpningen av denna förordning och underrätta kommissionen om resultatet av kontrollerna.
Datum för förordningens ikraftträdande.
Ändring 20 Artikel 9a (ny)
Artikel 9a
Sanktioner
Medlemsstaterna skall fastställa vilka påföljder som skall tillämpas om det i samband med genomförda kontroller framkommer att villkoren i denna förordning inte respekteras.
Dessa påföljder skall vara effektiva, proportionerliga och avskräckande.
Medlemsstaterna skall informera kommissionen om dessa åtgärder senast den ...*, samt så snabbt som möjligt om alla påföljande ändringar av dessa.
________
* Tolv månader efter det att av denna förordning har trätt i kraft.
2.
utgår
Kategori
X
: nötdjur på högst åtta månader.
A)
Kategori
V
: nötdjur på högst åtta månader.
Bokstavsbeteckning för kategorin:
X
.
Bokstavsbeteckning för kategorin:
V
.
Kategori
Y
: nötdjur på mer än åtta månader, men högst tolv månader.
B)
Kategori
Z
: nötdjur på mer än åtta månader, men högst tolv månader.
Bokstavsbeteckning för kategorin:
Y
.
Bokstavsbeteckning för kategorin:
Z
.
Kött från nötdjur i kategori
X
:
A)
Kött från nötdjur i kategori
V
:
Kött från nötdjur i kategori
Y
:
B)
Kött från nötdjur i kategori
Z
:
P6_TA(2007)0093
Fullgörande av flaggstatsförpliktelser ***I
A6-0058/2007
Europaparlamentets lagstiftningsresolution av den 29 mars 2007 om förslaget till Europaparlamentets och rådets direktiv om fullgörande av flaggstatsförpliktelser ( KOM(2005)0586 – C6-0062/2006 – 2005/0236(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2005)0586 ) Ännu ej offentliggjort i EUT.
,
–
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för transport och turism ( A6-0058/2007 ).
1.
Europaparlamentet godkänner kommissionens förslag såsom ändrat av parlamentet.
2.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om kommissionen har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
3.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
P6_TC1-COD(2005)0236
(Text av betydelse för EES)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande EUT C
318, 23.12.2006, s.
195.
,
med beaktande av Regionkommitténs yttrande EUT C
229, 22.9.2006, s.
38.
,
i enlighet med förfarandet i artikel 251 i fördraget
Europaparlamentets ståndpunkt av den 29 mars 2007.
, och
av följande skäl: (1)
Säkerheten inom
sjöfarten i gemenskapen,
för dem som tillhandahåller sjöfartstjänster, liksom
(2)
Inom den internationella sjöfarten har det genom antagandet av ett antal konventioner för vilka Internationella sjöfartsorganisationen (IMO) är depositarie skapats ett omfattande ramverk för att öka sjösäkerheten och skyddet av miljön mot föroreningar från fartyg.
(3)
I enlighet med Förenta nationernas havsrättskonvention från 1982 (UNCLOS) och de konventioner för vilka IMO är depositarie, skall stater som är parter i dessa instrument utfärda lagar och förordningar och vidta nödvändiga åtgärder för att sätta dessa instrument i kraft helt och fullt, i syfte att skydda människoliv till havs och miljön genom att garantera att de fartyg som är i trafik är lämpliga för den verksamhet de är avsedda för och bemannat med behörigt sjöfolk.
(4)
de befintliga instrumenten för sjöfolk till ett enda instrument.
Konventionen omfattar
och
så snart som det har trätt i kraft
.
(5)
IMO-konventionerna bör ges full effekt i gemenskapen genom att konventionernas bindande bestämmelser införlivas med gemenskapens lagstiftning, eftersom alla medlemsstater skall vara parter i IMO-konventionerna och därmed är skyldiga att uppfylla konventionsförpliktelserna i fråga om fartyg under deras flagg.
(6)
De bindande bestämmelserna måste genomföras tillsammans med den relevanta gemenskapslagstiftningen om säkerheten i fråga om fartyg, besättningar, passagerare och last, och om förebyggande av förorening från fartyg och arbetstider för sjöfolk.
(7)
Några medlemsstater som ännu inte har fullbordat anslutningsprocessen för vissa IMO-konventioner – till exempel 1988 års SOLAS-konvention, lastlinjeprotokollen, MARPOL-bilagorna IV och VI och bilagorna till vissa IMO-konventioner som uttryckligen citeras i gemenskapslagstiftningen – bör uppmanas att slutföra dessa förfaranden.
(8)
av den ...
om gemensamma regler och standarder för organisationer som utför inspektioner och utövar tillsyn av fartyg och för sjöfartsadministrationernas verksamhet i förbindelse därmed
EUT L ...
(9)
IMO-resolution A.847 (20) upphävdes genom IMO-resolution A.973 (24) om koden för genomförande av bindande IMO-instrument, som innehåller de bindande bestämmelser som skall genomföras av flaggstater.
(10)
(11)
IMO-konventionerna ger flaggstaterna rätt att undanta fartyg från tillämpningen av grundläggande bestämmelser för flaggstater enligt IMO-konventionerna och att tillämpa likvärdiga bestämmelser, och detta har inneburit att administrationerna efter eget gottfinnande kan fatta beslut om ett stort antal krav.
Det krävs visserligen en viss flexibilitet i samband med genomförandet av särskilda åtgärder, men
(12)
I artikel 12 i rådets direktiv 98/18/EG av den 17 mars 1998 om säkerhetsbestämmelser och säkerhetsnormer för passagerarfartyg EGT L 144, 15.5.1998, s.
6).
utan att det påverkar tillämpningen av harmoniserade tolkningar som antas av IMO, på liknande bestämmelser för andra typer av fartyg som omfattas av IMO-konventionerna.
(13)
Sjöfartsadministrationerna i medlemsstaterna bör kunna förlita sig på resurser som är tillräckliga för fullgörandet av sina flaggstatsförpliktelser i proportion till flottans storlek och art och som grundar sig på relevanta IMO-krav.
(14)
Minimikriterier för dessa resurser bör fastställas med utgångspunkt i medlemsstaternas praktiska erfarenhet.
(15)
Ett obligatoriskt genomförande av de förfaranden som rekommenderas av IMO i MSC/Circ.1140/MEPC/Circ.424 av den 20 december 2004 om "Överföring av fartyg mellan stater" bör stärka de bestämmelser om byte av flagg som behandlas i IMO-konventionerna och i gemenskapens lagstiftning om sjösäkerhet, och de bör i sjösäkerhetens intresse öka öppenheten i förhållandet mellan flaggstater.
(16)
Medlemsstaterna bör för fartyg under deras flagg tillämpa harmoniserade krav på flaggstatens certifiering och besiktning enligt de relevanta förfaranden och riktlinjer som återfinns i bilagan till IMO-församlingens resolution A.948 (23) om riktlinjer för besiktning inom ramen för det harmoniserade systemet för besiktning och certifiering.
(17)
En sträng och grundlig kontroll av de erkända organisationer som utför flaggstaternas uppgifter på medlemsstaternas vägnar, och som står i proportion till storleken på och arten av medlemsstaternas flottor bör leda till en förbättring av den övergripande kvaliteten på fartyg som seglar under medlemsstaternas flaggor.
(18)
Om flaggstatsinspektörerna uppfyller vissa minimikrav bör detta garantera likvärdiga villkor för sjöfartsadministrationerna och höja kvaliteten på fartyg som seglar under medlemsstaternas flaggor.
(19)
Medlemsstaterna har förpliktelser såsom flaggstater när det gäller utredningar av olyckor och tillbud där deras fartyg är inblandade.
(20)
Medlemsstaterna skall följa de särskilda regler vid utredningar av olyckor vid sjötransporter som finns fastställda i
EUT L ...
.
(21)
IMO:s principer för säkerhetsbesättning bör bli bindande för att bidra till att förbättra kvaliteten på fartyg som seglar under medlemsstaternas flaggor.
(22)
En databas med viktiga uppgifter om fartyg som seglar under medlemsstaternas flaggor och fartyg som lämnat en medlemsstats register bör förbättra öppenheten när det gäller en högkvalitativ flottas prestanda, bidra till en bättre kontroll av flaggstaternas förpliktelser och skapa likvärdiga villkor för sjöfartsadministrationer.
(23)
(24)
(25)
IMO:s frivilliga revisionsprogram följer den standardiserade modellen för ett kvalitetsledningssystem som inkluderar principer, kriterier, revisionsområden, metoder och förfaranden som är lämpliga för att bedöma om medlemsstaterna genomför och verkställer de förpliktelser och åtaganden som ingår i de bindande IMO-konventioner som de är parter i.
Denna revisionsprocess kan därför redan nu föras in i gemenskapens lagstiftning om sjösäkerhet.
(26)
En kvalitetscertifiering av administrativa förfaranden i enlighet med ISO eller motsvarande normer skulle dessutom leda till likvärdiga villkor för sjöfartsadministrationer.
(27)
(28)
för att skapa synergier mellan flaggstaterna bör främjas av kommissionen
och bör tillhandahålla incitament för att registrera fartyg i medlemsstaternas register
(29)
Den europeiska sjösäkerhetsbyrån som inrättades genom Europaparlamentets och rådets förordning (EG) nr 1406/2002 EGT L 208, 5.8.2002, s.
1.
Förordningen senast ändrad genom förordning (EG) nr
1891/2006 (EUT L 394, 30.12.2006, s.
1).
bör ge det stöd som krävs för att detta direktiv skall genomföras.
(30)
De åtgärder som är nödvändiga för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter EGT L 184, 17.7.1999, s.
genom beslut 2006/512/EG (EUT L 200, 22.7.2006, s.
11).
.
(31)
I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå dessa mål.
1.
Syftet med detta direktiv är att
a)
se till att medlemsstaterna effektivt och konsekvent uppfyller sina förpliktelser som flaggstater enligt IMO-konventionerna
b)
öka säkerheten och förhindra föroreningar från fartyg som för en medlemsstats
flagg
,
c)
skapa en mekanism för en harmoniserad tolkning av de åtgärder som fastställs i IMO-konventionerna, och som tidigare har överlåtits åt parternas gottfinnande.
2.
1.
Förordningen senast ändrad genom kommissionens förordning (EG) nr 93/2007 (EUT L 22, 31.1.2007, s.
12).
eller rådets direktiv 1999/63/EG EGT L 167, 2.7.1999, s.
33.
.
1.
I detta direktiv gäller följande definitioner:
a)
"IMO-konventioner": följande konventioner, med tillhörande protokoll och ändringar och därmed förknippade koder med bindande status, antagna inom ramen för Internationella sjöfartsorganisationen (IMO), i uppdaterad version:
i)
1974 års internationella konvention om säkerheten för människoliv till sjöss (SOLAS 74)
ii)
1966 års internationella lastlinjekonvention (LL 66)
iii)
1969 års internationella konvention om skeppsmätning (TONNAGE 69)
iv)
v)
1978 års internationella konvention angående normer för sjöfolks utbildning, certifiering och vakthållning (STCW)
vi)
1972 års konvention om internationella regler till förhindrande av kollisioner till sjöss (COLREG 72)
vii)
1991 års kod för säkerheten vid transport av timmer som däckslast
viii)
1965 års kod för säkerheten vid transport av fast gods i bulk (BC-koden).
b)
c)
.
d)
"fartyg": fartyg och farkoster som omfattas av en eller flera IMO-konventioner.
e)
"administration": de behöriga sjöfartsmyndigheterna i den stat vars flagg fartyget har rätt att föra.
f)
"kvalificerad flaggstatsinspektör": en offentligt anställd tjänsteman eller annan person som är vederbörligen bemyndigad av en medlemsstats behöriga myndighet att utföra besiktningar och inspektioner som hänför sig till certifikaten och som uppfyller de kvalifikations- och oberoendekriterier som anges i bilaga II.
g)
[
h)
"certifikat": konventionscertifikat enligt IMO-konventionerna.
2.
det föreskrivande förfarande som avses
1.
Medlemsstaterna skall bli parter i IMO-konventionerna och de särskilda IMO-konventionerna.
Denna förpliktelse gäller emellertid bara konventionerna i den version som gäller på dagen för detta direktivs ikraftträdande.
2.
Medlemsstater som på dagen för detta direktivs ikraftträdande ännu inte är parter i samtliga IMO-konventioner och de särskilda IMO-konventionerna skall inleda ratifikations- eller anslutningsförfarandena för konventionerna i fråga enligt sin nationella lagstiftning.
De skall senast nittio dagar efter det att detta direktiv har trätt i kraft meddela kommissionen vid vilket datum de förväntas deponera ratifikations- eller anslutningsinstrumentet för konventionerna hos Internationella sjöfartsorganisationens generalsekreterare.
3.
Varje medlemsstat skall inom sin administration tydligt fördela arbetsuppgifter som gäller utformning och vidareutveckling av strategier för fullgörande av flaggstaternas åligganden enligt IMO-konventionerna, och se till att administrationen har förmåga att på ett lämpligt sätt bidra till utfärdandet av nationell lagstiftning och tillhandahålla vägledning om dess genomförande och upprätthållande.
4.
I synnerhet
när det gäller internationell sjöfart skall medlemsstaterna fullt ut tillämpa de bindande bestämmelser om flaggstater som fastställs i IMO-konventionerna i enligt med de villkor och avseende de fartyg som avses i dessa, och ta vederbörlig hänsyn till bestämmelserna i flaggstatskoden (FSC) i bilaga I till detta direktiv.
5.
Medlemsstaternas skall fortlöpande förbättra de åtgärder som vidtas för att genomföra IMO-konventionerna.
Förbättringar skall göras genom att den nationella lagstiftningen tillämpas och upprätthålls strängt och effektivt, och genom en fortlöpande kontroll av att reglerna följs.
6.
i artikel 18.2
får åtgärder antas i syfte att
a)
utveckla harmoniserade förfaranden för tillämpning av dispenser och liknande i enlighet med IMO-konventionerna,
b)
fastställa harmoniserade tolkningar av frågor som i IMO-konventionerna har överlåtits åt administrationernas gottfinnande,
c)
1.
Varje medlemsstat skall se till att dess administration har lämpliga resurser som står i proportion till dess flottas storlek och art.
Resurserna skall
a)
säkerställa att kraven i IMO-konventionerna
b)
säkerställa
att olyckor utreds och att fastställda brister hanteras korrekt och vid lämplig tidpunkt,
c)
medlemsstaterna i egenskap av fördragsslutande parter
d)
inbegripa ett lämpligt antal kvalificerade personer för att kunna tillämpa och upprätthålla den nationella lagstiftningen för genomförande av IMO-konventionerna, inbegripet
kvalificerade inspektörer från flaggstaten för att utföra
utredningar
e)
inbegripa ett tillräckligt antal kvalificerade flaggstatsanställda för att kunna utreda fall då fartyg som har rätt att föra medlemsstatens flagg har hållits kvar av en hamnstat,
f)
inbegripa ett tillräckligt antal kvalificerade flaggstatsanställda för att kunna utreda fall då en hamnstat har ifrågasatt giltigheten hos ett certifikat eller ett intyg om erkännande, eller behörigheten hos personer som har certifikat eller intyg om erkännande utfärdade av eller på uppdrag av flaggstaten.
2.
flaggstatsinspektörer och utredare, samt vid händelse av incidenter och brister, även kuststaten övervakas, liksom den
3.
Varje medlemsstat skall utarbeta eller bibehålla en kapacitet för
tekniskt beslutsfattande som står i proportion till dess flottas storlek och art.
4.
Minimikrav för uppfyllandet av de förpliktelser som fastställs i punkterna 1 och 2 skall antas i enlighet med
1.
Innan ett fartyg registreras skall medlemsstaten kontrollera dess identitet, inbegripet, i lämpliga fall, IMO-numret, och andra uppgifter om fartyget, så att fartyget inte seglar under två eller flera staters flagg samtidigt.
Det skall styrkas att ett fartyg som tidigare seglat under en annan stats flagg har strukits ur den statens register, eller att den statens registreringsmyndighet har samtyckt till överföring av fartyget.
2.
Som en förutsättning för att
ett fartyg skall
Medlemsstaten skall vid behov
och under alla omständigheter om fartyget inte är nybyggt
kontakta den tidigare flaggstaten
och begära att den överlämnar nödvändiga handlingar och uppgifter
.
3.
Om en begäran lämnas av en medlemsstat till en annan medlemsstat skall den tidigare flaggstaten vara skyldig att överlämna de berörda handlingarna och uppgifterna i enlighet med Europaparlamentets och rådets förordning (EG) nr 789/2004 av den 21 april 2004 om överföring av lastfartyg och passagerarfartyg mellan register inom gemenskapen
EUT L 138, 30.4.2004, s.
19.
.
4
5
skall tillämpas utan att det påverkar tillämpningen av artikel 4 i förordning (EG) nr 789/2004.
1.
Medlemsstaterna skall vidta alla åtgärder som är nödvändiga för att se till att fartyg som har rätt att föra deras flagg följer internationella regler och normer.
Dessa åtgärder skall särskilt inbegripa följande:
a)
Fartyg skall förbjudas att lägga ut innan de kan gå till sjöss utan att bryta mot internationella regler och normer.
b)
Fartyg skall bli föremål för regelbundna inspektioner av att fartygets skick och besättning stämmer överens med de certifikat som finns ombord.
c)
Under de regelbundna inspektioner som avses i b skall inspektören
på lämpligt sätt och med nödvändiga medel
kontrollera att det sjöfolk som förordnats för fartyget är väl förtrogna med sina arbetsuppgifter och fartygets arrangemang, installationer, utrustning och förfaranden.
d)
e)
Den nationella lagstiftningen skall innehålla bestämmelser om påföljder som är tillräckligt stränga för att avskräcka fartyg från att överträda internationella regler och normer.
f)
Förfaranden skall – efter utredning – inledas mot fartyg som har överträtt internationella regler och normer, oavsett var överträdelsen begicks.
g)
Den nationella lagstiftningen skall innehålla bestämmelser om påföljder som är tillräckligt stränga för att avskräcka personer med certifikat eller intyg om erkännande utfärdade av eller på uppdrag av medlemsstaten från att överträda internationella regler och normer.
h)
Förfaranden skall – efter utredning – inledas mot personer med certifikat eller intyg om erkännande som har överträtt internationella regler och normer, oavsett var överträdelsen begicks.
2.
Medlemsstaterna skall
, i enlighet med Europaparlamentets och rådets direktiv 2002/59/EG av den 27 juni 2002 om inrättande av ett övervaknings- och informationssystem för sjötrafik i gemenskapen
EGT L 208, 5.8.2002, s.
10.
,
utarbeta och genomföra ett lämpligt program för kontroll och övervakning
av fartyg som för deras flagg för att, inte minst genom användning av gemenskapssystemet för informationsutbyte SafeSeaNet, i god tid och på ett uttömmande sätt kunna tillmötesgå en begäran om information och klargöranden från en hamn- eller kuststat vid händelse av olyckor eller brister
.
3.
Medlemsstaterna, eller erkända organisationer som agerar för deras räkning, skall utfärda eller erkänna certifikat för ett fartyg först efter att de har fastställt att fartyget uppfyller alla tillämpliga krav.
4.
Medlemsstaterna skall utfärda ett internationellt behörighetscertifikat eller intyg om erkännande till en person först efter att de har fastställt att personen uppfyller alla tillämpliga krav.
5.
Medlemsstaterna skall se till att deras fartyg har besiktigats i enlighet med relevanta förfaranden och riktlinjer inom ramen för det harmoniserade system för besiktning och certifiering som fastställs i bilagan till IMO-församlingens resolution A.948 (23) i uppdaterad version.
6.
När ett fartyg som för en medlemsstats flagg hålls kvar av en hamnstat skall flaggstaten vidta åtgärder i enlighet med vägledningen i bilaga III.
7.
Bilaga III får ändras i enlighet med
1.
Medlemsstater som anlitar erkända organisationer för
[
2.
Medlemsstater som omfattas av punkt 1 skall
ha möjlighet
att
fartyg som för deras flagg, i syfte att se till att fartygen uppfyller kraven i IMO-konventionerna och de nationella kraven.
3.
som avses i punkt 2
för fartyg som
a)
har varit registrerade i medlemsstaten i
mindre än
två år,
b)
har
hållits kvar
i enlighet med
rådets
direktiv 95/21/EG
EGT L 157, 7.7.1995, s.
1.
53).
eller
Europaparlamentets och rådets
[
om hamnstatskontroll] *
.
4.
[
5.
Medlemsstater som omfattas av punkt 1 skall också
a)
utfärda särskilda instruktioner till sina erkända organisationer som noga beskriver vilka åtgärder som skall vidtas om det visar sig att ett fartyg inte kan gå till sjöss utan fara för fartyget eller människor ombord, eller visar sig utgöra ett orimligt hot mot den marina miljön, och
b)
förse sina erkända organisationer med alla lämpliga instrument i nationell lagstiftning och tolkning av denna för att bestämmelserna i IMO-konventionerna skall träda i kraft, eller ange om administrationens normer i något avseende går utöver de som föreskrivs i konventionerna.
6.
kompletterande utredningar
skall fastställas i enlighet med
1.
Medlemsstaterna skall definiera och dokumentera ansvarsområden, befogenheter och inbördes förhållande för all flaggstatspersonal som leder, utför och kontrollerar arbete som avser och påverkar säkerheten och förhindrandet av förorening.
2.
Medlemsstaterna skall se till att personal som ansvarar för eller utför besiktningar, inspektioner och revisioner på fartyg och företag, uppfyller de minimikrav som fastställs i bilaga II.
3.
Medlemsstaterna skall se till att annan personal än den som avses i punkt 2 som assisterar vid uppfyllandet av flaggstatens förpliktelser har utbildning och får handledning i proportion till de arbetsuppgifter de har behörighet att utföra.
4.
Medlemsstaterna skall
på lämpligt sätt och med nödvändiga medel
fortlöpande utveckling av kunskaperna hos den personal som avses i punkterna 1–3
, och kontinuerligt uppdatera personalens kunskaper på det sätt som krävs för de arbetsuppgifter de har fått
i uppdrag eller är behöriga
att utföra.
5.
Flaggstaten skall utfärda
6.
7
och de skyldigheter
som följer av koden för utredning av olyckor och tillbud till sjöss, antagen av IMO genom resolution
A.849 (20), bifogad IMO församlingens resolution A.884 (21), i uppdaterad version.
, oavsett var olyckan eller föroreningstillfället ägde rum.
Medlemsstaterna skall se till att fartyg som för deras flagg har adekvat bemanning ur sjösäkerhetssynpunkt och tillämpar principerna för säkerhetsbesättning enligt IMO-församlingens resolution A.890 (21) om principerna för säkerhetsbesättning, i uppdaterad version, med beaktande av relevanta riktlinjer som åtföljer den resolutionen.
1.
Medlemsstaterna skall utveckla eller upprätthålla en fartygsdatabas för sin flotta med de viktigaste tekniska uppgifterna om varje fartyg och de uppgifter som anges i punkt 2, eller se till att de har direkt tillgång till en databas som innehåller sådana uppgifter.
Medlemsstaterna skall ge kommissionen rätt att
få antingen egen eller delad tillgång, efter behov, till databaserna för
deras
fartyg och möjlighet att hämta uppgifter från
och utbyta data med dem.
2.
skall innehålla följande:
a)
Enskilda uppgifter för varje registrerat fartyg.
i)
Uppgifter om fartygen (namn, IMO-nummer etc.)
, registreringsdatum och i förekommande fall det datum då det ströks ur registret
.
ii)
Namnet på de erkända organisationer som har deltagit i fartygets certifiering och klassificering
iii)
.
iv)
Namnet på det organ som har inspekterat fartyget enligt bestämmelserna för hamnstatskontroll, och inspektionsdatum.
v)
Resultatet av hamnstatskontrollerna (brister:
; kvarhållanden:
).
vi)
Information om olyckor.
vii)
Information om överträdelser av
IMO-konventionerna, särskilt
11.
.
b)
Allmänna uppgifter beträffande alla fartyg i dess register.
i)
Förteckning över och
namn på fartyg som har utgått ur registret under de föregående tolv månaderna
ii)
Antal årliga inspektioner av alla slag, uppdelade efter besiktningstyp, som utförts av den berörda flaggstaten eller för dess räkning.
3.
i artikel 18.2.
4.
De uppgifter som avses i punkt 2 skall omedelbart överlämnas i sin helhet till den nya flaggstaten om ett fartyg utgår ur registret och överförs till ett annat register.
1.
Medlemsstaterna skall årligen utvärdera sin prestationsnivå i fråga om genomförande av bestämmelserna i det här direktivet.
2.
Utvärderingen av flaggstaternas prestationsnivåer skall bland annat inbegripa kvarhållandefrekvens inom ramen för hamnstatskontrollen, resultaten av flaggstatsinspektionerna, olycksstatistik, kommunikations- och informationsflöden, statistik över årliga förluster exklusive konstruktiva totalförluster, och andra lämpliga indikatorer, i syfte att avgöra om personal, resurser och administrativa förfaranden är tillräckliga för att fullgöra flaggstatsförpliktelserna.
3.
En gemensam metod för utvärdering av flaggstaternas prestationsnivåer skall fastställas i enlighet med
4.
Rapporten skall kartlägga de huvudsakliga skälen till den låga prestationsnivån, och ange de fartygskategorier som har orsakat resultatet.
Rapporten skall också innehålla en åtgärdsplan för bristernas avhjälpande, som vid behov kan föreskriva kompletteringsbesiktningar; planen skall genomföras snarast möjligt.
1.
Varje medlemsstat skall se till att en oberoende revision av hur medlemsstaten följer detta direktiv genomförs inom tre år efter det att direktivet har trätt i kraft, och därefter med jämna mellanrum.
2.
Revisionens omfattning och metod skall fastställas i enlighet med
Revisioner som utförs enligt bestämmelserna i
IMO-resolution A.974 (24) skall
godkännas som revision enligt punkt 1 om villkoren i punkt 3 är uppfyllda.
Ett sådant godkännande påverkar inte eventuella ytterligare inspektioner som kommissionen gör eller låter göra för att kontrollera att gemenskapens sjöfartslagstiftning följs.
3.
Medlemsstater som genomgår revision skall se till
a)
att det också kontrolleras att de följer bestämmelserna i det här direktivet,
b)
att kommissionen får möjlighet att delta som observatör i IMO-revisionen, och
c)
att kommissionen omedelbart får tillgång till rapporten och information om vilka åtgärder som kommer att vidtas.
4.
a)
fastställas en tidtabell för genomförandet av revisioner enligt punkt 1, och
b)
fastställas villkor för offentliggörandet av revisionsresultaten.
5.
Vid behov skall
kommissionen i samarbete med medlemsstaterna
utarbeta rekommendationer och förslag för att förbättra
förfarandena och resultaten
i IMO:s revisionsprogram
i det fall som avses i
punkt 2.
1.
Varje medlemsstat skall utarbeta, genomföra och upprätthålla ett kvalitetsledningssystem för sin administration.
Kvalitetsledningssystemet skall certifieras i enlighet med ISO-standarderna 9001:2000 eller en likvärdig standard som minst uppfyller alla delar av ISO 9001:2000, och det skall granskas i enlighet med ISO:s riktlinjer 19011:2002 eller en likvärdig standard som uppfyller alla delar av ISO 19011:2002.
När det gäller dessa likvärdiga standarder skall kraven enligt Europaparlamentets och rådets direktiv 98/34/EG EGT L 204, 21.7.1998, s.
37.
Direktivet senast ändrad genom 2003 års anslutningsakt.
vara uppfyllda.
2.
Kvalitetsledningssystemet skall införas inom tre år från det att detta direktiv träder i kraft.
3.
Kvalitetsledningssystemet skall certifieras inom fyra år från det att detta direktiv träder i kraft.
4.
Hänvisningarna till ISO-standarder i punkt 1 får uppdateras i enlighet med
Före utgången av [2007] skall kommissionen överlämna en rapport till Europaparlamentet och rådet om möjligheterna att utarbeta ett samförståndsavtal
mellan Europeiska gemenskapen, medlemsstaterna och tredjeländer
som har åtagit sig att tillämpa koden för genomförande av bindande IMO-instrument
genom IMO-resolutionen A.973 (24),
och som samtycker till att granskas i enlighet med
IMO-resolution A.974 (24)
.
Artikel 16
Tillhandahållande
av uppgifter och
meddelanden
1.
de uppgifter som krävs enligt IMO-konventionerna.
2.
Medlemsstaterna skall årligen underrätta kommissionen om
a)
hur många inspektioner och revisioner de har genomfört i egenskap av flaggstater,
b)
c)
3.
En harmoniserad blankettmall för
de obligatoriska rapporter
som avses i punkt 2 i denna artikel får fastställas i enlighet med
4.
Efter det att
uppgifterna
från medlemsstaterna har kommit in skall kommissionen utarbeta en konsoliderad rapport om genomförandet av det här direktivet.
Rapporten skall överlämnas till Europaparlamentet och rådet.
Artikel 17
Artikel 18
1.
Kommissionen skall biträdas av den kommitté för sjösäkerhet och förhindrande av förorening från fartyg (COSS) som inrättats enligt artikel 3 i förordning (EG) nr 2099/2002.
2.
1.
Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den […].
De skall genast överlämna texterna till dessa bestämmelser till kommissionen tillsammans med en jämförelsetabell för dessa bestämmelser och bestämmelserna i detta direktiv.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs.
Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2.
Medlemsstaterna skall till kommissionen överlämna texten till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Utfärdat i ... den ...
På Europaparlamentets vägnar På rådets vägnar
Ordförande Ordförande
BILAGA I
FLAGGSTATSKODEN (FSC) DELARNA 1 OCH 2 AV KODEN FÖR GENOMFÖRANDE AV BINDANDE IMO-INSTRUMENT DEL 1 – GEMENSAMMA OMRÅDEN
Syfte
1.
Syftet med denna kod är att öka sjösäkerheten i hela världen och förbättra skyddet av den marina miljön.
2.
Varje administration kommer att betrakta denna kod med utgångspunkt i deras egen situation, och kommer bara att vara bundna i fråga om genomförandet av de instrument som avses i punkt 6 som de själva är parter till.
På grund av geografi och omständigheter kan en del stater spela en viktigare roll som flaggstat än som hamnstat eller kuststat, medan andra är viktigare som hamnstater eller kuststater än som flaggstater.
En sådan obalans minskar inte på något sätt förpliktelserna som flaggstat, hamnstat eller kuststat.
Strategi
3.
För att en stat skall uppfylla syftet med denna kod bör staten utarbeta en strategi som täcker följande frågor:
1)
Genomförande och upprätthållande av relevanta internationella bindande instrument.
2)
Beaktande av internationella rekommendationer.
3)
Fortlöpande granskning och kontroll av statens fullgörande av internationella förpliktelser.
4)
Uppbyggnad, upprätthållande och förbättring av den övergripande organisationsstrukturens prestationsnivå och kapacitet.
Vid genomförandet av strategin bör den vägledning som ges i denna kod följas.
Allmänt
4.
Enligt bestämmelserna i Förenta Nationernas havsrättskonvention av 1982 (UNCLOS) och IMO-konventionerna är administrationerna ansvariga för att utfärda lagar och författningar och för att vidta alla andra åtgärder som kan krävas för att dessa instrument skall bli helt och fullt tillämpliga, så att det kan garanteras att ett fartyg är i tillräckligt gott skick för att användas till sitt avsedda ändamål och har den kompetenta personal som är nödvändig med tanke på skyddet för människoliv till havs och den marina miljön.
5.
Staterna skall, då de vidtar åtgärder för att förhindra, begränsa och kontrollera föroreningar av den marina miljön, handla på sådant sätt att de ej direkt eller indirekt överför skada eller risk från ett område till ett annat eller omvandlar en form av förorening till en annan (artikel 195 i UNCLOS).
Tillämpningsområde
6.
De bindande IMO-instrument som tas upp i denna kod är
1)
1974 års internationella konvention om säkerheten för människoliv till sjöss, i dess ändrade lydelse (SOLAS 74),
2)
1978 års protokoll till 1974 års internationella konvention om säkerheten för människoliv till sjöss, i dess ändrade lydelse (SOLAS PROT 1978),
3)
1988 års protokoll till 1974 års internationella konvention om säkerheten för människoliv till sjöss, i dess ändrade lydelse ((SOLAS PROT 1988),
4)
1973 års internationella konvention till förhindrande av förorening från fartyg, i dess lydelse enligt 1978 års protokoll (MARPOL 73/78),
5)
1997 års protokoll till 1973 års internationella konvention till förhindrande av förorening från fartyg, i dess lydelse enligt 1978 års protokoll (MARPOL PROT 1997),
6)
1978 års internationella konvention angående normer för sjöfolks utbildning, certifiering och vakthållning, i dess ändrade lydelse (STCW),
7)
1966 års internationella lastlinjekonvention (LL 66),
8)
1988 års protokoll till 1966 års internationella lastlinjekonvention (LL PROT 1988),
9)
1969 års internationella konvention om skeppsmätning (TONNAGE 69),
10)
1972 års konvention om internationella regler till förhindrande av kollisioner till sjöss, i dess ändrade lydelse (COLREG 72),
liksom instrument som gjorts bindande genom dessa konventioner och protokoll.
En icke uttömmande förteckning över förpliktelser enligt ovanstående bindande instrument finns i bilagorna 1–4.
En förteckning över de relevanta instrumenten finns i bilaga 5 och en sammanfattning av ändringarna av de bindande instrument som avspeglas i koden finns i bilaga 6 Bilagorna kommer att läggas till vid MSC 80 (maj 2005).
Bara bilagorna 1, 2 och 5 berör flaggstatsförpliktelser.
.
Inledande åtgärder
7.
När ett nytt eller ändrat bindande IMO-instrument träder i kraft för en stat måste regeringen i den staten kunna genomföra och upprätthålla bestämmelserna med hjälp av lämplig nationell lagstiftning och skapa nödvändig infrastruktur för genomförande och upprätthållande.
Detta innebär att statens regering måste ha följande:
1)
Förmåga att utfärda lagar som skapar en i praktiken tillämplig jurisdiktion och kontroll i administrativa, tekniska och sociala frågor över fartyg som för statens flagg, och, särskilt, lägger den rättsliga grunden för utfärdande av allmänna villkor i fråga om registreringsmyndigheter och inspektioner av fartyg, säkerhetslagstiftning och lagstiftning om förhindrande av förorening för sådana fartyg, samt utfärdande av därmed förknippade bestämmelser.
2)
En rättslig grund för upprätthållande av statens nationella lagstiftning, inbegripet utrednings- och straffrättsliga förfaranden.
3)
En tillräckligt stor personal med sakkunskap i sjöfartsfrågor som kan bistå vid utformningen av nödvändig nationell lagstiftning och fullgöra statens förpliktelser, inbegripet rapportering i enlighet med de olika konventionerna.
8.
.
Informationsförmedling
9.
Staten bör meddela alla berörda parter om sin strategi enligt punkt 3, inbegripet uppgifter om den nationella lagstiftningen.
Protokoll
10.
Lämpliga protokoll bör upprättas och arkiveras för att visa att kraven har uppfyllts och att staten fungerar effektivt.
Protokollen bör vara läsliga, lätta att identifiera och åtkomliga.
Ett dokumenterat förfarande bör fastställas för att närmare ange vilka kontroller som krävs för identifiering, arkivering, skydd, åtkomst, förvaringstid och disponering i fråga om protokollen.
Förbättringar
11.
Staterna bör fortlöpande förbättra de åtgärder som vidtas för att genomföra de konventioner och protokoll som de har godtagit.
Förbättringarna bör göras genom att nationell lagstiftning tillämpas och upprätthålls strängt och effektivt, och genom en fortlöpande kontroll av att reglerna följs.
12.
Staterna bör stimulera en kultur som ger människor möjlighet att förbättra arbetet för sjösäkerhet och miljöskydd.
13.
Vidare bör staterna vidta åtgärder för att kartlägga och eliminera orsakerna till eventuella åsidosättanden för att förhindra att de upprepas, inbegripet
1)
granskning och analys av åsidosättanden,
2)
genomförande av nödvändiga korrigerande åtgärder, och
3)
granskning av de korrigerande åtgärder som har vidtagits.
14.
Staten skall besluta om åtgärder för att eliminera orsakerna till tänkbara åsidosättanden för att förhindra att de uppkommer.
DEL 2 – FLAGGSTATER
Genomförande
15.
För att flaggstaterna skall fullgöra deras ansvar och förpliktelser effektivt bör de
1)
med hjälp av nationell lagstiftning och vägledning bedriva en politik som bidrar till att genomföra och upprätthålla kraven i alla konventioner och protokoll om säkerhet och förhindrande av förorening som de är parter i, och
2)
inom sin administration fördela ansvaret för att vid behov uppdatera och ändra den antagna politiken på relevanta områden.
16.
Flaggstaterna bör upprätta resurser och förfaranden som gör det möjligt att förvalta ett program för säkerhet och miljöskydd som åtminstone bör bestå av följande:
1)
Administrativa instruktioner för genomförande av tillämpliga internationella regler och föreskrifter och utarbetande och spridning av nödvändiga nationella tolkningsföreskrifter.
2)
Resurser för att se till att kraven i IMO:s bindande instrument enligt punkt 6 följs, genom ett revisions- och inspektionsprogram som är oberoende av förvaltningsorgan som utfärdar föreskrivna certifikat eller relevant dokumentation och andra organ som staten har bemyndigat att utfärda sådana certifikat eller sådan dokumentation.
3)
Resurser för att se till att kraven i 1978 års STCW-konvention, i dess ändrade lydelse, följs.
Detta inbegriper bland annat att
3.
1 utbildning, behörighetsbedömning och certifiering av sjöfolk är i överensstämmelse med bestämmelserna i konventionen,
3.
2 certifikat och intyg om erkännande (s.k. påteckning) enligt konventionen ger en korrekt bild av sjöfolkets kompetens, och är utformade med lämplig STCW-terminologi och termer som är identiska med dem som används i eventuella dokument om säkerhetsbesättning som utfärdas för fartyget,
3.
3 opartiska utredningar kan göras när det har rapporterats att någon som har ett certifikat eller intyg om erkännande (s.k. påteckning) utfärdat av den parten har begått ett fel – genom handling eller underlåtenhet att handla – som kan utgöra ett direkt hot mot säkerheten för människor, egendom till sjöss eller den marina miljön,
3.
4 certifikat eller intyg om erkännande (s.k. påteckning) som har utfärdats av flaggstaten kan dras tillbaka eller upphävas tillfälligt eller slutgiltigt när det är motiverat och när det krävs för att förhindra bedrägeri,
3.
5 administrativa arrangemang, även för utbildnings-, bedömnings- och certifieringsverksamheter som bedrivs under en annan stats överinseende, är sådana att flaggstaten åtar sig ansvaret för att se till att befälhavare, befäl och annat sjöfolk som tjänstgör på fartyg som har rätt att föra dess flagg har den behörighet som krävs Regler I/2, I/9, I/10 och I/11 i 1978 års STCW-konvention, i dess ändrade lydelse.
.
4)
Resurser för att se till att olyckor utreds och att fartyg med konstaterade brister hanteras lämpligt och inom lämplig tid.
5)
Utarbetande, dokumentering och tillhandahållande av vägledning om de krav som återfinns i de relevanta bindande IMO-instrumenten, som administrationen finner tillfredsställande.
17.
Flaggstaterna skall se till att fartyg som har rätt att föra deras flagg har tillräcklig och effektiv bemanning, med beaktande av IMO:s principer för säkerhetsbesättning.
Delegering av behörighet
18.
Flaggstater som bemyndigar erkända organisationer att agera för deras räkning när det gäller besiktningar, inspektioner, utfärdande av certifikat och dokument, märkning av fartyg och annat arbete enligt IMO-konventionerna, skall reglera bemyndigandena i enlighet med regel XI-1/1 i SOLAS enligt följande:
1)
Flaggstaten skall verifiera att den erkända organisationen har tillräckliga resurser i fråga om teknik, ledarskap och forskning för att genomföra de arbetsuppgifter den anförtros, i enlighet med de minimistandarder för erkända organisationer som agerar för administrationens räkning som fastställs i den relevanta IMO-resolutionen Bihang I till resolution A.739 (18), Riktlinjer för bemyndigande av organisationer som agerar för administrationens räkning.
.
2)
Bemyndigandet skall grundas antingen på ett skriftligt avtal mellan administrationen och den erkända organisationen som minst innehåller de element som fastställs i den relevanta IMO-resolutionen Bihang II till resolution A.739 (18), Riktlinjer för bemyndigande av organisationer som agerar för administrationens räkning.
, eller ett likvärdigt bindande rättsligt arrangemang; avtalet kan grundas på mallen för avtal om bemyndigande av erkända organisationer som agerar för administrationens räkning MSC/Circ.710 – MEPC/Circ.307.
.
3)
Flaggstaten skall utfärda särskilda instruktioner som noga beskriver vilka åtgärder som skall vidtas om ett fartyg visar sig ha brister som gör att det inte kan gå till sjöss utan fara för fartyget eller människor ombord, eller visar sig utgöra ett orimligt hot mot den marina miljön.
4)
Flaggstaten skall förse den erkända organisationen med alla lämpliga instrument i nationell lagstiftning och tolkning av denna bestämmelserna i konventionerna skall träda i kraft, eller ange om administrationens normer i något avseende går utöver vad som föreskrivs i konventionerna.
5)
Flaggstaten skall ålägga den erkända organisationen att föra och arkivera protokoll ur vilka administrationen kan hämta data som kan vara till hjälp vid tolkningen av konventionskraven.
19.
Flaggstater som utnämner inspektörer för att göra besiktningar och inspektioner för deras räkning bör reglera sådana utnämningar på lämpligt sätt i enlighet med vägledningen i punkt 18, särskilt 18.3 och 18.4.
20.
Flaggstaten bör införa eller delta i ett tillsynsprogram med tillräckliga resurser för att övervaka och kommunicera med dess erkända organisationer för att se till att dess internationella förpliktelser uppfylls helt, genom att flaggstaten
1)
utövar sina befogenheter att genomföra kompletteringsbesiktningar för att se till att fartyg som har rätt att föra dess flagg följer bestämmelserna i bindande IMO-instrument,
2)
genomför kompletteringsbesiktningar när den anser att det behövs för att se till att fartyg som har rätt att föra dess flagg följer nationella bestämmelser som kompletterar kraven i IMO-konventionerna, och
3)
tillhandahåller personal som har goda kunskaper om flaggstatens och de erkända organisationernas regler och bestämmelser och kan övervaka de erkända organisationerna på platsen.
Upprätthållande av lagstiftningen
21.
Flaggstaterna bör garantera fullgörandet av deras internationella förpliktelser genom att vidta alla nödvändiga åtgärder för att se till att fartyg som har rätt att föra deras flagg och enheter och personer inom deras jurisdiktion följer internationella regler och normer.
Sådana åtgärder bör bland annat inbegripa följande:
1)
Fartyg som har rätt att föra flaggstatens flagg bör förbjudas att lägga ut innan fartyget kan gå till sjöss utan att bryta mot de krav som ställs i internationella regler och normer.
2)
Fartyg som har rätt att föra flaggstatens flagg bör bli föremål för regelbundna inspektioner av att fartygets skick och besättning stämmer överens med de certifikat som finns ombord.
3)
Under de regelbundna inspektioner som avses i punkt 2 bör inspektören se till att det sjöfolk som har förordnats för fartyget är väl förtrogna med
3.
1 sina arbetsuppgifter, och
3.
2 arrangemang, installationer, utrustning och förfaranden på fartyget.
4)
De bör se till att hela besättningen kan samordna sin verksamhet i en nödsituation och i fråga om arbetsuppgifter av central betydelse för säkerheten eller för förhindrande eller begränsning av förorening.
5)
Den nationella lagstiftningen bör innehålla bestämmelser om påföljder som är tillräckligt stränga för att avskräcka fartyg som har rätt att föra flaggstatens flagg från att överträda internationella regler och normer.
6)
Förfaranden bör – efter utredning – inledas mot fartyg som har rätt att föra flaggstatens flagg som har överträtt internationella regler och normer, oavsett var överträdelsen begicks.
7)
Den nationella lagstiftningen bör innehålla bestämmelser om påföljder som är tillräckligt stränga för att avskräcka personer med certifikat eller intyg om erkännande utfärdade av eller på uppdrag av flaggstaten från att överträda internationella regler och normer.
8)
Förfaranden bör – efter utredning – inledas mot personer med certifikat eller intyg om erkännande som har överträtt internationella regler och normer, oavsett var överträdelsen begicks.
22.
Flaggstaterna bör överväga att utarbeta och genomföra ett program för kontroll och övervakning för att
1)
olyckor skall kunna utredas snabbt och grundligt, med – i tillämpliga fall – rapport till IMO,
2)
statistiska data skall samlas in, så att problemområden kan kartläggas genom trendanalys, och
3)
brister och påstådda föroreningstillfällen som rapporteras av hamn- eller kuststater kan åtgärdas vid lämplig tidpunkt.
23.
Vidare bör flaggstaten
1)
se till att den nationella lagstiftningen garanterar att bindande IMO-instrument följs,
2)
tillhandahålla ett lämpligt antal kvalificerade personer för att kunna tillämpa och upprätthålla den nationella lagstiftning som avses i punkt 15.1, inbegripet personal som genomför utredningar och besiktningar,
3)
tillhandahålla ett tillräckligt antal kvalificerade flaggstatsanställda för att kunna utreda fall då fartyg som har rätt att föra dess flagg har hållits kvar av hamnstater,
4)
tillhandahålla ett tillräckligt antal kvalificerade flaggstatsanställda för att kunna utreda fall då en hamnstat har ifrågasatt giltigheten hos ett certifikat eller intyg om erkännande eller behörigheten hos personer som har certifikat eller intyg om erkännande utfärdat av eller på uppdrag av flaggstaten,
5)
se till att flaggstatsinspektörer och utredare utbildas, och att deras verksamhet övervakas.
24.
När en flaggstat får besked om att ett fartyg som har rätt att föra dess flagg har hållits kvar av en hamnstat bör flaggstaten se till att lämpliga korrigerande åtgärder vidtas så att fartyget omedelbart bringas i överensstämmelse med krav som ställs i tillämpliga internationella konventioner.
25.
En flaggstat eller en erkänd organisation som agerar för dess räkning bör utfärda eller erkänna ett internationellt certifikat för ett fartyg först efter det att den har fastställt att fartyget uppfyller alla tillämpliga krav.
26.
En flaggstat bör utfärda ett internationellt behörighetscertifikat eller intyg om erkännande till en person först efter det att de har fastställt att personen uppfyller alla tillämpliga krav.
Flaggstatsinspektörer
27.
Flaggstaten bör definiera och dokumentera ansvarsområden, befogenheter och inbördes förhållanden för all personal som leder, utför och kontrollerar arbete som avser och påverkar säkerheten och förhindrande av förorening.
28.
Personal som ansvarar för eller utför besiktningar, inspektioner och revisioner på fartyg och företag som omfattas av de relevanta bindande IMO-instrumenten bör minst ha följande kvalifikationer:
1)
Lämpliga kvalifikationer från en havs- eller sjöfartsinstitution och relevant erfarenhet till sjöss som fartygsbefäl med behörighet enligt STCW II/2 eller III/2, och bibehållna tekniska kunskaper om fartyg och handhavande av fartyg sedan behörighetscertifikatet erhölls, eller
2)
en teknisk eller naturvetenskaplig högskole- eller universitetsexamen eller motsvarande inom ett relevant ämnesområde som erkänns av staten.
29.
30.
31.
Dessutom bör sådan personal ha de lämpliga praktiska och teoretiska kunskaper om fartyg, handhavande av fartyg och bestämmelser i relevanta nationella och internationella instrument som krävs för att de skall kunna sköta sina arbetsuppgifter som flaggstatsinspektörer; dessa kunskaper skall ha inhämtats genom dokumenterade utbildningsprogram.
32.
Annan personal som assisterar vid sådant arbete bör ha utbildning och få handledning i proportion till de arbetsuppgifter de har behörighet att utföra.
33.
Relevant erfarenhet på området bör betraktas som en fördel; om personen saknar erfarenhet bör administrationen tillhandahålla lämplig praktisk utbildning.
34.
Flaggstaterna får ge inspektörsbehörighet åt personer som har genomgått ett formellt och detaljerat utbildningsprogram som ger den kunskapsnivå som krävs enligt punkterna 29–32.
35.
Flaggstaten bör ha infört ett dokumenterat system för kvalifikation av personal och fortlöpande uppdatering av deras kunskaper till en nivå som är lämplig med hänsyn till de arbetsuppgifter de är behöriga att utföra.
36.
Kvalifikationerna bör, beroende på vilka arbetsuppgifter som kommer i fråga, omfatta
1)
kunskap om tillämpliga nationella och internationella regler och föreskrifter för fartyg och fartygens företag, besättningar, last och handhavande,
2)
kunskap om de förfaranden som används vid besiktning, certifiering, kontroll, undersökning och övervakning,
3)
insikter i mål och syften med internationella och nationella instrument om sjösäkerhet och skydd av den marina miljön, och program som hänger samman med dessa,
4)
kunskaper om arbetsmetoderna ombord och i land, interna och externa,
5)
den nödvändiga yrkesmässiga kompetensen för att utföra arbetsuppgifterna väl och effektivt,
6)
säkerhetsmedvetenhet i alla situationer, också när det gäller den personliga säkerheten, och
7)
utbildning i eller erfarenhet av de olika arbetsuppgifter som skall utföras, och helst också i de funktioner som skall bedömas.
37.
Flaggstaten bör utfärda en identitetshandling som inspektören bär med sig under arbetet.
Flaggstaternas utredningar
38.
Sjöolyckor och föroreningstillfällen bör utredas.
Utredningar av olyckor bör göras av utredare med lämpliga kvalifikationer som är kompetenta i frågor som rör olyckan.
Flaggstaten bör vara beredd att ställa kvalificerade utredare till förfogande för detta ändamål, oavsett var olyckan eller föroreningstillfället ägde rum.
39.
Flaggstaten bör se till att de enskilda utredarna har praktiska kunskaper om och praktisk erfarenhet av de ämnesområden som ingår i deras normala arbetsuppgifter.
För att bistå enskilda utredare i deras arbete med frågor som ligger utanför deras normala uppdrag bör flaggstaten se till att lämplig expertis inom följande områden vid behov är lätt tillgänglig:
1)
Navigerings- och kollisionsregler.
2)
Flaggstatens bestämmelser om behörighetscertifiering.
3)
Havsföroreningarnas orsaker.
4)
Intervjuteknik.
5)
Bevisupptagning.
6)
Bedömning av den mänskliga faktorns inverkan.
40.
Alla olyckor som leder till personskador som kräver frånvaro från arbetet i tre dagar eller mer och alla dödsfall till följd av arbetsolyckor eller skador på flaggstatens fartyg bör utredas, och resultatet av utredningen offentliggöras.
41.
Fartygsolyckor bör utredas och rapporteras i enlighet med relevanta IMO-konventioner och de riktlinjer som har utarbetats av IMO Se koden för utredning av olyckor och tillbud till sjöss som antogs av IMO genom resolution A.849 (20), i dess lydelse enligt resolution A.884 (21).
.
Utredningsrapporten bör sändas till IMO tillsammans med flaggstatens iakttagelser i enlighet med de riktlinjer som avses ovan.
Utvärdering och granskning
42.
Flaggstaterna bör regelbundet utvärdera sin prestationsnivå i fråga om genomförandet av de administrativa metoder, förfaranden och resurser som krävs för att uppfylla deras förpliktelser enligt de konventioner som de är parter till.
43.
Utvärderingarna av flaggstaternas prestationsnivå kan bland annat inbegripa kvarhållandefrekvens inom ramen för hamnstatskontrollen, resultaten av flaggstatsinspektionerna, olycksstatistik, kommunikations- och informationsflöden, statistik över årliga förluster (exklusive konstruktiva totalförluster – CTL) och andra lämpliga indikatorer, i syfte att avgöra om personal, resurser och administrativa förfaranden är tillräckliga för att fullgöra flaggstatsförpliktelserna.
44.
Utvärderingarna kan inbegripa en regelbunden granskning av följande:
1)
Fartygsförluster och olycksfrekvenser, i syfte att kartlägga trender under utvalda tidsperioder.
2)
Antalet verifierade fall av kvarhållna fartyg i förhållande till flottans storlek.
3)
Antalet verifierade fall av inkompetens eller oegentligheter begångna av personer som har certifikat eller intyg om erkännande utfärdade av eller på uppdrag av flaggstaten.
4)
Vilka åtgärder som har vidtagits när hamnstater har rapporterat brister eller ingripanden.
5)
Utredningar av allvarliga olyckor och de lärdomar som kan dras av dessa.
6)
Ekonomiska, tekniska och andra resurser som tagits i anspråk.
7)
Resultatet av inspektioner, besiktningar och kontroller av fartygen i fartygsflottan.
8)
Utredningar av arbetsolyckor.
9)
Antalet incidenter och överträdelser enligt MARPOL 73/78, i dess ändrade lydelse.
10)
Antalet tillfälliga eller slutgiltiga indragningar av certifikat, intyg om erkännande, godkännanden m.m.
BILAGA II
MINIMIKRAV PÅ FLAGGSTATSINSPEKTÖRER (enligt artikel 8)
1.
Inspektörer skall vara bemyndigade av medlemsstatens behöriga myndighet att genomföra de besiktningar som avses i detta direktiv.
2.
Inspektörerna skall ha lämpliga teoretiska kunskaper om och praktisk erfarenhet av fartyg, handhavande av fartyg och relevant nationella och internationella krav.
Dessa kunskaper och erfarenheter skall ha inhämtats genom dokumenterade utbildningsprogram.
3.
Inspektörer skall ha minst något av följande:
1)
Lagstadgad examen
från en havs- eller sjöfartsinstitution
behörighet enligt STCW II/2 eller III/2.
2)
tre år, eller ett år kompletterat med två års praktik som fartygsinspektör hos en medlemsstats behöriga myndighet
.
3)
En relevant universitetsexamen eller motsvarande, och ha utbildats och godkänts på en skola för inspektörer och praktiserat som fartygsinspektör i minst två år hos en behörig
myndighet
.
4
.
5
6.
Inspektörer skall kunna kommunicera muntligt och skriftligt med sjöfolk på det språk som är vanligast till sjöss.
7.
, personligt eller familjemässigt
intresse
med anknytning till
det fartyg som besiktigas
icke-statliga organisationer som gör konventions- eller klassningsrelaterade besiktningar eller utfärdar certifikat för fartyg.
8
BILAGA III
VÄGLEDNING FÖR UPPFÖLJNING NÄR FARTYG HAR HÅLLITS KVAR AV EN HAMNSTAT (enligt artikel 6)
1.
NÄR EN HAMNSTAT HAR HÅLLIT KVAR ETT FARTYG
1
annan
hamnstat bör myndigheten se till att lämpliga korrigerande åtgärder vidtas så att fartyget bringas i överensstämmelse med tillämpliga regler och internationella konventioner.
Nedanstående åtgärder anses lämpliga, och listan förhindrar inte att åtgärder med liknande verkningar eller kompletterande åtgärder antas, förutsatt att de är förenliga med målen för och bestämmelserna i detta direktiv.
2.
OMEDELBARA ÅTGÄRDER
1.
Så snart flaggstaten får besked om kvarhållandet bör den kontakta företaget (med företag avses här ett företag enligt ISM-koden) och hamnstaten för att såvitt möjligt få alla närmare uppgifter om kvarhållandet.
2.
Mot bakgrund av de uppgifterna bör flaggstaten överväga vilka omedelbara åtgärder som krävs för att bringa fartyget i överensstämmelse.
Flaggstaten kan anse att vissa brister enkelt kan åtgärdas och godkännas av hamnstaten (exempelvis om en livbåt behöver service).
I så fall bör flaggstaten be hamnstaten bekräfta att bristerna har åtgärdats.
3.
en erkänd organisation, bör flaggstaten begära att en
särskild, kompletterande
inspektion utförs av någon av dess inspektörer, eller utse en inspektör från den erkända organisationen att göra en inspektion för dess räkning.
Inledningsvis bör denna inspektion koncentreras på de områden där hamnstaten har konstaterat brister.
Om inspektören från flaggstaten eller den erkända organisationen anser det nödvändigt kan inspektionen sedan utvidgas till en fullständig ombesiktning av de områden som omfattas av de relevanta konventionscertifikaten.
4.
Om den erkända organisationen har genomfört inspektionen enligt
punkt 3
bör organisationens inspektör rapportera till flaggstaten om vilka åtgärder som har vidtagits och om fartygets skick efter inspektionen, så att flaggstaten kan avgöra vilka eventuella ytterligare åtgärder som behövs.
5.
[
om hamnstatskontroll] bör flaggstaten ordna en ombesiktning av fartyget i fråga om de certifikat som gäller de områden där flaggstaten har noterat brister och andra områden där brister senare upptäcks.
Flaggstaten bör antingen genomföra denna besiktning själv eller begära en fullständig rapport från den erkända organisationens inspektör, och vid behov en bekräftelse på att en tillfredsställande besiktning har genomförts och alla brister åtgärdats.
När flaggstaten är nöjd med situationen bör den bekräfta för hamnstaten att fartyget uppfyller kraven i relevanta bestämmelser och internationella konventioner.
6.
När det gäller de allvarligaste överträdelserna av bestämmelser och internationella konventioner bör flaggstaten alltid skicka en egen inspektör, snarare än en inspektör från den erkända organisationen, för att genomföra eller övervaka de inspektioner och besiktningar som avses i
punkt 3–5.
7.
Utom i de fall som avses i
punkt 10
skall flaggstaten begära att korrigerande åtgärder vidtas av företaget så att fartyget bringas i överensstämmelse med tillämpliga bestämmelser och internationella konventioner innan fartyget tillåts lämna hamnen där det har hållits kvar (utöver de korrigerande åtgärder som hamnstaten har krävt).
Om inga sådana korrigerande åtgärder vidtas bör de berörda certifikaten dras in.
8.
Flaggstaten bör överväga i vilken utsträckning brister noterade av en hamnstat och upptäckta vid en flaggstatsinspektion eller flaggstatsbesiktning tyder på att fartygets och företagets säkerhetsorganisation inte fungerar.
Vid behov bör flaggstaten arrangera en ny revision av fartyget eller företaget och tillsammans med hamnstaten överväga om revisionen bör äga rum innan fartyget tillåts lämna den hamn där det har hållits kvar.
9.
Flaggstaten bör kontinuerligt stå i kontakt och samarbeta med hamnstaten för att bidra till att de brister som har konstaterats åtgärdas, och bör snarast möjligt besvara eventuella begäran om klargörande från hamnstaten.
10.
[
om hamnstatskontroll] tillåter fartyget att fortsätta till ett reparationsvarv bör flaggstaten kontakta hamnstaten för att bestämma på vilka villkor resan får äga rum och bekräfta dessa villkor skriftligen.
11.
Om fartyget inte uppfyller de villkor som avses i
punkt 10
eller inte anlöper det överenskomna reparationsvarvet bör flaggstaten omedelbart begära en förklaring från företaget och överväga att dra in fartygets certifikat.
Dessutom bör flaggstaten så snart det blir möjligt tilläggsbesiktiga fartyget.
12.
Om flaggstaten mot bakgrund av tillgängliga uppgifter anser att kvarhållandet är omotiverat bör den göra hamnstaten uppmärksam på detta och tillsammans med företaget överväga att överklaga beslutet i enlighet med hamnstatens bestämmelser.
3.
YTTERLIGARE ÅTGÄRDER
1.
Beroende på hur allvarliga de konstaterade bristerna är och vilka omedelbara åtgärder som har vidtagits bör flaggstaten också överväga att tilläggsbesiktiga fartyget efter det att kvarhållandet har upphört.
Denna besiktning bör inbegripa en bedömning av säkerhetsorganisationens effektivitet.
Ett riktmärke är att en tilläggsbesiktning bör göras inom [6] veckor efter det att flaggstaten fick besked om kvarhållandet.
Denna besiktning bör göras på företagets bekostnad.
Om flaggstaten planerar att genomföra en konventionsrelaterad besiktning inom [3] månader kan den skjuta upp besiktningen till dess.
2.
Vidare bör flaggstaten överväga om det bör genomföras en ny revision av det företag som är inblandat.
Flaggstaten skall också se över tidigare inspektionsrapporter om företagets andra fartyg, för att se om det finns några gemensamma nämnare när det gäller bristerna i det företagets flotta.
3.
Om fartyget har hållits kvar på goda grunder mer än en gång under de föregående 2 åren bör uppföljningen anses vara än mer angelägen, och i alla händelser bör flaggstaten tilläggsbesiktiga fartyget inom [4] veckor efter det att flaggstaten fick besked om kvarhållandet.
4.
[
om hamnstatskontroll] skall flaggstaten tilläggsbesiktiga fartyget och vidta alla nödvändiga åtgärder för att se till att företaget bringar fartyget i överensstämmelse med samtliga relevanta konventioner och bestämmelser.
När flaggstaten har försäkrat sig om att så har skett skall den skicka ett dokument som bekräftar detta till företaget.
5.
gemenskapsbestämmelser
och internationella konventioner bör flaggstaten överväga vilka ytterligare påföljder som kan krävas, inbegripet att stryka fartyget ur dess register.
6.
Efter fullbordande av de åtgärder som skall bringa fartyget i överensstämmelse
med internationella
konventioner
och gemenskapsbestämmelserna
bör flaggstaten skicka en rapport till IMO
och kommissionen, som, med avseende på IMO, skall utarbetas
i enlighet med regel 19 d i kapitel I i SOLAS 74, i dess ändrade lydelse och punkt 5.2 i IMO-resolution A.787 (19), i dess ändrade lydelse
4.
TILLÄGGSBESIKTNING
1.
En tilläggsbesiktning bör inbegripa en undersökning av nedan uppräknade områden som är tillräckligt grundlig för att flaggstatsinspektören skall vara säker på att fartyget, dess utrustning och dess besättning uppfyller alla krav i de bestämmelser och internationella konventioner som är tillämpliga:
Certifikat och dokument.
Skrovets struktur och utrustning.
Villkoren för fastställande av fribord.
Huvudmaskineri och viktiga system.
Renlighet i maskinutrymmena.
Livräddningsutrustning.
Brandsäkerhet.
Navigeringsutrustning.
Lasthanteringsutrustning.
Radioutrustning.
Elektrisk utrustning.
Förhindrande av förorening.
Bostads- och arbetsvillkor.
Bemanning.
Besättningens certifikat.
Passagerarsäkerhet.
Driftskrav, inbegripet kommunikation i besättningen, övningar, arbetet på bryggan och i maskinrummet och säkerhet.
2.
Den bör också inbegripa de relevanta punkterna för en utökad inspektion
enligt bilaga
Flaggstatsinspektörer bör inte avstå från att vid behov inbegripa funktionstester på exempelvis livräddningsfarkoster och deras sjösättningsanordningar, huvud- och hjälpmaskineri, lastluckor, huvudelsystem och system för länspumpning.
P6_TA(2007)0153
Multilateralt avtal om inrättande av ett gemensamt europeiskt luftrum
B6-0148/2007
Europaparlamentets resolution av den 25 april 2007 om förslaget till rådets beslut om ingående av det multilaterala avtalet mellan Republiken Albanien, Bosnien och Hercegovina, Republiken Bulgarien, Europeiska gemenskapen, Republiken Island, Republiken Kroatien, f.d. jugoslaviska republiken Makedonien, Konungariket Norge, Serbien och Montenegro, Rumänien och Förenta nationernas övergångsförvaltning i Kosovo om inrättandet av ett gemensamt europeiskt luftrum
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till rådet ( KOM(2006)0113 ) Ännu ej offentliggjort i EUT.
,
–
med beaktande av Europaparlamentets resolution av den 17 januari 2006 om fortsatt utveckling av EU:s luftfartspolitik gentemot länder utanför EU EUT C 287 E, 24.11.2006, s.
84.
,
–
A.
B.
B Rådet har antagit det provisoriska avtalet i enlighet med kommissionens förslag och detta avtal bör ännu ratificeras av alla avtalsslutande parter.
C.
Avtalet om ett gemensamt europeiskt luftrum är viktigt som ramavtal för att lösa luftfartsrelaterade frågor, särskilt med länderna på västra Balkan, Island och Norge, och det erbjuder en modell för framtida avtal av detta slag med andra tredjeländer.
Miljön
1.
Europaparlamentet anser att det är viktigt att avtalet om ett gemensamt europeiskt luftrum omfattar nuvarande och framtida gemenskapslagstiftning om utsläpp och andra åtgärder som minskar luftfartens miljökonsekvenser.
2.
Man bör välkomna det faktum att signatärstaterna accepterar att utsläpp från luftfarten i framtiden eventuellt kommer att inkluderas i systemen för handel med utsläppsrätter.
3.
Europaparlamentet betonar att avtalet är viktigt för att skapa förutsättningar för att utöka det gemensamma europeiska luftrummet (SES), så att det sträcker sig utanför EU:s medlemsstater.
Säkerhet
4.
Europaparlamentet understryker betydelsen av teknisk assistans och anslutningsförhandlingar bör därför uttryckligen betonas som medel för att få till stånd den konsensus med partner utanför EU och EES som är nödvändig för att uppnå detta mål.
5.
Europaparlamentet insisterar på att all gemenskapslagstiftning på området för säkerhet och Europaparlamentets och rådets förordning (EG) nr 1107/2006 av den 5 juli 2006 måste om rättigheter i samband med flygresor för personer med funktionshinder och personer med nedsatt rörlighet EUT L 204, 26.7.2006, s.
1.
skall inkluderas i den operationella bilagan till avtalet.
6.
Flygledningstjänster ingår i avtalet, vilket är viktigt för tillämpningen av bestämmelserna om SES, exempelvis dem för utvecklandet av gränsöverskridande luftrumsblock.
7.
Europaparlamentet välkomnar fördelarna med alla avtalsslutande parters ömsesidiga och konsekventa tillämpning av Europaparlamentets och rådets direktiv 2004/36/EG av den 21 april 2004 om säkerheten i fråga om luftfartyg från tredje land som använder flygplats i gemenskapen EUT L 143, 30.4.2004, s.
76.
Direktivet ändrat genom förordning (EG) nr 2111/2005 (EUT L 344, 27.12.2005, s.
15).
.
8.
Europaparlamentet påminner om att genomförandet av SES medför även flexibilitet i luftrummet som fordrar ett institutionaliserat samarbete mellan militära och civila myndigheter på flygledningsområdet.
Sociala frågor
9.
Europaparlamentet välkomnar den roll som Europeiska byrån för luftfartssäkerhet har för att fortbilda experter, utarbeta manualer och tillhandahålla teknisk rådgivning i partnerländerna samt bidra till att inrätta genomförandemekanismer.
10.
Europaparlamentet betonar att tillämplig gemenskapslagstiftning på området för sociala frågor skall respekteras vid genomförandet av avtalet.
11.
Europaparlamentet noterar att avtalet föreskriver tillämpning av rådets förordning (EEG) nr 3922/91 av den 16 december 1991 om harmonisering av tekniska krav och administrativa förfaranden inom området civil luftfart EGT L 373, 31.12.1991, s.
4.
Förordningen senast ändrad genom Europaparlamentets och rådets förordning (EG) nr 1900/2006 (EUT L 377, 27.12.2006, s.
176).
.
12.
Europaparlamentet noterar att åtagandena i avtalet skall genomföras snarast och en framstegsrapport skall läggas fram för Europaparlamentet senast den 31 december 2008.
13.
Europaparlamentet uppmanar kommissionen och rådet att se till att avtalet återspeglar dessa viktiga aspekter och att det inrättas en övervakningsmekanism i samband med genomförandeprocessen.
o
o o
14.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet och kommissionen.
P6_TA(2007)0301
Fastställande av en ny statistisk indelning av produkter efter näringsgren (CPA) ***I
A6-0242/2007
Europaparlamentets lagstiftningsresolution av den 10 juli 2007 om förslaget till Europaparlamentets och rådets förordning om fastställande av en ny statistisk indelning av produkter efter näringsgren (CPA) och om upphävande av förordning (EEG) nr 3696/93 ( KOM(2006)0655 – C6-0376/2006 – 2006/0218(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2006)0655 ) Ännu ej offentliggjort i EUT.
,
–
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för ekonomi och valutafrågor ( A6-0242/2007 ).
1.
Europaparlamentet godkänner kommissionens förslag såsom ändrat av parlamentet.
2.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
P6_TC1-COD(2006)0218
Europaparlamentets ståndpunkt fastställd vid första behandlingen den 10 juli 2007 inför antagandet av Europaparlamentets och rådets förordning (EG) nr .../2007 om fastställande av en ny statistisk indelning av produkter efter näringsgren (CPA) och om upphävande av rådets förordning (EEG) nr 3696/93
(Eftersom det nåddes en överenskommelse mellan parlamentet och rådet, motsvarar parlamentets ståndpunkt vid första behandlingen den slutliga rättsakten, förordning (EG) nr .../2007.)
P6_TA(2007)0343
Unionens framtida havspolitik
A6-0235/2007
Europaparlamentets resolution av den 12 juli 2007 om unionens framtida havspolitik: En europeisk vision för oceanerna och haven ( 2006/2299(INI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens grönbok "Unionens framtida havspolitik: En europeisk vision för oceaner och hav" ( KOM(2006)0275 ),
–
–
,
–
med beaktande av artikel 45 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för transport och turism och yttrandena från utskottet för miljö, folkhälsa och livsmedelssäkerhet, utskottet för industri, forskning och energi, fiskeriutskottet och utskottet för regional utveckling ( A6-0235/2007 ), och av följande skäl:
A.
B.
C.
D.
E.
F.
G.
H.
Uppskattningar i FN:s miljöprogram visar att cirka 80 procent av havsföroreningarna orsakas av landbaserade källor.
I.
J.
Stora fartyg för med sig stora mängder bunkrad olja under färden, och denna olja kan vid en olyckshändelse eller tillbud orsaka stora miljöskador och har redan orsakat stora skador, och möjligheterna är små att rätta till och gottgöra skadorna.
K.
Enligt officiella uppskattningar är 80 procent av de olyckshändelser som sker till sjöss direkt orsakade av den mänskliga faktorn.
L.
M.
Havsvattennivån har stigit och hotar därmed kustområden, deras befolkning och näringar som kustturism.
N.
De många olika havs- och kustverksamheterna kräver flexibel fysisk planering från medlemsstaternas och deras myndigheters sida.
O.
P.
Q.
Havsmotorvägarna hör sedan 2004 till de 30 mest prioriterade projekten inom ramen för TEN, men ännu har mycket få framsteg gjorts.
R.
S.
T.
U.
Havet och oceanerna spelar en viktig roll för produktionen av energi från alternativa energikällor och ökar energileveranssäkerheten.
V.
Det är nödvändigt att uppmärksamma den särskilda situationen för EU:s yttersta randområden och öar, framför allt när det gäller olaglig invandring, naturkatastrofer, transporter och dessa områdens bidrag till den biologiska mångfalden.
W.
En stor del av EU:s yttre gräns utgörs av hav, och övervakningen och skyddet av denna gräns innebär extra kostnader för kustmedlemsstaterna.
X.
Medelhavet och Svarta havet delas mellan EU-medlemsstaterna och tredjeländer som har mindre resurser att genomföra miljöbestämmelser och säkerhets- och skyddsåtgärder.
1.
2.
Europaparlamentet välkomnar en havspolitik som kräver att politik, åtgärder och beslut som rör havsfrågor skall integreras och som främjar bättre samordning, mer öppenhet och ökat samarbete mellan alla aktörer vars verksamhet påverkar Europas oceaner och hav.
3.
Europaparlamentet konstaterar att när ansvaret för politik och åtgärder som rör haven fördelas mellan EU:s myndigheter, nationella regeringar och regionala och lokala myndigheter bör de beslutsfattande organen på alla nivåer sträva efter ett mer samordnat synsätt som ser till att deras verksamhet på havsområdet tar full hänsyn till den höga graden av interaktion mellan dem.
4.
Europaparlamentet uppmanar kommissionen att beakta de olika rekommendationerna i den ovannämnda resolutionen av den 15 mars 2007 och framför allt att prioritera inrättandet av en administrativ enhet för öar inom kommissionen, för att kunna utveckla den sedan länge efterlysta sektorsövergripande strategin som skall hantera problemen i dessa områden och för att öarna skall ges en riktig plats i EU:s statistiska program i samband med den framtida havspolitiken.
5.
Klimatförändringarna är den största utmaningen för havspolitiken
6.
7.
Europaparlamentet betonar att EU måste inta en ledande och vägvisande ställning i kampen mot klimatförändringarna.
8.
Europaparlamentet betonar att kust- och havsbaserad vindkraft har en mycket stor utvecklingspotential och kan ge ett betydande bidrag till klimatskyddet och uppmanar därför kommissionen att vidta åtgärder genom att inrätta en stab eller samordningsenhet för vindkraft och genom att införa en handlingsplan för vindkraft.
9.
10.
11.
12.
Europaparlamentet insisterar på att man vid planering av utvecklingsprojekt längs med gemenskapens långa kust, såsom stadsutveckling, industrianläggningar, små och stora hamnar, fritidsanläggningar etc. uttryckligen måste beakta konsekvenserna av klimatförändringarna och de därmed sammanhängande höjningarna av havsnivån, inbegripet den ökade frekvensen och styrkan av stormar och den ökade höjden på vågorna.
13.
Europaparlamentet understryker vikten av en övergripande strategi, som exempelvis en strategi som syftar till en integrerad förvaltning av kustområdena, för att åtgärderna skall bli effektiva.
Den förbättrade europeiska sjöfarten med bättre europeiska fartyg
14.
15.
1).
16.
17.
18.
Europaparlamentet uppmanar kommissionen att stödja den europeiska varvsindustrin, som hela tiden är utsatt för illojal konkurrens från de asiatiska skeppsbyggarna, genom interventioner på WTO-nivå.
19.
Europaparlamentet välkomnar kommissionens arbetsdokument om hur arbetet med initiativet LeaderSHIP 2015 fortskrider ( KOM(2007)0220 ) och betonar särskilt framgången med det nya heltäckande synsättet på industripolitik som LeaderSHIP 2015 gick i bräschen för, som ett av de första sektorsvisa initiativen.
20.
Europaparlamentet betonar att bättre (gränsöverskridande) samordning och samarbete mellan hamnar, och en mer balanserad fördelning av ansvaret mellan EU:s hamnar i hög grad kan bidra till att undvika ohållbara landtransporter.
21.
22.
–
att fastställa utsläppsstandarder för kväveoxider för fartyg som använder hamnar i EU,
–
att utse Medelhavet och nordöstra Atlanten till övervakningsområden för utsläpp av svaveloxider (SECA-områden) enligt Marpolkonventionen,
–
att sänka den högsta tillåtna svavelhalten i marina bränslen som används av passagerarfartyg i SECA-områden från 1,5 procent till 0,5 procent,
–
att införa instrument som skatter eller avgifter på utsläpp av svaveldioxid eller kväveoxider från fartyg,
–
att uppmuntra differentierade avgifter i hamnar och farleder som gynnar fartyg med lägre utsläpp av svaveldioxid eller kväveoxider,
–
att uppmuntra fartyg att använda landström när de ligger i hamn,
–
ett EG-direktiv om kvaliteten på marina bränslen.
23.
24.
25.
11.
.
26.
Europaparlamentet erkänner kommissionens aktiviteter på området för fartygs- och sjösäkerhet efter fartygskatastroferna med "Erika" och "Prestige", vars viktigaste resultat är åtgärdspaketen om sjöfartssäkerhet.
27.
Europaparlamentet kräver eftertryckligen att rådet (transport) snabbt förbereder "det tredje sjösäkerhetspaketet" och fattar ett gemensamt beslut tillsammans med Europaparlamentet för att det inte skall uppstå en trovärdighetslucka.
28.
Europaparlamentet uppmanar kommissionen att förstärka alla åtgärder som rör civilt och straffrättsligt skadeståndsansvar vid olyckor eller tillbud, samtidigt som subsidiaritetsprincipen, kompetensfördelningen och det internationella regelverket måste respekteras.
29.
Europaparlamentet påminner om sin resolution av den 21 april 2004 om ökad sjösäkerhet EUT C 104 E, 30.4.2004, s.
730.
och kräver att kommissionen i nästa steg på ett bättre sätt tar hänsyn till den mänskliga faktorn.
30.
31.
32.
Europaparlamentet påminner kommissionen om kravet att så snart som möjligt lägga fram ett förslag till parlamentet och rådet för att kunna säkerställa att bunkerolja för bränsle i nya fartyg också lagras i säkrare tankar med dubbla skrov, eftersom frakt- och containerfartyg ofta har tung brännolja som bränsle i sina bränsleförråd i sådana mängder som ofta avsevärt överstiger mindre oljetankfartygs frakt.
Parlamentet anser att kommissionen, innan den lägger fram ett sådant förslag, först måste undersöka huruvida de befintliga IMO-regler som har fastställts i MEPC-resolution 141.54 är tillräckliga för att garantera säker transport av bunkerolja som används som bränsle.
33.
Europaparlamentet uppmanar kommissionen att skärpa övervakningen av tillämpningen av bestämmelserna om obligatorisk användning av dubbla skrov.
34.
35.
36.
Europaparlamentet uppmanar medlemsstaterna och den marina sektorns berörda parter att se över karriärplanerna och möjligheterna till livslångt lärande inom den marina sektorn, dels för att kunna använda förvärvade färdigheter och erfarenheter i praktiken, dels för att kunna införa system för att skifta mellan havs- och landbaserade yrken så att expertisen bevaras och karriärmöjligheterna blir attraktivare.
37.
38.
Europaparlamentet anser i likhet med vad som föreslås i ovannämnda grönbok att arbetsmarknadens parter bör se över det faktum att sjömän inte omfattas av sociala direktiv.
39.
Europaparlamentet framhåller att fiskare och sjömän undantas från många områden av sociallagstiftningen inom EU (exempelvis direktiv 98/59/EG EGT L 225, 12.8.1998, s.
16.
16.
om skydd för arbetstagares rättigheter vid överlåtelse av företag, verksamheter eller delar av företag eller verksamheter, direktiv 2002/14/EG EGT L 80, 23.3.2002, s.
29.
om inrättande av en allmän ram för information till och samråd med arbetstagare samt direktiv 96/71/EG om utstationering av arbetstagare i samband med tillhandahållande av tjänster EGT L 18, 21.1.1997, s.
Parlamentet uppmanar kommissionen att i nära samarbete med arbetsmarknadens parter granska dessa undantagsbestämmelser.
40.
41.
Europaparlamentet kräver att en europeisk kvalitetsmärkning för fartyg införs, i linje med IMO:s vita klassificeringslista, som motsvarar senaste säkerhetsstandarder och sociala villkor, vilket medför att dessa fartyg får preferensbehandling inom ramen för hamnstatskontrollen.
42.
43.
44.
45.
Europaparlamentet konstaterar att ett av huvudmålen med havspolitiken är att skapa förutsättningar som säkerställer hygien, säkerhet och komfort för de anställda inom fiskeindustrin, både för fiskarna själva och för dem som arbetar inom sektorer i tidigare och senare led av produktionskedjan.
46.
Europaparlamentet anser att i jämförelse med lagstiftning är begreppet företagens sociala ansvar av begränsat värde i samband med att bevara havsmiljön, och att en korrekt rättslig grund därför måste fortsätta att lägga till grund för gemenskapens program för att bevara miljön, vilket skall förstärkas med frivilliga åtgärder från de företag som önskar visa sitt ansvarsfulla beteende.
47.
48.
49.
50.
51.
Europaparlamentet begär att utbildning och information skall tillhandahållas genom insamling, analys och spridning av bästa praxis, tekniker, instrument för att övervaka tanktömning och innovativa åtgärder för att bekämpa oljeföroreningar och föroreningar av giftiga och farliga ämnen, och att man skall utveckla tekniska lösningar – med användning av inspektion och satellitbaserad övervakning – för att övervaka läckage som sker genom olyckshändelser eller med avsikt.
En bättre europeisk kustpolitik, inklusive bättre europeiska hamnar
52.
53.
54.
55.
56.
Europaparlamentet anser att det är mycket viktigt att utveckla system för tidig varning längs de områden längs de delar av Atlantens kuster som riskerar att drabbas av tsunamier.
57.
Europaparlamentet understryker hamnarnas grundläggande betydelse för kanaliseringen av den internationella handeln, som ekonomiska motorer, som skapare av arbetstillfällen i kustregioner, som marknadsplats för fisket och som viktiga säkerhetskontrollpunkter.
58.
51.
, så att de medlemsstater som utnyttjar möjligheten att bli befriade från skatt på bunkerolja, i enlighet med artikel 14 i direktivet, förpliktar att i samma utsträckning befria landbaserad elektricitet från skatt.
59.
Europaparlamentet kräver en översynav Europaparlamentets och rådets direktiv 2000/59/EG av den 27 november 2000 om mottagningsanordningar i hamn för fartygsgenererat avfall och lastrester
EGT L 332, 28.12.2000, s.
60.
61.
62.
63.
64.
40.
och tillämpliga internationella konventioner samt regelbunden övervakning och kontroll.
65.
66.
Europaparlamentet insisterar emellertid på att ett av huvudmålen för förvaltningen av kustområden måste vara att bevara havsmiljön snarare än att etablera några få förevisningsområden som tecken på åtgärder för bevarande, i synnerhet med beaktande av Europaparlamentets och rådets rekommendation 2002/413/EG av den 30 maj 2002 om genomförandet av en integrerad förvaltning av kustområden i Europa EGT L 148, 6.6.2002, s.
24.
.
67.
68.
69.
70.
71.
Europaparlamentet uppmuntrar inrättandet av nya nätverk för att genomföra projekt och verksamheter i form av partnerskap mellan den privata sektorn, frivilligorganisationer och lokala myndigheter och regioner i syfte att skapa ökad dynamik, innovation och effektivitet och att förbättra livskvaliteten i kustområdena.
72.
73.
74.
75.
76.
77.
3.
78.
Europaparlamentet uppmuntrar kommissionen att genomföra specifika, vetenskapliga, miljömässiga och socioekonomiska statistiska och andra undersökningar av havsregionerna, i syfte att övervaka och kontrollera vilka effekter utvecklingen av ekonomiska aktiviteter och idrotts- och fritidsaktiviteter har i dessa regioner.
79.
80.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att göra samtliga berörda parter delaktiga i alla steg i processen för att förbättra EU:s havspolitik, både vid genomförandet och verkställandet av befintlig lagstiftning och vid utarbetandet av nya initiativ.
Hållbar turism i kustområden
81.
82.
83.
Europaparlamentet understryker att avsaknaden av ändamålsenliga och jämförbara uppgifter är ett av nyckelproblemen när det gäller att erhålla tillförlitliga uppgifter om sysselsättningssituationen inom turismen i kustområden.
84.
85.
Europaparlamentet konstaterar att Europa är en favoritdestination för kryssningsfartyg och betonar att tillhandahållandet av tjänster bör organiseras på ett sätt som garanterar fri konkurrens, och att behovet av bättre infrastruktur på detta område måste tillfredsställas.
86.
87.
Europaparlamentet anser att EU:s Agenda 21 för en hållbar europeisk turism måste ta hänsyn till kustturismens – och öturismens – särdrag och lägga fram användbara initiativ och utbyta god praxis för att på ett effektivt sätt bekämpa sektorns säsongsbetonade karaktär, exempelvis utveckla turism för äldre människor.
88.
Europaparlamentet uppmanar kommissionen att lägga fram en hållbar maritim europeisk turismstrategi som följer ett integrerat politiskt tillvägagångssätt.
En hållbar maritim miljö
89.
Europaparlamentet påminner om sin resolution av den 14 november 2006 om en temainriktad strategi för skydd och bevarande av den marina miljön Antagna texter, P6_TA(2006)0486 .
och upprepar särskilt behovet av att
-
EU:s övergripande mål skall vara en hållbar användning av haven och att bevara de marina ekosystemen, vilket inbegriper en stark EU-politik om marint skydd som skall förhindra ytterligare förluster av den biologiska mångfalden och ytterligare försämring av den marina miljön,
-
införa en för hela gemensam EU-definition av god miljöstatus,
-
Europeiska miljöbyrån tillhandhåller regelbundna bedömningar av den marina miljön, vilket kräver förbättringar av den nationella insamlingen, rapporteringen och utbytet av uppgifter,
-
erkänna betydelsen av samråd på förhand, samordning och samarbete med angränsande länder vid antagande och genomförande av det kommande direktivet om en marin strategi.
90.
Europaparlamentet konstaterar att en sund havsmiljö utgör grunden för en hållbar utveckling inom EU:s sjöfartssektor och erinrar om EU:s åtagande att inbegripa miljöaspekterna i alla delar av gemenskapspolitiken.
91.
92.
93.
Europaparlamentet understryker med eftertryck behovet av att de kriterier som används för att definiera ett gott miljötillstånd är tillräckligt långtgående, eftersom dessa mål som hänför sig till kvalitet troligen kommer att vara styrande för åtgärdsprogrammen under lång tid framöver.
94.
Europaparlamentet anser vidare att åtgärder för att förbättra vattenkvaliteten måste vidtas snabbt och är därför bekymrat över den utsträckta tidsplan som föreslås i förslaget till direktiv om en marin strategi.
95.
Europaparlamentet begär med eftertryck att genomförandet av nätverket för marina skyddade områden skall påskyndas.
96.
97.
98.
Europaparlamentet anser att klusterkonceptet skulle kunna ha positiva effekter på havsmiljön om bevarande av livsmiljöer, kontroll av föroreningar och andra miljötekniker införlivas i utformningen och genomförandet av klustren från planeringsstadiet och framåt.
99.
Parlamentet betonar att alla system med marin fysisk planering på EU-nivå måste tillföra ett mervärde i förhållande till de nationella systemen och planerna, där sådana finns, och att de måste grunda sig på de marina regionerna och underregionerna i direktivet om en marin strategi och främja användningen av en ekosystembaserad strategi till marin förvaltning och målen med god miljöutveckling enligt direktivet om en marin strategi.
100.
Europaparlamentet noterar att uppnående av god miljöstatus också kräver att mänskliga verksamheter som utförs utanför ekologiskt känsliga områden skall regleras noga så att all eventuell negativ påverkan på havsmiljön minimeras.
Integrerad fiskeripolitik
101.
102.
103.
104.
Europaparlamentet uppmanar kommissionen att ta vederbörlig hänsyn till de goda erfarenheterna av lokala och regionala myndigheters förvaltning av fisket så att de kan tillämpas som modell inom andra regioner, speciellt de erfarenheter som omfattar en integrerad och hållbar förvaltning av havet genom ett förbud mot icke-selektiv fiskeutrustning, anpassning av fiskeflottornas storlek till befintliga resurser, kustplanering, reglering av turistaktiviteter såsom valskådning, utarbetande av förvaltningsplaner för områden inom Natura 2000-nätet och inrättande av skyddade områden.
105.
Europaparlamentet betonar att de regionala rådgivande nämndernas värdefulla rådgivande roll bör erkännas och nämnderna bör rådfrågas angående förvaltning av den marina miljön.
106.
107.
108.
109.
110.
111.
112.
113.
Europaparlamentet betonar vikten av att övervaka fisket på internationellt vatten, eftersom detta även påverkar fiskeresurserna inom EU:s exklusiva ekonomiska zoner.
Havsforskning, energi, teknik och innovation
114.
115.
116.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att utarbeta och genomföra ett mätprogram för havsbottnen och kustvattnen i Europa, för att på denna grund kunna utveckla en europeisk havsatlas.
117.
118.
119.
120.
121.
Europaparlamentet betonar - utöver det att skadliga metoder måste avskaffas - vikten av att utveckla sådan verksamhet utanför fisket som är förenlig med fiskesektorn genom att exempelvis uppmuntra planering av plattformar för energiproduktion eller vindturbiner som bidrar till att främja och bevara ett blomstrande ekosystem och därmed underlättar inrättandet av lek- och yngelområden för marina arter i områden där det råder fiskeförbud.
122.
123.
124.
Europaparlamentet anser mot bakgrund av den ovanligt snabba utvecklingen av avsaltningsanläggningar för havsvatten, som släpper ut tonvis med saltlösning och andra produkter i havet, att kommissionen bör inleda studier om dessa anläggningars inverkan på plankton och havsbotten samt på förändringar och mutationer i ekosystemet.
125.
126.
127.
Europaparlamentet påpekar att eftersom de yttersta randområdena i Atlanten och Indiska oceanen och ligger bra till för att observera fenomen som rör vädercykler och vulkanologi, och eftersom oceanografi, biologisk mångfald, miljökvalitet, förvaltning av naturresurser, energi och vatten, genetik, folkhälsa, hälsovetenskap, nya telekommunikationssystem och -tjänster i dessa territorier är favoritområden för europeisk forskning, bör man ta hänsyn till dessa regioner vid planeringen av framtida forsknings- och utvecklingsprogram.
128.
129.
En gemensam havspolitik
130.
131.
132.
133.
134.
135.
136.
Europaparlamentet anser att fullständigt genomförande i god tid av all gemenskapslagstiftning på miljöområdet (vilken omfattar bland annat ramdirektivet om vatten Europaparlamentets och rådets direktiv 2000/60/EG av den 23 oktober 2000 om upprättande av en ram för gemenskapens åtgärder på vattenpolitikens område (EGT L 327, 22.12.2000, s.
1).
, habitatdirektivet, fågeldirektivet, nitratdirektivet Rådets direktiv 91/676/EEG av den 12 december 1991 om skydd mot att vatten förorenas av nitrater från jordbruket (EGT L 375, 31.12.1991, s.
1).
, direktivet om marina bränslens svavelhalter Rådets direktiv 1999/32/EG av den 26 april 1999 om att minska svavelhalten i vissa flytande bränslen och om ändring av direktiv 93/12/EEG (EGT L 121, 11.5.1999, s.
13).
och direktivet om föroreningar förorsakade av fartyg och införandet av sanktioner för överträdelser) är absolut nödvändigt för att havsmiljöns kvalitet skall bevaras, och att kommissionen bör utöva de påtryckningar som behövs för att uppmuntra medlemsstaterna att uppnå detta, om nödvändigt även genom lagstiftningsåtgärder.
137.
138.
139.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att i anslutning till sin havspolitik genomföra grundliga undersökningar av de gamla ammunitionsförråd från tidigare krig som sänkts i de europeiska haven och den fara som dessa utgör för människor och miljön samt vidta eventuella säkrings- och/eller bärgningsåtgärder.
140.
141.
Europaparlamentet betonar att EU aktivt måste engagera sig i marin förvaltning på internationell nivå för att främja rättvisa konkurrensvillkor för marin ekonomi, utan att äventyra ambitionerna vad gäller de marina verksamheternas miljömässiga hållbarhet.
142.
143.
144.
i)
Säkerheten till sjöss och skydd av den marina miljön (bland annat övervakning av fisket), skydd mot terrorism, sjöröveri och sjöfartsbrottslighet samt mot olagligt, oreglerat och icke-rapporterat fiske.
ii)
Genomförandet av samordnade inspektioner av fisket och verkställandet av bestämmelser på samma sätt inom hela EU samt medlemsstaternas domstolars tillämpning av likadana sanktioner och påföljder.
iii)
145.
Europaparlamentet förväntar sig att den europeiska grannskapspolitiken ska ta hänsyn till EU:s havspolitik och nödvändigheten att samarbeta med EU:s grannländer när det gäller miljö, havsskydd och sjösäkerhet.
146.
147.
148.
149.
o
o o
150.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet och kommissionen samt till Europeiska ekonomiska och sociala kommittén och Regionkommittén.
P6_TA(2007)0362
Naturkatastrofer
B6-0323 , 0324 , 0325 och 0327/2007
Europaparlamentets resolution av den 4 september 2007 om naturkatastrofer
Europaparlamentet utfärdar denna resolution
–
med beaktande av artiklarna 2, 6 och 174 i EG-fördraget,
–
med beaktande av sina resolutioner av den 7 september 2006 om skogsbränder och översvämningar EUT C 305 E, 14.12.2006, s.
240.
, den 5 september 2002 om översvämningskatastrofen i Europa EUT C 272 E, 13.11.2003, s.
471.
, den 14 april 2005 om torkan i Portugal EUT C 33 E, 9.2.2006, s.
599.
, den 12 maj 2005 om torkan i Spanien EUT C 92 E, 20.4.2006, s.
414.
, den 8 september 2005 om naturkatastrofer (bränder och översvämningar) i Europa EUT C 193 E, 17.8.2006, s.
322.
och sina resolutioner av den 18 maj 2006 om naturkatastrofer (bränder och översvämningar) – jordbruksaspekter EUT C 297E, 7.12.2006, s.
363.
, – regionala utvecklingsaspekter EUT C 297 E 7.12.2006, s.
369.
och – miljöaspekter EUT C 297 E 7.12.2006, s.
375.
,
–
med beaktande av de två gemensamma utfrågningarna organiserade av utskottet för regional utveckling, utskottet för miljö, folkhälsa och livsmedelssäkerhet och utskottet för jordbruk och landsbygdens utveckling om en EU-strategi för naturkatastrofer (den 20 mars 2006) och om en europeisk civilskyddsstyrka: Europe Aid (den 5 oktober 2006),
–
med beaktande av rådets beslut 2001/792/EG, Euratom av den 23 oktober 2001 om inrättande av en gemenskapsindustri för att underlätta ett förstärkt samarbete vid biståndsinsatser inom räddningstjänsten EGT L 297, 15.11.2001, s.
7.
samt av det förväntade antagandet av rådets omarbetade beslut om gemenskapens räddningstjänstmekanism och parlamentets ståndpunkt av den 24 oktober 2006 om detsamma EUT C 313 E, 20.12.2006, s.
100.
,
–
med beaktande av kommissionens förslag till Europaparlamentets och rådets förordning om inrättande av Europeiska unionens solidaritetsfond ( KOM(2005)0108 ) och av parlamentets ståndpunkt av den 18 maj 2006 om detsamma EUT C 297 E, 7.12.2006, s.
331.
,
–
med beaktande av Michel Barniers rapport av den 9 maj 2006 om en europeisk civilskyddsstyrka: Europe Aid,
–
,
–
med beaktande av rådets beslut 2007/162/EG, Euratom av den 5 mars 2007 om inrättande av ett finansiellt instrument för civilskydd EUT L 71, 10.3.2007, s.
9.
,
–
med beaktande av slutsatserna från rådets (rättsliga och inrikes frågor) möte den 12–13 juni 2007 om stärkandet av övervaknings- och informationscentrets samarbetsförmåga inom ramen för gemenskapens räddningstjänstmekanism,
–
med beaktande av Kyotoprotokollet till Förenta nationernas ramkonvention om klimatförändringar (UNFCCC) av den 11 december 1997 och gemenskapens ratificering av Kyotoprotokollet den 4 mars 2002,
–
med beaktande av förordning (EG) nr 2152/2003 av den 17 november 2003 (Forest Focus-förordningen) EUT L 324, 11.12.2003, s.
1.
,
–
med beaktande av punkt 12 i ordförandeskapets slutsatser från Europeiska rådets möte i Bryssel den 15 och 16 juni 2006 om unionens förmåga att agera vid stora olyckor, kriser och katastrofer,
–
med beaktande av kommissionens meddelande om problemet med vattenbrist och torka i Europeiska unionen KOM(2007)0414 ,
–
A.
B.
C.
Enbart de förödande skogsbränderna som nyligen härjat i Grekland kostade mer än 60 människor livet och skadade många samt ledde till mer än 250 000 hektar nedbränd skog och snårskog, döda djur, ett stort antal förstörda hus och egendomar samt utplånade byar.
D.
E.
F.
G.
Naturkatastroferna får svåra ekonomiska och sociala konsekvenser för regionala ekonomier, produktiv verksamhet och turism.
H.
Det stora antalet skogsbränder i södra Europa under 2007 och deras omfattning beror på flera olika faktorer däribland klimatförändringar, otillräcklig och bristande skogsvård samt en kombination av naturliga orsaker och mänskligt slarv, men även brottslig verksamhet och en bristande tillämpning av lagar som förbjuder olaglig byggnation på nedbrunnen mark.
I.
EU måste erkänna särdragen hos naturkatastroferna (såsom torka och bränder) i Medelhavsområdet, samt anpassa sina instrument för förebyggande, forskning, riskhantering, civilskydd och solidaritet.
1.
Europaparlamentet uttrycker sitt djupa deltagande och sin starka solidaritet med anhöriga till dem som förlorat sina liv och med invånarna i de berörda områdena.
2.
Europaparlamentet betygar sin vördnad för de brandmän, andra fackmän och frivilliga som oförtröttligt arbetat och riskerat sina liv med att släcka bränder, rädda människor och begränsa de skador som uppstått till följd av sommarens naturkatastrofer och alla de enskilda medborgare som kämpat med att försöka rädda det som var deras livsuppehälle och den omgivande miljön.
3.
4.
Europaparlamentet uppmanar kommissionen att anslå särskilt ekonomiskt gemenskapsbistånd till stöd för återställandet av de regioner som har drabbats hårt, återskapa de drabbade områdenas produktionspotential, försöka återuppta arbetet med att skapa arbetstillfällen och vidta lämpliga åtgärder för att kompensera de sociala kostnader som följer av förlusten av arbetstillfällen och andra inkomstkällor.
5.
6.
7.
8.
9.
10.
11.
Europaparlamentet anser att de erfarenheter som man gjort under tidigare år och den senaste tiden understryker behovet av att öka gemenskapens förebyggande åtgärder, beredskap och insatser inom räddningstjänsten när det gäller skogsbränder och andra vilda bränder, och uppmanar med kraft kommissionen att ta ett initiativ i denna riktning.
12.
13.
14.
15.
16.
17.
18.
19.
Europaparlamentet betonar att det i samband med naturkatastrofer måste tas särskild hänsyn till funktionshindrades särskilda behov i alla åtgärder som vidtas med användning av räddningstjänstmekanismerna.
20.
21.
Europaparlamentet anser att det för att garantera ett långsiktigt skogs- och områdesskydd krävs en hållbar programplanering och tillämpning av regionala utvecklingsplaner och landsbygdsutvecklingsplaner som syftar till att minska avfolkningen av landsbygdsområden och som genererar nya diversifierade landsbygdsinkomster, särskilt för den yngre generationen, och som inrättar den nödvändiga moderniserade infrastruktur som främjar en hållbar turism och hållbara tjänster i landsbygdsområdena.
22.
23.
24.
Europaparlamentet uppmanar kommissionen att övervaka att alla katastrofmedel som medlemsstaterna ställt till förfogande används på ett korrekt, ändamålsenligt och effektivt sätt för att hantera följderna av naturkatastroferna och uppmanar medlemsstaterna att se till att gemenskapsstöd som använts på felaktigt sätt betalas tillbaka, exempelvis i samband med återbeskogningsprogram som inte fullföljts, och att se till att fastighetsregistren uppdateras.
25.
Europaparlamentet fördömer legalisering av olaglig byggverksamhet på skyddade områden och i områden där bygglov i allmänhet inte ges och uppmanar till att alla försök att minska skogsskyddet genom ändring av den grekiska konstitutionen (artikel 24) omedelbart stoppas.
26.
Europaparlamentet föreslår att det sänds en delegation från parlamentet till de länder som drabbats värst av den senaste tidens naturkatastrofer för att uttrycka parlamentets medkänsla med befolkningen, för att se hur allvarlig förstörelsen är när det gäller liv, egendomar, sociala nätverk, miljö och ekonomi och att dra nödvändiga slutsatser för att förebygga och svara på liknande extrema situationer inom EU i framtiden.
27.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen och till medlemsstaternas regeringar och parlament.
P6_TA(2007)0443
Utnyttjande av Europeiska fonden för justering för globaliseringseffekter
A6-0378/2007
Europaparlamentets resolution av den 23 oktober 2007 om förslaget till Europaparlamentets och rådets beslut om utnyttjande av Europeiska fonden för justering för globaliseringseffekter med tillämpning av punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning ( KOM(2007)0415 – C6-0323/2007 – 2007/2168(ACI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2007)0415 – C6-0323/2007 ),
–
med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning EUT C 139, 14.6.2006, s.
1.
, särskilt punkt 28,
–
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1927/2006 av den 20 december 2006 om upprättande av Europeiska fonden för justering för globaliseringseffekter EUT L 406, 30.12.2006, s.
1.
,
–
med beaktande av resultaten av trepartsöverläggningarna den 6 juli 2007 och budgetförlikningen den 13 juli 2007,
–
med beaktande av betänkandet från budgetutskottet och yttrandet från utskottet för sysselsättning och sociala frågor ( A6-0378/2007 ), och av följande skäl:
A.
Europeiska unionen har inrättat lämpliga lagstiftningsinstrument och budgetinstrument för att kunna ge kompletterande stöd till arbetstagare som sagts upp och som drabbats av effekterna av större strukturella förändringar i världshandelsmönstren, för att underlätta deras återanpassning på arbetsmarknaden.
B.
Europeiska unionens ekonomiska stöd till arbetstagare som sagts upp bör vara dynamiskt och ställas till förfogande så snabbt och effektivt som möjligt.
C.
.
1.
Europaparlamentet uppmanar de berörda institutionerna att vidta de åtgärder som krävs för att fonden snarast skall kunna tas i anspråk.
2.
Europaparlamentet godkänner det bifogade beslutet.
3.
4.
Europaparlamentet uppdrar åt talmannen att översända denna resolution, inklusive bilagan, till rådet och kommissionen.
BILAGA
EUROPAPARLAMENTETS OCH RÅDETS BESLUT
av den 23 oktober 2007
om utnyttjande av Europeiska fonden för justering för globaliseringseffekter med tillämpning av punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning EUT C 139, 14.6.2006, s.
1.
, särskilt punkt 28,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1927/2006 av den 20 december 2006 om upprättande av Europeiska fonden för justering för globaliseringseffekter EUT L 406, 30.12.2006, s.
1.
,
med beaktande av kommissionens förslag,
och av följande skäl:
(1)
Europeiska unionen har inrättat Europeiska fonden för justering för globaliseringseffekter ("fonden") för att erbjuda ytterligare stöd till uppsagda arbetstagare som drabbats av större strukturförändringar i de världshandelsmönstren och att stödja dem i deras återintegrering på arbetsmarknaden.
(2)
Det interinstitutionella avtalet av den 17 maj 2006 gör det möjligt att utnyttja medel från fonden inom det årliga taket på 500 miljoner EUR.
(3)
Förordning (EG) nr 1927/2006 innehåller bestämmelser för att utnyttja fonden.
(4)
Frankrike har ansökt om medel från fonden med anledning av två fall som gäller uppsägningar inom bilsektorn: Peugeot SA och Renault SA.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Europeiska unionens allmänna budget för 2007 ska ett totalt belopp om 3 816 280 belasta rubriken Europeiska fonden för justering för globaliseringseffekter.
Artikel 2
Detta beslut skall offentliggöras i
Europeiska unionens officiella tidning
.
Utfärdat i Strasbourg den 23 oktober 2007
P6_TA(2007)0631
Kvinnors rättigheter i Saudiarabien
B6-0526 , 0530 , 0534 , 0537 , 0539 och 0540/2007
Europaparlamentets resolution av den 13 december 2007 om kvinnors rättigheter i Saudiarabien
Europaparlamentet utfärdar denna resolution
–
med beaktande av att Saudiarabien ratificerade FN:s konvention om avskaffande av all slags diskriminering av kvinnor den 7 september 2000,
–
med beaktande av FN:s konvention mot tortyr och annan grym, omänsklig eller förnedrande behandling eller bestraffning, som Saudiarabien ratificerade den 23 september 1997,
–
med beaktande av att Saudiarabien är en signatärstat till konventionen om barnets rättigheter sedan den 26 januari 1996,
–
med beaktande av att Saudiarabien valdes in i FN:s nya människorättsråd i maj 2006,
–
med beaktande av sina tidigare resolutioner om Saudiarabien av den 18 januari 1996 EUT C 32, 5.2.1996, s.
98.
,
–
A.
Kvinnor i Saudiarabien utsätts alltjämt för många olika former av diskriminering i det privata och offentliga livet, drabbas ofta av sexuellt våld och möter enorma hinder i det straffrättsliga systemet.
B.
I oktober 2006 dömdes en 19-årig kvinna, känd som "Qatif-flickan", till 90 piskrapp efter en incident där hon befann sig ensam i en bil och samtalade med en man som inte var en nära anhörig, när hon plötsligt attackerades och utsattes för gruppvåldtäkt.
C.
Det är djupt bekymmersamt att domstolen i Qatif (Saudiarabien) i november 2007 ändrade domen och dömde henne till sex månaders fängelse och 200 piskrapp.
D.
En tjänsteman vid domstolen i Qatif har uppgett att kvinnans straff skärptes på Högsta domstolens inrådan eftersom hon försökt kompromettera och påverka rättsväsendet via media.
E.
F.
G.
H.
Runt två miljoner kvinnliga migrerande arbetstagare är anställda som hemarbetare i Saudiarabien, där de ofta utsätts för övergrepp av statliga myndigheter och privata arbetsgivare, bland annat genom fysisk och psykisk misshandel, lön som inte betalas ut, frihetsberövande utan åtal eller rättegång och till och med dödsstraff efter orättvisa rättsliga förfaranden.
I.
Särskilt noterbara är fallen med Rizana Nafeek, en srilankesisk hemarbetare som i juni 2007 dömdes till döden eftersom ett spädbarn som hon hade hand om vid 17 års ålder hade dött, samt de indonesiska hemarbetarna Siti Tarwiyah Slamet och Susmiyati Abdul Fulan, som i augusti 2007 misshandlades till döds av den familj som de var anställda hos, samtidigt som två andra sårades svårt.
J.
Signatärstaterna till internationella konventioner om mänskliga rättigheter (exempelvis konventionen om avskaffande av all slags diskriminering av kvinnor) är skyldiga att garantera lika rättigheter för kvinnor och män.
1.
Europaparlamentet kräver att Saudiarabiens regering vidtar ytterligare åtgärder för att upphäva begränsningarna av kvinnors rättigheter, som deras rätt att röra sig fritt och köra bil, deras möjligheter att ta en anställning, deras rättskapacitet och deras rätt att företrädas i rättsprocesser, samt att avskaffa all slags diskriminering av kvinnor i det privata och offentliga livet och främja deras deltagande i den ekonomiska, sociala och politiska sfären.
2.
Europaparlamentet beklagar det ovannämnda beslutet av domstolen i Qatif att straffa våldtäktsoffret och uppmanar de saudiska myndigheterna att upphäva domen och lägga ner alla anklagelser mot våldtäktsoffret.
3.
4.
Europaparlamentet anser att en medvetandehöjande kampanj om våld mot kvinnor i Saudiarabien, framför allt våld i hemmet, vore ett lika välkommet som brådskande initiativ.
5.
Europaparlamentet uppmanar myndigheterna att se över och tillämpa nationell arbetsrättslig lagstiftning för att ge hemarbetare samma skydd som arbetstagare i andra branscher och se till att det väcks åtal mot arbetsgivare som gör sig skyldiga till sexuella eller fysiska övergrepp eller arbetsrättsliga övergrepp som strider mot gällande nationell lagstiftning.
6.
Europaparlamentet uppmanar Saudiarabiens regering att se över alla mål mot minderåriga gärningsmän som dömts till döden, avskaffa dödstraffet för minderåriga gärningsmän samt införa ett moratorium för dödsstraff.
7.
Europaparlamentet uppmanar rådet och kommissionen att ta upp dessa frågor vid ministermötet i det gemensamma rådet mellan EU och Gulfstaternas samarbetsråd.
8.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, FN:s generalsekretariat, Saudiarabiens regering, generalsekreteraren för Islamiska konferensen samt generalsekreteraren för Gulfstaternas samarbetsråd.
P6_TA(2008)0023
Situationen i Egypten
B6-0023 , 0029 , 0032 , 0036 , 0039 och 0042/2008
Europaparlamentets resolution av den 17 januari 2008 om situationen i Egypten
Europaparlamentet utfärdar denna resolution
–
med beaktande av sina tidigare resolutioner om Europa–Medelhavspartnerskapet,
–
med beaktande av sin resolution av den 15 november 2007 om allvarliga händelser som äventyrar kristna samfunds och andra religiösa samfunds existens Antagna texter, P6_TA(2007)0542 .
,
–
med beaktande av Barcelonaförklaringen från november 1995,
–
med beaktande av kommissionens meddelande till rådet och Europaparlamentet av den 21 maj 2003 om stärkande av EU:s åtgärder för mänskliga rättigheter och demokratisering i samarbete med Medelhavsparterna – Strategiska riktlinjer ( KOM(2003)0294 ),
–
med beaktande av den första konferensen som anordnades av Europa–Medelhavsnätverket för mänskliga rättigheter i Kairo den 26 och 27 januari 2006,
–
med beaktande av FN-konventionen mot tortyr, grym omänsklig eller förnedrande behandling eller bestraffning från 1984,
–
med beaktande av EU:s riktlinjer om försvarare av mänskliga rättigheter,
–
med beaktande av artikel 19 i FN:s internationella konvention om medborgerliga och politiska rättigheter, som Egypten ratificerade 1982,
–
med beaktande av den internationella konventionen om avskaffande av all slags diskriminering av kvinnor,
–
med beaktande av det arbetsprogram som godkändes vid toppmötet mellan stats- och regeringscheferna i Barcelona i november 2005,
–
med beaktande av de slutsatser som antogs i Barcelona den 26 november 2005, vid den femte europeiska parlamentsordförandekonferensen,
–
med beaktande av de resolutioner som antogs vid sammanträdet för den parlamentariska församlingen för Europa–Medelhavet den 27 mars 2006 och det uttalande som församlingens ordförande gjorde,
–
med beaktande av sin resolution av den 19 januari 2006 om den europeiska grannskapspolitiken EUT C 287 E, 24.11.2006, s.
312.
,
–
A.
B.
C.
D.
De egyptiska myndigheterna har lovat att sätta stopp för fängslandet av journalister, men hittills har man inte uppfyllt detta löfte.
E.
Oppositionens presidentkandidat Ayman Nour avtjänar fortfarande det femåriga fängelsestraff som 2005 utdömdes efter en orättvis rättegång till följd av ett politiskt motiverat åtal, och hans hälsa blir allt sämre på grund av denna fängelsevistelse.
F.
G.
Kopterna, bahaierna, shiiterna, koranisterna och medlemmar av andra religiösa minoriteter lider fortfarande allvarliga nackdelar på grund av sekterisk isolering som innebär en beklaglig begränsning för dem.
1.
2.
3.
Europaparlamentet uppmanar den egyptiska regeringen att upphöra med alla former av trakasserier, inklusive rättsliga åtgärder, mot och gripanden av mediaarbetare samt människorättsförsvarare och aktivister i allmänhet som begär reformer, och att fullt ut respektera yttrandefriheten i enlighet med artikel 19 i FN:s internationella konvention om medborgerliga och politiska rättigheter.
4.
5.
6.
7.
8.
9.
10.
Europaparlamentet välkomnar Egyptens ansträngningar för att garantera säkerheten vid gränsen till Gaza, och uppmanar samtliga berörda parter att intensifiera kampen mot smuggling genom tunnlar in till Gazaremsan.
11.
12.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till Egyptens regering och parlament, kommissionen, regeringarna och parlamenten i medlemsstaterna och i de Medelhavsländer som undertecknat Barcelonadeklarationen samt till talmannen i den parlamentariska församlingen för Europa–Medelhavsområdet samt till rådet och kommissionen.
P6_TA(2008)0027
Statistik över vattenbruket ***I
A6-0001/2008
Europaparlamentets lagstiftningsresolution av den 31 januari 2008 om förslaget till Europaparlamentets och rådets förordning om inlämning av statistik över vattenbruket från medlemsstaterna ( KOM(2006)0864 – C6-0005/2007 – 2006/0286(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2006)0864 ),
–
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från fiskeriutskottet ( A6-0001/2008 ).
1.
Europaparlamentet godkänner kommissionens förslag såsom ändrat av parlamentet.
2.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om kommissionen har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
3.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
P6_TC1-COD(2006)0286
Europaparlamentets ståndpunkt fastställd vid första behandlingen den 31 januari 2008 inför antagandet av Europaparlamentets och rådets förordning (EG) nr .../2008 om inlämning av statistik över vattenbruket från medlemsstaterna och om upphävande av rådets förordning (EG) nr 788/96
(Eftersom det nåddes en överenskommelse mellan parlamentet och rådet, motsvarar parlamentets ståndpunkt vid första behandlingen den slutliga rättsakten, förordning (EG) nr .../2008.)
P6_TA(2008)0039
Installation av belysnings- och ljussignalanordningar på jordbruks- och skogsbrukstraktorer med hjul (kodifierad version) ***I
A6-0022/2008
Europaparlamentets lagstiftningsresolution av den 19 februari 2008 om förslaget till Europaparlamentets och rådets direktiv om installationen av belysnings- och ljussignalanordningar på jordbruks- och skogsbrukstraktorer med hjul (kodifierad version) ( KOM(2007)0192 – C6-0108/2007 – 2007/0066(COD) )
(Medbeslutandeförfarandet – kodifiering)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2007)0192 ),
–
med beaktande av artiklarna 251.2 och 95 i EG-fördraget, i enlighet med vilka kommissionen har lagt fram sitt förslag ( C6-0108/2007 ),
2.
,
–
med beaktande av artiklarna 80 och 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för rättsliga frågor ( A6-0022/2008 ).
1.
Europaparlamentet godkänner kommissionens förslag såsom anpassat till rekommendationerna från den rådgivande gruppen för de juridiska avdelningarna vid Europaparlamentet, rådet och kommissionen.
2.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
P6_TA(2008)0116
Stöd till små och medelstora företag som bedriver forskning och utveckling ***I
A6-0064/2008
Europaparlamentets lagstiftningsresolution av den 10 april 2008 om förslaget till Europaparlamentets och rådets beslut om gemenskapens deltagande i ett forsknings- och utvecklingsprogram som syftar till att stödja små och medelstora företag som bedriver forskning och utveckling och som inletts av flera medlemsstater ( KOM(2007)0514 – C6-0281/2007 – 2007/0188(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2007)0514 ),
–
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för industrifrågor, forskning och energi ( A6-0064/2008 ).
1.
Europaparlamentet godkänner kommissionens förslag såsom ändrat av parlamentet.
2.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om kommissionen har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
3.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
P6_TC1-COD(2007)0188
(Eftersom det nåddes en överenskommelse mellan parlamentet och rådet, motsvarar parlamentets ståndpunkt vid första behandlingen den slutliga rättsakten, beslut nr .../2008/EG.)
P6_TA(2008)0149
Ansvarsfrihet 2006: Europeiska byrån för återuppbyggnad
A6-0112/2008
1.
Europaparlamentets beslut av den 22 april 2008 om ansvarsfrihet för genomförandet av budgeten för Europeiska byrån för återuppbyggnad för budgetåret 2006 ( C6-0373/2007 – 2007/2048(DEC) )
Europaparlamentet fattar detta beslut
–
med beaktande av den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad för budgetåret 2006 EUT C 261, 31.10.2007, s.
13.
,
–
med beaktande av revisionsrättens rapport om den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad för budgetåret 2006, samt byråns svar EUT C 309, 19.12.2007, s.
40.
,
–
med beaktande av rådets rekommendation av den 12 februari 2008 (5843/2008 – C6-0084/2008 ),
–
med beaktande av EG-fördraget, särskilt artikel 276,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
Förordningen senast ändrad genom förordning (EG) nr 1525/2007 (EUT L 343, 27.12.2007, s.
9).
, särskilt artikel 185,
–
med beaktande av rådets förordning (EG) nr 2667/2000 av den 5 december 2000 om Europeiska byrån för återuppbyggnad EGT L 306, 7.12.2000, s.
7.
Förordningen senast ändrad genom förordning (EG) nr 1756/2006 (EUT L 332, 30.11.2006, s.
18).
, särskilt artikel 8,
–
med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002 EGT L 357, 31.12.2002, s.
72.
, särskilt artikel 94,
–
med beaktande av artikel 71 och bilaga V i arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för utrikesfrågor ( A6-0112/2008 ).
1.
Europaparlamentet beviljar ansvarsfrihet för den verkställande direktören för Europeiska byrån för återuppbyggnad avseende genomförandet av byråns budget för budgetåret 2006.
2.
Europaparlamentet redovisar sina iakttagelser i resolutionen nedan.
3.
Europaparlamentet uppdrar åt talmannen att översända detta beslut och den resolution som utgör en del av beslutet till direktören för Europeiska byrån för återuppbyggnad, rådet, kommissionen och revisionsrätten samt att se till att de offentliggörs i Europeiska unionens officiella tidning (L-serien).
2.
Europaparlamentets beslut av den 22 april 2008 om avslutande av räkenskaperna för Europeiska byrån för återupbyggnad för budgetåret 2006 ( C6-0373/2007 – 2007/2048(DEC) )
Europaparlamentet fattar detta beslut
–
med beaktande av den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad för budgetåret 2006 EUT C 261, 31.10.2007, s.
13.
,
–
med beaktande av revisionsrättens rapport om den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad för budgetåret 2006, samt byråns svar EUT C 309, 19.12.2007, s.
40.
,
–
med beaktande av rådets rekommendation av den 12 februari 2008 (5843/2008 – C6-0084/2008 ),
–
med beaktande av EG-fördraget, särskilt artikel 276,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
Förordningen senast ändrad genom förordning (EG) nr 1525/2007 (EUT L 343, 27.12.2007, s.
9).
, särskilt artikel 185,
–
med beaktande av rådets förordning (EG) nr 2667/2000 av den 5 december 2000 om Europeiska byrån för återuppbyggnad EGT L 306, 7.12.2000, s.
7.
Förordningen senast ändrad genom förordning (EG) nr 1756/2006 (EUT L 332, 30.11.2006, s.
18).
, särskilt artikel 8,
–
med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002 EGT L 357, 31.12.2002, s.
72.
, särskilt artikel 94,
–
med beaktande av artikel 71 och bilaga V i arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för utrikesfrågor ( A6-0112/2008 ).
1.
Europaparlamentet konstaterar att den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad är den som bifogats revisionsrättens årsrapport.
2.
Europaparlamentet godkänner avslutandet av räkenskaperna för Europeiska byrån för återuppbyggnad för budgetåret 2006.
3.
Europaparlamentet uppdrar åt talmannen att översända detta beslut till den verkställande direktören för Europeiska byrån för återuppbyggnad, rådet, kommissionen och revisionsrätten samt att se till att det offentliggörs i Europeiska unionens officiella tidning (L-serien).
3.
Europaparlamentets resolution av den 22 april 2008 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska byrån för återuppbyggnad för budgetåret 2006 ( C6-0373/2007 – 2007/2048(DEC) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad för budgetåret 2006 EUT C 261, 31.10.2007, s.
13.
,
–
med beaktande av revisionsrättens rapport om den slutliga årsredovisningen för Europeiska byrån för återuppbyggnad för budgetåret 2006, samt byråns svar EUT C 309, 19.12.2007, s.
40.
,
–
med beaktande av rådets rekommendation av den 12 februari 2008 (5843/2008 – C6-0084/2008 ),
–
med beaktande av EG-fördraget, särskilt artikel 276,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
Förordningen senast ändrad genom förordning (EG) nr 1525/2007 (EUT L 343, 27.12.2007, s.
9).
, särskilt artikel 185,
–
med beaktande av rådets förordning (EG) nr 2667/2000 av den 5 december 2000 om Europeiska byrån för återuppbyggnad EGT L 306, 7.12.2000, s.
7.
Förordningen senast ändrad genom förordning (EG) nr 1756/2006 (EUT L 332, 30.11.2006, s.
18).
, särskilt artikel 8,
–
med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002 EGT L 357, 31.12.2002, s.
72.
, särskilt artikel 94,
–
med beaktande av artikel 71 och bilaga V i arbetsordningen,
–
A.
Revisionsrätten har förklarat att den har uppnått en rimlig säkerhet om att räkenskaperna för budgetåret är tillförlitliga och att de underliggande transaktionerna är lagliga och korrekta.
B.
Den 24 april 2007 beviljade Europaparlamentet direktören för Europeiska byrån för återuppbyggnad ansvarsfrihet för genomförandet av detta organs budget för budgetåret 2005 EUT L 187, 15.7.2008, s.
182.
, och i sin resolution som åtföljde beslutet om ansvarsfrihet framförde parlamentet bland annat följande synpunkter:
–
–
Europaparlamentet noterade att revisionsrätten i sin rapport för 2004 hade upptäckt, i samband med en genomgång av de verksamheter som överlåtits på Förenta nationernas övergångsförvaltning i Kosovo (UNMIK), att byrån inte utövade vederbörlig finansiell kontroll vid betalningar och att den hade stora svårigheter när den skulle avsluta verksamheterna, främst på grund av att bokföringen för projekten var bristfällig och att utgifterna inte var tillräckligt styrkta.
Allmänna punkter som rör övergripande frågor för de decentraliserade EU-organen och som därmed också är av betydelse för varje enskilt organs ansvarsfrihetsförfarande
1.
Europaparlamentet noterar att totalbudgeten för de 24 byråer och satellitorgan som revisionsrätten granskat uppgick till 1 080,5 miljoner EUR 2006 (där den största är Europeiska byrån för återuppbyggnad med 271 miljoner EUR och den minsta är Europeiska polisakademien (Cepol) med 5 miljoner EUR).
2.
Europaparlamentet påpekar att de externa EU-organ som nu är föremål för revision och ansvarsfrihet inte bara omfattar traditionella tillsynsmyndigheter utan också genomförandeorgan som inrättats för att genomföra enskilda program och inom en snar framtid även kommer att omfatta gemensamma företag som inrättats som offentlig-privata partnerskap (gemensamma teknikinitiativ).
3.
Europaparlamentet noterar att antalet organ som är föremål för ansvarsfrihetsförfarandet från parlamentets sida har utvecklats enligt följande: Budgetåret 2000: 8, 2001: 10, 2002: 11, 2003: 14, 2004: 14, 2005: 16, 2006: 20 tillsynsmyndigheter och 2 genomförandeorgan (förutom 2 organ som visserligen granskas av revisionsrätten men som blir föremål för ett internt ansvarsfrihetsförfarande).
4.
Principiella överväganden
5.
Europaparlamentet begär att kommissionen ska ge tydliga förklaringar för följande faktorer innan ett nytt organ inrättas eller ett befintligt organ reformeras: typ av organ, organets mål, interna styrstrukturer, produkter, tjänster, huvudsakliga förfaranden, målgrupp, kunder och intressenter, formella relationer med externa aktörer, budgetansvar, ekonomisk planering och personal- och rekryteringspolitik.
6.
Europaparlamentet begär att varje organ ska styras av ett årligt prestationsavtal som formuleras av organet och det ansvariga generaldirektoratet och som ska innehålla de huvudsakliga målsättningarna för det kommande året med en finansieringsram och klara indikatorer för att mäta prestationerna.
7.
Detta bör inte begränsas till traditionella delar som ekonomisk förvaltning och korrekt användning av offentliga medel utan bör också omfatta administrativ effektivitet och ändamålsenlighet och bör inkludera en värdering av den ekonomiska förvaltningen för vart och ett av organen.
8.
9.
10.
11.
12.
13.
Framläggande av redovisningsuppgifter
14.
15.
Europaparlamentet noterar att kommissionens gällande instruktioner för verksamhetsrapporter inte uttryckligen kräver att organet ska utarbeta en revisionsförklaring, men många direktörer har ändå gjort det för 2006, och i ett fall med en mycket viktig reservation.
16.
Europaparlamentet påminner om punkt 41 i sin resolution av den 12 april 2005 Europaparlamentets resolution innehållande iakttagelser som åtföljer beslutet om ansvarsfrihet för direktören för Europeiska byrån för återuppbyggnad med avseende på genomförandet av byråns budget för budgetåret 2003 (EUT L 196, 27.7.2005, s.
61).
där organens direktörer uppmanas att hädanefter låta deras verksamhetsrapporter, som läggs fram tillsammans med ekonomiska och administrativa uppgifter, åtföljas av en revisionsförklaring om transaktionernas laglighet och korrekthet, liknande de förklaringar som undertecknas av kommissionens generaldirektörer.
17.
Europaparlamentet uppmanar kommissionen att ändra sina gällande instruktioner till organen i enlighet härmed.
18.
Europaparlamentet föreslår dessutom att kommissionen ska arbeta med organen för att skapa en harmoniserad modell som gäller för alla byråer och satellitorgan och där det görs en tydlig åtskillnad mellan
–
en årsrapport, som riktas till en allmän läsekrets, om organets verksamhet, arbete och resultat,
–
en ekonomisk årsredovisning och en rapport om genomförandet av budgeten,
–
en verksamhetsrapport liknande den som kommissionens generaldirektörer lämnar,
–
en revisionsförklaring som undertecknats av organets direktör, med reservationer och iakttagelser som denne anser att den ansvarsfrihetsbeviljande myndigheten lämpligen bör uppmärksamma.
Allmänna iakttagelser från revisionsrätten
19.
Europaparlamentet noterar revisionsrättens iakttagelser (punkt 10.29 i årsrapporten EUT C 273, 15.11.2007, s.
1.
) att kommissionens utbetalningar av bidrag från gemenskapsbudgeten inte bygger på tillräckligt motiverade uppskattningar av byråernas behov av likvida medel.
20.
Europaparlamentet noterar att i slutet av 2006 hade 14 byråer ännu inte infört redovisningssystemet ABAC (fotnot till punkt 10.31 i årsrapporten).
21.
Internrevision
22.
Internrevisorn rapporterar till varje organs styrelse och direktör.
23.
Europaparlamentet uppmärksammar följande reservation i internrevisorns verksamhetsrapport för 2006:
På grund av personalbrist är kommissionens internrevisor inte i stånd att ordentligt uppfylla den funktion som internrevisor för gemenskapens decentraliserade organ som denne ges i artikel 185 i budgetförordningen.
24.
Europaparlamentet noterar dock internrevisorns anmärkning i dennes verksamhetsrapport för 2006 att från och med 2007 har internrevisionsenheten fått extra personalresurser från kommissionen och alla tillsynsmyndigheter kommer att bli föremål för internrevision på årlig basis.
25.
26.
27.
När det gäller den interna revisionskapaciteten, särskilt i förhållande till mindre organ, noterar Europaparlamentet det förslag som internrevisorn gjorde inför parlamentets ansvariga utskott den 14 september 2006 om att mindre organ ska tillåtas att köpa in interrevisionstjänster från den privata sektorn.
Utvärdering av organ
28.
Europaparlamentet påminner om det gemensamma uttalandet från parlamentet, rådet och kommissionen Rådsdokument DS 605/1/07 Rev1.
som förhandlades fram vid medlingen inför Ekofinrådets budgetmöte den 13 juli 2007 där man efterlyser i) en förteckning på organ som kommissionen avser att utvärdera och xii) en förteckning på de organ som redan utvärderats, tillsammans med en sammanfattning av resultaten.
Disciplinära förfaranden
29.
Organen uppmanas att överväga att inrätta en gemensam disciplinnämnd för organen.
Förslag till interinstitutionellt avtal
30.
I den sammanfattande rapporten om kommissionens förvaltning 2006 (punkt 3.1, KOM(2007)0274 ) sägs att förhandlingarna sedermera avbröts, men att diskussioner om innehållet återupptogs i rådet i slutet av 2006.
31.
Europaparlamentet välkomnar därför kommissionens åtagande att lägga fram ett meddelande om framtiden för EU:s tillsynsmyndigheter under loppet av 2008.
Självfinansierade organ
32.
—
Kontoret för harmonisering inom den inre marknaden har likvida medel på 281 miljoner EUR Källa: Rapport om årsredovisningen för Kontoret för harmonisering inom den inre marknaden (varumärken och mönster) för budgetåret 2006 samt kontorets svar (EUT C 309, 19.12.2007, s.
141).
.
—
Gemenskapens växtsortsmyndighet har likvida medel på 18 miljoner EUR Källa: Rapport om årsredovisningen för Gemenskapens växtsortsmyndighet för budgetåret 2006 samt myndighetens svar (EUT C 309, 19.12.2007, s.
135).
.
Specifika punkter
33.
Europaparlamentet välkomnar byråns utmärkta bidrag till att utveckla och stärka stabiliteten i regionen genom sina olika program samt en sund förvaltning av programmet Cards.
34.
35.
I detta sammanhang upprepar Europaparlamentet sin begäran om att bli regelbundet informerat av kommissionen om överföringen av verksamheten från byrån till delegationerna.
36.
Europaparlamentet gratulerar byråns direktör och hans personal för det arbete som utförts under mycket svåra omständigheter och som i betydande grad har förbättrat bilden av EU och dess synlighet.
37.
Europaparlamentet anser att byrån inte bara har de system (logistik, IT och andra) för att snabbt genomföra stora stödinsatser i områden som genomgått konflikter utan också har visat prov på särskilt hög expertis och sakkunskap i återuppbyggnaden efter krig.
38.
39.
Europaparlamentet anser att ett nytt mandat för denna framgångsrika byrå skulle vara det effektivaste sättet att genomföra de nya uppgifter inom ramen för de externa åtgärderna som inte kan utföras av kommissionens avdelningar i Bryssel eller av kommissionens delegationer.
40.
41.
Europaparlamentet noterar revisionsrättens iakttagelse när det gäller budgetåret 2006 att även om genomförandegraden när det gäller budgeten var tillfredsställande, måste dock byrån uppmärksammas på den nivå av åtaganden som ännu ska ingås, vilket kommer att kräva särskild övervakning av programmen med tanke på att byråns mandat upphör i slutet av 2008.
42.
Europaparlamentet konstaterar vidare att revisionsrätten noterade att redovisningssystemet och internkontrollsystemet hade förbättrats jämfört med de föregående åren, särskilt i fråga om övervakningen av medel som förvaltas av externa organ och av genomförandet av upphandlingsförfaranden.
43.
Europaparlamentet påminner om att byrån har den i särklass största budgeten (2006: 271 miljoner EUR) av de organ som är föremål för ansvarsfrihetsförfarandet.
44.
Europaparlamentet konstaterar emellertid från byråns räkenskaper att de anslag som överfördes till 2007 uppgick till sammanlagt 678 miljoner EUR.
45.
Europaparlamentet uppmanar kommissionen att informera parlamentets behöriga utskott hur återstoden av outnyttjade anslag vid utgången av byråns mandat skall hanteras.
46.
Europaparlamentet noterar att byråns direktör undertecknade en revisionsförklaring utan reservationer den 30 maj 2007.
47.
Europaparlamentet konstaterar att internrevisionsenheten i slutet av 2004 genomförde en granskning av effektiviteten och ändamålsenligheten vid byråns fem arbetsorter och att en serie åtgärder vidtogs under 2006 av byråns ledning för att ta itu med de frågor som internrevisionsenheten tagit upp.
48.
Europaparlamentet uppmanar kommissionen att ändra byråns mandat när detta utlöper 2008 och omvandla byrån till ett organ för genomförande av särskilda externa EU-åtgärder, framför allt i regioner som just genomgått en krissituation.
P6_TA(2008)0188
Punktskattesats för öl från Madeira *
A6-0146/2008
Europaparlamentets lagstiftningsresolution av den 8 maj 2008 om förslaget till rådets beslut om tillstånd för Portugal att tillämpa en nedsatt punktskattesats för öl som produceras lokalt i den autonoma regionen Madeira ( KOM(2007)0772 – C6-0012/2008 – 2007/0273(CNS) )
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till rådet ( KOM(2007)0772 ),
–
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för regional utveckling och yttrandet från utskottet för jordbruk och landsbygdens utveckling ( A6-0146/2008 ).
1.
Europaparlamentet godkänner kommissionens förslag.
2.
Rådet uppmanas att underrätta Europaparlamentet om rådet har för avsikt att avvika från den text som parlamentet har godkänt.
3.
Rådet uppmanas att på nytt höra Europaparlamentet om rådet har för avsikt att väsentligt ändra kommissionens förslag.
4.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
P6_TA(2008)0215
Straffrättsliga påföljder till skydd för miljön ***I
A6-0154/2008
Europaparlamentets lagstiftningsresolution av den 21 maj 2008 om förslaget till Europaparlamentets och rådets förordning om straffrättsliga påföljder till skydd för miljön ( KOM(2007)0051 – C6-0063/2007 – 2007/0022(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2007)0051 ),
–
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för rättsliga frågor och yttrandena från utskottet för miljö, folkhälsa och livsmedelssäkerhet och utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor ( A6-0154/2008 ).
1.
Europaparlamentet godkänner kommissionens förslag såsom ändrat av parlamentet.
2.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om kommissionen har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
3.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
P6_TC1-COD(2007)0022
Europaparlamentets ståndpunkt fastställd vid första behandlingen den 21 maj 2008 inför antagandet av Europaparlamentets och rådets direktiv 2008/.../EG om skydd för miljön genom straffrättsliga bestämmelser
P6_TA(2008)0292
Saknade personer i Cypern - Uppföljning (artikel 131 i arbetsordningen)
A6-0139/2008
Europaparlamentets resolution av den 18 juni 2008 om saknade personer i Cypern – Uppföljning av Europaparlamentets resolution av den 15 mars 2007 ( 2007/2280(INI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av sin resolution av den 15 mars 2007 om saknade personer i Cypern EUT C 301 E, 13.12.2007, s.
243.
,
–
med beaktande av relevanta rapporter från FN:s generalsekreterare Särskilt den senaste om FN:s insats på Cypern (S/2008/353), kapitel IV.
och resolutioner från FN:s säkerhetsråd Särskilt resolution 1818(2008) av den 13 juni 2008.
och de internationella initiativ som tagits för att utreda vad som har hänt med de saknade personerna i Cypern Kommittén för saknade personer i Cypern: http://www.cmp-cyprus.org
,
–
med beaktande av avgörandena från Europeiska domstolen för de mänskliga rättigheterna (Europadomstolen) av den 10 maj 2001 Cypern mot Turkiet, nr 25781/94, ECHR 2001-IV.
och den 10 januari 2008 Varnava m.fl. mot Turkiet , nr 16064/90, 16065/90,16066/90, 16068/90, 16069/90, 16070/90, 16071/90, 16072/90 och 16073/90 (överklagande väntar på avgörande).
beträffande saknade personer i Cypern,
–
med beaktande av artikel 45 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor ( A6-0139/2008 ), och av följande skäl:
A.
Det besök som parlamentets föredragande gjort hos kommittén för saknade personer, på uppgrävningsplatserna, på det antropologiska laboratoriet – i vars arbete båda befolkningsgrupper deltar – och hos saknade personers familjer i Cypern hade uteslutande i syfte att undersöka det humanitära problem med de saknade personerna (grekcyprioter och turkcyprioter) som är kopplat till de anhörigas rätt att få veta vad som har hänt dessa personer.
B.
C.
Kommittén för saknade personer i Cypern har gjort framsteg sedan 2004 när det gäller uppgrävning och identifiering av kvarlevor och visar beslutsamhet att gå vidare i syfte att uppnå resultat som kan uppnås endast om dess kapacitet ökas, särskilt på fältet.
D.
Kommitténs projekt för uppgrävning, identifiering och återbördande av kvarlevor efter saknade personer har pågått sedan augusti 2006, och hittills har kvarlevorna efter 398 personer grävts upp, varav 266 har analyserats vid kommitténs antropologiska laboratorium i ett försök att göra sannolika identifieringar.
E.
F.
De första säkra identifieringarna gjordes i slutet av juni 2007, och fram till i dag har 91 kvarlevor efter personer som grävts upp inom ramen för kommitténs projekt identifierats genom denna process.
G.
Det största enskilda bidraget till kommittén för saknade personer, 1,5 miljoner EUR, täcker endast perioden fram till slutet av 2008 och ingår i EU:s ekonomiska stöd till den turkcypriotiska befolkningsgruppen.
H.
Det konstruktiva samarbetet mellan grekcypriotiska och turkcypriotiska medlemmar av kommittén för saknade personer, liksom det goda samarbetet mellan de blandade grek- och turkcypriotiska arbetslagen, både i laboratoriet och på fältet bör noteras.
1.
Europaparlamentet uppmanar de berörda parterna att fortsätta det ärliga och uppriktiga samarbetet för att snabbt slutföra nödvändiga utredningar om vad som hänt alla personer som saknas i Cypern och att ge full verkan åt avgörandet från Europadomstolen av den 10 maj 2001.
2.
Europaparlamentet uppmanar de berörda parterna och alla dem som har eller kan få tillgång till uppgifter eller bevis från personlig kunskap, arkiv, rapporter från slagfält eller register från interneringsanläggningar att ställa dessa uppgifter eller bevis till förfogande för kommittén för saknade personer i syfte att hjälpa till att påskynda dess arbete.
3.
Europaparlamentet anser att ytterligare ekonomiskt stöd bör anslås till kommittén för saknade personer för åren från och med 2009 och att det är nödvändigt att avsätta ett tilläggsbelopp på 2 miljoner EUR i Europeiska unionens allmänna budget för 2009.
4.
Europaparlamentet uppmanar rådet och kommissionen att enas om detta ytterligare ekonomiska bistånd för 2009, inte bara för att medge fortsatt arbete, utan även för att öka kapaciteten, särskilt på fältet, och göra det möjligt att anställa fler forskare och anskaffa mer utrustning.
5.
Europaparlamentet uppmanar medlemsstaterna att fortsätta med sitt hittillsvarande stöd.
6.
Europaparlamentet uppmanar utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor att fortsätta att följa upp frågan om saknade personer i Cypern och att avlägga årliga rapporter.
7.
Europaparlamentet bemyndigar parlamentets föredragande och utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor att vidta alla tänkbara åtgärder för att förmå alla berörda parter att uppriktigt och aktivt medverka i arbetet att utreda vad som har hänt var och en av de saknade personerna.
8.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, FN:s generalsekreterare, regeringarna och parlamenten i Cypern, Turkiet, Grekland och Förenade kungariket och till kommittén för saknade personer i Cypern.
P6_TA(2008)0386
Vissa frågor som rör motorfordonsförsäkring
A6-0249/2008
Europaparlamentets resolution av den 2 september 2008 om vissa frågor som rör motorfordonsförsäkring ( 2007/2258(INI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens rapport om vissa frågor som rör motorfordonsförsäkring ( KOM(2007)0207 ) (kommissionens rapport),
–
med beaktande av Europaparlamentets och rådets direktiv 2000/26/EG av den 16 maj 2000 om tillnärmning av medlemsstaternas lagar om ansvarsförsäkring för motorfordon (fjärde direktivet om motorfordonsförsäkring) EGT L 181, 20.7.2000, s.
65.
,
–
med beaktande av artikel 45 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för den inre marknaden och konsumentskydd och yttrandet från utskottet för rättsliga frågor ( A6-0249/2008 ),
A.
Den fria rörligheten för personer i EU har särskilt i samband med de två senaste utvidgningsrundorna och den motsvarande utökningen av Schengengruppen resulterat i en snabb ökning av både antalet personer och fordon som rör sig över nationsgränserna både i arbetsrelaterat syfte och i privat syfte.
B.
Den prioriterade frågan att skydda olycksdrabbade personer kräver en tydlig, precis och verkningsfull lagstiftning på området för motorfordonsförsäkringar på EU-nivå.
C.
I det fjärde direktivet om motorfordonsförsäkring uppmanades kommissionen att till Europaparlamentet och rådet rapportera om genomförandet av och effektiviteten hos de nationella sanktioner som införts när det gäller förfarandet med motiverat ersättningsanbud/motiverat svar samt om överensstämmelsen mellan dessa, och att lägga fram förslag om detta ansågs nödvändigt.
D.
I kommissionens rapport granskas de nationella sanktionsbestämmelserna, effektiviteten avseende mekanismen med skaderegleringsrepresentanten och den rådande tillgången till frivillig rättsskyddsförsäkring, som kan tecknas av personer som kan drabbas av trafikolyckor.
E.
F.
G.
Det krävs fortfarande ett klargörande av hur denna bestämmelse fungerar.
H.
Kommissionen måste ta fullständig hänsyn till utvidgningen när den genomför EU:s politik, i synnerhet den förhållandevis höga kostnaden för motorfordonsförsäkringar i de nya medlemsstaterna.
I.
Olika sanktionsbestämmelser avseende förfarandet med motiverat ersättningsanbud/motiverat svar har tillämpats i medlemsstaterna.
J.
Samråd med nationella myndigheter, även i de nya medlemsstaterna, har bekräftat att de gällande sanktionsbestämmelserna, där sådana finns, är adekvata och att tillämpningen av dem är verkningsfull i hela EU.
K.
En del medlemsstater har dock inte infört några särskilda sanktioner, utan där gäller bara försäkringsbolagets skyldighet att betala lagstadgad ränta på ersättningsbeloppet om det motiverade ersättningsanbudet/motiverade svaret inte föreligger inom tre månader.
L.
Systemet med skaderegleringsrepresentanter är förhållandevis välkänt i de flesta medlemsstater.
M.
I kommissionens samråd för att bedöma medborgarnas kännedom om systemet med skaderegleringsrepresentanter deltog endast medlemsstaterna och försäkringsbranschen och man lyckades inte på ett lämpligt sätt engagera medborgarna och konsumentorganisationerna, dvs. de aktörer som är mest intresserade av att systemet fungerar ordentligt.
N.
O.
Frågan om sådana skäliga rättegångskostnader bör täckas av tredje parts ansvarsförsäkring för motorfordon i alla medlemsstater är fortfarande öppen.
P.
En ansvarsförsäkring för motorfordon som täcker rimliga rättegångskostnader i alla medlemsstater bidrar emellertid till ett bättre skydd av de europeiska konsumenterna och ett större förtroende från deras sida.
Q.
R.
Obligatorisk täckning av rättegångskostnader borde öka konsumenternas förtroende för tredje parts ansvarsförsäkring för motorfordon, särskilt i fall då man söker ersättning för rättegångskostnader, eftersom konsumenterna i många nya medlemsstater aktar sig för höga rättegångskostnader, som skulle täckas genom en obligatorisk försäkring.
S.
En obligatorisk rättsskyddsförsäkring skulle innebära en ytterligare och mer komplex arbetsbörda för rättsväsendet, vilket skulle kunna försena biläggandet av tvister och medföra en högre andel oberättigade ersättningsanspråk.
T.
Tredje parts ansvarsförsäkring för motorfordon och rättsskyddsförsäkringen har olika mål och funktioner genom att tredje parts ansvarsförsäkring för motorfordon gör det möjligt för konsumenterna att hantera kostnaden för alla ersättningsanspråk som riktas mot dem till följd av en vägtrafikolycka, medan rättsskyddsförsäkringen täcker rättegångskostnaderna i samband med ersättningskrav mot tredje part till följd av en vägtrafikolycka.
U.
Allmänna kampanjer från nationella myndigheter, försäkringsbranschen och konsumentorganisationer är viktiga för att de nationella marknaderna ska utvecklas.
1.
Europaparlamentet välkomnar kommissionens rapport och betonar vikten av att låta alla berörda parter, särskilt konsumenterna, delta fullt ut och effektivt i samrådsprocessen i samband med utvecklingen av EU:s politik på detta område.
2.
Europaparlamentet begär därför att i synnerhet konsumentorganisationer som företräder skadelidande systematiskt ska delta i utvärderingsprocessen avseende effektiviteten hos de rådande systemen i medlemsstaterna.
3.
Europaparlamentet välkomnar denna efterhandsutvärdering av lagstiftningsåtgärderna, där syftet är att se till att bestämmelserna fungerar som avsett och att belysa alla oförutsedda felaktiga tillämpningar.
4.
Europaparlamentet betonar vikten av att öka konsumenternas förtroende för motorfordonsförsäkringarna när det gäller gränsöverskridande resor med motorfordon inom EU, särskilt för bilister från de gamla medlemsstaterna som färdas till destinationer i de nya medlemsstaterna och vice versa.
5.
Europaparlamentet anser att främjandet av befintliga och marknadsdrivna lösningar som skyddar konsumenterna stärker konsumenternas förtroende för motorfordonsförsäkringen.
6.
Europaparlamentet anser att medlemsstaterna även har ett ansvar för att deras nationella försäkringssystem fungerar väl i förhållande till EU-lagstiftning om förfarandet med motiverat ersättningsanbud/motiverat svar och rättegångskostnader som bekostas av skadelidande.
7.
Europaparlamentet uppmanar kommissionen att fortsätta att nära övervaka marknadsmekanismernas effektivitet och att regelbundet rapportera till parlamentet om denna.
8.
9.
Europaparlamentet understryker att arbetsrelationerna mellan kommissionen, de nationella myndigheterna, försäkringsbranschen och konsumenterna bör stärkas för att garantera ett oavbrutet tillhandahållande av korrekta uppgifter om de rådande tillsynssystemen.
10.
Europaparlamentet anser, i linje med EU:s allmänt etablerade synsätt när det gäller sanktioner, att subsidiaritetsprincipen bör tillämpas och att det inte finns något behov av harmonisering av de nationella sanktionsbestämmelserna.
11.
Europaparlamentet finner att nationella tillsynsmyndigheter har bättre förutsättningar att garantera högsta möjliga konsumentskydd på sina nationella marknader.
12.
Europaparlamentet rekommenderar därför med avseende på förfarandet med motiverat ersättningsanbud/motiverat svar att medlemsstaterna tillåts avgöra vilka sanktioner som ska vidtas och vilken typ av bestämmelser som är lämplig.
13.
Europaparlamentet uppmanar medlemsstaterna att garantera att deras påföljder, om tidsfristen på tre månader för att lämna ett motiverat svar eller ett motiverat ersättningsanbud på en ersättningsansökan inte respekteras, är effektiva.
14.
15.
Europaparlamentet upprepar betydelsen av att öka medborgarnas förtroende för systemet med skaderegleringsrepresentanten genom att främja detta med hjälp av allmänna kampanjer och andra lämpliga åtgärder.
16.
Europaparlamentet uppmanar medlemsstaterna och kommissionen att öka konsumenternas förtroende genom att främja lämpliga åtgärder som ökar kännedomen om och användningen av nationella centrum för försäkringsinformation, t.ex. krav på att försäkringsbolagens avtalsinformation ska innehålla kontaktuppgifter till informationscentrumet i den aktuella medlemsstaten.
17.
Europaparlamentet uppmanar dessutom medlemsstaterna att kräva att försäkringsbolagen, som ett led i förhandsinformationen om försäkringsavtal, förser konsumenterna med heltäckande information om hur systemet med skaderegleringsrepresentanten fungerar och om dess nytta för försäkringstagarna.
18.
Europaparlamentet uppmanar kommissionen att fortsätta att övervaka systemets funktion och att samordna och hjälpa till då detta behövs eller då nationella myndigheter ber om hjälp.
19.
Europaparlamentet anser dessutom, i förbindelse med tredje parts ansvarsförsäkring för motorfordon, att obligatorisk täckning av rättegångskostnader tydligt skulle minska viljan att bilägga tvister utanför domstol och eventuellt öka antalet domstolsförfaranden, vilket skulle leda till en omotiverad ökning av arbetsbördan för rättsväsendet och riskera att destabilisera den befintliga och framväxande marknaden för frivilliga rättsskyddsförsäkringar.
20.
Europaparlamentet anser därför att de negativa effekterna av att införa ett system med obligatorisk täckning av rättegångskostnader i tredje parts ansvarsförsäkring för motorfordon skulle vara större än de potentiella fördelarna.
21.
Europaparlamentet uppmanar kommissionen att tillsammans med medlemsstaterna vidta de ytterligare åtgärder som är nödvändiga för att öka kännedomen om rättsskyddsförsäkringar och andra försäkringar, särskilt i de nya medlemsstaterna, och inrikta sig på att informera konsumenterna om fördelarna med endera typen av försäkringsskydd.
22.
Europaparlamentet anser att de nationella tillsynsmyndigheternas roll i detta sammanhang är avgörande för genomförandet av bästa metoder från andra medlemsstater.
23.
Europaparlamentet uppmanar därför kommissionen att stärka konsumentskyddet främst genom att uppmana medlemsstaterna att uppmuntra sina nationella tillsynsmyndigheter och nationella försäkringsbolag att öka kännedomen om frivilliga rättsskyddsförsäkringar.
24.
Europaparlamentet anser att förhandsinformation om motorfordonsförsäkring även skulle kunna innehålla uppgifter om möjligheten att teckna rättsskyddsförsäkring.
25.
Europaparlamentet uppmanar medlemsstaterna att be nationella tillsynsmyndigheter och mellanhänder att informera kunderna om möjliga risker och om kompletterande frivilliga försäkringar som kan vara till nytta för dem, som t.ex. rättsskyddsförsäkring, assistansskydd och stöldförsäkring.
26.
Europaparlamentet uppmanar de medlemsstater som inte har infört alternativa tvistlösningssystem i samband med ersättningskrav att överväga att införa sådana system grundade på bästa metoder i andra medlemsstater.
27.
Europaparlamentet begär att kommissionen inte föregriper resultatet av den utredning som beställts om olika skadeståndsnivåer vid personskada i samband med antagandet av Rom II-förordningen Europaparlamentets och rådets förordning (EG) nr 864/2007 av den 11 juli 2007 om tillämplig lag för utomobligatoriska förpliktelser (EUT L 199, 31.7.2007, s.
40).
, eftersom utredningen kan komma att föreslå en försäkringsbaserad lösning och därav följande ändring av det fjärde direktivet om motorfordonsförsäkring.
28.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet och kommissionen.
P6_TA(2008)0411
Statskupp i Mauretanien
B6-0386 , 0392 , 0397 , 0398 , 0408 och 0409/2008
Europaparlamentets resolution av den 4 september 2008 om statskuppen i Mauretanien
Europaparlamentet utfärdar denna resolution
–
med beaktande av de uttalanden som efter statskuppen gjordes av Europaparlamentets talman, rådets ordförandeskap, den höge representanten för den gemensamma utrikes- och säkerhetspolitiken, kommissionen, FN:s säkerhetsråd, Afrikanska unionen (AU), Västafrikanska staters ekonomiska gemenskap (Ecowas) och Internationella organisationen för fransktalande länder (OIF),
–
med beaktande av det andra Mauretanienbesöket sedan statskuppen av Saïd Djinnit, FN:s generalsekreterares särskilde representant för Västafrika,
–
med beaktande av AU:s grundakt, som fördömer varje försök till maktövertagande genom våld,
–
A.
Den 6 augusti 2008 ägde en statskupp rum i Mauretanien, då landets president Sidi Mohamed Ould Cheikh Abdallahi störtades från makten av en grupp högt uppsatta generaler som han hade avskedat tidigare samma dag.
B.
Parlamentsvalen i november och december 2006, senatsvalet i januari 2007 och presidentvalet i mars 2007, då Sidi Mohamed Ould Cheikh Abdallahi valdes till president, bedömdes som rättvisa och öppna av internationella observatörer, däribland EU:s egna observatörer och särskilt de observatörsgrupper som skickats av Europaparlamentet, som på så vis stått som garant för att dessa val gått rätt till.
C.
D.
E.
F.
Det är glädjande att framsteg gjorts i fråga om flyktingars återvändande och att en lag som förbjuder slaveri i landet har antagits.
G.
H.
I.
Ett demokratiskt Mauretanien skulle vara en stabiliserande faktor i en annars ytterst bräcklig region: här finns å ena sidan GSPC (Groupe salafiste pour la prédication et le combat), som håller till i Sahara vid den nordöstra gränsen till Algeriet och Mali och som har blivit muslimska Maghrebs al-Qaida, och å andra sidan tuaregrebellerna.
J.
Den "författningsorder" i vilken juntan fastställer sina befogenheter och genom vilken juntan kan styra med hjälp av dekret har ingen rättslig grund.
1.
2.
Europaparlamentet kräver ett omedelbart frigivande av president Mohamed Ould Cheikh Abdallahi, premiärminister Yahya Ould Ahmed el-Waghef och andra regeringsmedlemmar som alltjämt sitter i husarrest på olika håll i landet.
3.
Europaparlamentet kräver att presidentens och parlamentets författningsenliga befogenheter respekteras fullt ut, vilket innebär att samstyret mellan president och parlament och maktdelningen mellan den verkställande och lagstiftande makten måste regleras med respekt för och inom ramen för konstitutionen, som kan ändras av hänsyn till stabiliteten endast om detta sker i enlighet med just konstitutionen och detta efter en omfattande debatt med samtliga politiska krafter.
4.
Europaparlamentet anser att en ärlig och uppriktig debatt mellan de viktigaste politiska krafterna bör bestämma vilka konstitutionella medel och metoder som ska användas för att få slut på krisen.
5.
6.
Europaparlamentet begär att de flyktingar som återvänt till Mauretanien ska kunna hävda sina rättigheter genom att få tillbaka de tillgångar de blivit av med.
7.
Europaparlamentet framhåller att det mauretanska folket, som redan är mycket hårt prövat av den ekonomiska krisen och livsmedelskrisen, inte får användas som gisslan i den kris som nu uppstått, och parlamentet uppmanar kommissionen att genomföra projekt till stöd för det civila samhället inom ramen för det europeiska instrumentet för demokrati och mänskliga rättigheter.
8.
9.
Europaparlamentet stöder AU:s ansträngningar att låta förnuftet leda fram till en lösning på krisen.
10.
Europaparlamentet uppmanar kommissionen att föra en politisk dialog i enlighet med artikel 8 i partnerskapsavtalet mellan medlemmarna i gruppen av stater i Afrika, Västindien och Stillahavsområdet, å ena sidan, och Europeiska gemenskapen och dess medlemsstater, å andra sidan, undertecknat i Cotonou den 23 juni 2000 EGT L 317, 15.12.2000, s.
3.
11.
Europaparlamentet uppmanar rådets ordförandeskap att fortsatt följa den politiska situationen i landet på nära håll, i nära samarbete med Afrikanska unionen, och att garantera säkerheten för EU-medborgare.
12.
Europaparlamentet vill att det snarast möjligt skickas en parlamentsdelegation som ska träffa sina mauretanska motsvarigheter och erbjuda hjälp för att landet ska kunna ta sig ur krisen.
13.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen och medlemsstaternas regeringar samt Afrikanska unionens institutioner, Västafrikanska staters ekonomiska gemenskap, OIF och FN:s säkerhetsråd.
P6_TA(2008)0440
Förfaranden vid domstolen (ändring av artikel 121)
A6-0324/2008
Europaparlamentets beslut av den 24 september 2008 om att ändra artikel 121 i Europaparlamentets arbetsordning om förfaranden vid domstolen ( 2007/2266(REG) )
Europaparlamentet fattar detta beslut
–
med beaktande av skrivelsen från ordföranden för utskottet för rättsliga frågor av den 26 september 2007,
–
med beaktande av artiklarna 201 och 202 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för konstitutionella frågor ( A6-0324/2008 ).
1.
Europaparlamentet beslutar att införa nedanstående ändring i arbetsordningen.
2.
Europaparlamentet påminner om att ändringen träder i kraft den första dagen under nästa sammanträdesperiod.
3.
Europaparlamentet uppdrar åt talmannen att för kännedom översända detta beslut till rådet och kommissionen.
Nuvarande lydelse
1
Europaparlamentets arbetsordning
3a.
Talmannen ska efter att ha hört ansvarigt utskott avge yttranden eller agera på parlamentets vägnar i domstolsförfaranden.
Om talmannen avser att avvika från det ansvariga utskottets rekommendation ska han eller hon informera utskottet om detta samt hänskjuta frågan till talmanskonferensen med angivande av sina skäl.
Om talmanskonferensen anser att parlamentet undantagsvis inte bör inkomma med inlagor eller skriftliga yttranden till domstolen i mål där giltigheten av en rättsakt som parlamentet antagit ifrågasätts, ska ärendet utan dröjsmål föreläggas kammaren.
I brådskande fall får talmannen vidta förebyggande åtgärder för att den berörda domstolens tidsfrister ska respekteras.
I sådana fall ska det förfarande som anges i denna punkt genomföras så snart som möjligt.
Tolkning:
P6_TA(2008)0469
IASCF
B6-0450/2008
Europaparlamentets resolution av den 9 oktober 2008 om den översyn av IASB:s offentliga redovisningsskyldighet och sammansättning som genomförts av IASCF – Förslag till förändring
Europaparlamentet utfärdar denna resolution
–
med beaktande av rådets slutsatser av den 8 juli 2008, angående IASB:s (International Accounting Standards Board) styrning,
–
1
,
–
med beaktande av Europaparlamentets resolution av den 24 april 2008 om internationella redovisningsstandarder (IFRS) och styrningen av International Accounting Standards Board (IASB) Antagna texter, P6_TA(2008)0183 .
,
–
med beaktande av kommissionens förordning (EG) nr 1358/2007 av den 21 november 2007 om ändring av förordning (EG) nr 1725/2003 om antagande av vissa redovisningsstandarder i enlighet med Europaparlamentets och rådets förordning (EG) nr 1606/2002, med avseende på den internationella redovisningsstandarden IFRS 8 EUT L 304, 22.11.2007, s.
9.
om rapportering för operativa segment, och parlamentets resolution av den 14 november 2007 om utkastet till kommissionens förordning Antagna texter, P6_TA(2007)0526 .
,
–
med beaktande av Europaparlamentets resolution av den 14 november 2007 om om utkastet till kommissionens förordning om ändring av förordning (EG) nr 809/2004 i fråga om redovisningsstandarder som tillämpas vid utarbetandet av historisk information i prospekt och om utkastet till kommissionens beslut om användningen bland värdepappersemittenter i tredjeland av information som utarbetats enligt internationellt godkända redovisningsstandarder Antagna texter, P6_TA(2007)0527 .
,
–
med beaktande av Europaparlamentets resolution av den 24 oktober 2006 om redovisningsstandarder som används av emittenter i tredjeländer och deras överensstämmelse med IFRS-standarderna i enlighet med förslaget till genomförandeåtgärder avseende prospektdirektivet och direktivet om insynskrav EUT C 313 E, 20.12.2006, s.
116.
, där de villkor som EU har fastställt för att nå konvergens och överensstämmelse mellan IFRS-standarderna och de amerikanska GAAP-standarderna anges,
–
med beaktande av IASCF:s rapport från juli 2008 "Översyn av stadgan – IASB:s offentliga redovisningsskyldighet och sammansättning – Förslag till förändring",
–
med beaktande av i rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter EGT L 184, 17.7.1999, s.
23.
,
–
A.
EU kräver att emittenter tillämpar internationella redovisningsstandarder i sina koncernredovisningar.
1.
Europaparlamentet noterar att IASCF har föreslagit att man ska inrätta en övervakningsgrupp, och anser att denna övervakningsgrupp bör få rekommendera kandidater till förvaltare/ombud samt ansvara för godkännandet av de utvalda förvaltarna/ombuden efter en överenskommen nomineringsprocess.
2.
3.
Europaparlamentet tvivlar på att det är lämpligt att inrätta en övervakningsgrupp i detta läge, innan andra fasen av samrådsprocessen rörande förnyelsen av IASB:s styrning har tagit sin början, och utan någon klar uppfattning om vilken förbindelse som bör upprättas mellan övervakningsgruppen och IASCF i den senares stadga.
4.
a)
den ansvariga ledamoten från kommissionen,
b)
ordföranden för kommittén för tillväxtekonomier inom den internationella organisationen för börstillsynsmyndigheter (IOSCO),
c)
ordföranden för den tekniska kommittén inom IOSCO (eller dess vice ordförande eller IOSCO:s utsedde ordförande, när IOSCO:s tekniska kommitté leds av ordföranden för en av EU:s börstillsynsmyndigheter, ledamoten från Japans Financial Service Agency eller ordföranden för USA:s Securities and Exchange Commission (SEC)),
d)
ledamoten från Japans Financial Service Agency,
e)
ordföranden för USA:s SEC, och
f)
ordföranden för Baselkommittén för banktillsyn.
5.
Europaparlamentet beklagar att man inte blev rådfrågad om inrättandet av en internationell rådgivningsgrupp för redovisningsfrågor.
6.
7.
8.
9.
10.
Europaparlamentet efterlyser en avsiktsförklaring mellan Europaparlamentet, rådet och kommissionen, som definierar hur lagstiftarna ska kopplas till övervakningsgruppens arbete, om en sådan grupp inrättas på detta stadium.
11.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, Europeiska centralbanken och Europeiska värdepapperstillsynskommittén samt medlemsstaternas regeringar och parlament.
P6_TA(2008)0603
Överföring av försvarsprodukter ***I
A6-0410/2008
Europaparlamentets lagstiftningsresolution av den 16 december 2008 om förslaget till Europaparlamentets och rådets direktiv om förenkling av villkoren för överföring av försvarsmateriel inom gemenskapen ( KOM(2007)0765 – C6-0468/2007 – 2007/0279(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2007)0765 ),
–
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för den inre marknaden och konsumentskydd och yttrandena från utskottet för utrikesfrågor och utskottet för industrifrågor, forskning och energi ( A6-0410/2008 ).
1.
Europaparlamentet godkänner kommissionens förslag såsom ändrat av parlamentet.
2.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om kommissionen har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
3.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
P6_TC1-COD(2007)0279
Europaparlamentets ståndpunkt fastställd vid första behandlingen den 16 december 2008 inför antagandet av Europaparlamentets och rådets direktiv 2009/.../EG om förenkling av villkoren för överföring av försvarsrelaterade produkter inom gemenskapen
(Eftersom det nåddes en överenskommelse mellan parlamentet och rådet, motsvarar parlamentets ståndpunkt vid första behandlingen den slutliga rättsakten, direktiv 2009/43/EG.)
P6_TA(2008)0616
Gränsöverskridande uppföljning av trafikförseelser ***I
A6-0371/2008
Europaparlamentets lagstiftningsresolution av den 17 december 2008 om förslaget till Europaparlamentets och rådets direktiv om att underlätta gränsöverskridande uppföljning av trafikförseelser ( KOM(2008)0151 – C6-0149/2008 – 2008/0062(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2008)0151 ),
–
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för transport och turism och yttrandet från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor ( A6-0371/2008 ).
1.
Europaparlamentet godkänner kommissionens förslag såsom ändrat av parlamentet.
2.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om kommissionen har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
3.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
P6_TC1-COD(2008)0062
2009/.../EG
om att underlätta gränsöverskridande uppföljning av trafikförseelser
(Text av betydelse för EES)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
,
,
med beaktande av europeiska datatillsynsmannens yttrande
9.
,
i enlighet med förfarandet i artikel 251 i fördraget
Europaparlamentets ståndpunkt av den 17 december 2008.
, och
av följande skäl: (1)
Europeiska unionen arbetar för att förbättra vägtrafiksäkerheten i syfte att minska antalet dödsolyckor, personskador och materiella skador.
För att nå detta syfte är det viktigt att konsekvent följa upp trafikförseelser som sätter vägtrafiksäkerheten på spel och utdöma påföljder för dem.
(2)
(3)
För att uppnå detta bör ett system med gränsöverskridande informationsutbyte införas.
(4)
Ett sådant system är särskilt värdefullt i samband med trafikförseelser som konstateras med automatisk utrustning och där trafiksyndarens identitet inte omedelbart kan fastställas, till exempel vid fortkörning eller rödljuskörning.
Det kan också med fördel användas för att följa upp trafikförseelser i fall då ett fordon har stoppats och det är nödvändigt att kontrollera fordonets registreringsuppgifter.
Detta gäller särskilt vid rattfylleri.
(5)
Detta system bör omfatta de trafikförseelser som är av störst risk för vägtrafiksäkerheten och som klassificeras som förseelser i alla medlemsstaternas lagstiftning.
Det bör därför omfatta fortkörning, rattfylleri, bristande bältesanvändning och rödljuskörning.
Kommissionen kommer att fortsätta att övervaka utvecklingen i
Europeiska unionen
.
(6)
(7)
För att kontrollsystemet ska vara effektivt bör det omfatta alla led mellan upptäckten av en förseelse och avsändandet av ett meddelande om trafikförseelse (utifrån en förlaga) till innehavaren av registreringsbeviset för fordonet i fråga.
När väl ett slutligt beslut har antagits,
kan
av den 24 februari 2005
om tillämpning av principen om ömsesidigt erkännande på bötesstraff EUT L 76, 22.3.2005, s.
.
Då nämnda rambeslut inte kan tillämpas, t.ex. då besluten om påföljd inte hänför sig till en brottslig handling, bör likväl andra åtgärder för verkställande av påföljder säkerställa att påföljderna är effektiva.
Det bör införas en minimistandard för meddelanden om trafikförseelse, inbegripet svarsblanketterna, och tillämpas mer kompatibla metoder för att sända dem så att den gränsöverskridande uppföljningen blir mer pålitlig och effektiv.
(8)
gemenskapsnät
.
(9)
31.
.
När gärningsmannen underrättas om trafikförseelsen bör denne följaktligen informeras om sin rätt att tillgå, rätta och radera uppgifter och om hur länge uppgifterna högst kan lagras på laglig väg.
(10)
De uppgifter som samlas in inom ramen för detta direktiv lagras endast tillfälligt och de får under inga omständigheter användas för andra ändamål än för vad som är nödvändigt för uppföljning av trafikförseelser.
Kommissionen och medlemsstaterna bör därför säkerställa att behandlingen av personuppgifter och förvaltningen av gemenskapens elektroniska nät gör det möjligt att undvika att de insamlade uppgifterna används för andra ändamål än uttryckliga trafiksäkerhetsändamål.
(11)
När det gäller trafikkontroller bör medlemsstaterna harmonisera sina metoder så att deras praxis blir jämförbar på EU-nivå.
Miniminormer för kontrollförfaranden bör således utvecklas i varje medlemsstat.
(12)
Den tekniska utrustning som används för trafiksäkerhetskontroller bör också harmoniseras i framtiden för att säkerställa konvergens mellan medlemsstaternas kontrollåtgärder.
Kommissionen bör föreslå en sådan teknisk harmonisering i samband med den översyn som föreskrivs i artikel 14
.
(13)
Kommissionen och medlemsstaterna bör vidta alla nödvändiga åtgärder för att informera och göra EU-medborgarna medvetna om genomförandet av detta direktiv.
Lämplig information om följderna av att bryta mot trafiksäkerhetsreglerna kan således ha en avskräckande effekt och därmed förhindra att trafikförseelser begås.
(14)
Kommissionen bör i framtiden inrikta sig på att underlätta gränsöverskridande uppföljning av trafikförseelser, särskilt när det gäller allvarliga trafikolyckor.
(15)
De åtgärder som är nödvändiga för att genomföra detta direktiv bör vidtas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter EGT L 184, 17.7.1999, s.
23. ║
.
(16)
(17)
dess
kan
gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget.
I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå
detta mål
.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
KAPITEL I
1.
Genom detta direktiv införs ett system för att underlätta gränsöverskridande uppföljning av följande trafikförseelser:
a)
Fortkörning
b)
Rattfylleri
c)
Bristande bältesanvändning
d)
Rödljuskörning
2.
I detta direktiv avses med
a)
"innehavare": den person som innehar registreringsbevis för fordonet i fråga
, inbegripet för motorcyklar
,
b)
"landet där förseelsen begicks": den medlemsstat där trafikförseelsen ägde rum,
c)
"bosättningsland": den medlemsstat där det fordon varmed trafikförseelsen begicks är registrerat,
d)
"behörig myndighet": den
enda kontaktpunkt i varje medlemsstat som är ansvarig för att underlätta genomförandet av detta direktiv
,
e)
"centralmyndighet": den myndighet som är ansvarig för att säkerställa uppgiftsskyddet i varje medlemsstat,
f)
"slutgiltigt administrativt beslut": ett slutgiltigt beslut som innebär att en finansiell påföljd måste betalas, och som inte utgör ett beslut enligt definitionen i artikel 1 i rambeslut 2005/214/RIF,
g)
"fortkörning": överskridning av de hastighetsbegränsningar som gäller i landet där förseelsen begicks för vägen eller fordonet i fråga,
h)
"rattfylleri": körning med en alkoholhalt i blodet som överskrider den högsta tillåtna promillegränsen i landet där förseelsen begicks,
i)
"bristande bältesanvändning": åsidosättande av kravet på bälte eller barnstol när det är obligatoriskt att använda sådan utrustning i enlighet med rådets direktiv 91/671/EEG Rådets direktiv 91/671/EEG av den 16 december 1991 om tillnärmning av medlemsstaternas lagstiftning om obligatorisk användning av bilbälten i fordon som väger mindre än 3,5 ton (EGT L 373, 31.12.1991, s.
26)║.
eller den nationella lagstiftningen i landet där förseelsen begicks,
j)
"rödljuskörning": körning mot rött trafikljus, i enlighet med den definition som ges i lagstiftningen för landet där förseelsen begicks.
Artikel 3
Riktlinjer för trafiksäkerheten i EU
1.
För att bedriva en trafiksäkerhetspolitik som syftar till en hög skyddsnivå för samtliga vägtrafikanter i Europeiska unionen, och med hänsyn till de mycket skiftande situationer som förekommer inom Europeiska unionen, ska medlemsstaterna, utan att detta påverkar mer restriktiv politik och lagstiftning, agera i syfte att tillhandahålla en minimiuppsättning riktlinjer för trafiksäkerhet inom tillämpningsområdet för detta direktiv.
För att uppnå detta mål ska kommissionen anta riktlinjer för vägsäkerhet inom hela EU i enlighet med det föreskrivande förfarande med kontroll som avses i artikel 13
.
2.
Dessa riktlinjer ska följa de miniminormer som fastställs i denna artikel
.
2.
När det gäller hastighet ska användningen av automatisk kontrollutrustning på motorvägar, landsvägar och stadsgator särskilt uppmuntras särskilt på avsnitt av vägnätet där antalet trafikolyckor till följd av fortkörning är högre än genomsnittet.
Syftet med de rekommendationer som antas inom ramen för dessa riktlinjer är att säkerställa antalet hastighetskontroller som sker med hjälp av automatisk utrustning ska öka med 30 % i de medlemsstater där antalet dödsfall i trafiken överstiger genomsnittet i unionen och minskningen av antalet dödsfall i trafiken sedan 2001 understiger genomsnittet i EU.
3.
När det gäller rattfylleri ska medlemsstaterna prioritera genomförandet av stickprov på platser och vid tillfällen då förseelser är vanligt förekommande och ökar risken för olyckor
.
Medlemsstaterna ska säkerställa att minst 30 % av förarna har kunnat kontrolleras varje år.
4.
När det gäller bältesanvändning ska medlemsstaterna genomföra intensiva kontroller i minst sex veckor under ett givet år i sådana medlemsstater där mindre än 70 % av väganvändarna använder bälte, särskilt på platser och vid tillfällen då förseelser är vanligt förekommande.
5.
När det gäller rödljuskörning ska användningen av automatisk kontrollutrustning framför allt i korsningar där förseelser är vanligt förekommande och där det inträffar fler olyckor än det genomsnittliga antalet olyckor till följd av rödljuskörning.
6.
Enligt riktlinjerna ska medlemsstaterna rekommenderas att utbyta god praxis och de medlemsstater som har kommit längst när det gäller automatiska kontroller ska särskilt uppmanas att ge tekniskt stöd till de medlemsstater som ber om detta.
KAPITEL II
BESTÄMMELSER SOM UNDERLÄTTAR GRÄNSÖVERSKRIDANDE UPPFÖLJNING
Artikel 4
Förfarande för informationsutbyte mellan medlemsstaterna
1.
2.
Den behöriga myndigheten i bosättningslandet ska omedelbart skicka följande information till den behöriga myndigheten i landet där förseelsen begicks:
a)
Märke och modell på fordonet med registreringsnumret i fråga.
b)
Namn, adress, födelseort och födelsedatum, om innehavaren av registreringsbeviset är en fysisk person.
c)
Namn och adress, om innehavaren av registreringsbeviset är en juridisk person.
3.
När det gäller behandling av personuppgifter och det fria flödet av sådana uppgifter ska informationsutbytet ske med iakttagande av direktiv 95/46/EG.
De behöriga myndigheterna i de andra medlemsstaterna ska inte lagra den information som översänds av landet där förseelsen begicks
Artikel 5
Ett elektroniskt nät
1.
Medlemsstaterna ska vidta alla nödvändiga åtgärder för att se till att informationsutbytet enligt
artikel 4
sker elektroniskt.
I detta syfte
2.
Gemensamma regler om genomförande av punkt 1 ska antas av kommissionen
senast
den dag som anges i
artikel 15.1
med kontroll
i
artikel 13
2
.
Dessa gemensamma regler ska omfatta särskilda bestämmelser om
a)
formatet för den information som utbyts,
b)
de tekniska förfarandena för det elektroniska informationsutbytet mellan medlemsstaterna
, med garantier för de översända uppgifternas säkerhet och konfidentialitet
,
c)
Artikel 6
Meddelande om trafikförseelse
1.
2.
relevanta uppgifter om trafikförseelsen.
bötesbeloppet
möjligheterna att bestrida grunderna för
utfärdandet av
3
4
.
Innehavaren ska genom meddelandet om trafikförseelse informeras om att ett svarsformulär måste fyllas i
inom en fastställd tidsfrist
de finansiella påföljderna
5
6
Detta ska inte tillämpas om det finns ett avtal mellan två eller flera medlemsstater för att lösa de problem som uppstår till följd av tillämpningen av denna artikel.
7
.
Meddelandet om trafikförseelse ska skickas till innehavaren på det eller de officiella språk i bosättningslandet som har uppgivits av landet.
8
.
Kommissionen får anpassa förlagan till meddelande om trafikförseelse för att ta hänsyn till den tekniska utvecklingen.
Åtgärder som syftar till att ändra mindre väsentliga
tekniska
.
2
.
9
Artikel 7
Uppföljning av trafikförseelser
1.
Om den finansiella påföljden inte betalas och möjligheterna att tillämpa de förfaranden som gäller vid tvist eller överklagan har uttömts, ska rambeslut 2005/214/RIF tillämpas på de finansiella påföljder som avses i artikel 1 i detta rambeslut.
2.
I sådana fall av betalningsvägran som de som avses i punkt 1, men där betalningsvägran avser finansiella påföljder som inte omfattas av tillämpningsområdet för nämnda rambeslut, ska den behöriga myndigheten i det land där förseelsen ägde rum översända det slutgiltiga beslutet till den behöriga myndigheten i bosättningslandet för verkställande av den finansiella påföljden.
Artikel 8
Erkännande och verkställande av finansiella påföljder
1.
a)
b)
Berörd part har inte informerats om sin rätt att överklaga och om tidsfristen för en sådan överklagan.
2.
Verkställandet av det beslut om en finansiell påföljd som fattats av behörig myndighet i bosättningslandet ska regleras av lagen i bosättningslandet på samma sätt som ett bötesstraff i detta land.
3.
Den behöriga myndigheten i landet där förseelsen ägde rum ska genast informera den behöriga myndigheten i bosättningslandet om varje beslut eller åtgärd som förhindrar genomförandet av beslutet.
Den behöriga myndigheten i bosättningslandet ska inställa genomförandet av beslutet, så snart den erhåller information från den behöriga myndigheten i landet där förseelsen ägde rum om ett sådant beslut eller en sådan åtgärd.
Artikel 9
Information från bosättningslandet
a)
b)
c)
Verkställandet av beslutet så snart detta har skett.
Artikel 10
Centralmyndigheter
1.
Varje medlemsstat ska utse en centralmyndighet som ska bistå vid tillämpningen av detta direktiv.
2.
Medlemsstaterna ska inom sex månader från och med att detta direktiv träder i kraft meddela kommissionen namn och adress till de myndigheter som utsetts i enlighet med denna artikel.
3.
Artikel 11
Rätt till tillgång, rättelse och radering
1.
Alla ska ha rätt att få tillgång till egna personuppgifter som registrerats i bosättningslandet och som har sänts över till den medlemsstat som begärt dem, utan att detta påverkar
2.
Alla berörda personer ska ha rätt att utan dröjsmål få oriktiga personuppgifter rättade och olagligt registrerade uppgifter raderade, utan att detta påverkar iakttagandet av de formella kraven i samband med den berörda medlemsstatens mekanismer för överklagan och prövning.
3.
Registrerade personer kan utöva rättigheterna i punkt 2 inför centralmyndigheten i sitt bosättningsland.
Artikel 12
Information till förarna i Europeiska unionen
1.
Medlemsstaterna ska vidta lämpliga åtgärder för att ge trafikanterna tillräcklig information om åtgärderna för tillämpning av detta direktiv.
Sådan information kan tillhandahållas av bl.a. trafiksäkerhetsorganisationer, icke-statliga organisationer som verkar på området för trafiksäkerhet eller klubbar.
2.
Kommissionen ska på sin hemsida offentliggöra en sammanfattning av de bestämmelser som gäller i medlemsstaterna och som omfattas av tillämpningsområdet för detta direktiv.
KAPITEL III
KOMMITTÉFÖRFARANDE
Artikel 13
Kommitté
1.
Kommissionen ska bistås av en kommitté för kontroller på området vägtrafiksäkerhet.
2
.
Artikel 14
Översyn och rapport
1.
Senast ...
*
Två år efter det att detta direktiv har trätt ikraft
.
2.
På grundval av denna rapport ska kommissionen granska möjligheterna att utvidga direktivets tillämpningsområde till att gälla andra trafikförseelser.
3.
I denna rapport ska kommissionen lägga fram förslag om en harmonisering av kontrollutrustningen på grundval av gemenskapskriterier och kontrollpraxis på trafiksäkerhetsområdet.
4.
I rapporten ska kommissionen dessutom utvärdera i vilken utsträckning medlemsstaterna frivilligt har genomfört de riktlinjer för vägsäkerhet inom hela EU som avses i artikel 3 och granska frågan om huruvida rekommendationer i dessa riktlinjer bör göras obligatoriska.
I lämpliga fall ska kommissionen lägga fram ett förslag om ändring av detta direktiv.
KAPITEL IV
SLUTBESTÄMMELSER
Artikel 15
Införlivande
1.
Medlemsstaterna ska sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa det här direktivet senast tolv månader efter det att direktivet träder i kraft.
De ska genast överlämna texterna till dessa bestämmelser till kommissionen tillsammans med en jämförelsetabell för dessa bestämmelser och bestämmelserna i detta direktiv.
När en medlemsstat antar dessa bestämmelser ska de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs.
Närmare föreskrifter om hur hänvisningen ska göras ska varje medlemsstat själv utfärda.
2.
Medlemsstaterna ska till kommissionen överlämna texten till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 16
Ikraftträdande
Detta direktiv träder i kraft dagen efter det att det har offentliggjorts i Europeiska unionens officiella tidning.
Artikel 17
Adressater
Detta direktiv riktar sig till medlemsstaterna.
Utfärdat i ║ den
På Europaparlamentets vägnar På rådets vägnar
Ordförande Ordförande
BILAGA
[Avsändarens namn, adress och telefonnummer] [Adressatens namn och adress]
meddelande om en trafikförseelse som begåtts i …….. [den medlemsstat där förseelsen ägde rum] [denna text återges på försättsbladet på alla officiella EU-språk] Sida 2
Den [datum ….. ] begicks en trafikförseelse med ett fordon med registreringsnummer ……….. av märket……., modell…….., vilken konstaterades av……………[namn på ansvarigt organ]
Du är registrerad som innehavare av registreringsbeviset för fordonet i fråga.
Förseelsen beskrivs närmare på sidan 3.
Bötesbeloppet för denna förseelse uppgår till ………euro/nationell valuta.
Betalningsfristen löper ut den ..............
Denna svarsblankett får översändas av [den behöriga myndigheten i landet där förseelsen begicks] till [den behöriga myndigheten i bosättningslandet] för verkställande av beslutet om påföljd.
INFORMATION
Detta ärende kommer att behandlas av den behöriga myndigheten i landet där förseelsen begicks.
Om ärendet inte lagförs, kommer ni att underrättas inom 60 dagar från det att myndigheten tagit emot svarsblanketten.
Om ärendet lagförs, kommer följande förfarande att tillämpas:
[Ifylles av landet där förseelsen begicks - redogörelse för vidare förfarande, inklusive närmare information om möjligheten att överklaga beslutet att lagföra ärendet och om förfarandet för detta.
Denna information ska under alla omständigheter omfatta namn och adress till myndigheten med ansvar för att följa upp ärendet, betalningsfrist, namn och adress till behörig instans för överklagan samt sista dag för överklagan].
___________________________________________________________________________ Sida 3 Beskrivning av förseelsen
a)
Registreringsnummer:
Registreringsland:
Märke och modell:
b)
Uppgifter om förseelsen
Ort, datum och tidpunkt för förseelsen:
Förseelsens art och rubricering:
fortkörning, rattfylleri, bristande användning av bälte eller barnstol, rödljuskörning Stryk det som ej är tillämpligt.
Detaljerad beskrivning av förseelsen:
Hänvisning till relevant lagstiftning:
Beskrivning av eller hänvisning till beviset för förseelsen:
c)
Uppgifter om den utrustning som användes för att konstatera förseelsen Ej tillämpligt om ingen utrustning använts.
Typ av utrustning för att konstatera fortkörning, rattfylleri, rödljuskörning eller bristande bältesanvändning1.
Specifikation av utrustningen:
Utrustningens identifieringsnummer:
Senaste kalibreringen giltig till och med:
d)
Resultat vid användningen av utrustningen:
[exemplet gäller fortkörning, andra förseelser läggs till:]
Högsta tillåtna hastighet:
Uppmätt hastighet:
Uppmätt hastighet efter avdrag av felmarginal:
Sida 4 Svarsblankett (ifylles med VERSALER, markera det riktiga alternativet)
A.
Förarens personuppgifter:
Körde du fordonet då förseelsen begicks
(ja/nej)
Om ja, fyll i uppgifterna nedan:
–
Efternamn och förnamn:
–
Födelseort och födelsedatum:
–
Körkortsnummer: ……, utställt den (datum): …….. i (ort):
–
Adress:
Om du inte körde fordonet då förseelsen begicks, kan du ange förarens identitet
(ja/nej)
Om ja, fyll i uppgifterna nedan avseende föraren:
–
Efternamn och förnamn:
–
Födelseort och födelsedatum:
–
Körkortsnummer: ……, utställt den (datum): …….. i (ort):
–
Adress:
B.
Frågor:
(1)
Är fordonet av märket …….. med registreringsnummer ……. registrerat i ert namn?
ja/nej
Om inte, ange vem som är innehavare av registreringsbeviset:
(efternamn, förnamn, adress)
(2)
Erkänner du dig skyldig till förseelsen?
ja/nej
(3)
Om inte,
och om du vägrar att ange förarens identitet,
förklara varför du anser att du inte är skyldig:
Den ifyllda blanketten skickas inom 60 dagar från och med datumet för detta meddelande till följande myndighet:
på följande adress:
▌
P6_TA(2009)0185
EIB:s och EBRD:s årsrapporter för 2007
A6-0135/2009
Europaparlamentet utfärdar denna resolution
–
med beaktande av Europeiska investeringsbankens (EIB) årsrapport för 2007,
–
med beaktande av årsrapporten från Europeiska banken för återuppbyggnad och utveckling (EBRD) för 2007,
–
med beaktande av artiklarna 9, 266 och 267 i EG-fördraget och protokoll nr 11 om EIB:s stadga,
–
med beaktande av avtalet om upprättande av Europeiska banken för återuppbyggnad och utveckling av den 29 maj 1990,
–
med beaktande av artiklarna 230 och 232 i EG-fördraget om EG-domstolens roll,
–
med beaktande av artikel 248 i EG-fördraget om revisionsrättens roll,
–
med beaktande av rådets beslut 2006/1016/EG av den 19 december 2006 om beviljande av en gemenskapsgaranti till Europeiska investeringsbanken mot förluster vid lån till och lånegarantier för projekt utanför gemenskapen EUT L 414, 30.12.2006, s.
95.
,
–
,
–
med beaktande av rådets beslut 2008/847/EG av den 4 november 2008 om berättigande för centralasiatiska länder till EIB-finansiering inom ramen för beslut 2006/1016/EG om beviljande av en gemenskapsgaranti till Europeiska investeringsbanken mot förluster vid lån till och lånegarantier för projekt utanför gemenskapen EUT L 301, 12.11.2008, s.
13.
,
–
med beaktande av rådets beslut 97/135/EG av den 17 februari 1997 om Europeiska gemenskapens tecknande av nya andelar kapital i Europeiska banken för återuppbyggnad och utveckling till följd av beslutet att fördubbla detta kapital EGT L 52, 22.2.1997, s.
15.
,
–
med beaktande av EBRD:s nuvarande översyn av kapitalresurserna (Capital Resources Review) från 2006 som omfattar perioden 2006−2010,
–
med beaktande av kommissionens rapport till Europaparlamentet och rådet om Europeiska gemenskapernas upp- och utlåning 2007 ( KOM(2008)0590 ),
–
med beaktande av sin resolution av den 22 april 2008 om Europeiska investeringsbankens årsrapport för 2006 Antagna texter, P6_TA(2008)0132 .
,
–
med beaktande av sin resolution av den 15 februari 2007 om EIB:s årsrapport för 2005 EUT C 287 E, 29.11.2007, s.
544.
,
–
med beaktande av sin resolution av den 16 januari 2003 om verksamheten vid Europeiska banken för återuppbyggnad och utveckling (EBRD) EUT C 38 E, 12.2.2004, s.
313.
,
–
med beaktande av Europarådets parlamentariska församlings resolution av den 24 juni 2008 om Europeiska banken för återuppbyggnad och utveckling som en stark partner för förändringen i övergångsländerna,
–
med beaktande av partnerskapsavtalet mellan medlemmarna i gruppen av stater i Afrika, Västindien och Stillahavsområdet å ena sidan, och Europeiska gemenskapen och dess medlemsstater å andra sidan, undertecknat i Cotonou den 23 juni 2000 EGT L 317, 15.12.2000, s.
3.
(Cotonou-avtalet),
–
med beaktande av den gemensamma förklaringen från rådet och företrädarna för medlemsstaternas regeringar församlade i rådet, Europaparlamentet och kommissionen om Europeiska unionens utvecklingspolitik – "Europeiskt samförstånd" EUT C 46, 24.2.2006, s.
1.
,
–
med beaktande av rådets slutsatser av den 14 maj 2008 om en investeringsram för västra Balkan: Att öka enhetligheten bland de nuvarande finansieringsinstrumenten för regionen i syfte att främja tillväxt och stabilitet,
–
med beaktande av kommissionens förslag av den 21 maj 2008 om en förordning om ändring av förordning (EG) nr 1638/2006 av den 24 oktober 2006 om fastställande av allmänna bestämmelser för upprättandet av ett europeiskt grannskaps- och partnerskapsinstrument ( KOM(2008)0308 ),
–
I-7141).
,
–
–
med beaktande av det avtal om samförstånd som undertecknades den 15 december 2006 mellan kommissionen, EIB och EBRD beträffande samarbete i Östeuropa och södra Kaukasus, Ryssland och Centralasien,
–
med beaktande av det avtal om samförstånd som undertecknades den 27 maj 2008 mellan kommissionen och Europeiska investeringsbanken om att främja samordningen av Europeiska unionens externa lånepolitik,
–
med beaktande av det avtal om deltagande i det europeiska centrumet för specialistkunskap på området för offentlig–privata partnerskap som undertecknades den 16 september 2008 mellan EIB, kommissionen och de nationella behöriga myndigheterna,
–
med beaktande av EIB:s verksamhetsplan för 2008–2010 som godkändes av bankens styrelse den 20 november 2007,
–
med beaktande av EIB:s offentliga samråd 2008 om dess förklaring om miljömässiga och sociala principer och standarder,
–
med beaktande av EBRD:s miljö- och socialpolitik som godkändes av styrelsen den 12 maj 2008,
–
med beaktande av EBRD:s politik för energiåtgärder som godkändes av styrelsen den 11 juli 2006,
–
med beaktande av EIB:s översyn av sin energipolitik som godkändes av styrelsen den 31 januari 2006,
–
med beaktande av EIB:s informationsmeddelande om förstärkta bidrag till EU:s energipolitik av den 5 juni 2007, som godkändes av styrelsen i juni 2007,
−
med beaktande av ordförandeskapets slutsatser från Europeiska rådets möte i Bryssel den 11-12 december 2008 om ekonomiska och finansiella frågor,
−
med beaktande av EIB:s rapport med titeln "Samråd med små och medelstora företag 2007/2008 – resultat och slutsatser", från maj 2008, och den efterföljande moderniseringen och förstärkningen av EIB-gruppens stöd till EU:s små och medelstora företag,
–
med beaktande av EIB:s förklaring om miljömässiga och sociala principer och standarder, av den 18 mars 2008,
−
med beaktande av rådets slutsatser från Ecofinrådet av den 7 oktober 2008 och den 2 december 2008 om EIB:s roll för stödet till små och medelstora företag,
−
med beaktande av kommissionens meddelande av den 29 oktober 2008 med titeln "Från finanskris till återhämtning: ram för åtgärder på EU-nivå" ( KOM(2008)0706 ),
−
med beaktande av kommissionens meddelande av den 26 november 2008 med titeln "En ekonomisk återhämtningsplan för Europa" ( KOM(2008)0800 ),
–
med beaktande av artikel 45 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för ekonomi och valutafrågor och yttrandet från budgetkontrollutskottet ( A6-0135/2009 ), och av följande skäl:
A.
EIB inrättades 1975 genom Romfördraget, och andelsägarna, det vill säga medlemsstaterna, har tecknat ett kapital som uppgår till 165 miljarder EUR.
B.
EIB har sedan 1963 genomfört transaktioner utanför gemenskapen till stöd för gemenskapens utrikespolitik.
C.
EBRD inrättades 1991 och dess andelsägare utgörs av 61 tredjeländer, Europeiska gemenskapen och EIB, som tillsammans har tecknat ett kapital som uppgår till totalt 20 miljarder EUR.
D.
Medlemsstaterna, Europeiska gemenskapen och EIB har tillsammans tecknat 63 procent av andelarna i EBRD.
E.
EIB:s lagstadgade mål är att genom att anlita kapitalmarknaderna och utnyttja egna medel bidra till en balanserad och störningsfri utveckling av den inre marknaden i gemenskapens intresse.
F.
Under den pågående finansiella oron och den enorma bristen på likviditet och krediter för företagen bör EIB spela en viktig roll i kommissionens och medlemsstaternas planer för den ekonomiska återhämtningen.
G.
EBRD:s lagstadgade mål är att genom att bidra till ekonomisk utveckling och återuppbyggnad gynna övergången till öppna marknadsorienterade ekonomier och att främja privata initiativ och företagaranda i de central- och östeuropeiska länder som bekänner sig till och som tillämpar principerna för demokratiskt flerpartisystem, pluralism och marknadsekonomi.
H.
EIB:s roll som utgivare av högt värderade AAA-obligationer för de internationella kapitalmarknaderna bör betonas och förstärkas.
I.
Enligt artikel 11 i avtalet om upprättandet av EBRD måste EBRD göra minst 60 procent av sina investeringar i den privata sektorn.
J.
Avtalet om upprättandet av EBRD föreskriver att styrelsen minst vart femte år ska företa en översyn av bankens kapital, och nästa översyn planeras äga rum 2010.
K.
En styrkommitté bestående av nio så kallade visa personer tillsattes den 1 oktober 2008 för att övervaka och sköta utvärderingen av halvtidsöversynen av EIB:s externa utlåningsmandat i enlighet med beslut 2006/1016/EG.
L.
Denna halvtidsöversyn bör göras i nära samråd med parlamentet, i enlighet med beslut 2006/1016/EC.
M.
I beslut 2006/1016/EG om EIB:s mandat för extern utlåning föreskrivs att lån till ett belopp av 25,8 miljarder EUR ska vara tillgängliga under perioden 2007−2013 fördelat på regioner enligt följande: föranslutningsländer, inklusive Kroatien och Turkiet, 8,7 miljarder EUR, Medelhavsländerna 8,7 miljarder EUR, Östeuropa, södra Kaukasus och Ryska federationen 3,7 miljarder EUR, Latinamerika 2,8 miljarder EUR, Asien 1 miljard EUR, och Republiken Sydafrika 0,9 miljarder EUR.
N.
De lån som EIB beviljat 2007 till stöd för EU:s politiska mål uppgick till 47,8 miljarder EUR, varav 41,4 miljarder EUR till länder i Europeiska unionen och Efta och 6,4 miljarder EUR till partner- och kandidatländer.
O.
EIB:s utlåningsverksamhet under 2007 utanför EU per geografiskt område såg ut på följande sätt: Asien och Latinamerika 925 miljoner EUR, Östeuropa, Södra Kaukasus, Ryssland och Centralasien 230 miljoner EUR, Medelhavsländerna 1 438 miljoner EUR, föranslutningsländer 2 870 miljoner EUR, AVS-länder 756 miljoner EUR och Sydafrika 113 miljoner EUR.
P.
EBRD:s årsomsättning uppgick under 2007 till 5,6 miljarder EUR och omfattade 353 projekt i 29 verksamhetsländer i Centraleuropa och de baltiska länderna Kroatien, Tjeckien, Estland, Ungern, Lettland, Litauen, Polen, Slovakien och Slovenien.
, sydöstra Europa Albanien, Bosnien och Hercegovina, Bulgarien, f.d. jugoslaviska republiken Makedonien, Montenegro, Rumänien och Serbien.
, västra OSS och Kaukasus Armenien, Azerbajdzjan, Vitryssland, Georgien, Moldavien och Ukraina.
, Ryssland och Centralasien Kazakstan, Kirgizistan, Mongoliet, Tadzjikistan, Turkmenistan och Uzbekistan.
.
Q.
EBRD: s investeringar i Ryssland ökade under 2007 till 2,3 miljarder EUR (det totala beloppet i Ryssland uppgick till 5,7 miljarder EUR) och omfattade 83 projekt och utgjorde 42 procent av EBRD:s årliga åtaganden (jämfört med 38 procent 2006).
R.
EBRD:s kapitalinvesteringar ökade under 2007 från 1 miljard EUR 2006 till 1,7 miljarder EUR 2007, och den del av EBRD:s årsomsättning som utgörs av eget kapital ökade från 20 procent 2006 till 30 procent 2007.
S.
T.
EIB har finansierat projekt i Turkiet sedan 1965 och investerat ungefär 10 miljarder EUR i alla viktiga sektorer av Turkiets ekonomi.
U.
I enlighet med Cotonou-avtalet ska EIB utöver att låna ut från det egna kapitalet även finansiera insatser i AVS-länderna med hjälp av ett riskbärande investeringsinstrument vars anslag kommer från Europeiska utvecklingsfonden.
V.
EIB:s finansieringsstrategi bör bidra till det allmänna målet att utveckla och befästa demokratin och rättsstatsprincipen samt att iaktta internationella miljöavtal i vilka gemenskapen eller dess medlemsstater är parter.
W.
Kommissionen, medlemsstaterna, partnerländerna i den europeiska grannskapspolitiken, de internationella finansinstituten och de europeiska regionala och bilaterala finansinstituten samarbetar för närvarande inom ramen för ett investeringsinstrument för grannskapspolitiken för ytterligare finansiering av infrastrukturprojekt, huvudsakligen avseende energi, transporter och miljö, i hela det område som omfattas av den europeiska grannskapspolitiken.
X.
EIB:s mål och verksamhet
1.
Europaparlamentet välkomnar EIB:s årsrapport för 2007, särskilt EIB:s finansieringsverksamhet i Europeiska unionen som inriktats på sex politiska prioriteringar (som säkerställer ekonomisk och social sammanhållning, genomförande av initiativet Innovation 2010, utveckling av transeuropeiska transport- och anslutningsnät, stöd till små och medelstora företag, skydd och förbättring av miljön samt hållbar, konkurrenskraftig och säker energi), och även genomförandet av EIB:s mandat för externa lån till tredjeländer.
2.
3.
Europaparlamentet noterar att EIB är det enda fördragsbaserade finansinstitutet och att majoriteten av dess verksamhet är koncentrerad till projekt i medlemsstaterna, samtidigt som banken också har en allt viktigare roll att spela i tredjeländer, i enlighet med beslut 2006/1016/EG.
4.
5.
6.
7.
8.
Parlamentet uppmanar med kraft EIB att i samband med bankens globala lån för stöd till små och medelstora företag förbättra övervakningen och säkerställa insyn när det gäller typen av lån och slutlig mottagare av dessa.
9.
När det gäller tillsynen av EIB
a)
påminner Europaparlamentet om att EIB, vars uppgifter är politiskt definierade, inte är föremål för den normalt förekommande tillsynen, och anser att tillsyn över EIB:s arbetsmetoder inte desto mindre är nödvändig,
b)
c)
välkomnar parlamentet EIB:s tekniska samarbete med de nationella tillsynsmyndigheterna i Luxemburg, men föreslår att samarbetet utvidgas,
d)
uppmanar parlamentet kommissionen och medlemsstaterna att undersöka om det är möjligt att göra en mer omfattande revidering av arrangemangen för tillsyn över EIB:s finansiella verksamhet, som skulle kunna genomföras av en framtida europeisk banktillsynsmyndighet, för att kontrollera att EIB:s finansiella situation är god, att dess resultat mäts exakt och att reglerna för god praxis inom yrket efterlevs.
10.
Europaparlamentet välkomnar utvecklingen och offentliggörandet under 2007 av EIB:s sektorsvisa operativa strategier i energi-, transport- och vattensektorerna som ett viktigt steg mot att öka insynen i EIB:s utlåningsverksamhet.
11.
Europaparlamentet välkomnar översynen av EIB:s offentlighetsstrategi för att beakta de relevanta bestämmelserna i Århusförordningen Europaparlamentets och rådets förordning (EG) nr 1367/2006 av den 6 september 2006 om tillämpning av bestämmelserna i Århuskonventionen om tillgång till information, allmänhetens deltagande i beslutsprocesser och tillgång till rättslig prövning i miljöfrågor på gemenskapens institutioner och organ (EUT L 264, 25.9.2006, s.
Parlamentet välkomnar offentliggörandet av EIB:s rapport för 2007 om utvärdering av verksamheten och uppmuntrar EIB att vidareutveckla avdelningen för utvärdering av verksamheten.
12.
13.
a)
administrativa förfaranden som utestänger företag som EIB eller andra multilaterala utvecklingsbanker funnit skyldiga till bedrägerier,
b)
en politik för att skydda personer som avslöjar missförhållanden, och
c)
en förstärkning av dess utredningsfunktion och av den därmed sammanhängande förebyggande och avslöjande rollen.
14.
15.
16.
17.
EBRD:s mål och verksamhet
18.
Europaparlamentet välkomnar EBRD:s årsrapport för 2007, särskilt den omständigheten att EBRD:s investeringsverksamhet inriktats på länder som befinner sig i ett tidigt skede eller i ett mellanskede av en övergångsperiod, och välkomnar de framsteg som gjorts när det gäller finansieringen av projekt inom ramen för bankens initiativ för hållbar energi, för vilka energiprojekt som är av intresse för EU bör prioriteras.
19.
Europaparlamentet konstaterar att EBRD främst är verksam i tredjeländer, men att det även i fortsättningen är viktigt med viss verksamhet i medlemsstaterna.
20.
Europaparlamentet konstaterar dessutom att mycket har förändrats sedan 1991 när det gäller EBRD:s roll i ett internationellt och regionalt sammanhang, och att EBRD:s mandat måste tillämpas i denna nya miljö i takt med att EBRD reagerar på marknadsförhållandena och flyttar sin verksamhet längre söder- och österut.
21.
Europaparlamentet konstaterar också att verksamhetsmiljön innebär allt större utmaningar eftersom företagsklimatet har blivit svårare på grund av att de lokala partnernas erfarenheter tenderar att minska och integritetsproblemen med tenderar att öka.
22.
Europaparlamentet anser att EBRD måste förbättra sitt tekniska stöd och sin rådgivningsverksamhet för att främja standarder för god förvaltning och se till att projekten förvaltas på lämpligt sätt på lokal nivå i EU:s grannskapsländer.
23.
Samarbete mellan EIB och EBRD och med andra internationella, regionala och nationella finansinstitut
24.
Europaparlamentet konstaterar att EIB och EBRD i allt större omfattning finansierar verksamhet i samma geografiska områden utanför Europeiska unionen, såsom i Östeuropa, södra Kaukasus, Ryssland, länderna i västra Balkan och inom en snar framtid även Turkiet.
25.
Europaparlamentet påpekar att i länder där båda bankerna bedriver verksamhet finns för närvarande tre olika typer av samarbete mellan EIB och EBRD: För östra Europa finns det ett avtal om samförstånd som EBRD ansvarar för och där gemensamma investeringar är den allmänna regeln, på västra Balkan har det skett en förskjutning från konkurrens eller parallell verksamhet till samarbete genom gemensamt utnyttjande av medlen, och nyligen, t.ex. när det gäller samarbetet i Turkiet, till ett avtal med utgångspunkt i särskilda gemensamma kompetensområden där huvudansvaret ska avgöras från fall till fall.
26.
27.
Europaparlamentet anser att EIB:s och EBRD:s verksamhet i de länder där båda är verksamma inte bör konkurrera, utan snarare komplettera varandra, att detta bör ske på grundval av varje banks komparativa fördelar, och att kunden inte bör drabbas av extra kostnad på grund av överlappningar.
28.
I syfte att uppnå ett bättre strukturerat samarbete mellan EIB och EBRD i länder med gemensam verksamhet rekommenderar därför Europaparlamentet
a)
att båda bankerna förbättrar sin funktionella arbetsfördelning för att öka specialiseringen och inrikta sig på sina respektive kompetenser och styrkor,
b)
att EIB specialiserar sig mer på finansieringen av mer storskaliga privata och offentliga infrastrukturer och projekt, inbegripet offentlig-privata partnerskapsinvesteringar samt utländska direktinvesteringar från EU-företag, och att EBRD specialiserar sig mer på småskaliga investeringar, institutionell uppbyggnad, privatiseringar, underlättande av handel, finansiella marknader och direkta kapitalinvesteringar för att främja normer för bolagsstyrning,
c)
att man definierar vilka typer av projekt, sektorer och produkter som är av potentiellt intresse för båda bankerna och där de skulle kunna bygga upp gemensamma kunskaps- och resurspooler, såsom finansiering av små och medelstora företag, främjande av investeringar för att bekämpa klimatförändringar, t.ex. uppmuntran av energi från förnybara källor och minskning av växthusgasutsläppen, och begär ett pragmatiskt tillvägagångssätt som anpassas till varje enskilt fall på de områden där det finns gemensamma intressen, och där en institution är huvudansvarig för varje samfinansieringsprojekt i syfte att undvika överlappningar, och att detta sker på grundval av ett ömsesidigt erkännande av förfaranden; i detta sammanhang måste projekt som stöds av EU motsvara EU:s standarder, till exempel när det gäller klimatskyddet eller de sociala rättigheterna, oavsett om det är EIB eller EBRD som är den ansvariga institutionen,
d)
att tydliga samarbetsmekanismer införs i båda institutionerna, både uppifrån och ned och på fältet,
e)
att båda bankerna lägger fram ett konkret förslag om ett mer konsekvent samarbete, som även omfattar en reflektion över gemensamma standarder, vilket är till fördel för andelsägarna, de berörda parterna och de mottagande länderna,
f)
att båda bankerna regelbundet rapporterar till kommissionen om samarbetet,
g)
att kommissionen avlägger en årlig rapport till parlamentet och rådet om bedömningen av resultaten av EIB:s och EBRD:s finansieringsverksamhet och dess effektivitet samt respektive banks bidrag till uppfyllandet av Europeiska unionens utrikespolitiska mål, och om det ömsesidiga samarbetet mellan bankerna och med andra finansinstitut, och
h)
att årliga utfrågningar av båda bankernas ordförande tillsammans med kommissionsledamoten med ansvar för ekonomiska och monetära frågor anordnas i parlamentet.
29.
30.
31.
32.
33.
Den globala oron på finansmarknaderna och konsekvenserna för EIB och EBRD
34.
35.
36.
37.
38.
Europaparlamentet uppmanar medlemsstaterna att till fullo utnyttja de instrument i form av riskkapital, globala lån och mikrokrediter som erbjuds genom EIB:s program och instrument.
39.
40.
Europaparlamentet uppmanar enträget kommissionen och EIB att tillsammans undersöka hur lånekrisen i den reala ekonomin kan bemästras med hjälp av nya innovativa finansiella instrument.
41.
Europaparlamentet välkomnar EBRD:s beslut att öka bankens årsomsättning 2009 med ca 20 procent till ca 7 miljarder EUR för att mildra den pågående finansiella och ekonomiska krisen, och konstaterar att hälften av de extra medlen på 1 miljard EUR 2009 är öronmärkta för Central- och Östeuropa.
42.
Europaparlamentet betonar att i den nuvarande situationen med snäva kreditvillkor framhävs de två bankernas roll både i och utanför Europeiska unionen, och uppmanar båda bankerna att hålla sina utfästelser gentemot tredjeländer, även i ekonomiskt svåra tider.
43.
44.
Europaparlamentet noterar med tillfredsställelse att EIB och EBRD har utsatts för den finansiella oron i ganska begränsad omfattning, även om EBRD redovisade sin första förlust 2008 under det här årtiondet till följd av nedgången på aktiemarknaderna.
Konsekvenserna av domstolens dom när det gäller EIB:s externa mandat
45.
Europaparlamentet välkomnar domstolens dom av den 6 november 2008 om den rättsliga grunden för beslut 2006/1016/EG.
46.
47.
48.
°
° °
49.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, Europeiska investeringsbanken, Europeiska banken för återuppbyggnad och utveckling samt medlemsstaternas regeringar och parlament.
P6_TA(2009)0289
Ansvarsfrihet 2007: Kommissionen
A6-0168/2009
1.
Europaparlamentets beslut av den 23 april 2009 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2007 - avsnitt III, kommissionen - verkställande organ ( SEK(2008)2359 – C6-0415/2008 – 2008/2186(DEC) )
Europaparlamentet fattar detta beslut
–
,
–
med beaktande av Europeiska gemenskapernas slutliga årsredovisning för budgetåret 2007 – Volym I ( SEK(2008)2359 – C6-0415/2008 ) EUT C 287, 10.11.2008, s.
1.
,
–
med beaktande av kommissionens årsrapporter till Europaparlamentet och rådet om uppföljningen av besluten om ansvarsfrihet 2006 ( KOM(2008)0629 och KOM(2008)0628 ) samt av de arbetsdokument från kommissionens tjänsteavdelningar som åtföljer dessa rapporter ( SEK(2008)2579 och SEK(2008)2580 ),
–
med beaktande av kommissionens meddelande med titeln "Sammanfattande rapport om kommissionens förvaltning 2007" ( KOM(2008)0338 ),
–
med beaktande av kommissionens årsrapport om de internrevisioner som genomförts under 2007, riktad till den myndighet som beviljar ansvarsfrihet ( KOM(2008)0499 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2008)2361 ),
–
med beaktande av kommissionens rapport om medlemsstaternas svar på revisionsrättens årsrapport 2006 ( KOM(2008)0112 ),
–
med beaktande av grönboken om det europeiska öppenhetsinitiativet som antogs av kommissionen den 3 maj 2006 ( KOM(2006)0194 ),
–
,
–
med beaktande av kommissionens meddelande om en färdplan för en integrerad ram för intern kontroll ( KOM(2005)0252 ),
–
med beaktande av kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2006)0009 ), kommissionens lägesrapport till rådet, Europaparlamentet och Europeiska revisionsrätten om kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2007)0086 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer rapporten ( SEK(2007)0311 ),
–
med beaktande av den första resultattavlan för genomförandet av kommissionens handlingsplan för en integrerad ram för intern kontroll, offentliggjord den 19 juli 2006 ( SEK(2006)1009 ), i enlighet med parlamentets begäran i resolutionen som åtföljde beslutet om ansvarsfrihet för budgetåret 2004,
–
med beaktande av revisionsrättens yttrande nr 6/2007 över medlemsstaternas årliga sammanfattningar, medlemsstaternas nationella förklaringar och nationella revisionsorgans revisionsarbete rörande EU-medel EUT C 216, 14.9.2007, s.
3.
,
–
med beaktande av kommissionens handlingsplan för att stärka kommissionens tillsynsfunktion vid delad förvaltning av strukturåtgärder ( KOM(2008)0097 ),
–
med beaktande av meddelandet från kommissionens ledamöter Danuta Hübner och Vladimír Špidla till kommissionen med en lägesrapport om genomförandet av handlingsplanen för att stärka kommissionens tillsynsfunktion vid delad förvaltning av strukturåtgärder ( SEK(2008)2756 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer detta meddelande ( SEK(2008)2755 ),
–
med beaktande av kommissionens rapport till Europaparlamentet, rådet och Europeiska revisionsrätten om kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2008)0110 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2008)0259 ),
–
med beaktande av revisionsrättens årsrapport om genomförandet av budgeten för budgetåret 2007 EUT C 286, 10.11.2008, s.
1.
och dess särskilda rapporter, samt de granskade institutionernas svar,
–
med beaktande av den revisionsförklaring om räkenskapernas tillförlitlighet och de underliggande transaktionernas laglighet och korrekthet som avges av revisionsrätten i enlighet med artikel 248 i EG-fördraget EUT C 287, 10.11.2008, s.
111.
,
–
med beaktande av kommissionens meddelande av den 16 december 2008 med titeln "Mot en samsyn på begreppet acceptabel risk" ( KOM(2008)0866 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer detta meddelande ( SEK(2008)3054 ),
–
med beaktande av rådets rekommendation av den 10 februari 2009 om beviljande av ansvarsfrihet för kommissionen för genomförandet av budgeten för budgetåret 2007 (5587/2009 – C6-0055/2009 ),
–
med beaktande av artiklarna 274, 275 och 276 i EG-fördraget samt artiklarna 179a och 180b i Euratomfördraget,
–
med beaktande av artikel 246 och följande artiklar om revisionsrätten i EG-fördraget,
–
med beaktande av internationella revisionsstandarder och internationella redovisningsstandarder, särskilt dem som avser den offentliga sektorn,
–
med beaktande av revisionsrättens internationella sakkunnighetsbedömning,
–
med beaktande av rådets förordning (EEG, Euratom, EKSG) nr 259/68 av den 29 februari 1968 om fastställande av tjänsteföreskrifter för tjänstemännen i Europeiska gemenskaperna och anställningsvillkor för övriga anställda i dessa gemenskaper EGT L 56, 4.3.1968, s.
1.
, särskilt avdelning V, kapitel 3 om pensioner och invaliditetspension och bilaga XII om genomförandebestämmelserna i artikel 83a i tjänsteföreskrifterna,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
, särskilt artiklarna 145, 146 och 147,
–
med beaktande av artikel 70 och bilaga V i arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet och yttrandena från övriga berörda utskott ( A6–0168/2009 ), och av följande skäl:
A.
I enlighet med artikel 274 i EG-fördraget ska kommissionen genomföra budgeten under eget ansvar i överensstämmelse med principerna för en sund ekonomisk förvaltning.
1.
Europaparlamentet beviljar kommissionen ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2007.
2.
Europaparlamentet redovisar sina iakttagelser i resolutionen nedan, som utgör en del av besluten om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2007, avsnitt III – kommissionen och genomförandeorgan.
3.
Europaparlamentet uppdrar åt talmannen att översända detta beslut och den resolution som utgör en del av beslutet till rådet, kommissionen, domstolen, revisionsrätten och Europeiska investeringsbanken samt till medlemsstaternas nationella och regionala revisionsorgan och att se till att de offentliggörs i Europeiska unionens officiella tidning (L-serien).
2.
Europaparlamentets beslut av den 23 april 2009 om ansvarsfrihet för genomförandet av budgeten för genomförandeorganet för utbildning, audiovisuella medier och kultur för budgetåret 2007 ( SEK(2008)2359 – C6-0415/2008 – 2008/2186(DEC) )
Europaparlamentet fattar detta beslut
–
,
–
med beaktande av Europeiska gemenskapernas slutliga årsredovisning för budgetåret 2007 – Volym I ( SEK(2008)2359 – C6-0415/2008 ) EUT C 287, 10.11.2008, s.
1.
,
–
med beaktande av den slutliga årsredovisningen för genomförandeorganet för utbildning, audiovisuella medier och kultur för budgetåret 2007 EUT C 278, 31.10.2008, s.
32.
,
–
med beaktande av kommissionens årsrapporter till Europaparlamentet och rådet om uppföljningen av besluten om ansvarsfrihet 2006 ( KOM(2008)0629 och KOM(2008)0628 ) samt av de arbetsdokument från kommissionens tjänsteavdelningar som åtföljer dessa rapporter ( SEK(2008)2579 och SEK(2008)2580 ),
–
med beaktande av kommissionens meddelande med titeln "Sammanfattande rapport om kommissionens förvaltning 2007" ( KOM(2008)0338 ),
–
med beaktande av kommissionens årsrapport om de internrevisioner som genomförts under 2007, riktad till den myndighet som beviljar ansvarsfrihet ( KOM(2008)0499 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2008)2361 ),
–
med beaktande av kommissionens rapport om medlemsstaternas svar på revisionsrättens årsrapport 2006 ( KOM(2008)0112 ),
–
med beaktande av grönboken om det europeiska öppenhetsinitiativet som antogs av kommissionen den 3 maj 2006 ( KOM(2006)0194 ),
–
,
–
med beaktande av kommissionens meddelande om en färdplan för en integrerad ram för intern kontroll ( KOM(2005)0252 ),
–
med beaktande av kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2006)0009 ), kommissionens lägesrapport till rådet, Europaparlamentet och Europeiska revisionsrätten om kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2007)0086 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2007)0311 ),
–
med beaktande av den första resultattavlan för genomförandet av kommissionens handlingsplan för en integrerad ram för intern kontroll, offentliggjord den 19 juli 2006 ( SEK(2006)1009 ), i enlighet med parlamentets begäran i resolutionen som åtföljde beslutet om ansvarsfrihet för budgetåret 2004,
–
med beaktande av revisionsrättens yttrande nr 6/2007 över medlemsstaternas årliga sammanfattningar, medlemsstaternas nationella förklaringar och nationella revisionsorgans revisionsarbete rörande EU-medel EUT C 216, 14.9.2007, s.
3.
,
–
med beaktande av kommissionens handlingsplan för att stärka kommissionens tillsynsfunktion vid delad förvaltning av strukturåtgärder ( KOM(2008)0097 ),
–
med beaktande av meddelandet från kommissionens ledamöter Danuta Hübner och Vladimír Špidla till kommissionen med en lägesrapport om genomförandet av handlingsplanen för att stärka kommissionens tillsynsfunktion vid delad förvaltning av strukturåtgärder ( SEK(2008)2756 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer detta meddelande ( SEK(2008)2755 ),
–
med beaktande av kommissionens rapport till Europaparlamentet, rådet och Europeiska revisionsrätten om kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2008)0110 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2008)0259 ),
–
med beaktande av revisionsrättens rapport om årsredovisningen för genomförandeorganet för utbildning, audiovisuella medier och kultur för budgetåret 2007 samt genomförandeorganets svar EUT C 311, 5.12.2008, s.
71.
,
–
med beaktande av den revisionsförklaring om räkenskapernas tillförlitlighet och de underliggande transaktionernas laglighet och korrekthet som avges av revisionsrätten i enlighet med artikel 248 i EG-fördraget EUT C 287, 10.11.2008, s.
111.
,
–
med beaktande av kommissionens meddelande av den 16 december 2008 med titeln "Mot en samsyn på begreppet acceptabel risk" ( KOM(2008)0866 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer detta meddelande ( SEK(2008)3054 ),
–
med beaktande av rådets rekommendation av den 10 februari 2009 om beviljande av ansvarsfrihet för genomförandeorganen för genomförandet av budgeten för budgetåret 2007 (5589/2009 – C6-0056/2009 ),
–
med beaktande av artiklarna 274, 275 och 276 i EG-fördraget samt artiklarna 179a och 180b i Euratomfördraget,
–
med beaktande av artikel 246 och följande artiklar om revisionsrätten i EG-fördraget,
–
med beaktande av internationella revisionsstandarder och internationella redovisningsstandarder, särskilt dem som avser den offentliga sektorn,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
, särskilt artiklarna 145, 146 och 147,
–
med beaktande av rådets förordning (EG) nr 58/2003 av den 19 december 2002 om stadgar för de genomförandeorgan som ansvarar för vissa uppgifter som avser förvaltningen av gemenskapsprogram EGT L 11, 16.1.2003, s.
1.
–
med beaktande av kommissionens förordning (EG) nr 1653/2004 av den 21 september 2004 om standardbudgetförordning för genomförandeorgan enligt rådets förordning (EG) nr 58/2003 om stadgar för genomförandeorgan som ansvarar för vissa uppgifter som avser förvaltning av gemenskapsprogram EUT L 297, 22.9.2004, s.
6.
–
med beaktande av kommissionens beslut 2005/56/EG av den 14 januari 2005 om inrättande av "Genomförandeorganet för utbildning, audiovisuella medier och kultur" för att förvalta gemenskapsprogram inom utbildning, audiovisuella medier och kultur enligt rådets förordning (EG) nr 58/2003 EUT L 24, 27.1.2005, s.
35.
,
–
med beaktande av artikel 70 och bilaga V i arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet och yttrandena från övriga berörda utskott ( A6–0168/2009 ), och av följande skäl:
A.
I enlighet med artikel 274 i EG-fördraget ska kommissionen genomföra budgeten under eget ansvar i överensstämmelse med principerna för en sund ekonomisk förvaltning.
1.
Europaparlamentet beviljar ansvarsfrihet för direktören för genomförandeorganet för utbildning, audiovisuella medier och kultur avseende genomförandet av genomförandeorganets budget för budgetåret 2007.
2.
Europaparlamentet redovisar sina iakttagelser i resolutionen nedan, som utgör en del av besluten om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2007, avsnitt III – kommissionen och genomförandeorgan.
3.
Europaparlamentet uppdrar åt talmannen att översända detta beslut om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2007, avsnitt III – kommissionen och den resolution som utgör en del av beslutet till direktören för genomförandeorganet för utbildning, audiovisuella medier och kultur, rådet, kommissionen, domstolen och revisionsrätten samt att se till att de offentliggörs i Europeiska unionens officiella tidning (L-serien).
3.
Europaparlamentets beslut av den 23 april 2009 om ansvarsfrihet för genomförandet av budgeten för genomförandeorganet för konkurrenskraft och innovation för budgetåret 2007 ( SEK(2008)2359 – C6-0415/2008 – 2008/2186(DEC) )
Europaparlamentet fattar detta beslut
–
,
–
med beaktande av Europeiska gemenskapernas slutliga årsredovisning för budgetåret 2007 – Volym I ( SEK(2008)2359 – C6-0415/2008 ) EUT C 287, 10.11.2008, s.
1.
,
–
med beaktande av den slutliga årsredovisningen för genomförandeorganet för konkurrenskraft och innovation för budgetåret 2007 EUT C 278, 31.10.2008, s.
29.
,
–
med beaktande av kommissionens årsrapporter till Europaparlamentet och rådet om uppföljningen av besluten om ansvarsfrihet 2006 ( KOM(2008)0629 och KOM(2008)0628 ) samt av de arbetsdokument från kommissionens tjänsteavdelningar som åtföljer dessa rapporter ( SEK(2008)2579 och SEK(2008)2580 ),
–
med beaktande av kommissionens meddelande med titeln "Sammanfattande rapport om kommissionens förvaltning 2007" ( KOM(2008)0338 ),
–
med beaktande av kommissionens årsrapport om de internrevisioner som genomförts under 2007, riktad till den myndighet som beviljar ansvarsfrihet ( KOM(2008)0499 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2008)2361 ),
–
med beaktande av kommissionens rapport om medlemsstaternas svar på revisionsrättens årsrapport 2006 ( KOM(2008)0112 ),
–
med beaktande av grönboken om det europeiska öppenhetsinitiativet som antogs av kommissionen den 3 maj 2006 ( KOM(2006)0194 ),
–
,
–
med beaktande av kommissionens meddelande om en färdplan för en integrerad ram för intern kontroll ( KOM(2005)0252 ),
–
med beaktande av kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2006)0009 ), kommissionens lägesrapport till rådet, Europaparlamentet och Europeiska revisionsrätten om kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2007)0086 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2007)0311 ),
–
med beaktande av den första resultattavlan för genomförandet av kommissionens handlingsplan för en integrerad ram för intern kontroll, offentliggjord den 19 juli 2006 ( SEK(2006)1009 ), i enlighet med parlamentets begäran i resolutionen som åtföljde beslutet om ansvarsfrihet för budgetåret 2004,
–
med beaktande av revisionsrättens yttrande nr 6/2007 över medlemsstaternas årliga sammanfattningar, medlemsstaternas nationella förklaringar och nationella revisionsorgans revisionsarbete rörande EU-medel EUT C 216, 14.9.2007, s.
3.
,
–
med beaktande av kommissionens handlingsplan för att stärka kommissionens tillsynsfunktion vid delad förvaltning av strukturåtgärder ( KOM(2008)0097 ),
–
med beaktande av meddelandet från kommissionens ledamöter Danuta Hübner och Vladimír Špidla till kommissionen med en lägesrapport om genomförandet av handlingsplanen för att stärka kommissionens tillsynsfunktion vid delad förvaltning av strukturåtgärder ( SEK(2008)2756 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer detta meddelande ( SEK(2008)2755 ),
–
med beaktande av kommissionens rapport till Europaparlamentet, rådet och Europeiska revisionsrätten om kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2008)0110 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2008)0259 ),
–
med beaktande av revisionsrättens rapport om årsredovisningen för genomförandeorganet för konkurrenskraft och innovation för budgetåret 2007 samt genomförandeorganets svar EUT C 311, 5.12.2008, s.
79.
,
–
med beaktande av den revisionsförklaring om räkenskapernas tillförlitlighet och de underliggande transaktionernas laglighet och korrekthet som avges av revisionsrätten i enlighet med artikel 248 i EG-fördraget EUT C 287, 10.11.2008, s.
111.
,
–
med beaktande av kommissionens meddelande av den 16 december 2008 med titeln "Mot en samsyn på begreppet acceptabel risk" ( KOM(2008)0866 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer detta meddelande ( SEK(2008)3054 ),
–
med beaktande av rådets rekommendation av den 10 februari 2009 om beviljande av ansvarsfrihet för genomförandeorganen för genomförandet av budgeten för budgetåret 2007 (5589/2009 – C6-0056/2009 ),
–
med beaktande av artiklarna 274, 275 och 276 i EG-fördraget samt artiklarna 179a och 180b i Euratomfördraget,
–
med beaktande av artikel 246 och följande artiklar om revisionsrätten i EG-fördraget,
–
med beaktande av internationella revisionsstandarder och internationella redovisningsstandarder, särskilt dem som avser den offentliga sektorn,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
, särskilt artiklarna 145, 146 och 147,
–
med beaktande av rådets förordning (EG) nr 58/2003 av den 19 december 2002 om stadgar för de genomförandeorgan som ansvarar för vissa uppgifter som avser förvaltningen av gemenskapsprogram EGT L 11, 16.1.2003, s.
1.
–
med beaktande av kommissionens förordning (EG) nr 1653/2004 av den 21 september 2004 om standardbudgetförordning för genomförandeorgan enligt rådets förordning (EG) nr 58/2003 om stadgar för genomförandeorgan som ansvarar för vissa uppgifter som avser förvaltning av gemenskapsprogram EUT L 297, 22.9.2004, s.
6.
–
85.
,
–
med beaktande av kommissionens beslut 2007/372/EG av den 31 maj 2007 om ändring av beslut 2004/20/EG för att ändra Exekutiva byrån för intelligent energi till genomförandeorganet för konkurrenskraft och innovation EUT L 140, 1.6.2007, s.
–
med beaktande av artikel 70 och bilaga V i arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet och yttrandena från övriga berörda utskott ( A6–0168/2009 ), och av följande skäl:
A.
I enlighet med artikel 274 i EG-fördraget ska kommissionen genomföra budgeten under eget ansvar i överensstämmelse med principerna för en sund ekonomisk förvaltning.
1.
Europaparlamentet beviljar ansvarsfrihet för direktören för genomförandeorganet för konkurrenskraft och innovation avseende genomförandet av genomförandeorganets budget för budgetåret 2007.
2.
Europaparlamentet redovisar sina iakttagelser i resolutionen nedan, som utgör en del av besluten om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2007, avsnitt III – kommissionen och genomförandeorgan.
3.
Europaparlamentet uppdrar åt talmannen att översända detta beslut om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2007, avsnitt III – kommissionen och den resolution som utgör en del av beslutet till direktören för genomförandeorganet för konkurrenskraft och innovation, rådet, kommissionen, domstolen och revisionsrätten samt att se till att de offentliggörs i Europeiska unionens officiella tidning (L-serien).
4.
Europaparlamentets beslut av den 23 april 2009 om ansvarsfrihet för genomförandet av budgeten för genomförandeorganet för folkhälsoprogrammet för budgetåret 2007 ( SEK(2008)2359 – C6-0415/2008 – 2008/2186(DEC) )
Europaparlamentet fattar detta beslut
–
,
–
med beaktande av Europeiska gemenskapernas slutliga årsredovisning för budgetåret 2007 – Volym I ( SEK(2008)2359 – C6-0415/2008 ) EUT C 287, 10.11.2008, s.
1.
,
–
med beaktande av den slutliga årsredovisningen för genomförandeorganet för folkhälsoprogrammet för budgetåret 2007 EUT C 278, 31.10.2008, s.
81.
,
–
med beaktande av kommissionens årsrapporter till Europaparlamentet och rådet om uppföljningen av besluten om ansvarsfrihet 2006 ( KOM(2008)0629 och KOM(2008)0628 ) samt av de arbetsdokument från kommissionens tjänsteavdelningar som åtföljer dessa rapporter ( SEK(2008)2579 och SEK(2008)2580 ),
–
med beaktande av kommissionens meddelande med titeln "Sammanfattande rapport om kommissionens förvaltning 2007" ( KOM(2008)0338 ),
–
med beaktande av kommissionens årsrapport om de internrevisioner som genomförts under 2007, riktad till den myndighet som beviljar ansvarsfrihet ( KOM(2008)0499 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2008)2361 ),
–
med beaktande av kommissionens rapport om medlemsstaternas svar på revisionsrättens årsrapport 2006 ( KOM(2008)0112 ),
–
med beaktande av grönboken om det europeiska öppenhetsinitiativet som antogs av kommissionen den 3 maj 2006 ( KOM(2006)0194 ),
–
,
–
med beaktande av kommissionens meddelande om en färdplan för en integrerad ram för intern kontroll ( KOM(2005)0252 ),
–
med beaktande av kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2006)0009 ), kommissionens lägesrapport till rådet, Europaparlamentet och Europeiska revisionsrätten om kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2007)0086 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2007)0311 ),
–
med beaktande av den första resultattavlan för genomförandet av kommissionens handlingsplan för en integrerad ram för intern kontroll, offentliggjord den 19 juli 2006 ( SEK(2006)1009 ), i enlighet med parlamentets begäran i resolutionen som åtföljde beslutet om ansvarsfrihet för budgetåret 2004,
–
med beaktande av revisionsrättens yttrande nr 6/2007 över medlemsstaternas årliga sammanfattningar, medlemsstaternas nationella förklaringar och nationella revisionsorgans revisionsarbete rörande EU-medel EUT C 216, 14.9.2007, s.
3.
,
–
med beaktande av kommissionens handlingsplan för att stärka kommissionens tillsynsfunktion vid delad förvaltning av strukturåtgärder ( KOM(2008)0097 ),
–
med beaktande av meddelandet från kommissionens ledamöter Danuta Hübner och Vladimír Špidla till kommissionen med en lägesrapport om genomförandet av handlingsplanen för att stärka kommissionens tillsynsfunktion vid delad förvaltning av strukturåtgärder ( SEK(2008)2756 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer detta meddelande ( SEK(2008)2755 ),
–
med beaktande av kommissionens rapport till Europaparlamentet, rådet och Europeiska revisionsrätten om kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2008)0110 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2008)0259 ),
–
med beaktande av revisionsrättens rapport om årsredovisningen för genomförandeorganet för folkhälsoprogrammet för budgetåret 2007 samt genomförandeorganets svar EUT C 311, 5.12.2008, s.
86.
,
–
med beaktande av den revisionsförklaring om räkenskapernas tillförlitlighet och de underliggande transaktionernas laglighet och korrekthet som avges av revisionsrätten i enlighet med artikel 248 i EG-fördraget EUT C 287, 10.11.2008, s.
111.
,
–
med beaktande av kommissionens meddelande av den 16 december 2008 med titeln "Mot en samsyn på begreppet acceptabel risk" ( KOM(2008)0866 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer detta meddelande ( SEK(2008)3054 ),
–
med beaktande av rådets rekommendation av den 10 februari 2009 om beviljande av ansvarsfrihet för genomförandeorganen för genomförandet av budgeten för budgetåret 2007 (5589/2009 – C6-0056/2009 ),
–
med beaktande av artiklarna 274, 275 och 276 i EG-fördraget samt artiklarna 179a och 180b i Euratomfördraget,
–
med beaktande av artikel 246 och följande artiklar om revisionsrätten i EG-fördraget,
–
med beaktande av internationella revisionsstandarder och internationella redovisningsstandarder, särskilt dem som avser den offentliga sektorn,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
, särskilt artiklarna 145, 146 och 147,
–
med beaktande av rådets förordning (EG) nr 58/2003 av den 19 december 2002 om stadgar för de genomförandeorgan som ansvarar för vissa uppgifter som avser förvaltningen av gemenskapsprogram EGT L 11, 16.1.2003, s.
1.
–
med beaktande av kommissionens förordning (EG) nr 1653/2004 av den 21 september 2004 om standardbudgetförordning för genomförandeorgan enligt rådets förordning (EG) nr 58/2003 om stadgar för genomförandeorgan som ansvarar för vissa uppgifter som avser förvaltning av gemenskapsprogram EUT L 297, 22.9.2004, s.
6.
–
med beaktande av kommissionens beslut 2004/858/EG av den 15 december 2004 om inrättandet av ett genomförandeorgan med namnet "Genomförandeorgan för folkhälsoprogrammet" för förvaltning av gemenskapsåtgärder inom folkhälsoområdet – med tillämpning av rådets förordning (EG) nr 58/2003 EGT L 369, 16.12.2004, s.
73.
,
–
med beaktande av artikel 70 och bilaga V i arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet och yttrandena från övriga berörda utskott ( A6–0168/2009 ), och av följande skäl:
A.
I enlighet med artikel 274 i EG-fördraget ska kommissionen genomföra budgeten under eget ansvar i överensstämmelse med principerna för en sund ekonomisk förvaltning.
1.
Europaparlamentet beviljar ansvarsfrihet för direktören för genomförandeorganet för folkhälsoprogrammet avseende genomförandet av genomförandeorganets budget för budgetåret 2007.
2.
Europaparlamentet redovisar sina iakttagelser i resolutionen nedan, som utgör en del av besluten om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2007, avsnitt III – kommissionen och genomförandeorgan.
3.
Europaparlamentet uppdrar åt talmannen att översända detta beslut om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2007, avsnitt III – kommissionen och den resolution som utgör en del av beslutet till direktören för genomförandeorganet för hälso- och konsumentfrågor (tidigare genomförandeorganet för folkhälsoprogrammet), rådet, kommissionen, domstolen och revisionsrätten samt att se till att de offentliggörs i Europeiska unionens officiella tidning (L-serien).
5.
Europaparlamentets beslut av den 23 april 2009 om avslutande av räkenskaperna avseende genomförandet av Europeiska unionens allmänna budget för budgetåret 2007, avsnitt III – kommissionen ( SEK(2008)2359 – C6-0415/2008 – 2008/2186(DEC) )
Europaparlamentet fattar detta beslut
–
,
–
med beaktande av Europeiska gemenskapernas slutliga årsredovisning för budgetåret 2007 – Volym I ( SEK(2008)2359 – C6-0415/2008 ) EUT C 287, 10.11.2008, s.
1.
,
–
med beaktande av kommissionens årsrapporter till Europaparlamentet och rådet om uppföljningen av besluten om ansvarsfrihet 2006 ( KOM(2008)0629 och KOM(2008)0628 ) samt av de arbetsdokument från kommissionens tjänsteavdelningar som åtföljer dessa rapporter ( SEK(2008)2579 och SEK(2008)2580 ),
–
med beaktande av kommissionens meddelande med titeln "Sammanfattande rapport om kommissionens förvaltning 2007" ( KOM(2008)0338 ),
–
med beaktande av kommissionens årsrapport om de internrevisioner som genomförts under 2007, riktad till den myndighet som beviljar ansvarsfrihet ( KOM(2008)0499 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2008)2361 ),
–
med beaktande av kommissionens rapport om medlemsstaternas svar på revisionsrättens årsrapport 2006 ( KOM(2008)0112 ),
–
med beaktande av grönboken om det europeiska öppenhetsinitiativet som antogs av kommissionen den 3 maj 2006 ( KOM(2006)0194 ),
–
,
–
med beaktande av kommissionens meddelande om en färdplan för en integrerad ram för intern kontroll ( KOM(2005)0252 ),
–
med beaktande av kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2006)0009 ), kommissionens lägesrapport till rådet, Europaparlamentet och Europeiska revisionsrätten om kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2007)0086 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2007)0311 ),
–
med beaktande av den första resultattavlan för genomförandet av kommissionens handlingsplan för en integrerad ram för intern kontroll, offentliggjord den 19 juli 2006 ( SEK(2006)1009 ), i enlighet med parlamentets begäran i resolutionen som åtföljde beslutet om ansvarsfrihet för budgetåret 2004,
–
med beaktande av revisionsrättens yttrande nr 6/2007 över medlemsstaternas årliga sammanfattningar, medlemsstaternas nationella förklaringar och nationella revisionsorgans revisionsarbete rörande EU-medel EUT C 216, 14.9.2007, s.
3.
,
–
med beaktande av kommissionens handlingsplan för att stärka kommissionens tillsynsfunktion vid delad förvaltning av strukturåtgärder ( KOM(2008)0097 ),
–
med beaktande av meddelandet från kommissionens ledamöter Danuta Hübner och Vladimír Špidla till kommissionen med en lägesrapport om genomförandet av handlingsplanen för att stärka kommissionens tillsynsfunktion vid delad förvaltning av strukturåtgärder ( SEK(2008)2756 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer detta meddelande ( SEK(2008)2755 ),
–
med beaktande av kommissionens rapport till Europaparlamentet, rådet och Europeiska revisionsrätten om kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2008)0110 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2008)0259 ),
–
med beaktande av revisionsrättens årsrapport om genomförandet av budgeten för budgetåret 2007 EUT C 286, 10.11.2008, s.
1.
och dess särskilda rapporter, samt de granskade institutionernas svar,
–
med beaktande av den revisionsförklaring om räkenskapernas tillförlitlighet och de underliggande transaktionernas laglighet och korrekthet som avges av revisionsrätten i enlighet med artikel 248 i EG-fördraget EUT C 287, 10.11.2008, s.
111.
,
–
med beaktande av kommissionens meddelande av den 16 december 2008 med titeln "Mot en samsyn på begreppet acceptabel risk" ( KOM(2008)0866 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer detta meddelande ( SEK(2008)3054 ),
–
med beaktande av rådets rekommendation av den 10 februari 2009 om beviljande av ansvarsfrihet för kommissionen för genomförandet av budgeten för budgetåret 2007 (5587/2009 – C6-0055/2009 ),
–
med beaktande av artiklarna 274, 275 och 276 i EG-fördraget samt artiklarna 179a och 180b i Euratomfördraget,
–
med beaktande av artikel 246 och följande artiklar om revisionsrätten i EG-fördraget,
–
med beaktande av internationella revisionsstandarder och internationella redovisningsstandarder, särskilt dem som avser den offentliga sektorn,
–
med beaktande av revisionsrättens internationella sakkunnighetsbedömning,
–
med beaktande av rådets förordning (EEG, Euratom, EKSG) nr 259/68 av den 29 februari 1968 om fastställande av tjänsteföreskrifter för tjänstemännen i Europeiska gemenskaperna och anställningsvillkor för övriga anställda i dessa gemenskaper EGT L 56, 4.3.1968, s.
1.
, särskilt avdelning V, kapitel 3 om pensioner och invaliditetspension och bilaga XII om genomförandebestämmelserna i artikel 83a i tjänsteföreskrifterna,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
, särskilt artiklarna 145, 146 och 147,
–
med beaktande av rådets förordning (EG) nr 58/2003 av den 19 december 2002 om stadgar för de genomförandeorgan som ansvarar för vissa uppgifter som avser förvaltningen av gemenskapsprogram EGT L 11, 16.1.2003, s.
1.
–
med beaktande av artikel 70 och bilaga V i arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet och yttrandena från övriga berörda utskott ( A6–0168/2009 ), och av följande skäl:
A.
I enlighet med artikel 275 i EG-fördraget är kommissionen behörig att redovisa räkenskaperna.
1.
Europaparlamentet godkänner avslutandet av räkenskaperna avseende genomförandet av Europeiska unionens allmänna budget för budgetåret 2007.
2.
Europaparlamentet redovisar sina iakttagelser i resolutionen nedan, som utgör en del av besluten om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2007, avsnitt III – kommissionen och genomförandeorgan.
3.
Europaparlamentet uppdrar åt talmannen att översända detta beslut till rådet, kommissionen, domstolen, revisionsrätten och Europeiska investeringsbanken samt till de nationella parlamenten och medlemsstaternas nationella och regionala revisionsorgan och att se till att de offentliggörs i Europeiska unionens officiella tidning (L-serien).
6.
Europaparlamentets resolution av den 23 april 2009 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2007, avsnitt III – kommissionen och genomförandeorgan ( SEK(2008)2359 – C6-0415/2008 – 2008/2186(DEC) )
Europaparlamentet utfärdar denna resolution
–
,
–
med beaktande av Europeiska gemenskapernas slutliga årsredovisning för budgetåret 2007 – Volym I ( SEK(2008)2359 – C6-0415/2008 ) EUT C 287, 10.11.2008, s.
1.
,
–
med beaktande av kommissionens årsrapporter till Europaparlamentet och rådet om uppföljningen av besluten om ansvarsfrihet 2006 ( KOM(2008)0629 och KOM(2008)0628 ) samt av de arbetsdokument från kommissionens tjänsteavdelningar som åtföljer dessa rapporter ( SEK(2008)2579 och SEK(2008)2580 ),
–
med beaktande av kommissionens meddelande med titeln "Sammanfattande rapport om kommissionens förvaltning 2007" ( KOM(2008)0338 ),
–
med beaktande av kommissionens årsrapport om de internrevisioner som genomförts under 2007, riktad till den myndighet som beviljar ansvarsfrihet ( KOM(2008)0499 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2008)2361 ),
–
med beaktande av kommissionens rapport om medlemsstaternas svar på revisionsrättens årsrapport 2006 ( KOM(2008)0112 ),
–
med beaktande av grönboken om det europeiska öppenhetsinitiativet som antogs av kommissionen den 3 maj 2006 ( KOM(2006)0194 ),
–
,
–
med beaktande av kommissionens meddelande om en färdplan för en integrerad ram för intern kontroll ( KOM(2005)0252 ),
–
med beaktande av kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2006)0009 ), kommissionens lägesrapport till rådet, Europaparlamentet och Europeiska revisionsrätten om kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2007)0086 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2007)0311 ),
–
med beaktande av den första resultattavlan för genomförandet av kommissionens handlingsplan för en integrerad ram för intern kontroll, offentliggjord den 19 juli 2006 ( SEK(2006)1009 ), i enlighet med parlamentets begäran i resolutionen som åtföljde beslutet om ansvarsfrihet för budgetåret 2004,
–
med beaktande av revisionsrättens yttrande nr 6/2007 över medlemsstaternas årliga sammanfattningar, medlemsstaternas nationella förklaringar och nationella revisionsorgans revisionsarbete rörande EU-medel EUT C 216, 14.9.2007, s.
3.
,
–
med beaktande av kommissionens handlingsplan för att stärka kommissionens tillsynsfunktion vid delad förvaltning av strukturåtgärder ( KOM(2008)0097 ),
–
med beaktande av meddelandet från kommissionens ledamöter Danuta Hübner och Vladimír Špidla till kommissionen med en lägesrapport om genomförande av handlingsplanen för att stärka kommissionens tillsynsfunktion vid delad förvaltning av strukturåtgärder ( SEK(2008)2756 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer detta meddelande ( SEK(2008)2755 ),
–
med beaktande av kommissionens rapport till Europaparlamentet, rådet och Europeiska revisionsrätten om kommissionens handlingsplan för en integrerad ram för intern kontroll ( KOM(2008)0110 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer denna rapport ( SEK(2008)0259 ),
–
med beaktande av revisionsrättens årsrapport om genomförandet av budgeten för budgetåret 2007 EUT C 286, 10.11.2008, s.
1.
och dess särskilda rapporter, samt de granskade institutionernas svar,
–
med beaktande av den revisionsförklaring om räkenskapernas tillförlitlighet och de underliggande transaktionernas laglighet och korrekthet som avges av revisionsrätten i enlighet med artikel 248 i EG-fördraget EUT C 287, 10.11.2008, s.
111.
,
–
med beaktande av kommissionens meddelande av den 16 december 2008 med titeln "Mot en samsyn på begreppet acceptabel risk" ( KOM(2008)0866 ) och det arbetsdokument från kommissionens tjänsteavdelningar som åtföljer detta meddelande ( SEK(2008)3054 ),
–
med beaktande av rådets rekommendation av den 10 februari 2009 om beviljande av ansvarsfrihet för kommissionen för genomförandet av budgeten för budgetåret 2007 (5587/2009 – C6-0055/2009 ),
–
med beaktande av rådets rekommendation av den 10 februari 2009 om beviljande av ansvarsfrihet för genomförandeorganen för genomförandet av budgeten för budgetåret 2007 (5589/2009 – C6-0056/2009 ),
–
med beaktande av artiklarna 274, 275 och 276 i EG-fördraget samt artiklarna 179a och 180b i Euratomfördraget,
–
med beaktande av artikel 246 och följande artiklar om revisionsrätten i EG-fördraget,
–
med beaktande av internationella revisionsstandarder och internationella redovisningsstandarder, särskilt dem som avser den offentliga sektorn,
–
med beaktande av revisionsrättens internationella sakkunnighetsbedömning,
–
med beaktande av rådets förordning (EEG, Euratom, EKSG) nr 259/68 av den 29 februari 1968 om fastställande av tjänsteföreskrifter för tjänstemännen i Europeiska gemenskaperna och anställningsvillkor för övriga anställda i dessa gemenskaper EGT L 56, 4.3.1968, s.
1.
, särskilt avdelning V, kapitel 3 om pensioner och invaliditetspension och bilaga XII om genomförandebestämmelserna i artikel 83a i tjänsteföreskrifterna,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
, särskilt artiklarna 145, 146 och 147 i denna,
–
med beaktande av rådets förordning (EG) nr 58/2003 av den 19 december 2002 om stadgar för de genomförandeorgan som ansvarar för vissa uppgifter som avser förvaltningen av gemenskapsprogram EGT L 11, 16.1.2003, s.
1.
–
med beaktande av artikel 70 och bilaga V i arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet och yttrandena från övriga berörda utskott ( A6–0168/2009 ), och av följande skäl:
A.
Enligt artikel 274 i EG-fördraget åligger ansvaret för genomförandet av gemenskapsbudgeten kommissionen, som ska genomföra budgeten i överensstämmelse med principerna för en sund ekonomisk förvaltning i samarbete med medlemsstaterna.
B.
C.
D.
Det verkar som om Europeiska gemenskapernas politiska makt över de gemenskapsbyråer som inte har genomförandeuppgifter, något som är en förutsättning för att deras budgetar ska konsolideras i gemenskapsbudgeten, utökas för varje år som går och deras plats i det politiska organisationsschemat för gemenskapens operativa strukturer blir allt svårare att skönja.
E.
Genomförandet av vissa av EU:s politikområden kännetecknas av "delad förvaltning" av gemenskapsbudgeten mellan kommissionen och medlemsstaterna, vilket innebär att omkring 80 procent av gemenskapsutgifterna förvaltas av medlemsstaterna.
F.
I sin resolution av den 24 april 2007 EUT L 187, 15.7.2008, s.
25.
om ansvarsfrihet för budgetåret 2005 ansåg Europarlamentet att varje medlemsstat måste kunna ta ansvar för de gemenskapsmedel som man tar emot, antingen genom en enda nationell förvaltningsförklaring eller genom flera förklaringar inom en nationell ram.
G.
I sin årsrapport om budgetåret 2007 underströk revisionsrätten i sin utvärdering av framstegen i införandet av en integrerad ram för intern kontroll att "EU-utgifternas karaktär innebär att risken för fel är störst hos den slutliga stödmottagaren" (punkt 1.47).
H.
De årliga sammanfattningar av revisioner och förklaringar från medlemsstaterna som finns tillgängliga på området för delad förvaltning i enlighet med punkt 44 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning EUT C 139, 14.6.2006, s.
I.
och revisionsrätten har förklarat att "alla kontrollsystem är en avvägning mellan å ena sidan kostnaden för att genomföra kontroller med den frekvens som fastställts, och å andra sidan den nytta dessa förfaranden innebär.
Inom gemenskapen handlar nyttan om att minska risken för att medel slösas bort, och att hålla risken för felaktigheter på en godtagbar nivå".
J.
I sin årsrapport 2007 ansåg revisionsrätten att "kontrollkostnaderna är en viktig fråga, både för EU:s budget och för medlemsstaterna" och att "balansen mellan kostnad och kvarstående risk när det gäller vissa utgiftsområden är av sådan betydelse att den bör godkännas på politisk nivå (det vill säga av budgetmyndigheten/den myndighet som beviljar ansvarsfrihet) i unionsmedborgarnas namn" (punkt 1.52 b och 1.52 c) och i punkt 2.42 c rekommenderade revisionsrätten att man skulle gå vidare med utvecklingen av begreppet tolererbar risk.
K.
I punkt 5 i slutsatserna från Ekofinrådets sammanträde den 8 november 2005 anges det att det att det är mycket viktigt att införa en integrerad ram för internkontroll och att förenkla lagstiftningen för kontrollerna och rådet uppmanade "kommissionen att bedöma kostnaden för kontroller per utgiftsområde".
L.
M.
Om det emellertid krävs en dialog mellan den externa revisorn (revisionsrätten) och det granskade organet (kommissionen) är det tveklöst upp till den externa revisorn att, i enlighet med de internationella revisionsstandarder som bör utgöra den övergripande ramen för budgetkontroll, bedöma de risker som får ligga till grund för valet av revisionsförfaranden.
N.
Dessutom beror kostnaderna för en kontroll inte bara på den godtagbara felfrekvensen utan även på komplexiteten i den granskade organisationen och kvaliteten på dess interna kontroll.
O.
P.
Q.
Det årliga förfarandet för att bevilja ansvarsfrihet ger parlamentet möjlighet att få direktkontakt med dem som har det främsta ansvaret för denna förvaltning och att mot bakgrund av resultaten av revisionsrättens granskning säkerställa en bättre förvaltning av EU:s utgifter för medborgarna och därmed skapa ett bättre beslutsunderlag.
R.
S.
I artikel 83 i förordning (EEG, Euratom, EKSG) nr 259/68 införs en kollektiv garanti från medlemsstaternas sida, vilket innebär att denna garanti kan inträda om en eller flera medlemsstater fallerar men detta betyder inte att gemenskaperna inte har en fordran gentemot de medlemsstater som ingått detta åtagande.
T.
2007 var det första året för genomförandet av instrumentet för utvecklingssamarbete.
U.
År 2007 var Europeiska året för lika möjligheter för alla, vilket riktade särskild uppmärksamhet på de olika former av diskriminering som kvinnor ofta möter.
V.
På grund av den bestående bristen på jämställdhet mellan män och kvinnor har användningen av budgetmedel olika effekter på dessa.
W.
Under nästa budgetförfarande bör rådet ta hänsyn till resultatet av och rekommendationerna i beslutet om ansvarsfrihet 2007 och stödja de reformförslag som syftar till att stärka medlemsstaternas ansvar i syfte att slutligt lösa de problem som revisionsrätten har påpekat i flera år.
X.
Kommissionen, rådet och parlamentet bör i samarbete med revisionsrätten fastställa som ett gemensamt mål att erhålla en positiv revisionsförklaring.
HUVUDSAKLIGA SLUTSATSER
1.
Europaparlamentet välkomnar de ytterligare framsteg som kommissionen och vissa av medlemsstaterna gjort mot en effektivare användning av gemenskapsmedel och den förbättrade övergripande kontrollen, vilket revisionsrätten påpekar i sin revisionsförklaring (DAS).
2.
3.
Europaparlamentet noterar att 2007 var det första året då fleråriga program från perioden 2000–2006 avslutades och att mycket medel återvanns.
4.
5.
6.
ÖVERGRIPANDE FRÅGOR
Revisionsförklaring (DAS)
7.
8.
Europaparlamentet välkomnar att revisionsrättens rapport visar att det inte finns några betydande fel i inkomster, administrativa utgifter, utgifter på området ekonomi och finans eller utgifter inom ramen för Europeiska garantifonden för jordbruket (EGFJ).
9.
Europaparlamentet konstaterar att situationen har förbättrats, särskilt i fråga om kontrollsystemen, men att detta inte är tillräckligt och att det går alltför långsamt.
Räkenskapernas tillförlitlighet
10.
11.
12.
Europaparlamentet förstår inte varför de tillgångar som Europeiska gemenskaperna har fått in i samband med Galileo-programmet inte redovisas i årsredovisningen.
13.
14.
Europaparlamentet begär att det när det saknas kapitalförbindelser bör göras en noggrann kontroll av att Europeiska gemenskapernas politiska inflytande i de organ som ingår i området för konsolideringen av räkenskaperna är förenligt med de villkor som anges i de internationella redovisningsstandarderna för den offentliga sektorn.
15.
Europaparlamentet uttrycker oro och tvivel kring möjligheten att utse högre tjänstemän "utanför kategori", såvida detta inte uttryckligen nämns i tjänsteförteckningen, under alla omständigheter i det sista steget av AD16, och uppmanar kommissionen att klarlägga möjligheterna enligt tjänsteföreskrifterna i ljuset av denna specifika budgetposition.
Lagligheten i de transaktioner som ligger till grund för räkenskaperna
16.
Europaparlamentet noterar med tillfredsställelse att det inte finns några väsentliga fel inom de områden där kommissionen har genomfört ändamålsenliga kontroll- och övervakningssystem (inkomster, åtaganden och betalningar när det gäller administrativa och andra utgifter samt ekonomi och finans) när det gäller lagligheten och korrektheten i de transaktioner som ligger till grund för räkenskaperna (kapitel 1 punkt IX i revisionsförklaringen).
17.
18.
Europaparlamentet uppmanar kommissionen att framför allt förstärka sin övervakning av de kontroller som delegerats till medlemsstaterna och att utfärda tydliga riktlinjer för att förhindra, identifiera och korrigera felaktigheter och kräver att kommissionen, när medlemsstaternas kontrollsystem är ineffektiva, vidtar alla åtgärder för att förmå medlemsstaterna att respektera sina förpliktelser och göra nödvändiga förbättringar, särskilt genom att ställa in betalningar och verkställa finansiella korrigeringar.
Budgetförvaltning – finansiella korrigeringar
19.
Europaparlamentet noterar att revisionsrätten konstaterar att jämfört med början av föregående programplaneringsperiod har utnyttjandet av åtaganden förbättrats tydligt under 2007, som är det första året av den nya programplaneringsperioden 2007–2013.
20.
Återvinningar
21.
22.
Europaparlamentet påpekar också att det är mycket viktigt att fatta beslut och vidta slutgiltiga korrigerande åtgärder för att utesluta utgifter som inte har verkställts i enlighet med gemenskapslagstiftningen ur gemenskapsfinansieringen och upprepar sitt krav på att det måste anges exakt vilken budgetrubrik och vilket år som de enskilda återvinningarna avser, i likhet med vad som görs för jordbruket och naturresurserna.
23.
24.
Europaparlamentet kräver med hänsyn till att problemen med återvinningar kvarstår att systemet utvärderas.
Uppskjutande av betalningar
25.
Europaparlamentet ger kommissionen sitt fulla stöd i dess stränga tillämpning av lagstiftningen om uppskjutande av betalningar och välkomnar de åtgärder som har vidtagits för att inga överföringar ska ske så länge kommissionen inte har fått absoluta garantier i fråga om tillförlitligheten i förvaltnings- och kontrollsystemet hos den medlemsstat som tar emot medlen i fråga.
Årliga sammanfattningar av revisioner, förklaringar som finns tillgängliga på området för delad förvaltning och nationella förvaltningsförklaringar
26.
27.
28.
I detta sammanhang begär Europaparlamentet att kommissionen analyserar de sammanfattningar som mottas 2009 i syfte att optimera deras mervärde när det gäller de garantier som ges för hur medlemsstaternas interna kontrollsystem fungerar.
29.
Europaparlamentet beklagar att kommissionen inte har följt parlamentets begäran i resolutionen av den 22 april 2008 om ansvarsfrihet för budgetåret 2006 EUT L 88, 31.3.2009, s.
25.
30.
31.
Kommissionen uppmanas att efter tre år utföra en fullständig utvärdering, med en analys av det mervärde som de årliga sammanfattningarna innebär för en sund ekonomisk förvaltning av EU-medel i medlemsstaterna, samt av graden av oberoende hos de berörda revisorerna.
32.
33.
Europaparlamentet välkomnar att några medlemsstater (Danmark, Nederländerna, Sverige och Storbritannien) har tagit initiativ till att anta en nationell förklaring om förvaltningen av gemenskapsmedel, men beklagar att majoriteten av de övriga medlemsstaterna trots detta initiativ motsätter sig införandet av en sådan förklaring och beklagar djupt att Belgien, Bulgarien, Tjeckien, Tyskland, Estland, Irland, Grekland, Spanien, Frankrike, Italien, Cypern, Lettland, Litauen, Luxemburg, Ungern, Malta, Österrike, Polen, Portugal, Rumänien, Slovenien, Slovakien och Finland ännu inte vidtar några åtgärder för att utveckla ett effektivt system för nationella förklaringar.
34.
Kontrollsystem
Handlingsplanen för en integrerad ram för intern kontroll
35.
Europaparlamentet noterar med tillfredsställelse de framsteg som har gjorts i genomförandet av handlingsplanen, att majoriteten av åtgärderna har vidtagits och att de flesta brister som tas upp i handlingsplanen har åtgärdats.
36.
Europaparlamentet uttrycker sin oro över revisionsrättens upprepade kritik av den bristande kvaliteten på kontrollerna i medlemsstaterna och noterar bekymrat klagomålen från mottagare och nationella kontrollinstanser om antalet kontroller och om avgifterna.
37.
Europaparlamentet noterar även med oro mottagarnas kritik av antalet manualer, handböcker, arbetsdokument och deltaganderegler som ska tillämpas på stöd och begär att dessa dokument konsolideras och att en diskussion bör föras med parlamentet för att förenkla dessa tillämpningsföreskrifter.
38.
39.
40.
Europaparlamentet beklagar att genomförandet av åtgärd 4 i handlingsplanen för en integrerad ram för intern kontroll, som gäller införandet av ett interinstitutionellt initiativ om de grundprinciper som ska beaktas i fråga om acceptabla risker i underliggande transaktioner, kommer att försenas.
41.
Europaparlamentet påminner också om vikten i detta sammanhang av att genomföra åtgärd 10 i handlingsplanen som syftar till att göra en "analys av kostnaderna för kontrollerna", med tanke på behovet "att uppnå en lämplig balans mellan kostnaderna för och nyttan med kontroller".
42.
Europaparlamentet förväntar sig också att generaldirektoratens årliga verksamhetsrapporter återigen kommer att innehålla uppgifter om kvaliteten på kontrollerna i medlemsstaterna och om deras förbättringar och kräver att kommissionen ska klassificera samtliga utbetalande och attesterande organ.
43.
Europaparlamentet uppmanar kommissionen att regelbundet lägga fram utvärderingar av det integrerade interna kontrollsystemet och kräver att de årliga verksamhetsrapporterna och den sammanfattande rapporten på ett ännu bättre sätt omfattar kommissionens tjänsteavdelningars och medlemsstaternas system för den delade förvaltningen, särskilt när det gäller den tekniska kvaliteten och de etiska övervägandena, t.ex. i fråga om de nationella revisionsmyndigheternas oberoende.
44.
Europaparlamentet uppmanar kommissionen att göra en mer fullständig och uttömmande utvärdering av kostnaderna för de resurser som läggs på kontrollsystem per utgiftsområde och att göra detta för samtliga av EU:s utgiftsområden, precis som parlamentet har begärt i sina resolutioner om beviljande av ansvarsfrihet under föregående år, och med tanke på begreppet "att uppnå resultat".
45.
46.
Europaparlamentet anser att denna jämförande analys bör överlämnas till parlamentet, rådet och revisionsrätten i slutet av 2009 eller i början av 2010 och att den bör ligga till grund för en interinstitutionell dialog om den godtagbara felfrekvensen.
47.
Europaparlamentet konstaterar att även om begreppet tolererbar risknivå (acceptabel risk för fel) är grundläggande för den integrerade ramen för intern kontroll som revisionsrätten måste beakta när den utfärdar sin revisionsförklaring i enlighet med revisionsrättens yttrande nr 4/2006 över förslaget till rådets förordning om ändring av förordning (EG, Euratom) nr 1605/2002 EUT C 273, 9.11.2006, s.
2.
, har det ännu inte definierats hur denna tolererbara risknivå ska fastställas.
Acceptabel risk för fel
48.
49.
Europaparlamentet beklagar att kommissionen i sitt meddelande förklarar att den har svårigheter med att få in tillräckligt tillförlitliga uppgifter från medlemsstaterna och anser att denna bedömning skadar EU:s framtoning.
50.
Europaparlamentet tvivlar på tillförlitligheten i uppgifterna som medlemsstaterna lämnar och uppmanar kommissionen att samla in sifferuppgifter på nytt, med tekniskt stöd från revisionsrätten, och att göra en fördjupad analys så snart som effekterna av bestämmelserna för perioden 2007–2013 blir synliga och att översända denna analys till parlamentet och rådet före utgången av 2011.
51.
Europaparlamentet anser att det är ytterst viktigt och samtidigt mycket komplicerat att fastställa en tolererbar risknivå och att denna nivå bör hänga nära samman med en fördjupad undersökning av kostnadseffektiviteten i kommissionens och medlemsstaternas kontrollsystem för vart och ett av gemenskapens utgiftsområden.
52.
Med tanke på hur viktigt det är att fortsätta att analysera kostnader och fördelar av kontroller uppmanar Europaparlamentet kommissionen att med tekniskt stöd från revisionsrätten göra en fördjupad analys av områdena för forskning, yttre förbindelser och administrativa utgifter och att leverera en rapport om detta före utgången av 2010.
53.
Europaparlamentet anser att beloppet för de EU-medel som går förlorade på grund av felaktigheter också bör beaktas när en godtagbar felfrekvens fastställs.
54.
Europaparlamentet anser att det behövs konkreta förslag om hur förvaltningen och kontrollen av gemenskapsmedlen kan förbättras och rentav harmoniseras i vissa fall och föreslår att parlamentet vid nästa budgetförfarande ger kommissionen de resurser som krävs för att genomföra en undersökning.
55.
Europaparlamentet uppmanar kommissionen att utan dröjsmål överlämna sina förslag till hur målet om en positiv revisionsförklaring ska kunna uppnås.
Öppenhet
56.
57.
Europaparlamentet beklagar att dess begäran om en ny uppförandekod för ledamöter av kommissionen, vilken skulle förbättra och tydligare definiera deras individuella och kollektiva politiska ansvar och redovisningsskyldighet för sina beslut och för tjänsteavdelningarnas genomförande av politiken, inte hörsammats.
58.
Europaparlamentet påminner återigen om kommissionens ansvar för att säkerställa att uppgifter om mottagare av EU-finansiering är fullständiga, sökbara och jämförbara, och beklagar att detta mål ännu inte har uppnåtts.
59.
Europaparlamentet påminner återigen om vikten av fullständig öppenhet och offentlighet när det gäller personal vid kommissionsledamöternas kabinett som inte har rekryterats enligt personalföreskrifterna.
60.
61.
EUT L 340, 6.12.2006, s.
5.
.
62.
Europaparlamentet påminner kommissionen om att en fullständig och lättåtkomlig databas med uppgifter om alla slutmottagare av gemenskapsfinansiering bör vara tillgänglig och öppen för en bredare publik före nästa val till Europaparlamentet.
Budgetförordning
63.
Europaparlamentet noterar med tillfredsställelse att den förenkling som gjordes vid den senaste revideringen av förordning (EG, Euratom) nr 1605/2002 har gett de önskade effekterna för offentliga upphandlingar.
64.
65.
Europaparlamentet uppmanar kommissionen att på ett mycket tidigt stadium konsultera andra institutioner som omfattas av förordning (EG, Euratom) nr 1605/2002.
Europeiska byrån för bedrägeribekämpning (Olaf)
66.
Europaparlamentet noterar med oro arbetsvillkoren för Olaf och uppmanar kommissionen att se till att Olaf får direkt tillgång till kommissionens databaser när det uppstår behov i samband med en undersökning för att det ska vara möjligt att inleda och administrera undersökningar utan dröjsmål.
67.
68.
69.
70.
SEKTORSSPECIFIKA FRÅGOR
Egna medel
71.
72.
Europaparlamentet påminner om punkt 93 i sin ovannämnda resolution av den 24 april 2007 om ansvarsfrihet för 2005 där parlamentet förutsätter att FISIM automatiskt kommer att inkluderas i beslutet om egna medel, för beräkning av egna medel från BNI, eftersom kommissionen i sitt förslag till rådets beslut om systemet för Europeiska gemenskapernas egna medel ( KOM(2006)0099 ) inte gjorde någon reservation om begränsningar i detta hänseende.
73.
Europaparlamentet konstaterar att inte heller rådet gjorde någon minsta reservation om begränsningar för FISIM, i enlighet med kommissionens förslag (KOM (2006) 0099), i samband med antagandet av beslut 2007/436/EG, Euratom av den 7 juni 2007 om systemet för Europeiska gemenskapernas egna medel EUT L 163, 23.6.2007, s.
Parlamentet förväntar sig därför att beräkningen av Europeiska gemenskapernas egna medel, i och med att det nya beslutet träder i kraft, retroaktivt från och med den 1 januari 2007 ska göras på grundval av BNI-uppgifter som beaktar FISIM, och att det på denna grundval görs nya beräkningar av hittillsvarande och framtida betalningar från medlemsstaterna.
Jordbruk och naturresurser
74.
75.
76.
Europaparlamentet konstaterar emellertid att revisionsrätten drar slutsatsen att det integrerade systemet för förvaltning och kontroll fortfarande är ändamålsenligt för att begränsa risken för oriktiga utgifter förutsatt att systemet genomförs på rätt sätt och att riktiga och tillförlitliga uppgifter registreras för de betalningar inom systemet med samlat gårdsstöd som baseras på tilldelade stödrättigheter (punkt 5.20 och 5.21 i årsrapporten 2007).
77.
Europaparlamentet är dock oroat över revisionsrättens kritik i fråga om feltolkningar av bestämmelser i lagstiftningen och över slutsatsen att alla de fel som uppstår under flera års tid kommer att leda till en betydande ackumulerad effekt om de inte korrigeras och uppmanar kommissionen att så snart som möjligt vidta lämpliga åtgärder, som åtminstone bör innebära en förenkling av politikområdet och ett klarare och konsekventare kontrollsystem, för att korrigera dessa fel och att informera parlamentet om de vidtagna åtgärderna i slutet av 2009.
78.
79.
Europaparlamentet noterar med oro de stora svagheter som revisionsrätten avslöjar i kontrollsystemen i flera medlemsstater när det gäller landsbygdsutvecklingen till följd av att vissa villkor för stödberättigande inte är tillräckligt tydligt definierade i den nationella lagstiftningen och att reglerna ofta är komplicerade, vilket påverkar kvaliteten i kontrollerna negativt.
80.
81.
Europaparlamentet uppmanar medlemsstaterna att i samarbete med kommissionen omedelbart intensifiera sina kontroller, särskilt av att stödmottagarna uppfyller villkoren för att få stöd, och uppmanar kommissionen att så snart som möjligt förtydliga och förenkla dessa villkor.
82.
Europaparlamentet beklagar att revisionsrätten även för år 2007 har konstaterat samma inneboende begränsningar i systemet för granskning och godkännande, t.ex. att besluten om överensstämmelse grundar sig på retroaktivitet och flerårighet och det faktum att det inte finns någon giltig koppling mellan de belopp som återbetalats på detta sätt och de faktiska belopp som betalats ut på felaktiga grunder (punkt 5.47 i årsrapporten 2007).
83.
Europaparlamentet anser att efter flera år med samma allvarliga kritik från revisionsrätten om samma problem måste kommissionen lägga fram förslag för att reformera systemet så att det blir möjligt att göra tydliga och giltiga kopplingar mellan återbetalade belopp och de belopp som betalats ut på felaktiga grunder och att i så hög grad som möjligt säkerställa att kostnaderna för de finansiella korrigeringarna bärs av de slutliga stödmottagarna och inte av skattebetalarna, och att schablonkorrigeringar ska tillämpas på medlemsstater som inte respekterar sina förpliktelser.
Fiskestöd
84.
Europaparlamentet välkomnar att utvalda medlemsstater har offentliggjort namnen på stödmottagarna, namnen på de aktuella projekten och storleken på den offentliga finansieringen (på gemenskapsnivå och nationell nivå) på kommissionens webbplats som också innehåller länkar till medlemsstaternas informationskällor.
85.
1).
.
86.
Europaparlamentet välkomnar kommissionens förslag till rådets förordning om införande av ett kontrollsystem i gemenskapen för att säkerställa att bestämmelserna i den gemensamma fiskeripolitiken efterlevs ( KOM(2008)0721 ), vilket syftar till att göra det rättsligt möjligt att skjuta upp eller minska ekonomiskt stöd till medlemsstater som inte tillämpar bestämmelserna i den gemensamma fiskeripolitiken på ett korrekt sätt.
87.
Europaparlamentet begär dock att kommissionen också föreslår att medlemsstater som inte tillämpar bestämmelserna i den gemensamma fiskeripolitiken på ett korrekt sätt inte heller ska kunna dra fördel av partnerskapsavtal om fiske.
88.
Europaparlamentet begär att kommissionen inför gemenskapslagstiftning som utesluter alla fartygsägare som begått allvarliga överträdelser (enligt rådets förordning (EG) nr 1447/1999 Rådets förordning (EG) nr 1447/1999 av den 24 juni 1999 om att upprätta en förteckning över sådana beteenden som utgör allvarliga överträdelser av den gemensamma fiskeripolitikens bestämmelser (EGT L 167, 2.7.1999, s.
5).
från gemenskapsstöd från Europeiska fiskerifonden och/eller från utnyttjande av partnerskapsavtal om fiske.
89.
Europaparlamentet uppmanar kommissionen att se till att gemenskapsstödet inte används till modernisering av sådana flottsegment som har överkapacitet.
90.
Europaparlamentet påminner kommissionen om dess åtaganden inom ramen för strategin för hållbar utveckling, vilken godkändes av Europeiska rådet vid mötet i Göteborg i juni 2001 och reviderades av Europeiska rådet vid mötet i Wien i juni 2006, att avveckla miljöskadligt stöd och att senast 2008 presentera en färdplan med sektorsvisa reformer av dessa stöd med syftet att eliminera dem.
Sammanhållning
91.
Europaparlamentet noterar med stor oro revisionsrättens beräkning att minst 11 procent av det totala belopp som ersatts inte borde ha ersatts när det gäller strukturpolitiska projekt.
92.
Europaparlamentet konstaterar att kommissionen inte ifrågasätter denna andel på 11 procent.
93.
Europaparlamentet konstaterar att det antal kontroller som revisionsrätten genomfört förefaller lågt i förhållande till antalet betalningar till slutmottagarna (till exempel för sammanhållningspolitiken har revisionsrätten enligt punkt 6.21 i årsrapporten 2007 kontrollerat 180 delbetalningar av flera hundratusentals betalningar till slutmottagare), men konstaterar att denna revisionsmetod överensstämmer med internationella revisionsstandarder enligt de synpunkter som lagts fram i rapporten International Peer Review of the European Court of Auditors som gjorts av en grupp erfarna finans- och effektivitetsrevisorer från de högsta nationella revisionsorganen i Österrike, Kanada, Norge och Portugal.
94.
Visserligen uppskattar Europaparlamentet förbättringarna i den samlade bedömningen av systemen för övervakning och kontroll i revisionsrättens årsrapport, men beklagar ändå att systemen för förvaltning och kontroll på såväl medlemsstatsnivå som kommissionens övervakningsnivå inte är tillräckligt effektiva för att begränsa felfrekvensen, trots kommissionens fortsatta ansträngningar, och uppmanar kommissionen att rapportera till parlamentet i början av 2010 om de ytterligare åtgärder som har genomförts under 2009 samt om de inledande effekterna av åtgärderna i den ovan nämnda handlingsplanen.
95.
Europaparlamentet noterar med stor oro att utnyttjandet av regionalfonden och Sammanhållningsfonden uppnådde oacceptabelt låga nivåer, och uppmanar kommissionen att fortsätta revisionsförfarandet och att genast förenkla gällande förordningar.
96.
97.
Europaparlamentet uppmanar även kommissionen att göra en bedömning av sammanhållningspolitikens positiva effekter per medlemsstat och lägga fram en rapport till parlamentet om det mervärde som politiken medför på EU-nivå.
98.
99.
100.
101.
102.
103.
Europaparlamentet uppmanar kommissionen, som har det slutliga ansvaret för en god finansiell förvaltning av gemenskapens medel, att strikt tillämpa gemenskapsbestämmelserna om uppskjutande av betalningar när en medlemsstat inte lämnar de begärda garantierna.
104.
105.
106.
107.
108.
109.
110.
Europaparlamentet betonar att den felnivå som redovisas i rapporten från revisionsrätten inte nödvändigtvis hänför sig till bedrägerier och uppmanar därför kommissionen och revisionsrätten att härvidlag göra en klar åtskillnad i framtida dokument.
111.
Inre politik
112.
Europaparlamentet beklagar att revisionsrätten anser att samma problem kvarstår som under föregående år avseende de områden som kommissionen förvaltar direkt (brister i ersättningen av kostnader, komplexa bestämmelser och avsaknad av en effektiv sanktionsmekanism) och uppmanar kommissionen att fortsätta sina insatser för att förenkla och ytterligare förtydliga de regler som gäller för program med delade kostnader.
Forskning
113.
Europaparlamentet välkomnar utvecklingen på området för forskning och teknisk utveckling där den årliga felfrekvensen minskat från 8,03 procent 2006 till 2,39 procent 2007, vilket utgör en stor bedrift som visar att kommissionens forskningsansvariga enheter, i nära samarbete med budgetkontrollutskottet och revisionsrätten, varit framgångsrika i att genomföra rekommendationerna från 2005 års ansvarsfrihetsförfarande.
114.
Europaparlamentet konstaterar att systemet med revisionsintyg under 2007 fick ned felfrekvensen till 2,5 procent för projekt inom det sjätte ramprogrammet, i jämförelse med 4,06 procent för projekt inom det femte ramprogrammet som inte ingår i systemet med revisionsintyg.
115.
Europaparlamentet välkomnar det arbetsdokument från kommissionens tjänsteavdelningar ( SEK(2008)3054 ) som innehåller en första analys av bland annat kontrollkostnaderna för generaldirektoratet för forskning och generaldirektoratet för informationssamhället och medier för att väcka nytt liv i den interinstitutionella diskussionen i syfte att åstadkomma ett gemensamt avtal om den godtagbara felfrekvensen på området för EU:s forskningspolitik.
116.
Europaparlamentet uppmanar kommissionen att fortsätta att uppfylla de ersättningsmöjligheter som fastställs i det sjunde ramprogrammet, särskilt genom att ytterligare analysera huruvida det sjunde ramprogrammets bestämmelser om förfarande för schablonersättningar är lämpliga, och att informera parlamentets behöriga utskott i samband med halvtidsöversynen om hur man har bidragit till att förenkla bestämmelserna för betalningsmottagarna samt om nödvändiga förbättringar av systemet.
117.
118.
119.
Med syftet att förenkla de administrativa rutinerna och bidragsansökningarna vill Europaparlamentet påminna om sin begäran om en enda kontaktpunkt för stödmottagarna för frågor i samband med ramprogrammet, och som har behörighet att fatta beslut i dessa ärenden.
120.
Europaparlamentet begär att kommissionen, som en förutsättning för rättssäkerheten, avstår från att räkna om årsredovisningarna för projekt inom det sjätte ramprogrammet som redan har godkänts och avslutats av kommissionen, genom att tillämpa nya tolkningar av vilka kostnader som är stödberättigade enligt de allmänna villkoren (bilaga II) i det sjätte ramprogrammets standardkontrakt.
121.
122.
123.
Eftersom kommissionens revisionsstrategi omfattar kostnaderna för ett ramprogram under en fyraårsperiod, medan revisionsrätten ska utarbeta rapporter på årsbasis, uppmanar Europaparlamentet revisionsrätten att lägga fram fleråriga tabeller där de finansiella effekterna av de felaktigheter som konstaterats under revisionsrättens revisionsarbete presenteras på ett sätt som stämmer överens med kommissionens kontrollmetod.
Miljö, folkhälsa och livsmedelssäkerhet
124.
Europaparlamentet anser att de övergripande genomförandenivåerna för budgetens utgiftskategorier miljö, folkhälsa och livsmedelssäkerhet är tillfredsställande.
125.
Europaparlamentet betonar att den övergripande budgetgenomförandenivån på 94,6 procent för miljö, folkhälsa och livsmedelssäkerhet är ett tillfredsställande resultat med tanke på att 2007 var det första året i den nya budgetramen 2007–2013 och ett år som kännetecknades av antagandet och ikraftträdandet av nya program på politikområdet miljö.
126.
127.
Europaparlamentet uppmanar kommissionen att utveckla ytterligare stöd till sökande inom fleråriga program, särskilt genom att erbjuda sökande särskild utbildning och utarbeta användarvänliga riktlinjer.
128.
Europaparlamentet välkomnar ansträngningarna att göra anbudsinfordringar mer fokuserade och att ge mer stöd till sökande, särskilt inom folkhälsoprogrammen, så att man kan undvika att projektansökningar lämnas in som uppenbarligen inte kan komma ifråga för stöd eller som är av dålig kvalitet, men noterar att ytterligare insatser behövs för att situationen ska bli tillfredsställande.
129.
130.
Europaparlamentet betonar att administrativa och finansiella bestämmelser i förordning (EG, Euratom) nr 1605/2002 inte får leda till onödiga förseningar för beviljandet av bidrag eller urvalet av projekt som ska finansieras och uppmanar kommissionen att fortsätta sina ansträngningar att förbättra administrativa förfaranden som påverkar genomförandet av åtagande- och betalningsbemyndiganden.
Inre marknaden och konsumentskydd
131.
Europaparlamentet välkomnar iakttagelserna i revisionsrättens rapport, som ger en rättvis bedömning av politiken för den inre marknaden, tullpolitiken och konsumentskyddspolitiken.
132.
133.
134.
135.
136.
Transport och turism
137.
- 933 578 000 EUR som åtagandebemyndiganden och 369 665 000 EUR som betalningsbemyndiganden för transeuropeiska transportnät (TEN-T).
- 15 348 000 EUR som åtaganden och 14 500 000 EUR som betalningar för transportsäkerhet.
- 56 890 000 EUR som åtaganden och 10 425 000 EUR som betalningar för Marco Polo-programmet.
- 113 631 000 EUR som åtaganden och 114 716 000 EUR i betalningar för transportbyråerna och övervakningsmyndigheten för GNSS.
- 6 000 000 EUR i åtaganden och 6 578 000 EUR i betalningar för transportsäkerhet, inbegripet pilotprojekt för säkerhet inom det transeuropeiska vägnätet.
138.
Europaparlamentet välkomnar att både åtagandebemyndiganden och betalningsbemyndiganden för TEN-T-projekt fortsättningsvis utnyttjas i hög grad, nästan till 100 procent vardera, och uppmanar medlemsstaterna att se till att adekvat finansiering görs tillgänglig ur de nationella budgetarna för att matcha detta gemenskapsåtagande.
139.
140.
Europaparlamentet noterar med tillfredsställelse att till följd av reaktionerna på revisionsrättens särskilda rapport nr 6/2005 om det transeuropeiska transportnätet EUT C 94, 21.4.2006, s.
1.
141.
Europaparlamentet noterar med tillfredsställelse att revisionsrättens analys av interna kontrollstandarder med en direkt koppling till de underliggande transaktionernas laglighet och korrekthet visar att generaldirektoratet för energi och transport uppfyller de grundläggande kraven.
Kultur och utbildning
142.
Europaparlamentet konstaterar att revisionsrätten i sin årsrapport 2007 uttalar sig om den felfrekvens som den har upptäckt på politikområdet för utbildning och kultur (punkt 9.11 och bilaga 9.1, en felprocent på mellan 2 procent och 5 procent), men inte ger någon förklaring angående arbetssättet hos de olika nationella organen och genomförandeorganen och inte heller angående kvaliteten i deras arbete eller varför denna organisation ska räknas med.
143.
Europaparlamentet uppmanar revisionsrätten att i sin nästa årsrapport göra en mer ingående analys av frågan om effektivitet och förekomsten av olika organ på området för utbildnings- och kulturpolitik.
144.
145.
146.
Parlamentet uppmanar kommissionen att harmonisera förklaringarna och att hålla parlamentet och revisionsrätten informerade om hur harmoniseringsarbetet fortskrider.
147.
148.
Europaparlamentet beklagar att vissa nationella myndigheter och organ inte uppfyller sina skyldigheter, vilket har lett till att kommissionen har skickat officiella påminnelseskrivelser, och ger kommissionen sitt fulla stöd när det gäller att skjuta upp utbetalningarna av bidrag i de fall slutrapporter saknas.
149.
150.
Europaparlamentet ser med tillfredsställelse på att antalet sena betalningar på utbildnings- och kulturområdet minskat och förväntar sig att kommissionen fortsätter sina ansträngningar att minska dem ytterligare.
151.
Europaparlamentet hoppas att det kontrollsystem som generaldirektoratet för kommunikation upprättade i slutet av 2007 kommer att göra det onödigt att lämna en reservation om dess budgetförvaltning i framtiden, vilket var fallet för budgetåret 2007.
152.
Europaparlamentet begär mer information från kommissionen om inrättandet av administrativa strukturer i medlemsstaterna för att medverka i vänortsverksamhet, särskilt behovet av sådana strukturer, kostnaderna i samband härmed och deras syfte.
153.
Medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor
154.
155.
156.
Europaparlamentet beklagar att beskrivningarna av medlemsstaternas system för övervakning och kontroll av fonden för de yttre gränserna lämnades till kommissionen först under det sista kvartalet 2007, vilket fick till följd att kommissionen inte kunde bedöma medlemsstaternas system före utgången av 2007.
Kvinnors rättigheter och jämställdhet mellan kvinnor och män
157.
158.
Europaparlamentet upprepar sin begäran till kommissionen om att jämställdhet ska betraktas som ett ständigt prioriterat mål under budgetplaneringen, i enlighet med principen om integrering av ett jämställdhetsperspektiv i budgeten, vilket parlamentet begärde i sin resolution av den 3 juli 2003 om gender budgeting — att utarbeta offentliga budgetar utifrån ett genusperspektiv EUT C 74 E, 24.3.2004, s.
746.
, och beklagar att kommissionens genomförbarhetsstudie om ärendet i fråga har försenats.
159.
Europaparlamentet beklagar att revisionsrättens årsrapport om genomförandet av budgeten för 2007 inte innehåller upplysningar om huruvida budgeten framgångsrikt bidragit till att främja jämställdhet.
160.
Europaparlamentet föreslår att revisionsrätten inkluderar jämställdhetsaspekter i sina årsrapporter och särskilda rapporter, särskilt relevant information om åtgärder för integrering av principen om icke-diskriminering mellan män och kvinnor och om tillgången till könsspecifika uppgifter.
Externa åtgärder
161.
Europaparlamentet noterar med stor oro att revisionsrätten framför samma kritik som föregående år, framför allt i fråga om utbetalningar på slutlig stödmottagarnivå.
162.
Europaparlamentet påpekar att bistånd till tredjeland i princip inte berördes av den senaste revideringen av förordning (EG, Euratom) nr 1605/2002 och kräver en översyn av avdelning IV "Externa åtgärder" i förordning (EG, Euratom) nr 1605/2002 för att anpassa den bättre till de särskilda marknads- och stödvillkoren på detta område.
163.
multi donor trust fond
) när den deltar i dessa fonder.
164.
165.
166.
Europaparlamentet konstaterar att denna uppskattning enligt den information som lämnats av kommissionen endast omfattar en del av de sammanlagda kostnaderna för de humanitära insatser som finansieras av ECHO eftersom kostnaderna för de kontroller som genomförs av de humanitära organisationerna och som ingår i totalkostnaderna för bidragsavtalen också finansieras av ECHO.
167.
Europaparlamentet konstaterar att utifrån hypotesen att kontrollkostnaderna utgörs av tre stora kategorier – kostnaderna för de kontroller som kommissionens tjänsteavdelningar utför vid huvudkontoret och vid delegationerna, kostnaderna för externa revisioner av kommissionen och kostnaderna för verifiering av utgifterna genom revisioner som beställs av mottagarna – uppskattar kommissionen att kontrollkostnaderna för fonder som förvaltas av byrån för samarbete, EuropeAid, under 2007 uppgick till omkring 120 000 000 EUR.
168.
Europaparlamentet uppmanar revisionsrätten att i sin nästa årsrapport ta hänsyn till detta i sina beräkningar och uttala sig om denna uppskattning och om kostnadseffektiviteten i dessa kontrollsystem med hänsyn till de särskilda egenskaperna och begränsningarna hos EU:s yttre åtgärder.
169.
Europaparlamentet beklagar att kommissionen betalade ut ett budgetstöd till Kenya precis efter valet den 27 december 2007, vilket gav intrycket av att den valde sida i diskussionen om valets legitimitet.
och förväntar sig att kommissionen tar hänsyn till den.
170.
171.
172.
Europaparlamentet uppmanar kommissionen att ytterligare förbättra, och mer noggrant definiera, de villkor och resultatindikatorer som används för att betala ut budgetstöd till tredjeländer, så att man tillhandahåller klara, otvetydiga och mätbara bedömningskriterier, i förekommande fall med en specifik tidtabell.
173.
174.
Europaparlamentet ser fram emot konkreta resultat av tillämpningen av nya direktiv för utgiftskontroller via externa revisioner som genomförs på initiativ av stödmottagarna eller kommissionen.
175.
Europaparlamentet tar del av revisionsrättens särskilda rapport nr 5/2007 om kommissionens förvaltning av Cardsprogrammet EUT C 285, 27.11.2007, s.
176.
Europaparlamentet förväntar sig att regelbundet informeras om de åtgärder som kommissionen vidtar för att genomföra den viktiga utfästelsen om stöd till Georgiens återhämtning efter konflikten och framtida utveckling vid den internationella givarkonferens som hölls i Bryssel den 22 oktober 2008.
177.
Europaparlamentet uppmanar återigen kommissionen att regelbundet lägga fram konkreta åtgärder för parlamentet för att ytterligare öka EU:s ansvar för och kontroll över sina externa åtgärder i deras geografiska sammanhang, i enlighet med principerna om effektivitet, ansvar och synlighet.
Icke-statliga organisationer
178.
Europaparlamentet noterar de icke-statliga organisationernas roll och växande antal i förvaltningen av gemenskapsmedlen, och uppmanar kommissionen att utvärdera hur effektivt driftsstödet till de icke-statliga organisationernas huvudkontor i Bryssel är och att strikt tillämpa den princip om gradvis nedtrappning av driftsstödet som fastslås i budgetförordningen.
179.
Europaparlamentet uppmanar kommissionen att senast i slutet av 2009 sammanställa en fullständig förteckning över alla frivilligorganisationer som har mottagit gemenskapsmedel.
Utveckling
180.
Europaparlamentet noterar att revisionsrätten än en gång har konstaterat att ECHO bör förbättra sin revisionsstrategi genom att garantera en bättre täckning av transaktioner vid verkställande organ och mer specifikt på fältnivå när det gäller alla typer av partner (punkt 8.33 f i årsrapporten 2007).
181.
Europaparlamentet uppmuntrar kommissionen i dess målsättning sedan 2007 att varje projekt ska besökas minst en gång av en expert, såvida det inte på grund av säkerhetsförhållanden eller svårtillgänglighet är omöjligt, så att humanitära biståndsspecialister permanent befinner sig på plats för att underlätta och maximera effekterna av de humanitära insatser som finansieras av kommissionen, oavsett vilket land eller region det rör sig om.
182.
Europaparlamentet anser att kommissionen när projekten genomförs måste se till att de bestämmelser som antogs tillsammans med FN i april 2007 om rapportering tillämpas strikt och att de finansiella rapporterna utformas i enlighet med dessa bestämmelser.
183.
Europaparlamentet är medvetet om riskerna med otillräckliga kontroller på plats i områden som är svårtillgängliga eller där det humanitära biståndets neutralitet inte respekteras och att dessa risker i viss mån är förknippade med biståndsmålen för humanitära behov och det som brukar kallas "bortglömda kriser".
184.
Europaparlamentet noterar också att enligt den årliga verksamhetsrapporten från ECHO 2007 har kommissionens humanitära bistånd i Irak uteslutande genomförts via Röda korsets internationella kommitté inom sektorerna för vattenskydd och rening till ett sammanlagt belopp av 7 800 000 EUR.
185.
186.
187.
Europaparlamentet betonar att inom utbildningen måste prioritet ges till inskrivning av barn från grupper som är svåra att nå i länder med kritiska millennieutvecklingsmålsindikatorer, särskilt barn med funktionshinder.
188.
Europaparlamentet uppmanar med kraft kommissionen att prioritera stöd till partnerländer för att utveckla parlamentarisk kontroll- och revisionskapacitet, särskilt när biståndet tillhandahålls via budgetstöd och kommissionen uppmanas också att regelbundet rapportera om de framsteg som gjorts.
189.
190.
191.
41).
Föranslutningsstrategin
Samarbets- och kontrollmekanismen
192.
Europaparlamentet påminner om att kommissionen för första gången efter en anslutning av nya medlemsstater har inrättat en samarbets- och kontrollmekanism för Rumänien och Bulgarien för att åtgärda "brister när det gäller reformen av rättsväsendet och kampen mot korruption och organiserad brottslighet och att övervaka framstegen på dessa områden" ( KOM(2008)0063 ) och undrar hur effektiv och relevant denna mekanism är samt hur tillförlitliga uppgifterna till den myndighet som beviljar ansvarsfrihet är.
193.
EU-medel i Bulgarien och Rumänien
194.
Europaparlamentet konstaterar att 650 000 000 EUR har ställts till Bulgariens förfogande mellan 2004 och 2007 inom ramen för gemenskapsprogrammet för ekonomiskt stöd till länder i Central- och Östeuropa (Phareprogrammet), 226 000 000 EUR inom ramen för det särskilda föranslutningsprogrammet för jordbruket och landsbygdens utveckling (Sapard), 440 500 000 EUR inom ramen för det strukturpolitiska föranslutningsinstrumentet (Ispa) och att omkring 1 346 500 000 EUR har ställts till Rumäniens förfogande mellan 2004 och 2007 inom ramen för Phareprogrammet, 526 300 000 EUR inom Sapard och 1 040 500 000 EUR inom Ispa.
195.
Europaparlamentet påminner om att revisionsrätten redan i sin särskilda rapport 4/2006 om investeringsprojekt inom Phareprogrammet i Bulgarien och Rumänien EUT C 174, 26.7.2006, s.
1.
konstaterade ett flertal problem i förvaltningen av EU-medlen, bl.a. i form av oriktigheter i anbudsförfarandena och utgifternas stödberättigande, avyttring av kapitalvaror och bristande administrativ kapacitet.
196.
Europaparlamentet noterar också med oro att budgetkontrollutskottet inte fick tillfredsställande information om bristernas omfattning inom de fastställda tidsfristerna av den kommissionsledamot som har ansvar för utvidgningen.
197.
198.
Europaparlamentet är medvetet om att bristen på tillförlitliga kontrollsystem och förvaltningsproblemen innebär risker för de europeiska bidragsgivarnas pengar, välkomnar de insatser som har gjorts under tiden för att lösa problemen och uppmanar medlemsstaterna att fortsätta vidta alla åtgärder som krävs för att uppfylla sina skyldigheter inför EU.
199.
200.
201.
Europaparlamentet anser att kommissionen inte på ett tillräckligt seriöst sätt har hanterat frågan om Rumäniens och Bulgariens kapacitet att tillgodogöra sig medlen på jordbruks- och sammanhållningsområdena, och att kommissionens uttalanden och åtgärder i detta sammanhang var missledande, inte enbart för parlamentet utan även för Bulgariens och Rumäniens regeringar, och att de var ett av skälen till att dessa länder förlorade medel.
202.
Europaparlamentet uppmanar kommissionen att hålla parlamentet underrättat om de praktiska konsekvenserna av arbetet med de rättsliga reformerna och kampen mot korruptionen och begär att det i framstegsrapporterna införs kriterier för att mäta framstegen på dessa områden.
203.
Europaparlamentet anser att EU:s institutioner bör tillämpa nolltolerans när det gäller missbruk av EU-medel, bedrägerier och korruption och uppmanar kommissionen att se till att belopp som har betalats ut oriktigt verkligen återvinns.
204.
Europaparlamentet uppmanar även Olaf att överlämna resultatet av sina pågående undersökningar i medlemsstaterna till parlamentet.
205.
206.
Mot bakgrund av den senaste lägesrapporten och bakslagen vad gäller korruptionsbekämpningen begär Europaparlamentet att från gemenskapsmedel i Rumänien och om vilka åtgärder som vidtagits vad gäller korruptionsbekämpningen och vilka resultat detta har gett, under perioden fram till den 15 juli 2009.
Turkiet, Kroatien, Serbien, f.d. jugoslaviska republiken Makedonien, Kosovo och övriga länder på västra Balkan
207.
208.
209.
210.
Europaparlamentet uppmanar revisionsrätten att utarbeta en särskild rapport om effektiviteten i de kontrollsystem som kommissionen har infört för de medel som Kosovo har fått från EU samt deras verkan när det gäller att förebygga bedrägerier och att kontrollera att finansieringen fullt ut har omfattats av de villkor som fastställts i avtalen för de berörda programmen, inbegripet bestämmelserna i föranslutningsinstrumentet Rådets förordning (EG) nr 1085/2006 av den 17 juli 2006 om upprättande av ett instrument för stöd inför anslutningen (EUT L 210, 31.7.2006, s.
82).
och i förordning (EG, Euratom) nr 1605/2002.
211.
Europaparlamentet föreslår att kommissionen kräver att Kosovos regering visar upp ett revisionsintyg från landets revisionsrätt i fråga om EU:s medel och särskilt dem som har använts i budgeten.
212.
Administrativa utgifter
213.
Europaparlamentet konstaterar med tillfredsställelse att revisionsrättens granskning inte har avslöjat några väsentliga fel som påverkar lagligheten och korrektheten i de administrativa utgifterna.
Europaskolor
214.
Europaparlamentet förväntar sig att kommissionen ser till att Belgiens och Storbritanniens regeringar åtar sig att fullgöra sina skyldigheter enligt gällande avtal mellan regeringarna – för Belgiens del att snarast färdigställa en fjärde eller rent av en femte europaskola, för Storbritanniens del att avdela tillräckligt många lärare – samt att den gällande antagningspolicyn för skolorna i Berkendael/Laeken ses över, så att långa och oacceptabla restider för barnen kan undvikas.
Decentraliseringens effekter för personalen
215.
Europaparlamentet noterar med tillfredsställelse att kommissionen på parlamentets begäran har genomfört en undersökning av personalresurserna 2007 ( SEK(2007)0530 ) i fråga om den administrativa verksamheten.
216.
217.
218.
Frågor i samband med gemenskapens fastighetsinfrastruktur
219.
Europaparlamentet beklagar kommissionens bristande öppenhet i fråga om förvaltningen av de 61 byggnader som den disponerar i Bryssel och om utvecklingen av dess fastighetsbestånd.
220.
Europaparlamentet uppmanar kommissionen att underrätta det om alla nya projekt avseende fastighetsbeståndet innan sådana beslut fattas, samt att regelbundet informera parlamentets budgetkontrollutskott om alla initiativ och nya beslut om fastighetsprojekt, inklusive förberedande arbeten och anbudsförfaranden för vilka det föreslås att inrätta en kommitté för anbudsförfaranden med företrädare för parlamentet.
221.
Europaparlamentet uppmanar Olaf att informera parlamentet om upptäckta fall av bedrägerier inom ramen för fastighetspolitiken och att undersöka eventuella intressekonflikter.
222.
Europaparlamentet uppmanar kommissionen att genomföra en revision av fastighetsförvaltningen, inte bara för kommissionen utan för Europeiska gemenskapernas samtliga institutioner och att undersöka möjligheten till en gemensam fastighetsförvaltning.
Följdåtgärder i samband med beviljandet av ansvarsfrihet
223.
Europaparlamentet beklagar att kommissionen i Europeiska gemenskapernas årsredovisning för 2007 EUT C 287, 10.11.2008, s.
9.
SLUTSATSER OM REVISIONSRÄTTENS SÄRSKILDA RAPPORTER
Del I: ärskild rapport nr 6/2007 om det tekniska biståndets ändamålsenlighet vid kapacitetsutveckling
224.
Europaparlamentet anser att tekniskt bistånd och andra former av externt bistånd, som fortfarande i stor utsträckning styrs av givarna, ofta är ineffektivt och ohållbart och omedelbart behöver reformeras, bl.a. genom att främja lokalt egenansvar, effektivare samordning av resurser mellan medlemsstaterna på EU-nivå och internationell nivå och genom att se till att det avsätts tillräckligt med tid för att genomföra projekt.
225.
226.
227.
228.
Europaparlamentet beklagar att upphävandeklausulen, som möjliggör ett påskyndat upphandlingsförfarande, knappt används av kommissionen och uppmanar den att använda denna möjlighet klokt för att förbättra tidplanen för genomförandet av tekniska biståndsinsatser.
229.
230.
12.
och beslut 2008/969/EG, Euratom av den 16 december 2008 om systemet för tidig varning som ska användas av kommissionens utanordnare och genomförandeorgan EUT L 344, 20.12.2008, s.
125.
231.
Parlamentet uppmanar därför kommissionen att se till att dessa åtaganden snabbt uppfylls på grundval av den strategiska dialog som förutses inom ramen för de arbetsområden som diskuterades i Accra och efter Accra och åtgärderna inom arbetsplanen (axel 1, särskilt åtgärd 20).
232.
Europaparlamentet uppmanar kommissionen att i så stor utsträckning som möjligt följa sina öppenhetsinitiativ och att ta hänsyn till parlamentets resolution av den 19 februari 2008 om öppenhet i ekonomiska frågor Antagna texter, P6_TA(2008)0051 .
och rekommenderar att det inrättas en databas som ger en översikt över tekniska biståndsuppdrag och resultat som går att använda i kommande tekniska biståndsuppdrag och för att förhindra dubbelarbete.
Del II: Särskild rapport nr 1/2008 om förfarandena för utredning och utvärdering av större investeringsprojekt under programperioderna 1994–1999 och 2000–2006
233.
234.
Europaparlamentet uppmanar kommissionen att avlägga fullständiga rapporter om tillämpningen i praktiken av n+2- och n+3-bestämmelserna för större projekt, eftersom vissa länder har försökt "kringgå" ERUF-bestämmelserna (närmare bestämt n+2-bestämmelsen) genom att slå samman ett antal projekt så att deras totalsumma hamnar precis under tröskelvärdet för större projekt och sedan invänta att kommissionen fattar ett beslut om att upphäva n+2-bestämmelsen för projektet i fråga.
235.
236.
237.
238.
Del III: ärskild rapport nr 2/2008 om bindande klassificeringsbesked
239.
Europaparlamentet insisterar på att kommissionen måste anstränga sig för att snarast åtgärda de återstående problemen och svagheterna eftersom de kan leda till inkomstförluster för EU i form av traditionella egna medel.
240.
Europaparlamentet noterar kommissionens svar att den moderniserade tullkoden, som antogs 2008 Europaparlamentets och rådets förordning (EG) nr 450/2008 av den 23 april 2008 om fastställande av en tullkodex för gemenskapen (Moderniserad tullkodex) (EUT L 145, 4.6.2008, s.
1).
, kommer att innebära att de bindande klassificeringsbeskeden blir obligatoriska för innehavaren, uppdateringsarbetet för ordlistan kommer att fortsätta och att användargränssnittet finns tillängligt på samtliga officiella EU-språk.
241.
Europaparlamentet uppmanar kommissionen att se till att konflikter i fråga om tullklassificering blir lösta inom de tidsfrister som fastställs i gemenskapslagstiftningen och senast inom fem månader, och uppmanar dessutom kommissionen att med hänsyn till eventuella förluster av egna medel utöka personalen som arbetar med de bindande klassificeringsbeskeden och klassificering till 4 personer och se till att dessa även utför fler riskanalyser och mer noggrant kontrollerar medlemsstaternas bidrag till systemet, eventuella fall av missbruk av anstånd och fall där aktörer ser sig om efter de mest fördelaktiga bindande klassificeringsbeskeden.
242.
Europaparlamentet uppmanar kommissionen att informera det före utgången av 2009 om alla åtgärder som har vidtagits på grundval av revisionsrättens iakttagelser och om deras genomförande.
Del IV: Särskild rapport nr 3/2008 om Europeiska unionens solidaritetsfond: hur snabb, effektiv och flexibel är den?
243.
Europaparlamentet välkomnar revisionsrättens överlag positiva bedömning av kommissionens resultat i fråga om Europeiska unionens solidaritetsfond.
244.
Europaparlamentet konstaterar att kritiken i fråga om "snabbhet" inte enbart kan hänföras till kommissionens förvaltning av fonden eftersom problemen ofta är förknippade med brister i medlemsstaternas förvaltning, t.ex. när det gäller kvaliteten i den information som de sökande lämnar in.
245.
Europaparlamentet konstaterar också att det i sin ståndpunkt av den 18 maj 2006 EUT C 297 E, 7.12.2006, s.
331.
ställde sig positivt till förslaget till Europaparlamentets och rådets förordning om inrättande av Europeiska unionens solidaritetsfond ( KOM(2005)0108 ) som innehåller enklare och tydligare kriterier för att kunna aktivera fonden snabbare och som rådet hittills inte har gått vidare med.
Del V: Särskild rapport nr 4/2008 om genomförandet av mjölkkvoter i de medlemsstater som anslöt sig till Europeiska unionen den 1 maj 2004
246.
7).
som minskar kontrollprocenten till 1 procent för producenter vars produktion understiger 5 000 kilo.
247.
Europaparlamentet anser att kommissionen inom ramen för den delade förvaltningen måste fortsätta att ta alla de initiativ som krävs för att säkerställa en effektiv övervakning av införandet och förvaltningen av systemet med mjölkkvoter.
248.
Europaparlamentet uppmanar de behöriga nationella myndigheterna att på grundval av en riskanalys upprätta en kontrollplan för varje tolvmånadersperiod och att utföra kontroller under och efter kvotåret men senast 18 månader efter aktuellt regleringsår.
249.
Europaparlamentet anser att kommissionen i förenklingssyfte bör uppmana de nya medlemsstaterna att se till att den allmänna principen enligt vilken all saluförd mjölk ska bokföras efterlevs.
250.
Europaparlamentet uppmanar kommissionen att uppmana de nya medlemsstaterna att förbättra underhållet av databaserna i enlighet med revisionsrättens begäran i sin rapport och att undvika onödiga kontroller.
251.
Europaparlamentet uppmanar kommissionen att fortsätta att utvärdera utvecklingen inom mjölksektorn, särskilt vad avser dess marknad, producenternas situation och konsekvenserna av den fysiska planeringen och detta inom ramen för de utvärderingsrapporter som ska läggas fram före den 31 december 2010 och före den 31 december 2012 enligt den politiska överenskommelsen från november 2008 om "hälsokontrollen" av den gemensamma jordbrukspolitiken.
252.
Europaparlamentet uppmanar kommissionen att följa samtliga rekommendationer från revisionsrätten i fråga om denna "hälsokontroll" och att särskilt inrikta sina överväganden om vilka justeringar som kan göras av den gemensamma organisationen av marknaden för mjölk och systemet för mjölkkvoter på följande punkter:
a)
Kompletterande åtgärder och övergångsåtgärder i regioner där små producenter fortfarande är i stor majoritet.
b)
Behovet för mjölkproducenter att ha ett stabilt regelverk och tydliga utvecklingsmöjligheter som uppmuntrar dem att göra nödvändiga investeringar för att säkerställa verksamhetens bärkraftighet.
Del VI: Särskild rapport nr 5/2008 om unionens tillsynsmyndigheter: att uppnå resultat
253.
Europaparlamentet välkomnar revisionsrättens särskilda rapport och rekommenderar kraftfullt kommissionen att beakta de brister som identifierats i rapporten och vidta åtgärder i enlighet med revisionsrättens rekommendationer.
254.
255.
Europaparlamentet uppmanar kommissionen att införa ett operativt kontrollsystem för EU:s organ som möjliggör intern överföring av bästa praxis och metoder och som omfattar en uppsättning av såväl generella som specifika utvärderingsindikatorer.
256.
Europaparlamentet uppmanar kommissionen att ta fram riktlinjer för att förbättra planering, kontroll, utformning av rapporter och utvärdering av organens verksamhet och att fullt ut genomföra begreppet väntade resultat som införs genom förordning (EG, Euratom) nr 1605/2002 och rambudgetförordningen för organen Kommissionens förordning (EG, Euratom) nr 2343/2002 av den 23 december 2002 om rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002 med budgetförordning för Europeiska gemenskapernas allmänna budget (EUT L 357, 31.12.2002, s.
72).
.
Del VII: Särskild rapport nr 6/2008 om Europeiska kommissionens återanpassningsstöd efter tsunamin och orkanen Mitch
257.
Europaparlamentet uppmanar kommissionen att dra alla slutsatser som krävs av erfarenheterna efter orkanen Mitch och tsunamin för att förbättra framtida insatser och råder kommissionen att spela en aktiv roll på internationell nivå för att åtgärda de systemiska svagheterna i de internationella resurserna för katastrofinsatser.
258.
Europaparlamentet uppmanar kommissionen att särskilt uppmärksamma följande frågor i sina framtida återanpassningsinsatser: att garantera att finansieringen bygger på behoven, att säkerställa att den drabbade befolkningen – inklusive fattiga, kvinnor och barn – står i centrum för hjälpinsatserna och att se till att detaljerad och korrekt information om resultatet av biståndet finns tillgänglig för bidragsgivarna i givarländerna och de drabbade länderna.
259.
Europaparlamentet uppmanar de nationella revisionsorganen och revisionsrätten att förstärka samarbetet för att utreda, revidera och utvärdera användningen av biståndsmedlen vid naturkatastrofer.
260.
Europaparlamentet uppmanar kommissionen att revidera sin förteckning över icke-statliga organisationer för att utesluta de organisationer som den saknar förtroende för och att utforma en upphandlingspolicy för att förhindra att dessa icke-statliga organisationer förskingrar medel.
261.
Europaparlamentet uppmanar dessutom kommissionen att göra EU:s bistånd tillräckligt synligt utan att för den skull äventyra den övergripande effektiviteten och rättvisemålen.
262.
Europaparlamentet uppmanar FN, Röda korset, Röda halvmånen och alla andra givare att enas om en detaljerad ram för kontroll och revision för att
a)
intensifiera och förbättra den övergripande kontrollen över insamlade medel,
b)
undanröja dubbelarbete eller fragmentering av kontrollförfaranden och minska sina kostnader.
263.
Europaparlamentet förväntar sig att kommissionen inte bara godtar revisionsrättens rekommendationer utan även anger att de kommer att genomföras inom en snar framtid.
264.
Europaparlamentet anser också att det är nödvändigt att kommissionen i fråga om humanitärt bistånd ser till att kriterierna för biståndseffektivitet respekteras så som de fastställs i Parisförklaringen om biståndseffektivitet.
265.
Europaparlamentet uppmanar kommissionen att fastställa en realistisk och konkret tidsgräns för hur länge medlen ska finnas tillgängliga för att motivera mottagarländerna att genomföra de godkända projekten i tid.
266.
Europaparlamentet anser att humanitärt bistånd bör erbjudas utan politiska villkor vid naturkatastrofer, men anser ändå att kommissionen bör kräva av mottagarländerna att
a)
möjligheten att nå offren inte begränsas,
b)
biståndet är undantaget från skatter, tullavgifter och alla andra skattepålagor,
c)
viseringar för personal från internationella biståndsorgan inte fördröjs eller avslås,
d)
stödmottagarna inte tvingas betala för donerade varor och tjänster (eller att sådana intäkter i sin helhet återinvesteras i återuppbyggnaden).
267.
Europaparlamentet uppmanar kommissionen att överväga att avbryta biståndet om ovannämnda principer inte följs.
Del VIII: Särskild rapport nr 7/2008 om programmet "Intelligent energi - Europa 2003–2006"
268.
Europaparlamentet välkomnar revisionsrättens seriösa arbete och dess slutsatser som innehåller visst beröm men även kritik av hur kommissionen och Exekutiva byrån för intelligent energi har förvaltat programmet Intelligent energi – Europa (IEE-programmet) 2003-2006 och uppskattar byråns, revisionsrättens och parlamentets nära och framtidsinriktade samarbete med parlamentet.
269.
Europaparlamentet drar slutsatsen av revisionsrättens analys att kostnader som bärs av stödmottagarna (för att utarbeta förslag och rapporter) är ganska höga och även om parlamentet förstår att dessa kostnader skiljer sig från rent administrativa kostnader förordar det att även dessa beaktas och minskas i enlighet med principerna för bättre lagstiftning.
270.
Europaparlamentet anser att revisionsrättens slutsatser också kan vara användbara för andra genomförandeorgan och ser fram emot revisionsrättens kommande särskilda rapport om genomförandeorganen.
271.
Del IX: Särskild rapport nr 8/2008 – Är tvärvillkoren ändamålsenliga?
272.
Europaparlamentet anser att målet med rådets förordning (EG) nr 1782/2003 Rådets förordning (EG) nr 1782/2003 av den 29 september 2003 om upprättande av gemensamma bestämmelser för system för direktstöd inom den gemensamma jordbrukspolitiken och om upprättande av vissa stödsystem för jordbrukare (EUT L 270, 21.10.2003, s.
273.
Europaparlamentet anser att regelverket för tvärvillkor bör förenklas genom att begränsas till de huvudsakliga jordbruksverksamheter som man vill förbättra och genom att förväntade resultat, krav och normer specificeras.
274.
275.
276.
277.
Europaparlamentet uppmanar kommissionen att lägga fram förslag senast i samband med budgetöversynen och nästa reform av den gemensamma jordbrukspolitiken.
278.
Europaparlamentet uppmanar revisionsrätten att rapportera om hur tvärvillkoren uppfylls i sin årsrapport (revisionsförklaring).
Del X: Särskild rapport nr 9/2008 – EU-stödets ändamålsenlighet på området för frihet, säkerhet och rättvisa i Vitryssland, Moldavien och Ukraina
279.
Europaparlamentet uppmanar kommissionen att göra en fullständig analys av anledningarna till bristerna och avsaknaden av resultat i vissa projekt i Vitryssland, Moldavien och Ukraina och att förbättra planeringen, förvaltningen och kontrollen av EU-medel i dessa länder.
280.
Europaparlamentet kräver att kommissionen ska fortsätta att styra EU-medlen mot de särskilda prioriteringarna för Vitryssland, Moldavien och Ukraina med hänsyn till framstegen i föregående projekt.
281.
Europaparlamentet uppmanar kommissionen att öka flexibiliteten i gemenskapens finansieringsförfaranden, vilket skulle göra det möjligt att justera projekthandlingar, riktmärken och mål för att avspegla förändringar i ländernas ekonomiska och politiska situation.
282.
Europaparlamentet kräver att kommissionen säkerställer hållbarheten i EU-finansierade projekt genom att tydligt definiera mottagarregeringens åtaganden vid slutet av projektet.
283.
Europaparlamentet beklagar att gemenskapsmedlen inte har varit tillräckligt ändamålsenliga i fall där det, trots att det förekom tillkortakommanden i projektförvaltningen, beviljades bidrag till samma kontraktspart för nya projekt, och uppmanar därför kommissionen att fastställa tydliga kriterier för att välja kontraktsparter och för att undvika att en otillfredsställande förvaltning av gemenskaps medel upprepas.
284.
Europaparlamentet rekommenderar att kommissionen ska förbättra sin kommunikation med regeringarna i Vitryssland, Moldavien och Ukraina, och och vidta lämpliga åtgärder för att uppmuntra och bistå medlemsstaterna i att inrätta och utöva effektiv samordning mellan givarna.
285.
Europaparlamentet uppmuntrar kommissionen att i högre grad inrikta sig på en effektiv lagföring i kampen mot organiserad brottslighet och att undersöka möjligheten att öka allmänhetens delaktighet i korruptionsbegränsningspolitiken genom att stödja det civila samhällets organisationer i frågor som berör domarkårens oberoende och god samhälssstyrning.
Del XI: Särskild rapport nr 11/2008 om förvaltningen av Europeiska unionens stöd till offentlig lagring av spannmål
286.
Europaparlamentet håller med revisionsrätten om att kommissionen bör ta hänsyn till lagerlokalernas geografiska läge och framför allt spannmålspartiernas kvalitet när den fastställer det lägsta avyttringspriset.
287.
För att förbättra budgetprocessen uppmanar Europaparlamentet kommissionen att öka insynen i kostnader för verksamheter som inte är direkt relaterade till interventionslagring av spannmål och föreslår därför att stödkomponenten i programmen, som stödet till de sämst ställda eller till bioetanolindustrin, fördelas direkt till de berörda verksamheterna.
288.
Europaparlamentet uppmanar medlemsstaterna och kommissionen att utvärdera kostnaderna för kontroller på området för offentlig lagring av spannmål, och uppmanar kommissionen att skapa större incitament för medlemsstaterna att minska lagren och kapitalkostnaderna för sina interventioner och att sälja sina lager vid bästa möjliga tidpunkt.
289.
290.
Europaparlamentet stöder revisionsrättens uppfattning att inspektioner på plats för att kontrollera kostnadsuppgifter från medlemsstaternas utbetalande organ skulle vara användbara, men betonar emellertid att det måste garanteras att kontrollkraven är kostnadseffektiva.
291.
P6_TA-PROV(2009)0375
Europeiska flyktingfonden för perioden 2008–2013 (ändring av beslut nr 573/2007/EG) ***I
A6-0280/2009
Europaparlamentets lagstiftningsresolution av den 7 maj 2009 om förslaget till Europaparlamentets och rådets beslut om ändring av beslut nr 573/2007/EG om inrättande av Europeiska flyktingfonden för perioden 2008–2013 och om avskaffande av finansieringen av vissa gemenskapsåtgärder samt om nya gränser för högsta tillåtna finansiering ( KOM(2009)0067 – C6-0070/2009 – 2009/0026(COD) )
(Medbeslutandeförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2009)0067 ),
–
–
med beaktande av artikel 51 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor och yttrandet från budgetutskottet ( A6-0280/2009 ).
1.
Europaparlamentet godkänner kommissionens förslag.
2.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om kommissionen har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
3.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
som ersätter resolutionsförslagen från grupperna:
PPE ( B7‑0041/2010 )
ALDE ( B7‑0040/2010 )
Verts/ALE ( B7‑0055/2010 )
ECR ( B7‑0054/2010 )
GUE/NGL ( B7‑0053/2010 )
EFD ( B7‑0051/2010 )
om brott mot de mänskliga rättigheterna i Kina, särskilt fallet Liu Xiaobo
Tunne Kelam
,
Mario Mauro
,
Laima Liucija Andrikienė
,
Cristian Dan Preda
,
Bernd Posselt
,
Filip Kaczmarek
,
Eija-Riitta Korhola
,
Monica Luisa Macovei
,
Jean-Pierre Audy
,
László Tőkés
,
Elżbieta Katarzyna Łukacijewska
för PPE-gruppen
Renate Weber
,
Frédérique Ries
,
Ramon Tremosa i Balcells
,
Marielle De Sarnez
för ALDE-gruppen
Heidi Hautala
,
Barbara Lochbihler
,
Helga Trüpel
,
Philippe Lamberts
,
Daniel Cohn-Bendit
för Verts/ALE-gruppen
Charles Tannock
för ECR-gruppen
Marie-Christine Vergiat
,
Gabriele Zimmer
för GUE/NGL-gruppen
Fiorello Provera
för EFD-gruppen
Edward McMillan-Scott
PE432.888v01-00 } PE432.889v01-00 } PE432.899v01-00 } PE432.901v01-00 } PE432.902v01-00 } PE432.903v01-00 } RC1 Europaparlamentets resolution om brott mot de mänskliga rättigheterna i Kina, särskilt fallet Liu Xiaobo
Europaparlamentet utfärdar denna resolution
– med beaktande av sina tidigare resolutioner om Kina, i synnerhet av den 13 december 2007 om toppmötet EU/Kina och om EU–Kina-dialogen om mänskliga rättigheter och av den 26 november 2009 om minoriteters rättigheter och tillämpningen av dödsstraff,
– med beaktande av sin resolution av den 6 september 2007 om hur dialogerna och samråden om mänskliga rättigheter fungerar med tredjeländer,
– med beaktande av ordförandeskapets uttalande för EU av den 19 december 2008 om Charta 2008 och arresteringen av människorättsaktivister,
– med beaktande av toppmötet mellan EU och Kina i Prag 2009,
– med beaktande av ordförandeskapets uttalanden för EU av den 26 juni 2009 och den 14 december 2009 om åtalet mot Liu Xiaobo,
– med beaktande av EU–Kina-seminariet den 18–19 november 2009 och EU–Kina-dialogen om mänskliga rättigheter den 20 november 2009,
– med beaktande av ordförandeskapets uttalande för EU av den 29 december 2009 om avrättningen av Akmal Shaikh,
A. Liu Xiaobo, en framstående människorättsaktivist och akademiker samt medförfattare till Charta 2008, blev den 8 december 2008 på hemlig ort i Peking föremål för en form av häktning som kan användas i upp till sex månader utan att åtal väcks.
E. Liu Xiaobos hustru samt personal från ett dussintal olika ambassader i Peking begärde tillstånd att observera rättegången men nekades tillträde till rättegångssalen.
F. Domen har rönt omfattande kritik från inhemska Internetbloggare, internationella medborgargrupper samt utländska regeringar, och den har även överklagats av Liu Xiaobo.
G. Tjeckiens förre president Václav Havel nekades tillträde till Kinas ambassad i Prag när han ville vädja om frigivning av Liu Xiaobo.
H. De kinesiska myndigheterna hörsammade inte de upprepade kraven från EU och en av dess medlemsstater om att dödsdomen mot Akmal Shaikh skulle omvandlas.
I. För några dagar sedan erkände för första gången en kinesisk tjänsteman att Gao Zhiseng, en kristen människorättsaktivist som nominerats till Nobels fredspris, försvunnit.
J. I december 2009 ägde andra människorättsbrott rum i Kina, exempelvis trakasserier mot medlemmar av människorättsforumet Guizhou, som skulle hindras från att genomföra planerade aktiviteter med anledning av människorättsdagen, samt våld och misshandel av den frihetsberövade Qi Choghuai, reporter och tidigare chef för Fazhi Morning Posts redaktion i Shandong.
L. I april 2009 lämnade Kina in ett dokument till FN som syftade till att stärka landets kandidatur avseende medlemskap i människorättsrådet och enligt vilket Kina förbinder sig att främja och skydda det kinesiska folkets mänskliga rättigheter och grundläggande friheter.
M. Den 13 januari 2010 tillkännagav Google sin avsikt att avbryta samarbetet med den kinesiska Internetcensuren med anledning av de sofistikerade cyberattacker mot företagets datorsystem som man misstänkte hade sitt ursprung i Kina och som delvis var riktade mot människorättsaktivisters Gmail-konton.
Europaparlamentet uppmanar enträget Kina att säkerställa respekten för de mänskliga rättigheterna och grundläggande friheterna och kräver att landet ratificerar den internationella konventionen om medborgerliga och politiska rättigheter.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till unionens höga representant för utrikes frågor och säkerhetspolitik, Europeiska rådets ordförande, kommissionen samt Kinas president, premiärminister och nationella folkkongress.
som ersätter resolutionsförslagen från följande grupper:
Verts/ALE ( B7‑0413/2010 )
PPE ( B7‑0429/2010 )
S&D ( B7‑0430/2010 )
ALDE ( B7‑0431/2010 )
GUE/NGL ( B7‑0432/2010 )
om ikraftträdandet av konventionen mot klustervapen och EU:s roll
Elmar Brok
,
José Ignacio Salafranca Sánchez-Neyra
,
Michael Gahler
,
Arnaud Danjean
för PPE-gruppen
Adrian Severin
,
Roberto Gualtieri
,
Ana Gomes
,
María Muñiz De Urquiza
för S&D-gruppen
Johannes Cornelis van Baalen
,
Elizabeth Lynne
,
Sonia Alfano
för ALDE-gruppen
Ulrike Lunacek
,
Raül Romeva i Rueda
,
Barbara Lochbihler
,
Reinhard Bütikofer
för Verts/ALE-gruppen
Sabine Lösing
,
Willy Meyer
,
Helmut Scholz
,
Nikolaos Chountis
,
Takis Hadjigeorgiou
,
Kyriacos Triantaphyllides
för GUE/NGL-gruppen
PE442.011v01-00 } PE442.027v01-00 } PE442.028v01-00 } PE442.029v01-00 } PE442.030v01-00 } RC1 Europaparlamentets resolution om ikraftträdandet av konventionen mot klustervapen och EU:s roll
Europaparlamentet utfärdar denna resolution,
– med beaktande av konventionen om klustervapen som antogs av 107 länder vid den diplomatiska konferensen i Dublin den 19–30 maj 2008,
– med beaktande av att FN:s generalsekreterare i ett meddelande av den 30 maj 2008 uppmuntrade staterna att så snart som möjligt underteckna och ratificera detta viktiga avtal och sade att han ser fram emot att det kommer att träda i kraft inom kort,
A. Konventionen mot klustervapen har stått öppen för undertecknande sedan den 3 december 2008, först i Oslo och därefter vid FN:s högkvarter i New York, och den kommer att träda i kraft den första dagen i den sjätte månaden efter det att den har ratificerats av 30 stater, det vill säga den 1 augusti 2010.
B. I konventionen mot klustervapen definieras klustervapen som vapen som är utformade för att sprida eller släppa explosiva substridsdelar, som var och en väger mindre än 20 kg, och innefattar dessa explosiva substridsdelar.
C. Konventionen mot klustervapen kommer att förbjuda användning, tillverkning, lagring och överföring av klustervapen, och förbudet kommer att avse vapenkategorin.
D. Enligt konventionen mot klustervapen måste de undertecknande staterna förstöra de klustervapen som de har i lager.
E. Konventionen om klustervapen fastställer nya humanitära normer rörande stöd till offer, och ålägger de berörda staterna att avlägsna alla rester av odetonerade klustervapen som ligger kvar efter konflikter.
G. Fram till dags dato har tjugo EU-medlemsstater undertecknat konventionen mot klustervapen och elva har ratificerat den, medan sju varken har undertecknat eller ratificerat den.
H. När konventionen mot klustervapen träder i kraft den 1 augusti 2010 kommer det att bli besvärligare att ansluta sig till konventionen, eftersom staterna måste ansluta sig till konventionen i en process som består av ett steg.
I. Stödet från flertalet av EU-medlemsstaterna, interparlamentariska initiativ och ett stort antal organisationer i det civila samhället har på ett avgörande sätt bidragit till att Osloprocessen kunde resultera i konventionen mot klustervapen.
J. Om alla 27 EU-medlemsstater undertecknar och ratificerar konventionen mot klustervapen innan den träder i kraft den 1 augusti 2010 skulle detta bli en stark politisk signal till stöd för en värld utan klustervapen och för EU:s mål i kampen mot spridning av vapen som dödar urskillningslöst.
Europaparlamentet berömmer de stater som har undertecknat och ratificerat konventionen, vilka också har antagit ett moratorium mot användning, tillverkning och överföring av klustervapen samt förstört sina lager av dessa vapen.
Europaparlamentet uppmanar alla stater att delta i det första mötet mellan de undertecknande staterna, vilket kommer att hållas den 8–12 november 2010 i Vientiane i Laos, landet med världens största koncentration av odetonerade klusterbomber.
Europaparlamentet uppmanar rådet och kommissionen att införa förbudet mot klustervapen som en standardklausul i avtal med tredjeländer vid sidan av standardklausulen om icke-spridning av massförstörelsevapen.
13.
Europaparlamentet uppmanar EU:s medlemsstater, rådet och kommissionen att vidta åtgärder för att hindra tredjeländer från att förse icke-statliga aktörer med klustervapen.
som ersätter resolutionsförslagen från grupperna:
EFD ( B7‑0518/2010 )
S&D ( B7‑0519/2010 )
ALDE ( B7‑0520/2010 )
Verts/ALE ( B7‑0521/2010 )
PPE ( B7‑0523/2010 )
om den europeiska strategin för ekonomisk och social utveckling i bergsregioner, öregioner och glesbefolkade regioner
Lambert van Nistelrooij
,
Maurice Ponga
,
Marie-Thérèse Sanchez-Schmid
,
Nuno Teixeira
,
Rosa Estaràs Ferragut
,
Eleni Theocharous
,
Danuta Maria Hübner
,
Jean-Pierre Audy
,
Antonio López-Istúriz White
,
Veronica Lope Fontagné
för PPE-gruppen
Constanze Angela Krehl
,
Georgios Stavrakakis
,
Marita Ulvskog
,
Saïd El Khadraoui
,
Kriton Arsenis
,
Teresa Riera Madurell
,
Maria Badia i Cutchet
för S&D-gruppen
Riikka Manner
,
Ramona Nicole Mănescu
,
Pat the Cope Gallagher
,
Giommaria Uggias
,
Anneli Jäätteenmäki
,
Hannu Takkula
,
Carl Haglund
,
Niccolò Rinaldi
för ALDE-gruppen
François Alfonsi
för Verts/ALE-gruppen
Bairbre de Brún
,
Marisa Matias
för GUE/NGL-gruppen
Fiorello Provera
,
Lorenzo Fontana
för EFD-gruppen
PE446.607v01-00 } PE446.609v01-00 } PE446.610v01-00 } PE446.611v01-00 } PE446.613v01-00 } RC1 Europaparlamentets resolution om den europeiska strategin för ekonomisk och social utveckling i bergsregioner, öregioner och glesbefolkade regioner
Europaparlamentet utfärdar denna resolution
– med beaktande av avdelning XVIII i fördraget om Europeiska unionens funktionssätt och särskilt artikel 174,
– med beaktande av de förordningar som reglerar strukturfonderna för perioden 2007–2013,
– med beaktande av rådets beslut av den 6 oktober 2006 om gemenskapens strategiska riktlinjer för sammanhållningen EUT L 291, 21.10.2006, s.
11.
,
– med beaktande av sin resolution av den 2 september 2003 om regioner med strukturella nackdelar (öar, bergsområden och glesbygder) inom ramen för sammanhållningspolitiken och de institutionella perspektiven EUT C 76 E, 25.3.2004, s.
111.
,
– med beaktande av Regionkommitténs yttrande av den 7 juli 2005 om översynen av riktlinjerna för nationellt regionalstöd,
– med beaktande av sin resolution av den 15 mars 2007 om öarna och naturliga och ekonomiska hinder inom ramen för regionalpolitiken EUT C 301 E, 13.12.2007, s.
244.
,
– med beaktande av kommissionens meddelande av den 6 oktober 2008 med titeln ”Grönbok om territoriell sammanhållning – Att omvandla territoriell mångfald till styrka” ( KOM(2008)0616 ),
– med beaktande av kommissionens arbetsdokument ”Regions 2020 – an assessment of future challenges for EU regions” (Regioner 2020 – En bedömning av de framtida utmaningarna för EU:s regioner) ( SEK(2008)2868 ),
– med beaktande av sin resolution av den 24 mars 2009 om grönboken om den territoriella sammanhållningen och en lägesanalys av debatten om den framtida reformen av sammanhållningspolitiken Antagna texter, P6_TA(2009)0163 .
,
– med beaktande av kommissionens meddelande av den 25 juni 2009 om den sjätte rapporten om ekonomisk och social sammanhållning ( KOM(2009)0295 ),
– med beaktande av kommissionens meddelande av den 31 mars 2010 med titeln ”Sammanhållningspolitiken: Strategirapport 2010 om genomförandet av programmen 2007‑2013” ( KOM(2010)0110 ),
– med beaktande av artikel 110.4 i arbetsordningen, och av följande skäl:
2.
4.
Europaparlamentet begär att man fastställer en särskild europeisk integrerad och flexibel politisk ram, med rättsliga och finansiella konsekvenser, så att bergsregioner, öregioner och glesbefolkade regioner kan behandlas med utgångspunkt i deras gemensamma drag, samtidigt som vederbörlig hänsyn tas både till deras olika förutsättningar och till proportionalitetsprincipen.
Parlamentet anser att öregionernas situation bör tas upp inom sammanhållningspolitiken, inte bara via regionalpolitiken, utan också med hjälp av annan EU-politik som har en klar territoriell inverkan på utvecklingen i dessa regioner.
Parlamentet anser vidare att en europeisk politisk ram för bergsregioner, öregioner och glesbefolkade regioner kan ha det mervärde som behövs för att dessa regioners permanenta nackdelar ska kunna övervinnas och utvecklingsmodellen för dem anpassas utgående från deras resurser.
Ett vertikalt angreppssätt, där alla myndighetsnivåer deltar och där subsidiaritetsprincipen beaktas, är nämligen nödvändigt för att dessa regioner ska kunna slå in på den rätta vägen för hållbar utveckling och för att man samtidigt ska kunna beakta andra viktiga sektorer i regionen.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att se till att bergsregioner, öregioner och glesbefolkade regioner också i fortsättningen omfattas av särskilda föreskrifter, även inom den nya budgetplanen och under nästa programplaneringsperiod.
Europaparlamentet uppmanar medlemsstaterna att fullt ut utnyttja det europeiska grannskapsinstrumentet i bergsregioner, glesbefolkade regioner och öregioner, för att de ska kunna dra nytta av de resurser som finns tillgängliga över gränserna.
som ersätter resolutionsförslagen från grupperna:
EFD ( B7‑0637/2010 )
S&D ( B7‑0638/2010 )
ALDE ( B7‑0640/2010 )
ECR ( B7‑0642/2010 )
Verts/ALE ( B7‑0643/2010 )
PPE ( B7‑0644/2010 )
om Tibet – planer på att göra kinesiskan till huvudsakligt undervisningsspråk
Elmar Brok
,
José Ignacio Salafranca Sánchez-Neyra
,
Thomas Mann
,
Mario Mauro
,
Cristian Dan Preda
,
Bernd Posselt
,
Laima Liucija Andrikienė
,
Csaba Sógor
,
Filip Kaczmarek
,
Lena Kolarska-Bobińska
,
Róża Gräfin von Thun und Hohenstein
,
Eija-Riitta Korhola
,
Monica Luisa Macovei
,
Elena Băsescu
,
Tunne Kelam
,
Bogusław Sonik
,
Sari Essayah
,
Martin Kastler
för PPE-gruppen
Véronique De Keyser
,
Lidia Joanna Geringer de Oedenberg
för S&D-gruppen
Marietje Schaake
,
Niccolò Rinaldi
,
Graham Watson
,
Ramon Tremosa i Balcells
,
Frédérique Ries
,
Leonidas Donskis
,
Renate Weber
,
Edward McMillan-Scott
,
Sarah Ludford
,
Antonyia Parvanova
,
Kristiina Ojuland
,
Marielle De Sarnez
,
Sonia Alfano
för ALDE-gruppen
Heidi Hautala
,
Eva Lichtenberger
,
Raül Romeva i Rueda
,
François Alfonsi
,
Frieda Brepoels
,
Catherine Grèze
för Verts/ALE-gruppen
Charles Tannock
,
Michał Tomasz Kamiński
,
Konrad Szymański
,
Tomasz Piotr Poręba
,
Marek Henryk Migalski
,
Ryszard Czarnecki
,
Adam Bielan
,
Roberts Zīle
för ECR-gruppen
Fiorello Provera
för EFD-gruppen
PE450.473v01-00 } PE450.474v01-00 } PE450.476v01-00 } PE450.478v01-00 } PE450.479v01-00 } PE450.480v01-00 } RC1 Europaparlamentets resolution om Tibet – planer på att göra kinesiskan till huvudsakligt undervisningsspråk
Europaparlamentet utfärdar denna resolution
– med beaktande av sina tidigare resolutioner om Kina och Tibet, särskilt resolutionen av den 10 april 2008 om Tibet,
A. Respekten för de mänskliga rättigheterna, identitets-, kultur- och religionsfrihet, är en grundläggande princip för Europeiska unionen och prioriteras inom Europeiska unionens utrikespolitik.
B. Folkrepubliken Kina har uttryckt en önskan om harmoniska etniska relationer mellan alla 56 etniska minoriteter.
G. Överallt inom den autonoma regionen Tibet håller tibetanskan på att inom lågstadie-, högstadie- och gymnasieundervisningen successivt ersättas av kinesiska och för det mesta går det inte att få tag på officiella handlingar på tibetanska.
H. Omläggningarna i undervisningspolitiken skulle begränsa tibetanskans användning i skolorna, eftersom alla läroböcker och ämnen skulle vara på mandarinkinesiska, med undantag för undervisningen i tibetanska och engelska.
I. Folkrepubliken Kina röstade den 13 september 2007, tillsammans med 142 andra länder, för att godkänna FN:s förklaring om ursprungsfolkens rättigheter, i vars 14 artikel det framför allt står att ”ursprungsfolken har rätt att inrätta och övervaka sitt utbildningsväsen samt inrättningar som bedriver utbildning på deras egna språk, på ett sätt som är lämpligt utgående från deras kulturbetingade metoder för undervisning och lärande.”
J. Till följd av kinesiskans dominans blir personer med universitets- och högskoleexamen i de tibetanska områdena alltmer oroliga inför sina utsikter att få arbete eftersom, såsom det stod i en framställning som undertecknats av lärare och elever, de flesta eleverna och studenterna i Tibet aldrig vistats i en kinesiskspråkig omgivning och därför inte kan kommunicera på kinesiska.
Europaparlamentet noterar oron över försöken att få tibetanskan att framstå som mindre värd och betonar att tibetanskan måste vara inhemskt språk för att den tvåspråkiga undervisningen ska lyckas.
Europaparlamentet uppmanar de kinesiska myndigheterna att göra allt för att minska de språkliga och kulturella nackdelar som tibetaner drabbas av när de söker arbete i städerna, låt vara att detta bör göras på sådant sätt att det inte blir till skada för det tibetanska språket och den tibetanska kulturen.
Europaparlamentet uppmanar än en gång Kina att ratificera Internationella konventionen om medborgerliga och politiska rättigheter och beklagar den ofta diskriminerande behandlingen av etniska och religiösa minoriteter i Kina.
som ersätter resolutionsförslagen från grupperna:
S&D ( B7‑0347/2011 )
ALDE ( B7‑0348/2011 )
PPE ( B7‑0357/2011 )
Verts/ALE ( B7‑0358/2011 )
ECR ( B7‑0359/2011 )
om toppmötet mellan EU och Ryssland
Elmar Brok
,
José Ignacio Salafranca Sánchez-Neyra
,
Ria Oomen-Ruijten
,
Ioannis Kasoulides
,
Alojz Peterle
,
Tunne Kelam
,
Cristian Dan Preda
,
Jacek Saryusz-Wolski
,
Inese Vaidere
,
Vytautas Landsbergis
,
Arnaud Danjean
,
Krzysztof Lisek
,
Michael Gahler
,
Paweł Zalewski
,
Nadezhda Neynsky
,
Zuzana Roithová
,
Andrzej Grzyb
,
Joachim Zeller
,
Giovanni La Via
för PPE-gruppen
Hannes Swoboda
,
Véronique De Keyser
,
Knut Fleckenstein
,
Kristian Vigenin
,
Pino Arlacchi
,
Mitro Repo
för S&D-gruppen
Kristiina Ojuland
,
Leonidas Donskis
,
Marielle De Sarnez
,
Ivo Vajgl
,
Graham Watson
,
Ramon Tremosa i Balcells
,
Anneli Jäätteenmäki
,
Marietje Schaake
,
Edward McMillan-Scott
för ALDE-gruppen
Charles Tannock
,
Ryszard Antoni Legutko
,
Marek Henryk Migalski
,
Paweł Robert Kowal
,
Konrad Szymański
,
Ryszard Czarnecki
,
Geoffrey Van Orden
,
Tadeusz Cymański
för ECR-gruppen
Rebecca Harms
,
Heidi Hautala
,
Werner Schulz
för Verts/ALE-gruppen
PE465.652v01-00 } PE465.653v01-00 } PE465.662v01-00 } PE465.663v01-00 } PE465.664v01-00 } RC1 Europaparlamentets resolution om toppmötet mellan EU och Ryssland
Europaparlamentet utfärdar denna resolution
– med beaktande av det befintliga avtalet om partnerskap och samarbete mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Ryska federationen, å andra sidan EGT L 327, 28.11.1997, s.
1.
, och de förhandlingar som inleddes 2008 om ett nytt avtal mellan EU och Ryssland, samt det partnerskap för modernisering som inleddes 2010,
– med beaktande av det gemensamma mål som EU och Ryssland angav i ett gemensamt uttalande den 31 maj 2003 efter det elfte toppmötet mellan EU och Ryssland som hölls i Sankt Petersburg om att skapa ett gemensamt ekonomiskt område, ett gemensamt område med frihet, säkerhet och rättvisa, ett gemensamt område för samarbete kring yttre säkerhet och ett gemensamt område för forskning och utbildning, vilket även ska inbegripa kulturella aspekter (”de fyra gemensamma områdena”),
– med beaktande av sina tidigare betänkanden och resolutioner om Ryssland och förbindelserna mellan EU och Ryssland, särskilt resolutionerna av den 17 februari 2011 om rättsstatsprincipen Antagna texter, P7_TA-PROV(2011)0066 .
, av den 17 juni 2010 om toppmötet mellan EU och Ryssland Antagna texter, P7_TA(2010)0234 .
, av den 12 november 2009 inför toppmötet mellan EU och Ryssland i Stockholm den 18 november 2009 Antagna texter, P7_TA(2009)0064 .
, av den 17 september 2009 om morden på människorättsaktivister i Ryssland Antagna texter, P7_TA(2009)0022 .
och av den 17 september 2009 om de externa aspekterna av en tryggad energiförsörjning Antagna texter, P7_TA(2009)0021 .
,
– med beaktande av människorättssamrådet mellan EU och Ryssland och dess senaste möte den 4 maj 2011,
– med beaktande av de avtal som undertecknades och de gemensamma uttalanden som gjordes vid toppmötet mellan EU och Ryssland i Rostov-na-Donu den 31 maj–1 juni 2010,
– med beaktande av EU:s höga representant Catherine Ashtons uttalande av den 24 maj 2011 om målet mot Michail Chodorkovskij och Platon Lebedev,
– med beaktande av den gemensamma förklaring som medordförandena för den parlamentariska samarbetskommittén EU-Ryssland utfärdade i Sochi den 18 maj 2011,
– med beaktande av dagordningen för det toppmöte mellan EU och Ryssland som ska hållas i Nizjnij Novgorod den 9–10 juni 2011,
– med beaktande av artikel 110.4 i arbetsordningen, och av följande skäl:
2.
4.
Europaparlamentet hoppas att toppmötet kommer att bidra till att lösa de sista frågorna om Rysslands anslutning till WTO, efter det att EU och Ryssland i december 2010 ingått ett bilateralt avtal för att landet ska kunna gå med i organisationen.
Parlamentet upprepar sitt stöd för Rysslands anslutning till WTO, som kommer att skapa enhetliga förutsättningar för företagsvärlden på båda sidor och underlätta och avreglera handeln i den globala ekonomin.
Europaparlamentet uppmanar Ryssland att respektera de avtal det undertecknat, uppfylla alla åtaganden i sexpunktsavtalet om vapenvila och omedelbart dra tillbaka sina styrkor från de ockuperade georgiska territorierna Sydossetien och Abchazien till de ställningar som rådde före konflikten samt garantera tillträde för Europeiska unionens övervakningsuppdrag (EUMM) till dessa territorier.
som ersätter resolutionsförslagen från grupperna:
S&D ( B7‑0048/2012 )
PPE ( B7‑0049/2012 )
ALDE ( B7‑0051/2012 )
ECR ( B7‑0054/2012 )
om avtalet mellan EU och Marocko om ömsesidiga liberaliseringsåtgärder angående jordbruksprodukter och fiskeriprodukter
Cristiana Muscardini
,
Daniel Caspary
,
Elisabeth Jeggle
för PPE-gruppen
Véronique De Keyser
,
Bernd Lange
,
David Martin
,
Vital Moreira
för S&D-gruppen
Metin Kazak
,
George Lyon
för ALDE-gruppen
Robert Sturdy
för ECR-gruppen
PE479.474v01-00 } PE479.475v01-00 } PE479.477v01-00 } PE479.480v01-00 } RC1 Europaparlamentets resolution om avtalet mellan EU och Marocko om ömsesidiga liberaliseringsåtgärder angående jordbruksprodukter och fiskeriprodukter
Europaparlamentet utfärdar denna resolution
– med beaktande av Barcelonaförklaringen av den 28 november 1995 som inrättade ett partnerskap mellan EU och länderna i södra Medelhavsområdet,
– med beaktande av Europa-Medelhavsavtalet om upprättande av en associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Konungariket Marocko, å andra sidan,
– med beaktande av rådets beslut av den 14 oktober 2005 om bemyndigande av förhandlingar med Marocko om ömsesidiga liberaliseringsåtgärder angående handel med jordbruksprodukter, bearbetade jordbruksprodukter, fisk och fiskeriprodukter,
– med beaktande av rådets beslut av den 14 december 2011 om bemyndigande av förhandlingar med Egypten, Jordanien, Marocko och Tunisien för att upprätta djupgående och omfattande frihandelsområden som en del i de befintliga Europa–Medelhavsavtalen om associering med dessa länder,
– med beaktande av det gemensamma meddelandet från kommissionen till Europeiska rådet, Europaparlamentet, rådet, Europeiska ekonomiska och sociala kommittén samt Regionkommittén av den 8 mars 2011 om ett partnerskap för demokrati och delat välstånd med södra medelhavsområdet, ( KOM(2011)0200 ),
– med beaktande av det gemensamma meddelandet från kommissionen till Europeiska rådet, Europaparlamentet, rådet, Europeiska ekonomiska och sociala kommittén samt Regionkommittén av den 25 maj 2011 om en ny respons på ett grannskap i förändring, ( KOM(2011)0303 ),
– med beaktande av sin resolution av den 25 november 2010 om företagens sociala ansvar vid internationella handelsavtal ( 2009/2201(INI) ) Antagna texter, P7_TA(2010)0446 .
,
– med beaktande av artikel 110.4 i arbetsordningen, och av följande skäl:
2.
Parlamentet anser att Marocko har gjort betydande framsteg för att befästa demokratin genom att reformera sin konstitution och genomföra rättvisa val.
3.
Avtalet
4.
Med tanke på jordbrukssektorns betydelse och inflytande i Marocko, särskilt när det gäller att skapa sysselsättning, betonar Europaparlamentet avtalets viktiga roll för landets ekonomiska utveckling och politiska stabilitet eftersom det erbjuder nya exportmöjligheter till EU, som är den största marknaden för marockanska produkter.
Parlamentet anser att avtalet också kommer att innebära möjligheter för EU:s jordbrukssektor, i synnerhet för bearbetade livsmedel.
Parlamentet påpekar att EU:s exportörer så småningom kommer att dra nytta av att man slopar de marockanska importtullarna för 70 procent av jordbruks- och fiskeriprodukterna, en åtgärd som beräknas medföra besparingar på 100 miljoner euro om året i tullavgifter när denna åtgärd väl genomförts fullt ut.
Parlamentet påminner vidare om att EU och Marocko har enats om en tvistlösningsmekanism som ger båda parter rätt till domstolsprövning om den andra parten inte respekterar villkoren i avtalet.
Parlamentet uppmanar därför kommissionen att lägga fram en bedömning av konsekvenserna för europeiska producenter, och särskilt för jordbrukarnas inkomster, och att ge parlamentet regelbunden information.
Parlamentet efterlyser garantier för att de ökade tullkvoterna enligt avtalet kommer att regleras av EU på lämpligt sätt och att det inte kommer att bli några missförstånd om de bestämmelser som reglerar systemet med ingångspriser.
Parlamentet påpekar att inga formella klagomål har framförts till Olaf sedan 2005.
I detta sammanhang noterar parlamentet förslagen att göra de bestämmelser som reglerar genomförandet av systemet med ingångspriser förenliga med gemenskapens tullkodex som en del i den senaste reformen av den gemensamma jordbrukspolitiken.
Europaparlamentet anser att avtalet innehåller särskilda institutionella arrangemang och mekanismer, exempelvis samarbete i syfte att undvika störningar på marknaderna, expertgrupper som inrättats av kommissionen tillsammans med tredjeländer, bland annat Marocko, underutskottet för jordbrukshandel som inrättats inom ramen för förvaltningen av associeringsavtal, informationsutbyte om strategier och produktion samt säkerhetsklausulen enligt artikel 7 i protokollet.
9.
Europaparlamentet betonar att tillträde till EU:s inre marknad bör bero på om vissa sanitära, fytosanitära och miljömässiga krav är uppfyllda och välkomnar den positiva rapport från Kontoret för livsmedels- och veterinärfrågor som kom 2011.
Parlamentet välkomnar den betydelse sanitära och fytosanitära åtgärder tillmäts i avtalet och vill se att tekniskt bistånd blir en central punkt i förhandlingarna om ett djupgående och omfattande frihandelsavtal.
Kommissionen uppmanas att främja överensstämmelse i åtgärder och kontroller mellan Marocko och Europeiska unionen på området för miljö- och livsmedelssäkerhetsnormer, i syfte att garantera rättvis konkurrens mellan de två marknaderna.
Parlamentet vill se fortsatt EU-stöd för förbättrade produktionsmetoder genom utbyte av bästa praxis, och för Marockos ansträngningar på området för vattenskydd.
Det finns dock fortfarande utrymme för förbättringar i fråga om förenings- och mötesfrihet samt barnarbete.
Parlamentet anser att bestämmelserna i de djupgående och omfattande frihandelsavtalen bör omfatta stöd för tillämpning av ILO:s konventioner, ratificering av ännu inte undertecknade centrala ILO-konventioner (t.ex. konventionen angående föreningsfrihet och skydd för organisationsrätten (nr 87)) samt initiativ rörande företagens sociala ansvar inom ramen för kapitlet om hållbar utveckling.
P7_TA(2009)0029
Effekterna av den globala finansiella och ekonomiska krisen på utvecklingsländerna
B7-0078/2009
Europaparlamentets resolution av den 8 oktober 2009 om effekterna av den globala finansiella och ekonomiska krisen på utvecklingsländerna och utvecklingssamarbetet
Europaparlamentet utfärdar denna resolution
–
med beaktande av G20-toppmötet i London den 2 april 2009 och dess förklaring om en global plan för återhämtning och reform,
–
med beaktande av FN:s millenniedeklaration av den 8 september 2000, i vilken världssamfundet gemensamt fastställde kriterier, bland annat för att utrota fattigdom och svält, i de s.k. millennieutvecklingsmålen,
–
med beaktande av rapporten från Världsbanken och Internationella valutafonden med titeln "Global Monitoring Report 2009: A Development Emergency" som offentliggjordes i april 2009,
–
med beaktande av Världsbankens rapport med titeln "Global Development Finance: Charting a Global Recovery 2009" som offentliggjordes i juni 2009,
–
med beaktande av FN:s konferens om finanskrisen och den ekonomiska krisen i världen och dess följder för utvecklingen, och FN:s generalförsamlings bekräftelse av resultatet av konferensen genom resolution 63/303 av den 9 juli 2009,
–
med beaktande av kommissionens meddelande av den 8 april 2009 om att hjälpa utvecklingsländerna att hantera krisen ( KOM(2009)0160 ),
–
med beaktande av slutsatserna från rådets (allmänna frågor och yttre förbindelser) möte den 18-19 maj 2009 om att hjälpa utvecklingsländerna att hantera krisen,
–
med beaktande av sin resolution av den 14 mars 2006 om den internationella valutafondens strategiska översyn EUT C 291 E, 30.11.2006, s.
118.
,
–
med beaktande av professor Ngaire Woods studie om det internationella gensvaret på den globala krisen och reformen av de globala finans- och stödstrukturerna En studie som beställts av utredningsavdelningen vid Europaparlamentets generaldirektorat för EU-extern politik och som kommer att offentliggöras.
,
–
med beaktande av konferensen om innovativ finansiering i Paris den 28–29 maj 2009 och den internationella konferensen om utvecklingsfinansiering i Doha den 28 november–2 december 2008.
–
med beaktande av rapporten med titeln "Impact of the Crisis on African Economies – Sustaining Growth and Poverty Reduction" av den 17 mars 2009 från den kommitté av Afrikanska finansministrar och centralbankschefer som fått i uppdrag att övervaka krisen,
–
med beaktande av frågan till kommissionen av den 3 september 2009 om effekterna av den globala finansiella och ekonomiska krisen på utvecklingsländerna och utvecklingssamarbetet ( O-0088/2009 – B7-0209/2009 ),
–
1.
Europaparlamentet betonar att trots att utvecklingsländerna inte förorsakade den globala finansiella och ekonomiska krisen så drabbas de oproportionerligt av den med en dramatisk nedgång i tillväxt och sysselsättning, negativa effekter på handelsbalansen och betalningsbalansen, en kraftig minskning av det privata nettokapitalinflödet och utländska direktinvesteringar, begränsad tillgång till kredit- och handelsfinansiering, minskade penningförsändelser från migranter, stora och häftiga svängningar i växelkurserna, kollapsade reserver, ökad instabilitet och fallande råvarupriser samt minskade inkomster från turism.
2.
Europaparlamentet stöder FN:s generalsekreterare Ban Ki Moons åsikt att den globala finanskrisen har gett upphov till en utvecklingskris som äventyrar och i vissa fall upphäver de med möda uppnådda framstegen när det gäller fattigdom, svält och mödra- och barnadödlighet, samt i fråga om grundskoleutbildning, jämställdhet och tillgång till rent dricksvatten och acceptabla sanitära förhållanden, vilket riskerar att medföra att millennieutvecklingsmålen, särskilt de som rör hälsa, inte kan uppnås.
3.
4.
Europaparlamentet understryker att många utvecklingsländer anser att samtliga av deras källor till utvecklingsfinansiering påverkats av krisen och att de inte kommer att kunna trygga de med möda uppnådda ekonomiska vinsterna utan omfattande stöd utifrån.
5.
Europaparlamentet uppmanar EU att vidta åtgärder för att utrota problemen med skatteparadis, skatteflykt och olaglig kapitalflykt i utvecklingsländerna och efterfrågar därför en ny bindande internationell överenskommelse som tvingar transnationella företagskoncerner att automatiskt uppge vilka vinster de gjort och vilka skatter de betalat i varje land i syfte att säkerställa insynsvänlighet med avseende på vad de betalar i varje utvecklingsland där de är verksamma.
6.
Europaparlamentet noterar G20-ledarnas erkännande av sitt kollektiva ansvar för att minska de sociala följderna av krisen för att minimera långvariga förluster för den globala potentialen, deras bekräftande av redan ingångna åtaganden om stöd och deras löften om nya resurser, inbegripet 50 000 miljoner USD för att stödja det sociala skyddet, öka handeln och skydda utvecklingen i låginkomstländerna som en del i en betydande ökning av krisstödet i utvecklingsländerna och mer resurser för socialt skydd i de fattigaste länderna.
7.
Europaparlamentet välkomnar G8-ledarnas beslut från toppmötet i Aquila (Italien) i juli 2009 om att ge 20 000 miljoner USD i stöd till utveckling av landsbygden och livsmedelssäkerhet.
8.
Europaparlamentet oroas över att de ekonomiska resurser som utlovats kanske inte kommer att räcka till eller inte riktas mot de fattigaste länderna eller befolkningsgrupperna samt över att resurserna kanske inte kommer att sättas in tillräckligt snabbt och på ett tillräcklig flexibelt sätt för att åstadkomma de förbättringar som krävs i utvecklingsländerna.
9.
Europaparlamentet stöder G8-ledarnas begäran om att genomföra en internationell översyn av strategierna för att uppnå millennieutvecklingsmålen under 2010.
10.
Europaparlamentet noterar de ökade anslagen till Internationella valutafonden och andra internationella finansiella institutioner.
11.
12.
13.
Europaparlamentet beklagar att Världsbanken har lämnats att reagera på krisen i huvudsak genom sina egna befintliga resurser och instrument, trots att ett effektivt svar på krisen skulle kräva en ny och stor resurstilldelning och trots G20-ledarnas löften om att tillhandahålla resurser till socialt skydd för de fattigaste länderna, inbegripet genom investeringar för att trygga livsmedelsförsörjningen på lång sikt och genom frivilliga bilaterala bidrag till Världsbankens sårbarhetsram (Vulnerability Framework), inbegripet krisinstrumentet för infrastruktur (Infrastructure Crisis Facility) och fonden för omedelbara sociala åtgärder (Rapid Social Response Fund).
14.
Europaparlamentet anser att den främsta prioriteringen helt enkelt bör vara att stödja strategier som minskar fattigdomen och som samtidigt innebär att skattebetalarnas pengar utnyttjas på bästa sätt, och som styrs av en insikt om det absoluta människovärdet hos alla människor i utvecklingsländerna.
15.
16.
17.
18.
19.
20.
21.
22.
Europaparlamentet påpekar att man upprepade gånger har begärt att Europeiska utvecklingsfonden ska ingå i gemenskapsbudgeten så att en demokratisk kontroll av fondens användningsområden kan säkerställas.
23.
24.
Europaparlamentet framhåller att omfattningen av det officiella utvecklingsbiståndet inte räcker till för att, med den snabbhet som krävs vid kris i denna storleksordning, möta de avsevärt utökade behoven i utvecklingsländerna som krisen förorsakat, och uppmanar kommissionen och medlemsstaterna att stå fast vid sina internationella åtaganden och fortsätta att bidra till uppnåendet av millennieutvecklingsmålen.
25.
Europaparlamentet betonar att samstämmigheten mellan EU:s handels-, budget-, klimat-, och utvecklingspolitik måste öka.
26.
Europaparlamentet rekommenderar därför att avtalen om ekonomiskt partnerskap används som ett instrument för att möta utvecklingsbehoven genom att AVS-länderna ges en handelsfördel och genom att uppnåendet av millennieutvecklingsmålen främjas, samtidigt som AVS-länderna tillåts lämna känsliga produkter och sektorer, såsom investeringar och tjänster, utanför förhandlingarna.
27.
Europaparlamentet framhåller, mot bakgrund av detta, att avtalen om ekonomiskt partnerskap måste tjäna som instrument för att främja regional integration och lyfta ekonomierna i AVS-länderna, att löftena om finansiering måste uppfyllas.
28.
Europaparlamentet understryker att Europeiska investeringsbanken (EIB) måste engagera sig på ett mer aktivt och öppet sätt som en föregångare när det gäller utvecklingen av nya finansieringsmekanismer.
29.
Europaparlamentet uppmanar med kraft kommissionen att inta en ledande roll för att snabbt stärka dessa mekanismer, inbegripet krediter på mikro- och mesonivå, särskilt för att sårbara grupper som kvinnor och jordbrukare ska kunna erbjudas möjligheter till finansiering.
30.
Europaparlamentet uppmanar EU att se till att lämpliga globala regleringsbestämmelser införs, så att man förhindrar att ytterligare en finanskris inträffar.
31.
Europaparlamentet uppmanar medlemsstaterna att iaktta och uppfylla sina åtaganden om offentligt utvecklingsbistånd.
32.
Europaparlamentet understryker hur viktigt det är ur utvecklingssynpunkt att politiken inom områden som ekonomi, handel, miljö och jordbruk är samstämmig, så att man förhindrar att den globala finansiella och ekonomiska krisen får ännu allvarligare konsekvenser för utvecklingsländerna.
33.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, medlemsstaterna, FN:s organisationer, Internationella valutafonden och Världsbanken samt till Internationella valutafondens och Världsbankens styrelseledamöter från EU:s medlemsstater, och G20-länderna.
P7_TA(2009)0042
Avtal EG/Mauritius om undantag från viseringskravet för kortare vistelser *
A7-0019/2009
Europaparlamentets lagstiftningsresolution av den 20 oktober 2009 om förslaget till rådets beslut om ingående av avtalet mellan Europeiska gemenskapen och Republiken Mauritius om undantag från viseringskravet för kortare vistelser ( KOM(2009)0048 – C7-0015/2009 – 2009/0012(CNS) )
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
–
med beaktande av förslaget till rådets beslut ( KOM(2009)0048 ),
–
–
–
–
med beaktande av betänkandet från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor ( A7-0019/2009 ).
1.
Europaparlamentet godkänner ingåendet av avtalet.
2.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen samt regeringarna och parlamenten i medlemsstaterna och Republiken Mauritius parlamentets ståndpunkt.
P7_TA(2009)0057
De institutionella aspekterna av inrättandet av den europeiska avdelningen för yttre åtgärder
A7-0041/2009
Europaparlamentets resolution av den 22 oktober 2009 om de institutionella aspekterna av inrättandet av den europeiska avdelningen för yttre åtgärder ( 2009/2133(INI) )
Europaparlamentet utfärdar denna resolution
–
–
med beaktande av förklaring nr 15 om artikel 27 i fördraget om Europeiska unionen, en förklaring som är bifogad slutakten från den regeringskonferens som antog Lissabonfördraget,
–
25.
,
–
med beaktande av sin resolution av den 5 september 2000 om den gemensamma EU-diplomatin EGT C 135, 7.5.2001, s.
69.
,
–
med beaktande av sin resolution av den 14 juni 2001 om kommissionens meddelande om utveckling av tjänsten för yttre representation EGT C 53 E, 28.2.2002, s.
390.
,
–
med beaktande av sin resolution av den 26 maj 2005 om de institutionella aspekterna av inrättandet av en europeisk avdelning för yttre åtgärder EUT C 117 E, 18.5.2006, s.
232.
,
–
med beaktande av det seminarium som anordnades av parlamentets utskott för konstitutionella frågor den 10 september 2008,
–
med beaktande av artikel 48 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för konstitutionella frågor och yttrandena från utskottet för utrikesfrågor och utskottet för utveckling ( A7-0041/2009 ), och av följande skäl:
A.
Den europeiska avdelningen för yttre åtgärder (European External Action Service, EEAS) har en mycket viktig roll att spela för att EU:s yttre förbindelser ska bli mer samstämda och effektivare, och för att de ska ges större uppmärksamhet.
B.
EEAS är en konsekvens av tre nyheter som införs genom Lissabonfördraget: Man kommer att välja en ständig ordförande för Europeiska rådet som ska representera unionen utåt på stats- och regeringschefsnivå; Europeiska rådet kommer, efter godkännande av kommissionens ordförande, att utse unionens höga representant för utrikes frågor och säkerhetspolitik, som kommer att vara kommissionens vice ordförande med ansvar för yttre förbindelser (kommissionens vice ordförande/den höga representanten); unionen blir uttryckligen en juridisk person, vilket ska ge unionen fullständig handlingsfrihet i internationella sammanhang.
C.
D.
EU:s roll som global aktör har ökat i betydelse de senaste årtiondena och det behövs ett nytt arbetssätt om EU ska kunna agera gemensamt och möta de globala utmaningarna på ett samstämt, konsekvent och effektivt sätt.
E.
F.
Inrättandet av EEAS måste bidra till att undvika dubbelarbete, ineffektivitet och slöseri med resurser i samband med unionens yttre åtgärder.
G.
EEAS bör ha till uppgift att framhäva EU:s roll som utvecklingsländernas viktigaste partner, och bör härvidlag bygga vidare på de starka förbindelser som EU har etablerat med utvecklingsländerna.
H.
Lissabonfördraget anger uttryckligen att utvecklingssamarbete är ett självständigt politikområde med specifika mål, jämställt med andra uttryck för EU:s utrikespolitik.
I.
I förklaring nr 15 om artikel 27 i fördraget om Europeiska unionen slog medlemsstaternas regeringar fast att kommissionens vice ordförande/den höga representanten, kommissionen och medlemsstaterna skulle inleda det förberedande arbetet med EEAS så snart Lissabonfördraget undertecknats.
J.
K.
L.
Så snart Lissabonfördraget har trätt i kraft kommer rådet, på förslag från kommissionens vice ordförande/den höga representanten och efter att ha hört parlamentet och ha erhållit kommissionens godkännande, att fastställa EEAS organisation och verksamhet.
M.
Ett antal principfrågor som rör utformningen av EEAS bör lösas i tillräckligt god tid för att avdelningen ska kunna inleda sitt arbete så snart som möjligt efter att kommissionens vice ordförande/den höga representanten har utsetts.
N.
Eftersom parlamentet kommer att höras om inrättandet av den europeiska avdelningen för yttre åtgärder, och med tanke på budgetkonsekvenserna, är en konkret dialog med parlamentet i ett tidigt skede av avgörande betydelse för att EEAS ska kunna inleda sin verksamhet på ett effektivt sätt och tillförsäkras nödvändiga ekonomiska resurser.
1.
2.
3.
Europaparlamentet uppmanar kommissionen, rådet, medlemsstaterna och den tillträdande kommissionens vice ordförande/höga representant att göra ett tydligt åtagande om att, tillsammans med parlamentet, nå en omfattande, ambitiös och gemensam plan för inrättandet av EEAS.
4.
5.
Europaparlamentet påminner om att EEAS måste garantera att Europeiska unionens stadga om de grundläggande rättigheterna tillämpas fullt ut i fråga om alla aspekter av EU:s yttre åtgärder i enlighet med Lissabonfördragets anda och syfte.
6.
Europaparlamentet bekräftar följande principer och uppmanar kommissionen att, då den i fortsättningen utarbetar sina förslag, insistera på att dessa principer följs i enlighet med Lissabonfördragets anda och syfte och med beaktande av konventets överläggningar:
a)
b)
c)
d)
e)
f)
EEAS måste se till att Europaparlamentet har kontaktpersoner i EU:s delegationer som ansvarar för samarbetet med parlamentet (till exempel genom att upprätthålla parlamentets kontakter i tredjeländer).
7.
a)
b)
Kommissionens vice ordförande/den höga representanten bör vara EEAS tillsättningsmyndighet, detta för att säkerställa dels att instruktionerna för de olika tjänsterna utformas i enlighet med de befogenheter som fördraget föreskriver, dels att kommissionens vice ordförande/den höga representanten är den som beslutar om anställning, befordran och avgång från tjänst.
c)
d)
I analogi med tidigare bestämmelser Till exempel artikel 6 i kommissionens beslut 1999/352/EG, EKGS, Euratom av den 28 april 1999 om inrättande av en europeisk byrå för bedrägeribekämpning (OLAF) (EGT L 136, 31.5.1999, s.
20).
bör ansvaret för att sköta tillsättningsmyndighetens administrativa uppgifter i samband med anställning av EEAS personal och för att genomföra de beslut som kommissionens vice ordförande/den höga representanten fattar i fråga om anställning, befordran, förlängning eller avgång från tjänst tillfalla ett lämpligt generaldirektorat inom kommissionen.
e)
Utstationering av personal till EEAS från medlemsstaternas nationella diplomattjänster bör ses som en integrerad del av karriärstigen inom dessa tjänster.
f)
g)
I och med att EEAS inrättas måste Interinstitutionella avtalet om budgetdisciplin och sund ekonomisk förvaltning Interinstitutionellt avtal mellan Europaparlamentet, rådet och kommissionen av den 17 maj 2006 om budgetdisciplin och sund ekonomisk förvaltning (EUT C 139, 14.6.2006, s.
1).
justeras, i enlighet med punkt 4 och avsnitt II, del G i avtalet.
1).
) bör respekteras fullt ut.
h)
Vid eventuell frånvaro bör kommissionens vice ordförande/den höga representanten från fall till fall och med hänsyn tagen till de uppgifter som är aktuella för tillfället besluta vem som ska ersätta honom eller henne.
8.
9.
Europaparlamentet anser att
a)
EEAS bör ledas av en generaldirektör som är ansvarig inför kommissionens vice ordförande/den höga representanten, och denna generaldirektör bör kunna företräda kommissionens vice ordförande/den höga representanten i vissa fall,
b)
EEAS bör delas in i ett antal direktorat som ska ansvara för var sin geostrategiskt viktiga del av unionens yttre förbindelser och med ytterligare direktorat som ansvarar för frågor som rör säkerhet och försvarspolitik, civil krishantering, multilaterala och horisontella frågor, bland annat mänskliga rättigheter och administrativa frågor,
c)
EEAS bör strukturera samarbetet mellan landsenheter i Bryssel och unionens delegationer (ambassader) i tredjeländer i frågor som rör de olika direktoraten.
d)
varken rådet eller Europeiska rådet bör ha mer än en avdelning för yttre åtgärder.
11.
Europaparlamentet anser att beslutet som ska fastställa EEAS organisation och verksamhet också bör slå fast att unionens ambassader i tredjeländer vid behov och utifrån tillgängliga resurser måste ge alla som tillhör någon EU-institution logistiskt och administrativt stöd.
12.
122).
med parlamentet, särskilt beträffande tillgång till känslig information och andra frågor som är relevanta för ett smidigt interinstitutionellt samarbete.
13.
14.
15.
Europaparlamentet uppmanar kommissionens vice ordförande/den höga representanten att lägga fram ett förslag till beslut om EEAS organisation och arbetssätt och därvid ta hänsyn till riktlinjerna i denna resolution.
Parlamentet avser att anta en detaljerad ståndpunkt om det förslaget i enlighet med artikel 27.3 i fördraget om Europeiska unionen enligt Lissabonfördragets formulering, och att i samband med budgetförfarandet undersöka de finansiella aspekterna.
Parlamentet rekommenderar emellertid att man når en politisk överenskommelse med parlamentet i samtliga frågor i ett tidigt skede för att undvika att man förlorar värdefull tid på politiska debatter om hur EEAS ska utformas efter att Lissabonfördraget trätt i kraft.
16.
Europaparlamentet uppmanar kommissionen att samtycka till det förslag som kommissionens vice ordförande/den höga representanten lägger fram endast om det till övervägande del följer riktlinjerna i denna resolution eller om man enhälligt kommer fram till en annan kompromisslösning genom interinstitutionella kontakter där parlamentet deltagit.
17.
Europaparlamentet är fast beslutet att be den tillträdande kommissionens vice ordförande att ta ställning i de frågor som tas upp i denna resolution då han eller hon sammanträder med det behöriga utskottet för utfrågningen i samband med förfarandet för utnämningen av den nya kommissionen.
18.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet och kommissionen.
P7_TA(2009)0076
Ändring av bilagorna II och III till Ospar-konventionen *
A7-0051/2009
Europaparlamentets lagstiftningsresolution av den 24 november 2009 om förslaget till rådets beslut om godkännande, på Europeiska gemenskapens vägnar, av ändringarna av bilagorna II och III till konventionen för skydd av den marina miljön i Nordostatlanten (Ospar-konventionen) gällande lagring av koldioxidströmmar i geologiska formationer ( KOM(2009)0236 – C7-0019/2009 – 2009/0071(CNS) )
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
–
med beaktande av förslaget till rådets beslut ( KOM(2009)0236 ),
–
–
–
–
med beaktande av betänkandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A7-0051/2009 ).
1.
Europaparlamentet godkänner förslaget till rådets beslut med de ändringar som gjorts i bilagorna II och III till konventionen.
2.
Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen samt regeringarna och parlamenten i Belgien, Danmark, Finland, Frankrike, Irland, Island, Luxemburg, Nederländerna, Norge, Portugal, Schweiz, Spanien, Storbritannien, Sverige och Tyskland parlamentets ståndpunkt.
Kommissionens förslag
Ändring
Ändring 1
Förslag till rådets beslut
Skäl 4a (nytt)
(4a)
Gemenskapen har nyligen antagit Europaparlamentets och rådets direktiv 2009/31/EG av den 23 april 2009 om geologisk lagring av koldioxid
1
__________
1
EUT L 140, 5.6.2009, s.
114.
Ändring 2
Förslag till rådets beslut
Skäl 4b (nytt)
(4b)
Delad behörighet mellan gemenskapen och medlemsstaterna, tillsammans med principen om enhetlighet vid företrädandet av gemenskapen på det internationella planet, talar för att gemenskapen och de av medlemsstaterna som är fördragsslutande parter i konventionen gemensamt ska deponera sina instrument för godkännande av ändringarna.
Ändring 3
Förslag till rådets beslut
De medlemsstater som är fördragsslutande parter i konventionen ska anstränga sig att vidta nödvändiga åtgärder för att deponera sina handlingar för ratifikation eller godkännande samtidigt med Europeiska gemenskapens och övriga medlemsstaters och i möjligaste mån inte senare än den 1 juni 2010.
P7_TA(2009)0104
Laos och Vietnam
B7-0157 , 0177 , 0178 och 0179/2009
Europaparlamentets resolution av den 26 november 2009 om situationen i Laos och Vietnam
Europaparlamentet utfärdar denna resolution
–
med beaktande av det femtonde toppmötet för Sydostasiatiska nationers förbund (Asean) den 23–25 oktober 2009,
–
med beaktande av att Aseans mellanstatliga kommission för mänskliga rättigheter invigdes den 23 oktober 2009,
–
med beaktande av EU:s årsrapport om de mänskliga rättigheterna 2008,
–
med beaktande av de pågående förhandlingarna om det nya partnerskaps- och samarbetsavtalet mellan EU och Vietnam och de samtal om mänskliga rättigheter som EU och Vietnams regering för med varandra två gånger om året,
–
med beaktande av sina tidigare resolutioner om Laos, framför allt resolutionen av den 15 november 2001 om de godtyckliga arresteringarna och den politiska situationen i Laos EUT C 140 E, 13.6.2002, s.
577.
och resolutionen av den 1 december 2005 om situationen för de mänskliga rättigheterna i Kambodja, Laos och Vietnam EUT C 285 E, 22.11.2006, s.
129.
,
–
med beaktande av samarbetsavtalet av den 1 december 1997 mellan Europeiska unionen och Demokratiska folkrepubliken Laos, som baseras på respekt för demokratiska principer och grundläggande mänskliga rättigheter sådana de fastställs i FN:s allmänna förklaring om de mänskliga rättigheterna,
–
Vietnam
A.
Den vietnamesiska regeringen har vägrat att efterleva många rekommendationer som utfärdades i samband med den allmänna återkommande utvärderingen som FN:s råd för mänskliga rättigheter genomförde mellan maj och september 2009, och som var avsedda att förbättra landets resultat på området för mänskliga rättigheter.
B.
I Vietnam sitter i dagsläget hundratals människor fängslade på grund av sin religiösa eller politiska övertygelse, till exempel montagnard-kristna, en katolsk präst, en mennonitisk pastor, medlemmar av Cao Dai-religionen och Hoa Hao-buddister.
C.
D.
Många anser att attacken mot klostret kan kopplas till det tiopunktsförslag om religiösa reformer som Thich Nhat Hanh lade fram för Vietnams president Nguyen Minh Triet 2007.
E.
F.
G.
H.
Flera samvetsfångar, till exempel Nguyen Van Ly, Le Thi Cong Nhan och Nguyen Binh Thanh, som alla dömts för att ha spridit "propaganda mot regeringen i Socialistiska republiken Vietnam", har nekats korrekt läkarvård i fängelset fastän deras hälsotillstånd kräver att de omedelbart läggs in på sjukhus.
I.
Eftersom det inte finns några egentliga människorättsorganisationer, tar kyrkliga ledare ofta på sig rollen att försvara de mänskliga rättigheterna och kämpa för mer tolerans och demokratiska principer.
J.
Laos
K.
Den 25 september 2009 ratificerade Demokratiska folkrepubliken Laos den internationella konventionen om medborgerliga och politiska rättigheter, i vilken t.ex. människors rätt till trosfrihet, föreningsfrihet, yttrandefrihet, tryckfrihet, rätt att demonstrera och politiska rättigheter garanteras.
L.
Nästan en månad efter den tionde årsdagen av "studentrörelsen" 26 oktober 1999 som startades av studenter och lärare i Vientiane, hålls fortfarande de främsta ledarna för rörelsen, Thongpaseuth Keuakoun, Seng-Aloun Phengphanh, Bouavanh Chanmanivong och Kèochay, i hemlig fångenskap, och enligt rapporter har Khamphouvieng Sisa-At avlidit i fängelse under oklara omständigheter.
M.
N.
O.
P.
Vietnam
1.
2.
3.
Europaparlamentet ber rådet och kommissionen att inom ramen för de pågående förhandlingarna om det nya partnerskaps- och samarbetsavtalet med Vietnam inkludera en bindande och otvetydig klausul om mänskliga rättigheter och demokrati, tillsammans med en mekanism som möjliggör dess tillämpning, för att få ett slut på de systematiska kränkningarna av demokratiska och mänskliga rättigheter.
4.
Europaparlamentet begär att all förföljelse och alla trakasserier ska upphöra, och att nunnor och munkar ska tillåtas att utöva buddism i enlighet med traditionerna inom den buddistiska Thich Nhat Hanh-gemenskapen i Bat Nha och på andra platser.
5.
Europaparlamentet kräver Thich Quang Dos ovillkorliga frigivning och återupprättande av Vietnams enade buddistkyrka och dess dignitärer.
6.
Europaparlamentet uppmanar regeringen att inrätta en oberoende nationell människorättskommission som ska samla in och utreda alla anklagelser om tortyr och andra former av maktmissbruk av tjänstemän, inklusive anställda inom säkerhetspolisen, och att inleda förfaranden för att avskaffa dödsstraffet.
7.
Europaparlamentet uppmanar Vietnams regering, med tanke på landets roll som medlem i FN:s säkerhetsråd, att utfärda stående inbjudningar till FN:s särskilda rapportörer, särskilt till dem som arbetar med yttrandefrihet, religionsfrihet, tortyr, människorättsaktivister och våld mot kvinnor och till FN:s arbetsgrupp för godtyckliga frihetsberövanden.
Laos
8.
Europaparlamentet välkomnar att Laos regering har ratificerat den internationella konventionen om medborgerliga och politiska rättigheter och uppmanar de laotiska myndigheterna att fullständigt respektera innehållet i konventionen, att utan dröjsmål harmonisera Laos lagstiftning med konventionens bestämmelser och att tillämpa bestämmelserna enligt internationella normer, särskilt när det gäller yttrande-, förenings- och trosfrihet.
9.
Europaparlamentet upprepar sin begäran om att ledarna för studentrörelsen "26 oktober 1999" och alla samvetsfångar som sitter fängslade i Laos ska släppas fria, och parlamentet ger sin EU-delegation i Vientiane ansvaret att följa upp ärendet.
10.
Europaparlamentet uppmanar Laos myndigheter att ovillkorligen släppa alla de människor som arresterades under försöket till fredlig demonstration den 2 november 2009.
11.
12.
Europaparlamentet uppmanar kommissionen att noggrant övervaka situationen för hmong lao-gruppen och regeringens program för etniska minoriteter.
13.
Europaparlamentet upprepar sin begäran till Laos myndigheter att utforma och så snabbt som möjligt genomföra alla de reformer som krävs för att införa demokrati i landet, garantera den politiska oppositionens rätt att yttra sig inom fredliga ramar och att se till att internationellt övervakade flerpartival kan genomföras snart, så att landet kan nå nationell försoning.
Allmänt
14.
15.
Europaparlamentet uppmanar rådet och kommissionen att genomföra en noggrann utvärdering av hur politiken för demokrati och mänskliga rättigheter tillämpats i Laos och Vietnam sedan partnerskaps- och samarbetsavtalen undertecknades, och att rapportera till parlamentet.
o
o o
16.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, medlemsstaternas regeringar och parlament, Laos och Vietnams regeringar och parlament, Aseans sekretariat, FN:s högkommissarie för mänskliga rättigheter och FN:s generalsekreterare.
P7_TA(2009)0107
Utnyttjande av Europeiska fonden för justering för globaliseringseffekter Sverige/Volvo - Österrike/Steiermark - Nederländerna/Heijmans
A7-0079/2009
Europaparlamentets resolution av den 16 december 2009 om förslaget till Europaparlamentets och rådets beslut om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning ( KOM(2009)0602 – C7-0254/2009 – 2009/2183(BUD) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2009)0602 – C7-0254/2009 ),
–
med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning EUT C 139, 14.6.2006, s.
1.
(IIA av den 17 maj 2006), särskilt punkt 28,
–
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1927/2006 av den 20 december 2006 om upprättande av Europeiska fonden för justering för globaliseringseffekter EUT L 406, 30.12.2006, s.
1.
,
–
med beaktande av betänkandet från budgetutskottet och yttrandet från utskottet för sysselsättning och sociala frågor ( A7-0079/2009 ), och av följande skäl:
A.
Europeiska unionen har inrättat lagstiftningsinstrument och budgetinstrument för att kunna ge kompletterande stöd till arbetstagare som blivit arbetslösa till följd av genomgripande strukturförändringar inom världshandeln och för att underlätta deras återinträde på arbetsmarknaden.
B.
Unionens ekonomiska stöd till arbetstagare som har blivit uppsagda bör vara dynamiskt och ges så snabbt och effektivt som möjligt, i enlighet med Europaparlamentets, rådets och kommissionens gemensamma uttalande, som antogs vid medlingsmötet den 17 juli 2008, och med vederbörlig hänsyn till IIA av den 17 maj 2006 när det gäller antagandet av beslut rörande fondens utnyttjande.
C.
Sverige, Österrike och Nederländerna har ansökt om stöd med anledning av uppsägningarna inom bilsektorn i Sverige EGF/2009/007 SE/Volvo.
och Österrike EGF/2009/009 AT/Steiermark.
och inom byggsektorn i ett företag, Heijmans N.V., i Nederländerna EGF/2009/011 NL/Heijmans N.V.
.
D.
Ansökningarna uppfyller kriterierna för berättigande till stöd enligt förordningen om upprättande av Europeiska fonden för justering för globaliseringseffekter.
1.
Europaparlamentet uppmanar de berörda institutionerna att vidta de åtgärder som krävs för att Europeiska fonden för justering för globaliseringseffekter snarast ska kunna tas i anspråk.
2.
Europaparlamentet erinrar om institutionernas åtagande att säkerställa ett smidigt och snabbt förfarande för antagandet av beslut om utnyttjande av fonden, i syfte att tillhandahålla ett tidsbegränsat och individuellt stöd av engångskaraktär för att hjälpa arbetstagare som har blivit uppsagda till följd av globaliseringen.
3.
4.
5.
6.
Europaparlamentet påminner kommissionen om att den i samband med utnyttjandet av fonden inte systematiskt ska överföra betalningsbemyndiganden från Europeiska socialfonden, eftersom Europeiska fonden för justering för globaliseringseffekter inrättades som ett enskilt och specifikt instrument med egna mål och tidsfrister.
7.
Europaparlamentet erinrar om att en utvärdering av hur Europeiska fonden för justering för globaliseringseffekter fungerar och vilket mervärde den skapar bör göras inom ramen för den allmänna bedömningen av programmen och andra instrument som skapats genom IIA av den 17 maj 2006, i samband med budgetöversynen av den fleråriga budgetramen 2007–2013.
8.
Europaparlamentet godkänner det beslut som bifogas denna resolution.
9.
Europaparlamentet uppmanar kommissionen att hädanefter, för varje enskild ansökan som inkommer, lägga fram ett separat förslag om att godkänna att fonden utnyttjas.
10.
Europaparlamentet uppdrar åt talmannen att underteckna detta beslut tillsammans med rådets ordförande och att se till att beslutet offentliggörs i Europeiska unionens officiella tidning.
11.
Europaparlamentet uppdrar åt talmannen att översända denna resolution, inklusive bilagan, till rådet och kommissionen.
BILAGA
EUROPAPARLAMENTETS OCH RÅDETS BESLUT
om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av fördraget om upprättandet av Europeiska gemenskapen och fördraget om Europeiska unionens funktionssätt,
med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning EUT C 139, 14.6.2006, s.
1.
, särskilt punkt 28,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1927/2006 av den 20 december 2006 om upprättande av Europeiska fonden för justering för globaliseringseffekter EUT L 406, 30.12.2006, s.
1.
av följande skäl:
(1)
Europeiska fonden för justering för globaliseringseffekter upprättades för att ge kompletterande stöd till arbetstagare som drabbats av konsekvenserna av större strukturella förändringar i världshandelsmönstren, för att hjälpa dem att återintegrera sig på arbetsmarknaden.
(2)
Tillämpningsområdet för fonden har utvidgats för ansökningar om stöd från fonden som inges från och med den 1 maj 2009 och omfattar nu stöd till arbetstagare som har blivit uppsagda som en direkt följd av den globala finansiella och ekonomiska krisen.
(3)
Det interinstitutionella avtalet av den 17 maj 2006 gör det möjligt att använda medel från fonden upp till ett högsta belopp på 500 miljoner EUR per år.
(4)
Sverige ingav den 5 juni 2009 en ansökan om stöd från fonden på grund av uppsägningar i bilsektorn.
(5)
Österrike ingav den 9 juli 2009 en ansökan om stöd från fonden på grund av uppsägningar i bilsektorn.
(6)
Nederländerna ingav den 4 augusti 2009 en ansökan om stöd från fonden på grund av uppsägningar i byggsektorn.
(7)
Fonden bör alltså tas i anspråk för att tillhandahålla ekonomiskt stöd med anledning av de ansökningar som ingivits av Sverige, Österrike och Nederländerna.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Europeiska fonden för justering för globaliseringseffekter ska tas i anspråk för att tillhandahålla beloppet 15 931 423 EUR i åtagandebemyndiganden och betalningsbemyndiganden i Europeiska unionens allmänna budget för budgetåret 2009.
Artikel 2
Utfärdat i Strasbourg den
På Europaparlamentets vägnar
På rådets vägnar
P7_TA(2010)0012
ERUF: Stödberättigande åtgärder avseende bostäder för marginaliserade grupper ***I
A7-0048/2009
Europaparlamentets lagstiftningsresolution av den 10 februari 2010 om förslaget till Europaparlamentets och rådets förordning (EU) nr .../2010 om ändring av förordning (EG) nr 1080/2006 om Europeiska regionala utvecklingsfonden vad gäller stödberättigade bostadsinsatser till förmån för marginaliserade befolkningsgrupper ( KOM(2009)0382 – C7-0095/2009 – 2009/0105(COD) )
(Ordinarie lagstiftningsförfarandet: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2009)0382 ),
–
–
med beaktande av meddelandet från kommissionen till Europaparlamentet och rådet "Konsekvenser av Lissabonfördragets ikraftträdande för pågående interinstitutionella beslutsförfaranden" ( KOM(2009)0665 ),
–
–
med beaktande av artikel 55 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för regional utveckling ( A7-0048/2009 ).
1.
Europaparlamentet antar nedanstående ståndpunkt vid första behandlingen.
2.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om kommissionen har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
3.
Europaparlamentet uppdrar åt talmannen att översända parlamentets ståndpunkt till rådet, kommissionen och de nationella parlamenten.
P7_TC1-COD(2009)0105
Europaparlamentets ståndpunkt fastställd vid första behandlingen den 10 februari 2010 inför antagandet av Europaparlamentets och rådets förordning (EU) nr .../2010 om ändring av förordning (EG) nr 1080/2006 om Europeiska regionala utvecklingsfonden vad gäller stödberättigande för bostadsinsatser till förmån för marginaliserade befolkningsgrupper
(Eftersom det nåddes en överenskommelse mellan parlamentet och rådet, motsvarar parlamentets ståndpunkt den slutliga rättsakten, förordning (EU) nr 437/2010.)
P7_TA(2010)0022
De viktigaste målen inför partskonferensen för Cites-konventionen
B7-0069/2010
Europaparlamentets resolution av den 10 februari 2010 om EU:s strategiska mål inför det femtonde mötet i partskonferensen för konventionen om internationell handel med utrotningshotade arter av vilda djur och växter (Cites), avsett att hållas i Doha (Qatar) den 13–25 mars 2010
Europaparlamentet utfärdar denna resolution
–
med beaktande av det kommande femtonde mötet i partskonferensen för konventionen om internationell handel med utrotningshotade arter av vilda djur och växter (Cites), avsett att hållas den 13–25 mars 2010 i Doha, Qatar,
–
med beaktande av frågorna av den 2 december 2009 till kommissionen och rådet om de viktigaste målen inför konferensen för parterna till Cites i Doha den 13–25 mars 2010 ( O-0145/2009 – B7-0003/2010 , O-0146/2009 – B7-0004/2010 ),
–
A.
Cites är det mest omfattande naturvårdsavtal som finns för att förhindra att vilda djur och växter överexploateras på grund av internationell handel, med 175 parter till konventionen, däribland EU:s 27 medlemsstater.
B.
De huvudsakliga orsakerna till utarmningen av jordens biologiska mångfald är människors användning av naturresurser, förstörelse av livsmiljöer, klimatförändringar, överexploatering av vilda arter och olaglig handel med vilda djur och växter.
C.
I vetenskapliga rapporter förutsägs det att klimatförändringen kommer att driva på förlusten av biologisk mångfald och förvärra situationen för de utrotningshotade arterna.
D.
E.
Allmänhetens medvetenhet i konsumtionsländerna har varit och fortsätter att vara avgörande för kontrollen av tjuvskyttet och den illegala internationella handeln med utrotningshotade arter av vilda djur och växter.
F.
Olaglig skogsavverkning kan innebära handel med växtarter upptagna i Cites-förteckningarna, och i förslaget till Europaparlamentets och rådets förordning om fastställande av skyldigheter för aktörer när det gäller utsläppande på marknaden av trä och träprodukter bör man se till att effektiva åtgärder vidtas för att lösa problemet med olaglig skogsavverkning.
G.
Den olagliga handeln försvårar allvarligt de världsomfattande strävandena efter hållbarhet inom utveckling och miljö, undergräver goda styrelseformer och underlättar spridning av smittsamma sjukdomar.
H.
I.
Furstendömet Monaco har lagt fram ett förslag om att införa blåfenad tonfisk i bilaga I till Cites-konventionen för att tillfälligt stoppa den internationella kommersiella handeln med arten.
J.
ICCATS (Internationella kommissionen för bevarande av tonfisk i Atlanten) vetenskapliga kommitté uppskattade vid sitt sammanträde den 21–23 oktober 2009 att det nuvarande lekande beståndets biomassa är lägre än 15 procent av vad den var innan fisket började, och bekräftade därmed att blåfenad tonfisk uppfyller detta kriterium för att föras in i bilaga I till Cites-konventionen.
K.
Sillhaj (håbrand) och pigghaj är mycket känsliga för överfiske och behöver lång tid för att återhämta sig på grund av sina biologiska egenskaper (långsam tillväxt, sen könsmognad, låg reproduktionskapacitet, lång livslängd och lång tid mellan generationerna).
L.
Dessa arter måste föras in i bilaga II till Cites-förordningen för att garantera att framtida internationell handel tryggas genom ett fiske som förvaltas hållbart och registreras korrekt, och som inte är skadligt för bevarandestatusen för det vilda bestånd som fisket utnyttjar.
M.
I konferensresolution 9.24 till Cites-konventionen anges att arter som är eller kan komma att bli föremål för handel, och som visar en markant nedgång i de vilda bestånden som härrör från eller kan beräknas utifrån att livsmiljöns areal eller kvalitet har minskat, ska föras in i bilaga I till Cites-konventionen.
N.
O.
Cites-parterna enades under det fjortonde mötet i partskonferensen (CoP 14) om att det inte skulle läggas fram några ytterligare förslag om handel med elfenben under en tidsperiod på minst nio år.
P.
Q.
R.
Vid CoP 14 antogs beslut 14.69, i vilket samtliga Cites-parter uppmanas att se till att asiatiska stora kattdjur föds upp i fångenskap endast om detta tjänar naturvårdsändamål, och i beslutet anges att tigrar inte bör avlas för att man ska kunna handla med delar av dem eller produkter av dessa.
S.
I de nyligen antagna rekommendationerna från Katmandu betonades vikten av att de internationella brottsbekämpande organen, såsom Interpol, Världstullorganisationen (WCO), FN:s drog- och brottsbekämpningsbyrå (UNODC) och Cites, ökar sin delaktighet i kampen mot naturvårdsbrott, och man begärde att dessa organs avdelningar för miljöbrott ska förstärkas i detta syfte.
T.
1.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att tillämpa försiktighetsprincipen som ledande princip i fråga om samtliga beslut om arbetsdokument och förslag till införande i listor och att även ta hänsyn till principen om att användaren betalar samt till ett ekosystembaserat synsätt och hävdvunna naturvårdsprinciper.
2.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att se till att inga beslut som syftar till att förstärka samordningen mellan Cites och andra konventioner om biologisk mångfald undergräver Cites ställning som internationellt naturvårdsavtal eller dess rigorösa naturvårdsåtgärder.
3.
Europaparlamentet motsätter sig kraftfullt slutna omröstningar och är besviket över att Cites stående kommitté inte lagt fram förslag för att förhindra möjligheten att använda slutna omröstningar i Cites beslutsprocesser.
Blåfenad tonfisk
4.
–
Möjlighet att ändra kommissionens förordning (EG) nr 865/2006 om tillämpningsföreskrifter för rådets förordning (EG) nr 338/97 om skyddet av arter av vilda djur och växter genom kontroll av handeln med dem, i syfte att införa ett allmänt undantag för handeln inom gemenskapen för att säkra ett varaktigt kustnära icke-industriellt fiske.
–
Ett EU-finansierat stöd till de sjömän och skeppsredare som berörs av detta beslut.
–
Förstärkta kontroller och sanktioner i kampen mot illegalt, icke rapporterat och oreglerat fiske (IUU).
5.
Europaparlamentet uppmanar kommissionen att ge ekonomisk ersättning till fiskesektorn, som kan komma att påverkas om blåfenad tonfisk införs i bilaga I till Cites-konventionen, för att slå vakt om sektorns ekonomiska bärkraft.
Hajar
6.
Europaparlamentet välkomnar varmt det förslag som lagts fram av Sverige på medlemsstaternas vägnar om att de två hajarterna sillhaj eller håbrand
(Lamna nasus)
och pigghaj
(Squalus acanthias)
7.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att stödja Förenta staternas förslag att ta upp de fem hajarterna flerhornig hammarhaj
(Sphyrna lewini)
, stor hammarhaj
(Sphyrna mokarran)
, hammarhaj
(Sphyrna zygaena)
, högfenad haj
(Carcharhinus plumbeus)
och mörkhaj
(Carcharhinus obscurus)
i bilaga II till Cites-konventionen.
8.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att stödja Förenta staternas förslag att ta upp årfenshaj
(Carcharhinus longimanus)
i bilaga II till Cites-konventionen.
Isbjörn
9.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att stödja Förenta staternas förslag att överföra isbjörn
(Ursus maritimus)
från konventionens bilaga II till dess bilaga I.
Elefanter och elfenben
10.
Europaparlamentet uppmanar med kraft kommissionen och medlemsstaterna att förkasta följande:
-
Förslaget från Tanzania och Zambia om att afrikansk elefant
(Loxondonta africana)
ska överföras från konventionens bilaga I till dess bilaga II i syfte att tillåta handel.
-
Samtliga förslag om att överföra afrikansk elefant från konventionens bilaga I till dess bilaga II, åtminstone till den tidpunkt då en verklig bedömning kan göras av konsekvenserna av engångsförsäljningen i november 2008 från Botswana, Namibia, Sydafrika och Zimbabwe, eftersom alltmer pekar på att den olagliga och organiserade handeln över hela Afrika ökar.
11.
Europaparlamentet uppmanar med kraft kommissionen och medlemsstaterna att stödja förslaget från Kenya, Ghana, Liberia, Mali, Sierra Leone, Togo, Kongo och Rwanda om att införa en not gällande afrikansk elefant som förhindrar alla framtida förslag om handel med elfenben eller om att föra över elefantpopulationer från bilaga I till Cites-konventionen till bilaga II, under minst 20 år efter engångsförsäljningen i november 2008.
12.
Europaparlamentet uppmanar de parter till Cites-konventionen som gynnades av engångsförsäljningen av elfenben från statsägda lager att ge ekonomiska bidrag till fonden för afrikanska elefanter för att stärka initiativ mot tjuvskytte och efterlevnaden av reglerna.
13.
Europaparlamentet uppmuntrar till ett bredare och öppnare samråd med samtliga stater som omfattas av elefanternas utbredningsområde för att överväga åtgärder gällande överförande av afrikansk elefant från konventionens bilaga I till dess bilaga II och efterföljande engångsförsäljningar.
14.
Europaparlamentet uppmuntrar till att kraftfullare metoder utarbetas för att övervaka den olagliga handeln med elfenben, och anser att ett brett spektrum av aktörer bör göras delaktiga i utarbetandet.
Tigrar och asiatiska stora kattdjur
15.
Europaparlamentet välkomnar EU:s förslag om att stärka konferensresolution 12.5 till Cites-konventionen om asiatiska stora kattdjur.
16.
17.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att stödja ansträngningarna att minska efterfrågan på de asiatiska stora kattdjurens delar eller produkter av dessa hos sin egen befolkning och i andra länder.
Övriga arter
18.
Europaparlamentet uppmanar med eftertryck kommissionen och medlemsstaterna att ställa sig bakom följande förslag:
–
Införande av
Corallium spp.
och
Paracorallium spp.
i bilaga II till Cites-konventionen, enligt det förslag som lagts fram av Sverige på medlemsstaternas vägnar.
–
Införande av
Bulnesia sarmientoi
i bilaga II till Cites-konventionen, i överensstämmelse med förslaget från Argentina.
–
Överförande av afrikansk dabbagam
(Uromastyx ornata)
från konventionens bilaga II till dess bilaga II, i överensstämmelse med förslaget från Israel.
–
Införande av iransk bergssalamander (
Neurergus kaiseri
) i bilaga I till Cites-konventionen, i överensstämmelse med förslaget från Iran.
–
Införande av leguanarterna
och
C. melanosterna
i bilaga II till Cites-konventionen, i överensstämmelse med förslaget från Honduras.
–
Införande av rödögda trädgrodor (
Agalychnis spp.
) i bilaga II till Cites-konventionen, i överensstämmelse med förslaget från Honduras och Mexico.
–
Införande av leguanarten
Ctenosaura palearis
i bilaga II till Cites-konventionen, i överensstämmelse med förslaget från Guatemala.
–
Införande av
Aniba rosaeodora
i bilaga II till Cites-konventionen, i överensstämmelse med förslaget från Brasilien.
–
Införande av
Dynastes satanas
i bilaga II till Cites-konventionen, i överensstämmelse med förslaget från Madagaskar.
–
Införande av fröna från
Beccariophoenix madagascariensis
i bilaga II till Cites-konventionen, i överensstämmelse med förslaget från Madagaskar.
–
Införande av fröna från
Dypsis decaryi
i bilaga II till Cites-konventionen, i överensstämmelse med förslaget från Madagaskar.
19.
Europaparlamentet välkomnar och stöder förslaget från Madagaskar om växter och arter av växtfröer som ska införas i förteckningen.
20.
Europaparlamentet uppmanar med eftertryck kommissionen och medlemsstaterna att avvisa följande förslag:
–
Strykningen av rödlo (
Lynx rufus
) från bilaga II till Cites-konventionen.
–
Överföringen av Moreletkrokodil (
Crocodylus moreletti
) från Cites-konventionens bilaga I till dess bilaga II (förslag från Belize och Mexiko).
–
Överföringen av de egyptiska populationerna av Nilkrokodil (
Crocodylus niloticus
) från Cites-konventionens bilaga I till dess bilaga II (förslag från Egypten).
21.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att avvisa Förenta staternas och Mexikos förslag om att stryka
Euphorbia misera
från bilaga II till Cites-konventionen.
22.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att förstärka det internationella samarbetet vid genomförandet av Cites-konventionen.
23.
24.
25.
26.
27.
Saiga tatarica tatarica
) och de tillhörande besluten i saigaantilopens utbredningsstater.
Parlamentet föreslår också att Cites-parterna ska uppmuntra de branscher som konsumerar horn från saigaantilopen att bidra till bevarandeåtgärder på plats för att återställa vilda populationer.
28.
29.
Europaparlamentet uppmanar med eftertryck kommissionen och medlemsstaterna att stödja insatserna inom Cites för att bekämpa illegalt, oreglerat och orapporterat fiske av napoleonfisk (
Cheilinus undulates
).
30.
o
o........o
31.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, parterna till Cites och Cites-sekretariatet.
P7_TA(2010)0104
Ansvarsfrihet för 2008: Europeiska kemikaliemyndigheten
A7-0089/2010
1.
Europaparlamentets beslut av den 5 maj 2010 om ansvarsfrihet för genomförandet av budgeten för Europeiska kemikaliemyndigheten för budgetåret 2008 ( C7-0202/2009 – 2009/2131(DEC) )
Europaparlamentet fattar detta beslut
–
med beaktande av den slutliga årsredovisningen för Europeiska kemikaliemyndigheten för budgetåret 2008,
–
med beaktande av revisionsrättens rapport om årsredovisningen för Europeiska kemikaliemyndigheten för budgetåret 2008, samt myndighetens svar EUT C 304, 15.12.2009, s.
33.
,
–
med beaktande av rådets rekommendation av den 16 februari 2010 (5827/2010 – C7-0061/2010 ),
–
med beaktande av artikel 276 i EG-fördraget och artikel 319 i fördraget om Europeiska unionens funktionssätt,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
, särskilt artikel 185,
–
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 EUT L 396, 30.12.2006, s.
1.
, särskilt artikel 97,
–
med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002 EGT L 357, 31.12.2002, s.
72.
, särskilt artikel 94,
–
med beaktande av artikel 77 i och bilaga VI till arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A7-0089/2010 ).
1.
Europaparlamentet beviljar ansvarsfrihet för den verkställande direktören för Europeiska kemikaliemyndigheten avseende genomförandet av myndighetens budget för budgetåret 2008.
2.
Europaparlamentet redovisar sina iakttagelser i resolutionen nedan.
3.
Europaparlamentet uppdrar åt talmannen att översända detta beslut och den resolution som utgör en del av beslutet till den verkställande direktören för Europeiska kemikaliemyndigheten, rådet, kommissionen och revisionsrätten samt att se till att de offentliggörs i Europeiska unionens officiella tidning (L-serien).
2.
Europaparlamentets beslut av den 5 maj 2010 om avslutande av räkenskaperna för Europeiska kemikaliemyndigheten för budgetåret 2008 ( C7-0202/2009 – 2009/2131(DEC) )
Europaparlamentet fattar detta beslut
–
med beaktande av den slutliga årsredovisningen för Europeiska kemikaliemyndigheten för budgetåret 2008,
–
med beaktande av revisionsrättens rapport om årsredovisningen för Europeiska kemikaliemyndigheten för budgetåret 2008, samt myndighetens svar EUT C 304, 15.12.2009, s.
33.
,
–
med beaktande av rådets rekommendation av den 16 februari 2010 (5827/2010 – C7-0061/2010 ),
–
med beaktande av artikel 276 i EG-fördraget och artikel 319 i fördraget om Europeiska unionens funktionssätt,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
, särskilt artikel 185,
–
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 EUT L 396, 30.12.2006, s.
1.
, särskilt artikel 97,
–
med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002 EGT L 357, 31.12.2002, s.
72.
, särskilt artikel 94,
–
med beaktande av artikel 77 i och bilaga VI till arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A7-0089/2010 ).
1.
Europaparlamentet godkänner avslutandet av räkenskaperna för Europeiska kemikaliemyndigheten för budgetåret 2008.
2.
Europaparlamentet uppdrar åt talmannen att översända detta beslut till den verkställande direktören för Europeiska kemikaliemyndigheten, rådet, kommissionen och revisionsrätten samt att se till att det offentliggörs i Europeiska unionens officiella tidning (L serien).
3.
Europaparlamentets resolution av den 5 maj 2010 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av budgeten för Europeiska kemikaliemyndigheten för budgetåret 2008 ( C7-0202/2009 – 2009/2131(DEC) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av den slutliga årsredovisningen för Europeiska kemikaliemyndigheten för budgetåret 2008,
–
med beaktande av revisionsrättens rapport om årsredovisningen för Europeiska kemikaliemyndigheten för budgetåret 2008, samt myndighetens svar EUT C 304, 15.12.2009, s.
33.
,
–
med beaktande av rådets rekommendation av den 16 februari 2010 (5827/2010 – C7-0061/2010 ),
–
med beaktande av artikel 276 i EG-fördraget och artikel 319 i fördraget om Europeiska unionens funktionssätt,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
, särskilt artikel 185,
–
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 EUT L 396, 30.12.2006, s.
1.
, särskilt artikel 97,
–
med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i rådets förordning (EG, Euratom) nr 1605/2002 EGT L 357, 31.12.2002, s.
72.
, särskilt artikel 94,
–
med beaktande av artikel 77 i och bilaga VI till arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet och yttrandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet ( A7-0089/2010 ).
A.
Revisionsrätten har förklarat att den har uppnått en rimlig säkerhet om att räkenskaperna för budgetåret 2008 är tillförlitliga och att de underliggande transaktionerna är lagliga och korrekta.
B.
År 2008 var myndighetens första verksamhetsår.
1.
Europaparlamentet noterar att myndigheten 2008 finansierades av ett bidrag från gemenskapen på 62 200 000 EUR i enlighet med artikel 185 i den allmänna budgetförordningen och i mindre utsträckning av avgifter som industrin erlägger vid registrering av kemikalier i enlighet med Reach-förordningen (Europaparlamentets och rådets förordning (EG) nr 1907/2006 av den 18 december 2006 om registrering, utvärdering, godkännande och begränsning av kemikalier (Reach) och om inrättande av en europeisk kemikaliemyndighet).
Verksamhetsresultat
2.
Europaparlamentet anser att myndigheten spelar en roll som kommissionen inte är i stånd att spela och att den till fullo utför sitt arbete i enlighet med unionens strategiska prioriteringar samt att dess verksamhet kompletterar andra byråers.
3.
Europaparlamentet noterar synpunkterna i den externa utvärderingen av EU:s decentraliserade byråer som kommissionen beställde 2009, i vilken det fastslås att målen och verksamheterna i det fleråriga arbetsprogrammet är förenliga med myndighetens mandat och att resultaten är användbara och av hög kvalitet och dessutom uppnås i tid.
4.
Europaparlamentet betonar dock att myndigheten skulle kunna dra nytta av att utveckla feedbackförfaranden och en starkare fokusering på kunderna.
5.
6.
Europaparlamentet noterar att det i förordning (EG) nr 1907/2006 om inrättande av myndigheten fastställs att den ska ses över vart tionde år.
Budgetförvaltning och ekonomisk förvaltning
7.
8.
9.
Parlamentet konstaterar att de likvida medlen uppgick till 18 747 210,75 EUR den 31 december 2008.
Parlamentet uppmanar kommissionen att undersöka vilka möjligheter det finns att se till att den behovsinriktade förvaltning av likvida medel som avses i artikel 15.5 i förordning (EG, Euratom) nr 2343/2002 till fullo tillämpas och vilka ändringar som krävs för att på lång sikt hålla myndighetens likvida medel på en så låg nivå som möjligt.
Personalresurser
10.
11.
12.
Internrevision
13.
Europaparlamentet konstaterar att 2008 var det första år då internrevisionstjänsten (IAS) gjorde en undersökning vid myndigheten och att en riskbedömning genomfördes i juli 2008 för att fastställa revisionsprioriteringarna och IAS revisionsplan för de kommande tre åren.
14.
o
o o
15.
Europaparlamentet hänvisar när det gäller andra övergripande iakttagelser som utgör en del av beslutet om ansvarsfrihet till sin resolution av den 5maj 2010 Antagna texter, P7_TA(2010)0139 .
om verksamhetsresultat, ekonomisk förvaltning och kontroll av byråerna.
P7_TA(2010)0201
Öppenhet och finansiering inom regionalpolitiken
A7-0139/2010
Europaparlamentets resolution av den 15 juni 2010 om öppenhet och finansiering inom regionalpolitiken ( 2009/2232(INI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av fördraget om Europeiska unionens funktionssätt, i synnerhet artiklarna 174–178,
–
med beaktande av rådets förordning (EG) nr 1083/2006 av den 11 juli 2006 om allmänna bestämmelser för Europeiska regionala utvecklingsfonden, Europeiska socialfonden och Sammanhållningsfonden EUT L 210, 31.7.2006, s.
25.
,
–
med beaktande av kommissionens förordning (EG) nr 1828/2006 av den 8 december 2006 om tillämpningsföreskrifter för rådets förordning (EG) nr 1083/2006 om allmänna bestämmelser för Europeiska regionala utvecklingsfonden, Europeiska socialfonden och Sammanhållningsfonden och för Europaparlamentets och rådets förordning (EG) nr 1080/2006 om Europeiska regionala utvecklingsfonden EUT L 371, 27.12.2006, s.
1.
,
–
med beaktande av rådets förordning (EG) nr 284/2009 av den 7 april 2009 om ändring av förordning (EG) nr 1083/2006 om allmänna bestämmelser för Europeiska regionala utvecklingsfonden, Europeiska socialfonden och Sammanhållningsfonden vad gäller vissa bestämmelser om den ekonomiska förvaltningen EUT L 94, 8.4.2009, s.
10.
,
–
med beaktande av Europaparlamentets och rådets förordning (EG) nr 397/2009 av den 6 maj 2009 om ändring av förordning (EG) nr 1080/2006 om Europeiska regionala utvecklingsfonden vad gäller stödberättigande för investeringar i energieffektivitet och förnybar energi i bostäder EUT L 126, 21.5.2009, s.
3.
,
–
med beaktande av Europaparlamentets beslut av den 22 april 2008 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2006, avsnitt III –kommissionen
EUT L 88, 31.3.2009, s.
23.
,
–
med beaktande av Europaparlamentets beslut av den 23 april 2009 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2007, avsnitt III – kommissionen
EUT L 255, 26.9.2009, s.
,
–
med beaktande av sin resolution av den 19 februari 2008 om öppenhet i ekonomiska frågor EUT C 184 E, 6.8.2009, s.
1.
,
–
med beaktande av sin resolution av den 21 oktober 2008 om styrelseformer och partnerskap på nationell och regional grundval samt på projektbasis inom regionalpolitiken Antagna texter, P6_TA(2008)0492 .
,
–
,
–
med beaktande av Europaparlamentets undersökning med titeln ’Initiativet om öppenhet i fråga om uppgifter och konsekvenserna för sammanhållningspolitiken’,
–
med beaktande av kommissionens grönbok av den 3 maj 2006 om Europeiska öppenhetsinitiativet ( KOM(2006)0194 ),
–
med beaktande av kommissionens meddelande av den 21 december 2009 med titeln ’Tjugonde årsrapporten om genomförandet av strukturfonderna (2008)’ ( KOM(2009)0617 ),
–
med beaktande av artikel 48 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för regional utveckling ( A7-0139/2010 ), och av följande skäl:
A.
B.
Enligt systemet för delad förvaltning hanteras informationen om mottagare av EU-medel på medlemsstatsnivå, men i frånvaro av en särskild skyldighet inom EU och en stark ’styrning’ från kommissionens sida skiljer sig graden av offentligt tillhandahållande av sådan information avsevärt åt mellan medlemsstaterna, vilket gör det svårt att göra jämförelser inom EU.
C.
Informationen om mottagarna av EU-finansiering gör det möjligt för allmänheten att delta i en meningsfull debatt om hur offentliga medel används, vilket är nödvändigt för fungerande demokratier.
D.
Det har inte upprättats någon koppling mellan öppenhetsinitiativet och de mer reglerade och tvingande ekonomiska kontrollerna och revisionerna.
E.
F.
G.
Tanken om insyn måste gå hand i hand med förenklingen av tilldelningsförfarandet för strukturfonderna.
1.
Europaparlamentet anser att insyn i sammanhållningspolitiken och dess programplaneringsperiod, fördelning av kostnader och tillgång till information för möjliga mottagare av medel från strukturfonderna är nödvändiga villkor för att man ska kunna uppfylla sammanhållningspolitikens övergripande mål, och att insyn därför bör införas som en sektorsövergripande princip inom sammanhållningspolitikens programplaneringsförfaranden och i beslutsprocessen.
Information om mottagare av sammanhållningsfinansiering
2.
3.
4.
5.
6.
Vad beträffar programmen inom ramen för det europeiska territoriella samarbetet vill Europaparlamentet att alla mottagare och inte bara de viktigaste förtecknas.
7.
Europaparlamentet understryker att en fullständig efterlevnad av öppenhetskraven är nödvändig och att detta bör uppnås genom lämpliga bestämmelser, bättre vägledning, en varningsmekanism och sanktioner, som en sista utväg i fall då kraven inte efterlevs.
Insyn och delad förvaltning
8.
9.
10.
11.
12.
13.
14.
Europaparlamentet uppmanar kommissionen att granska användningen av de ökade förskottsbetalningar som medlemsstaterna mottagit i enlighet med förenklingarna från 2009, som infördes genom förordning (EG) nr 1083/2006.
15.
16.
Europaparlamentet uppmanar revisorerna att anta ett strängare förhållningssätt avseende kommunikations- och informationskrav, inbegripet ’uthängning’ – i synnerhet om en statlig aktör är inblandad – och användandet av finansiella justeringar vid konstaterade bedrägerifall.
17.
Europaparlamentet välkomnar kommissionens och revisionsrättens insatser för att samordna sina revisionsmetoder.
Insyn och partnerskap
18.
19.
20.
Europaparlamentet uppmanar kommissionen att ge mer vägledning om hur partnerskapsklausulen ska tillämpas i de rådande programmen och efterlyser tillräckligt tvingande bestämmelser om partnerskap i framtida lagtexter, i synnerhet när det gäller regionala och lokala myndigheters delaktighet, dvs. valda organ som är oumbärliga partner i hela den här processen.
21.
Förbättring av insynen i samband med EU-finansiering av större projekt
22.
23.
Europaparlamentet kräver att information om stora projekt som godkänts eller inlämnats för godkännande under programperioden 2007–2013 ska offentliggöras retroaktivt på Internet.
24.
Europaparlamentet föreslår att det ska fastslås under vilka omständigheter oanvända medel får återanvändas och vilket ansvar den institution som beslutar om omfördelning av sådana medel har.
o
o o
25.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet och kommissionen.
P7_TA(2010)0405
Utnyttjande av Europeiska fonden för justering för globaliseringseffekter: Drenthe huvudgrupp 18 från Nederländerna
A7-0321/2010
Europaparlamentets resolution av den 23 november 2010 om förslaget till Europaparlamentets och rådets beslut om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning (ansökan EGF/2009/030 NL/ Drenthe huvudgrupp 18 från Nederländerna) ( KOM(2010)0531 – C7-0310/2010 – 2010/2226(BUD) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2010)0531 – C7-0310/2010 ),
–
med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning EUT C 139, 14.6.2006, s.
1.
, särskilt punkt 28,
–
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1927/2006 av den 20 december 2006 om upprättande av Europeiska fonden för justering för globaliseringseffekter EUT L 406, 30.12.2006, s.
1.
,
–
med beaktande av skrivelsen från utskottet för sysselsättning och sociala frågor,
–
med beaktande av betänkandet från budgetutskottet ( A7-0321/2010 ), och av följande skäl:
A.
Europeiska unionen har inrättat lagstiftningsinstrument och budgetinstrument för att kunna ge kompletterande stöd till arbetstagare som blivit arbetslösa till följd av genomgripande strukturförändringar inom världshandeln och för att underlätta deras återinträde på arbetsmarknaden.
B.
Tillämpningsområdet för fonden har utvidgats för ansökningar om stöd från fonden som inges från och med den 1 maj 2009 och omfattar nu stöd till arbetstagare som har blivit uppsagda som en direkt följd av den globala finansiella och ekonomiska krisen.
C.
Unionens ekonomiska stöd till arbetstagare som har blivit uppsagda bör vara dynamiskt och ges så snabbt och effektivt som möjligt, i enlighet med Europaparlamentets, rådets och kommissionens gemensamma uttalande, som antogs vid förlikningsmötet den 17 juli 2008, och med vederbörlig hänsyn till bestämmelserna i det interinstitutionella avtalet av den 17 maj 2006 om antagandet av beslut rörande fondens utnyttjande.
D.
Nederländerna har ansökt om ekonomiskt bidrag från fonden till följd av 140uppsägningar vid två företag som är verksamma inom sektorn Nace rev2 huvudgrupp 18 (Grafisk produktion och reproduktion av inspelningar) i Nuts II-regionen Drenthe.
E.
Ansökan uppfyller kriterierna för berättigande till stöd enligt förordningen om upprättande av Europeiska fonden för justering för globaliseringseffekter.
1.
Europaparlamentet uppmanar de berörda institutionerna att vidta de åtgärder som krävs för att Europeiska fonden för justering för globaliseringseffekter snarast ska kunna tas i anspråk.
2.
3.
4.
5.
Europaparlamentet välkomnar det faktum att kommissionen i samband med utnyttjandet av Europeiska fonden för justering för globaliseringseffekter föreslagit en alternativ källa till betalningsbemyndiganden utöver oanvända medel från Europeiska socialfonden, efter många påminnelser från Europaparlamentet om att Europeiska fonden för justering för globaliseringseffekter inrättades som ett separat särskilt instrument med egna mål och tidsfrister och att tillbörliga budgetposter för överföringar därför måste fastställas.
6.
7.
Europaparlamentet påminner om att en utvärdering av hur Europeiska fonden för justering för globaliseringseffekter fungerar och vilket mervärde den skapar bör göras inom ramen för den allmänna bedömningen av programmen och andra instrument som skapats genom det interinstitutionella avtalet av den 17 maj 2006, i samband med halvtidsöversynen av den fleråriga budgetramen 2007–2013.
8.
Europaparlamentet välkomnar det nya formatet för kommissionens förslag, där det i motiveringsdelen läggs fram tydliga och detaljerade uppgifter om ansökan med en analys av kriterier för stödberättigande och en förklaring av orsakerna till att ansökan godkänts, vilket ligger i linje med parlamentets krav.
9.
Europaparlamentet godkänner det bifogade beslutet.
10.
Europaparlamentet uppdrar åt talmannen att tillsammans med rådets ordförande underteckna beslutet och se till att det offentliggörs i Europeiska unionens officiella tidning.
11.
Europaparlamentet uppdrar åt talmannen att översända denna resolution med bilaga till rådet och kommissionen.
BILAGA
EUROPAPARLAMENTETS OCH RÅDETS BESLUT
av den
om utnyttjande av Europeiska fonden för justering för globaliseringseffekter i enlighet med punkt 28 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning (ansökan EGF/2009/030 NL/ Drenthe huvudgrupp 18 från Nederländerna)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av fördraget om Europeiska unionens funktionssätt,
med beaktande av det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning EUT C 139, 14.6.2006, s.
1.
, särskilt punkt 28,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1927/2006 av den 20 december 2006 om upprättande av Europeiska fonden för justering för globaliseringseffekter EUT L 406, 30.12.2006, s.
1.
av följande skäl:
(1)
Europeiska fonden för justering för globaliseringseffekter (nedan kallad fonden) inrättades för att ge kompletterande stöd till arbetstagare som blivit arbetslösa till följd av de genomgripande strukturförändringar som skett inom världshandeln på grund av globaliseringen och för att underlätta deras återinträde på arbetsmarknaden.
(2)
Tillämpningsområdet för fonden har utvidgats, och från och med den 1 maj 2009 är det möjligt att söka stöd för åtgärder som riktas till arbetstagare som har blivit uppsagda som en direkt följd av den globala finansiella och ekonomiska krisen.
(3)
Det interinstitutionella avtalet av den 17 maj 2006 gör det möjligt att använda medel från fonden upp till ett belopp på högst 500 miljoner EUR per år.
(4)
Nederländerna lämnade den 30 december 2009 in en ansökan om medel från fonden med anledning av uppsägningar vid två företag som är verksamma inom huvudgrupp 18 (Grafisk produktion och reproduktion av inspelningar) enligt Nace rev2, i Nuts II-regionen Drenthe (NL13), och kompletterade ansökan med ytterligare uppgifter fram till den 6 maj 2010.
Ansökan uppfyller villkoren för fastställande av det ekonomiska stödet enligt artikel 10 i förordning (EG) nr 1927/2006.
Kommissionen föreslår därför att ett belopp på 453 632 EUR ska anslås.
(5)
Fonden bör därför utnyttjas för att bevilja det ekonomiska stöd som Nederländerna ansökt om.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Europeiska fonden för justering för globaliseringseffekter ska belastas med 453 632 EUR i åtagande- och betalningsbemyndiganden ur Europeiska unionens allmänna budget för 2010.
Artikel 2
På Europaparlamentets vägnar På rådets vägnar
Ordförande Ordförande
P7_TA(2010)0426
Civilrättsliga, handelsrättsliga, familjerättsliga och internationella privaträttsliga aspekter av handlingsplanen för att genomföra Stockholmsprogrammet
A7-0252/2010
Europaparlamentets resolution av den 23 november 2010 om civilrättsliga, handelsrättsliga, familjerättsliga och internationella privaträttsliga aspekter av handlingsplanen för att genomföra Stockholmsprogrammet ( 2010/2080(INI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av artiklarna 67 och 81 i fördraget om Europeiska unionens funktionssätt,
–
med beaktande av kommissionens meddelande av den 10 juni 2009 med titeln ”Ett område med frihet, säkerhet och rättvisa i allmänhetens tjänst” ( KOM(2009)0262 ), i vilket kommissionen redogör för sina prioriteringar för området med frihet, säkerhet och rättvisa för 2010–2014, kommissionens utvärdering av Haagprogrammet och handlingsplanen ( KOM(2009)0263 ) och den därtill hörande resultattavlan för genomförande ( SEK(2009)0765 ) samt bidrag från de nationella parlamenten, det civila samhället och EU-byråer och EU-organ,
–
med beaktande av dokumentet från rådets ordförandeskap av den 2 december 2009 med titeln ”Stockholmsprogrammet – Ett öppet och säkert Europa i medborgarnas tjänst och för deras skydd” (17024/09),
–
med beaktande av sin resolution av den 25 november 2009 om Stockholmsprogrammet EUT C 285 E, 21.10.2010, s.
12.
,
–
med beaktande av kommissionens meddelande av den 20 april 2010 med titeln ”Handlingsplan för att genomföra Stockholmsprogrammet” ( KOM(2010)0171 ),
–
med beaktande av sin resolution av den 17 juni 2010 om rättslig utbildning – Stockholmsprogrammet Antagna texter, P7_TA(2010)0242 .
,
–
med beaktande av artikel 48 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för rättsliga frågor och yttrandena från utskottet för internationell handel, utskottet för den inre marknaden och konsumentskydd ( A7-0252/2010 ), och av följande skäl:
A.
Området med frihet, säkerhet och rättvisa är ett gemensamt ansvarsområde för unionen och medlemsstaterna.
B.
C.
D.
E.
Om vi ser tillbaka på vad som har uppnåtts inom ramen för området med frihet, säkerhet och rättvisa kan vi konstatera att i första hand harmoniseringen av internationella privaträttsliga bestämmelser har gått framåt i snabb takt.
F.
Vidare finns det fall av harmonisering eller tillnärmning som lämpar sig för vissa områden där en standardisering är önskvärd, om inte nödvändig, till exempel på konsumentskyddsområdet, men där detta utnyttjas i begränsad utsträckning inom ramen för området med frihet, säkerhet och rättvisa.
G.
Utarbetandet av en europeisk avtalsrätt kommer att vara en av de viktigaste uppgifterna inom ramen för området med frihet, säkerhet och rättvisa under de kommande åren, och detta arbete kan komma att resultera i en så kallad 28:e civilrättslig ordning som ett alternativ till det traditionella sättet att åstadkomma en harmonisering av lagstiftning på specifika områden.
H.
I.
J.
K.
L.
Detta utgör unionens verkliga styrka och samtidigt en utmaning för området med frihet, säkerhet och rättvisa och bör inte uppfattas som oförenligt med utvecklingen av och undervisningen i en verklig europeisk rättskultur.
M.
Beslutsamheten i ingressen till Lissabonfördraget att ”lägga grunden till en allt fastare sammanslutning mellan de europeiska folken” förutsätter en minskning av den verkliga och upplevda klyftan mellan EU, dess lagstiftning och medborgarna.
N.
Unionslagstiftningen måste vara i medborgarnas tjänst, inte minst på områden som rör familjerätt och civilståndsfrågor.
O.
Kommissionen måste säkerställa att handlingsplanen för Stockholmsprogrammet verkligen återspeglar enskilda individers och företags, och särskilt små och medelstora företags, behov av mer Europa (vad gäller rörlighet, anställningsrättigheter, näringslivets behov och lika möjligheter), och samtidigt främja rättssäkerhet och tillgång till snabb och effektiv rättslig prövning.
P.
I detta sammanhang måste allt mer vikt läggas vid att förenkla rättsapparaten och rättssystemet och skapa tydligare och mer tillgängliga förfaranden, samtidigt som hänsyn tas till behovet av att minska kostnaderna, särskilt i det rådande ekonomiska klimatet.
Q.
1.
Europaparlamentet lyckönskar kommissionen till dess förslag till handlingsplan.
2.
Europaparlamentet anser icke desto mindre att det är hög tid att fundera över den framtida utvecklingen inom området med frihet, säkerhet och rättvisa, och uppmanar kommissionen att initiera en ingående diskussion med alla berörda parter, däribland domare och andra yrkesutövare inom rättsväsendet.
3.
4.
Europaparlamentet uppmanar kommissionen att i samråd med parlamentet vidta åtgärder med anledning av parlamentets resolution av den 17 juni 2010 om juridisk utbildning.
5.
Europaparlamentet understryker på nytt behovet av att utnyttja alla till buds stående medel för att främja en europeisk rättskultur, särskilt genom juridisk utbildning och fortbildning.
6.
7.
Europaparlamentet konstaterar att befintliga inrättningar och nätverk för nationell utbildning bör utgöra den motor som för utvecklingen av en gemensam europeisk rättskultur framåt med tanke på att de vid medlemsstaternas genomförande av unionslagstiftningen befinner sig i främsta leden och att de har direktkontakt med ländernas domstolar och rättsväsende och även en djup förståelse av de olika medlemsstaternas rättskulturer och behov på detta område.
8.
9.
10.
11.
12.
13.
14.
15.
Parlamentet uppmanar med kraft kommissionen att svara på dess resolution av den 1 februari 2007 EUT C 250 E, 25.10.2007, s.
16.
Europaparlamentet välkomnar grönboken av den 1 juli 2010 om politiska alternativ för främjande av en europeisk avtalsrätt för konsumenter och företag och stöder kommissionens ambitiösa initiativ till en europeisk avtalsrättsakt som kan tillämpas frivilligt av avtalsparterna( KOM(2010)0348 ).
17.
Europaparlamentet betonar vikten av gränsöverskridande rättsliga prövningar när det gäller att lösa fall av bedrägerier och vilseledande affärsmetoder som har sitt ursprung i en medlemsstat och drabbar enskilda medborgare, icke-statliga organisationer och små och medelstora företag i andra medlemsstater.
18.
Europaparlamentet uppmärksammar sin resolution av den 10 mars 2009 om samarbete mellan medlemsstaternas domstolar i fråga om bevisupptagning i mål och ärenden av civil eller kommersiell natur EUT C 87 E, 1.4.2010, s.
21.
19.
20.
Europaparlamentet anser att sådana initiativ blir allt viktigare med tanke på konjunkturnedgången.
21.
Europaparlamentet uppmanar kommissionen att utan dröjsmål arbeta vidare med dessa initiativ och att fokusera på möjligheten att inrätta en självständig europeisk mekanism för insyn i och/eller frysning av tillgångar i gränsöverskridande fall.
22.
Europaparlamentet understryker att detta område får betydande finansiella och ryktesmässiga konsekvenser, och uppmuntrar därför till en preventiv användning av alternativa tvistelösningsförfaranden.
23.
Europaparlamentet anser att konsolideringen av lagstiftningen, genom de medel som fastställs i detta betänkande, med säkerhet bör leda till en utveckling och förstärkning av de ekonomiska och yrkesmässiga förbindelserna och därmed bidra till arbetet med att skapa en verklig inre marknad.
24.
25.
Europaparlamentet betonar att Stockholmsprogrammet syftar till att skapa ett europeiskt område med frihet, säkerhet och rättvisa som garanterar medborgarna grundläggande rättigheter, inklusive rätt till fri företagsamhet, för att företagarandan inom de olika sektorerna av ekonomin ska kunna utvecklas.
26.
Europaparlamentet ger sitt helhjärtade stöd till kommissionens målsättning att anta lagstiftning som medför minskade affärs- och transaktionskostnader, särskilt för små och medelstora företag.
27.
28.
29.
30.
31.
32.
33.
34.
35.
1).
36.
37.
38.
39.
40.
41.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen och medlemsstaternas regeringar och parlament.
P7_TA(2011)0013
Internationella adoptioner i Europeiska unionen
B7-0029 , 0030 , 0036 , 0037 och 0038/2011
Europaparlamentets resolution av den 19 januari 2011 om internationella adoptioner i Europeiska unionen
Europaparlamentet utfärdar denna resolution
–
med beaktande av FN:s konvention om barnets rättigheter, som antogs av FN:s generalförsamling den 20 november 1989, i synnerhet artikel 21,
–
med beaktande av 1967 års europeiska konvention om adoption av barn,
–
med beaktande av konventionen om skydd av barn och samarbete vid internationella adoptioner (undertecknad i Haag den 29 maj 1993) och av Europeiska konventionen om utövandet av barns rättigheter, antagen den 25 januari 1996 (ETS nr 160),
–
med beaktande av artikel 24 i Europeiska unionens stadga om de grundläggande rättigheterna,
–
–
med beaktande av sin resolution av den 12 december 1996 om förbättrad lagstiftning och förbättrat samarbete mellan medlemsstaterna beträffande adoption av minderåriga EGT C 20, 20.1.1997, s.
176.
,
–
med beaktande av sin resolution av den 16 januari 2008 om en EU-strategi för barnets rättigheter EUT C 41 E, 19.2.2009, s.
24.
,
–
A.
Varje barns välmående och tryggandet av barns intressen är ytterst viktigt, och skyddet av barns rättigheter är ett av EU:s mål.
B.
Adoptioner hör till medlemsstaternas behörighetsområde, och det är medlemsstaterna som genomför de relevanta förfarandena i enlighet med barnens intressen.
C.
Det finns gällande konventioner om skyddet av barn och föräldrars ansvar, närmare bestämt 1967 års europeiska konvention om adoptioner av barn som syftar till att närma medlemsstaternas lagstiftning i fall där adoptionen innebär att barnet flyttas från ett land till ett annat, och 1993 års konvention om skydd av barn och samarbete vid internationella adoptioner (Haagkonventionen).
D.
Alla EU:s medlemsstater har undertecknat Haagkonventionen.
E.
Betydande framsteg har kunnat göras till följd av Haagkonventionen.
F.
I FN:s konvention om barnets rättigheter och i Haagkonvention beskrivs familjen som den grundläggande enheten i samhället och den naturliga miljön för barns utveckling och välfärd i de allra flesta fall och som förstahandsval när det gäller omvårdnad av barn.
G.
Om familjen, dvs. förstahandsvalet, inte kan ta hand om barnen, bör adoption vara ett av de naturliga andrahandsval som kan komma i fråga, medan omhändertagande på institution bör vara den absolut sista lösningen.
H.
Barn som växer upp i otrygghet är ett allvarligt problem inom Europa, särskilt otryggheten bland övergivna barn och barn som växer upp på institutioner, och detta problem måste verkligen tas på största allvar.
I.
Kränkningar av barns rättigheter, våld mot barn och människohandel med barn för adoption, prostitution, olagligt arbete, tvångsäktenskap, gatutiggeri eller andra olagliga syften är fortfarande ett problem inom EU.
J.
Det är viktigt att barns rätt att leva i en familj tryggas och att man ser till att barn inte tvingas bo på barnhem under långa perioder.
K.
1.
Europaparlamentet begär att man undersöker möjligheten att på EU-nivå samordna de strategier som är kopplade till instrumentet för internationella adoptioner, i enlighet med de internationella konventionerna, för att förbättra hjälpen från informationstjänster, förberedandet av adoptioner mellan länder, handläggningen av internationella adoptionsansökningar och uppföljningen efter en adoption, med tanke på att alla internationella konventioner om skydd av barns rättigheter erkänner föräldralösa och övergivna barns rätt att leva i en familj och få skydd.
2.
Europaparlamentet uppmanar kommissionen att ta hänsyn till hur de nationella systemen fungerar på EU-nivå.
3.
Europaparlamentet anser att när så är möjligt och om det är till barnets bästa, ska en adoption i första hand ske i barnets ursprungsland där möjliga alternativ skulle kunna vara en familjehemslösning, så som en fosterfamilj eller annat boende, eller ett omhändertagande hos en familj inom ramen för internationell adoption, och att placering på institution bör användas bara som en tillfällig lösning.
4.
Europaparlamentet understryker att det vid internationella adoptioner är den nationella lagstiftningen i adoptivföräldrarnas ursprungsland som måste tillämpas i fråga om skyddet av barnets rättigheter på lång sikt.
5.
Europaparlamentet uppmanar medlemsstaterna och kommissionen att i samarbete med Haagkonferensen, Europarådet och barnorganisationer ta fram en ram för att garantera insyn i och effektiva bedömningar av utvecklingen när det gäller övergivna och adopterade barn, även barn som genomgått internationell adoption, samt att samordna sina insatser för att förhindra människohandel med barn i adoptionssyfte.
6.
Europaparlamentet uppmanar alla EU:s institutioner att spela en aktivare roll i och utöva påtryckning vid Haagkonferensen och på så sätt sträva efter att förbättra, effektivisera och underlätta internationella adoptionsförfaranden och få bort onödig byråkrati, och samtidigt åta sig att trygga rättigheterna för barn från tredjeländer.
7.
Europaparlamentet uppmanar de behöriga nationella myndigheterna att regelbundet rapportera till ursprungsmedlemsstaten om vad som händer med de barn som genomgått internationell adoption.
8.
Europaparlamentet uppmanar medlemsstaterna att uppmärksamma de psykiska, känslomässiga och sociala/utbildningsrelaterade följder som det kan få om ett barn flyttas från sitt ursprungsland samt att erbjuda stöd till adoptivföräldrarna och adoptivbarnet.
9.
Europaparlamentet uppmanar medlemsstaterna att i synnerhet uppmärksamma barn med särskilda behov, exempelvis barn med medicinska behov och barn med funktionshinder.
10.
11.
Europaparlamentet uppmanar EU:s institutioner och medlemsstater att engagera sig aktivt för att bekämpa människohandel med barn i adoptionssyfte.
12.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till Europeiska rådets ordförande, rådet, kommissionen och Haagkonferensen samt till medlemsstaternas regeringar och parlament.
P7_TA-PROV(2011)0112
Utnämning av den verkställande direktören för Europeiska försäkrings- och tjänstepensionsmyndigheten (EIOPA)
B7-0221/2011
Europaparlamentets resolution av den 24 mars 2011 om utnämningen av verkställande direktör för Europeiska tillsynsmyndigheten (Europeiska försäkrings- och tjänstepensionsmyndigheten)
Europaparlamentet utfärdar denna resolution
–
med beaktande av skrivelsen av den 10 mars 2011 från Europeiska tillsynsmyndigheten (Europeiska försäkrings- och tjänstepensionsmyndigheten),
–
48.
,
–
med beaktande av det faktum att utskottet för ekonomi och valutafrågor vid sitt sammanträde den 17 mars 2011 hörde den kandidat som valts ut av styrelsen för Europeiska tillsynsmyndigheten (Europeiska försäkrings- och tjänstepensionsmyndigheten),
–
med beaktande av artikel 120 i arbetsordningen, och av följande skäl:
A.
1.
Europaparlamentet ger sitt samtycke till utnämningen av Carlos Montalvo till verkställande direktör för Europeiska tillsynsmyndigheten (Europeiska försäkrings- och tjänstepensionsmyndigheten).
2.
Europaparlamentet uppdrar åt talmannen att vidarebefordra denna resolution till Europeiska tillsynsmyndigheten (Europeiska försäkrings- och tjänstepensionsmyndigheten).
P7_TA-PROV(2011)0162
Ansvarsfrihet för budgetåret 2009 – Europeiska datatillsynsmannen
A7-0117/2011
1.
Europaparlamentets beslut av den 10 maj 2011 om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2009, avsnitt IX – Europeiska datatillsynsmannen ( C7-0219/2010 – 2010/2150(DEC) )
Europaparlamentet fattar detta beslut
–
,
–
med beaktande av Europeiska unionens slutliga årsredovisning för budgetåret 2009 ( SEK(2010)0963 – C7-0219/2010 ) EUT C 308, 12.11.2010, s.
1.
,
–
med beaktande av Europeiska datatillsynsmannens årsrapport om internrevisioner som genomförts under 2009,
–
med beaktande av revisionsrättens årsrapport om genomförandet av budgeten för budgetåret 2009, samt de granskade institutionernas svar EUT C 303, 9.11.2010, s.
1.
,
–
med beaktande av förklaringen om räkenskapernas tillförlitlighet och de underliggande transaktionernas laglighet och korrekthet som avges av revisionsrätten i enlighet med artikel 287 i fördraget om Europeiska unionens funktionssätt EUT C 308, 12.11.2010, s.
129.
,
–
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
, särskilt artiklarna 50, 86, 145, 146 och 147,
–
med beaktande av artikel 77 och bilaga VI i arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet ( A7-0117/2011 ).
1.
Europaparlamentet beviljar Europeiska datatillsynsmannen ansvarsfrihet för genomförandet av budgeten för budgetåret 2009.
2.
Europaparlamentet redovisar sina iakttagelser i resolutionen nedan.
3.
Europaparlamentet uppdrar åt talmannen att översända detta beslut och den resolution som utgör en del av beslutet till rådet, kommissionen, domstolen, revisionsrätten, Europeiska ombudsmannen och Europeiska datatillsynsmannen samt att se till att de offentliggörs i Europeiska unionens officiella tidning (L-serien).
2.
Europaparlamentets resolution av den 10 maj 2011 med de iakttagelser som utgör en del av beslutet om ansvarsfrihet för genomförandet av Europeiska unionens allmänna budget för budgetåret 2009, avsnitt IX – Europeiska datatillsynsmannen ( C7-0219/2010 – 2010/2150(DEC) )
Europaparlamentet utfärdar denna resolution
–
,
–
med beaktande av Europeiska unionens slutliga årsredovisning för budgetåret 2009 ( SEK(2010)0963 – C7-0219/2010 ) EUT C 308, 12.11.2010, s.
1.
,
–
med beaktande av Europeiska datatillsynsmannens årsrapport om internrevisioner som genomförts under 2009, riktad till den myndighet som beviljar ansvarsfrihet,
–
med beaktande av revisionsrättens årsrapport om genomförandet av budgeten för budgetåret 2009, samt de granskade institutionernas svar EUT C 303, 9.11.2010, s.
1.
,
–
med beaktande av förklaringen om räkenskapernas tillförlitlighet och de underliggande transaktionernas laglighet och korrekthet som avges av revisionsrätten i enlighet med artikel 287 i fördraget om Europeiska unionens funktionssätt EUT C 308, 12.11.2010, s.
129.
,
–
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
, särskilt artiklarna 50, 86, 145, 146 och 147,
–
med beaktande av artikel 77 och bilaga VI i arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet ( A7-0117/2011 ).
1.
Europaparlamentet noterar att Europeiska ombudsmannen under 2009 hade tillgång till åtagandebemyndiganden som sammanlagt uppgick till 7 miljoner EUR (2008: 5,3 miljoner EUR 2006: 4,1 miljoner EUR.
), med en utnyttjandegrad på 81,44 procent, vilket är lägre än genomsnittet för de övriga institutionerna (97,69 procent).
2.
Europaparlamentet konstaterar att revisionsrätten under utarbetandet av årsrapporten för budgetåret 2009 genomförde en fördjupad bedömning av gransknings- och kontrollsystemen i domstolen, Europeiska ombudsmannen och Europeiska datatillsynsmannen som omfattade en granskning av ett ytterligare urval av betalningstransaktioner avseende personalresurser och andra administrativa utgifter.
3.
Europaparlamentet noterar att revisionsrätten fann att de uppgifter som Europeiska datatillsynsmannen förfogade över för att garantera att tillägg som fastställs i tjänsteföreskrifterna för tjänstemännen i Europeiska gemenskaperna EGT L 56, 4.3.1968, s.
1.
4.
Europaparlamentet stöder revisionsrättens förslag om att Europeiska datatillsynsmannens personal bör uppmanas att med jämna mellanrum visa upp handlingar som styrker deras personliga situation, och anser att Europeiska datatillsynsmannen bör förbättra sitt system för övervakning och kontroll av dessa handlingar vid lämplig tidpunkt.
5.
6.
Europaparlamentet noterar revisionsrättens uppgift att Europeiska datatillsynsmannen inte hade infört ett system för efterhandskontroll vid behov, såsom krävs enligt budgetförordningen, och att det enligt de normer för internkontroll som antagits av Europeiska datatillsynsmannen inte krävs att undantag till de ekonomiska standardförfarandena registreras på vederbörligt sätt i ett centralt register.
7.
8.
9.
Europaparlamentet noterar att revisionsrätten i sin årsrapport angav att revisionen inte ledde till några väsentliga iakttagelser när det gäller Europeiska datatillsynsmannen.
10.
11.
Europaparlamentet påminner, på grundval av det administrativa samarbetsavtalet mellan generalsekreterarna för kommissionen, parlamentet och rådet, som undertecknades tillsammans med Europeiska datatillsynsmannen den 7 december 2006 för ytterligare en period på tre år från och med den 16 januari 2007, om att den administrativa hanteringen av alla Europeiska datatillsynsmannens tjänsteresor sköts av kommissionens utbetalningsbyrå, och om att utvärderingen (som i själva verket genomförts av kommissionens internrevisor, i egenskap av datatillsynsmannens tjänst för internrevision på grundval av det administrativa samarbetsavtalet), har visat att detta system för internkontroll fungerar och är effektivt samt att det gav en rimlig säkerhet när det gäller Europeiska datatillsynsmannens uppnående av sina mål.
12.
Europaparlamentet välkomnar den årliga publiceringen av vilka ekonomiska intressen som institutionens ledamöter har (Europeiska datatillsynsmannen och den biträdande datatillsynsmannen), i vilken arvoderade tjänster eller verksamheter och deklarerad yrkesverksamhet redovisas.
13.
Europaparlamentet begär att Europeiska datatillsynsmannen i sin kommande verksamhetsrapport (budgetåret 2010) inkluderar ett kapitel med en detaljerad redovisning av uppföljningen under året av parlamentets tidigare beslut avseende ansvarsfriheten.
P7_TA-PROV(2011)0163
Ansvarsfrihet för 2009: EU-byråernas verksamhetsresultat, ekonomiska förvaltning och kontroll
A7-0149/2011
Europaparlamentets resolution av den 10 maj 2011 om ansvarsfrihet för 2009: EU-byråernas verksamhetsresultat, ekonomiska förvaltning och kontroll 2010/2271(DEC)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens rapport till Europaparlamentet av den 15 oktober 2008 om uppföljningen av besluten om ansvarsfrihet 2006 ( KOM(2008)0629 ) och det åtföljande arbetsdokumentet från kommissionen ( SEK(2008)2579 ),
–
med beaktande av kommissionens meddelande av den 11 mars 2008 ’EU:s tillsynsmyndigheter – mot en gemensam ansats’ ( KOM(2008)0135 ),
–
med beaktande av sin resolution av den 5 maj 2010 om ansvarsfrihet 2008: byråernas verksamhetsresultat, ekonomiska förvaltning och kontroll EUT L 252, 25.9.2010, s.
241.
,
–
med beaktande av rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget EGT L 248, 16.9.2002, s.
1.
,
–
med beaktande av kommissionens förordning (EG, Euratom) nr 2343/2002 EGT L 357, 31.12.2002, s.
72.
av den 19 november 2002 med rambudgetförordning för de gemenskapsorgan som avses i artikel 185 i förordning (EG, Euratom) nr 1605/2002, särskilt artikel 96,
–
med beaktande av revisionsrättens särskilda rapport nr 5/2008 ’Unionens tillsynsmyndigheter: att uppnå resultat’,
–
om årsredovisningarna för de decentraliserade byråerna för budgetåret 2009,
–
med beaktande av den undersökning som offentliggjordes den 7 april 2009 om lämpligheten och möjligheten av att inrätta gemensamma stödtjänster för EU-byråer,
–
med beaktande av sin förklaring av den 18 maj 2010 om unionens insatser när det gäller att bekämpa korruption Antagna texter, P7_TA(2010)0176 .
,
–
med beaktande av artikel 77 och bilaga VI i arbetsordningen,
–
med beaktande av betänkandet från budgetkontrollutskottet ( A7-0149/2011 ), och av följande skäl:
A.
Denna resolution innehåller för varje byrå, i den mening som avses i artikel 185 i förordning (EG, Euratom) nr 1605/2002, de övergripande iakttagelserna i samband med besluten om ansvarsfrihet enligt artikel 96 i förordning (EG, Euratom) nr 2343/2002 och artikel 3 i bilaga VI i parlamentets arbetsordning.
B.
Antalet byråer har ökat på ett sätt som saknar motstycke under de senaste åren, vilket har gjort det möjligt att lägga ut vissa av kommissionens uppgifter på externa organ.
C.
Efter antagande av ovannämnda meddelande från kommissionen av den 11 mars 2008 har parlamentet, rådet och kommissionen på nytt börjat arbeta med projektet att utforma en gemensam ram för gemenskapsbyråerna och 2009 bildat en interinstitutionell arbetsgrupp för byråer.
D.
Den interinstitutionella arbetsgruppen sammanträdde för tredje gången på politisk nivå den 10 november 2010 och diskuterade följande punkter: kriterier för inrättandet av nya organ, valet av säte för organen och avtalet om säte, styrelsernas sammansättning, förfarandena för utnämning av direktörer, utvärdering och resultat, det fleråriga programmet samt administrativt stöd.
E.
Revisionsrätten planerar också att överväga organens resultat och lägga fram en särskild rapport om kostnadsriktmärkning för unionens byråer i slutet av 2011.
F.
Unionens bidrag till decentraliserade byråer har ökat drastiskt mellan 2000 och 2011.
G.
I Europaparlamentets förklaring av den 18 maj 2010 om unionens insatser när det gäller att bekämpa korruption uppmanas kommissionen och EU:s relevanta organ att vidta alla nödvändiga åtgärder och tillhandahålla tillräckliga resurser för att garantera att EU-medel inte blir föremål för korruption, och att tillämpa avskräckande straffpåföljder i de fall där korruption och bedrägeri konstaterats.
I.
GEMENSAMMA UTMANINGAR NÄR DET GÄLLER EKONOMISK FÖRVALTNING
Överförda och förfallna driftsanslag
1.
2.
3.
Likviditetsförvaltning
4.
Brister i upphandlingsförfarandena
5.
Europaparlamentet är återigen bekymrat över revisionsrättens konstaterande att flera byråer hade brister i sina upphandlingsförfaranden.
6.
7.
Europaparlamentet uppmanar i detta avseende byråerna att
–
förbättra insynen i uppskattningar och ansvar för projekt,
–
förstärka sitt upphandlingsgodkännande i finansieringsbeslut och på arbetsprogramsnivå,
–
säkerställa en uttömmande redovisning av undantag i sina årliga verksamhetsrapporter,
–
säkerställa adekvat uppföljning av potentiella regelbrott,
–
utveckla och rapportera om efterhandskontroller.
8.
Europaparlamentet uppmuntrar dessutom byråerna att utarbeta och därefter regelbundet aktualisera en heltäckande tabell som beskriver deras ekonomiska flöden och de ekonomiska och operativa aktörernas skyldigheter.
9.
Europaparlamentet uppmanar alla byråer att på sina respektive webbplatser offentliggöra en förteckning över alla avtal som tilldelats under åtminstone de senaste tre åren och uppmanar kommissionen att fortsätta att göra denna information mer tillgänglig och slutligen integrera den i sitt system för finansiell öppenhet.
10.
Handläggning av bidrag
11.
Europaparlamentet anser att det är viktigt att byråerna förbättrar sin handläggning av bidrag genom att
–
genomföra kontroller på plats hos bidragsmottagare,
–
främja standardiserade enhetskostnader per kategori i stället för bidrag som bygger på ersättning för stödberättigande kostnader,
–
tydligt beskriva, informera om och övervaka aktörernas förpliktelser,
–
tillhandahålla en verksamhetsplan som godkänts av alla aktörer.
II.
GEMENSAMMA UTMANINGAR NÄR DET GÄLLER PERSONAL
Rekryteringsförfaranden
12.
–
Det finns inga bevis för att urvalskriterierna och de tröskelvärden som kandidaterna måste uppfylla för att bli kallade till skriftliga prov eller intervjuer har fastställts innan utvärderingsprocessen inleds.
–
Rekryteringsförfarandena är otillräckligt dokumenterade.
–
Interna och externa kandidater behandlas ojämlikt i rekryteringsförfarandet.
–
Begränsad konkurrens.
13.
Europaparlamentet anser att man bör inrätta ett system för dubbelkontroll mellan byråerna, så att man upptäcker om en person gjort sig skyldig till tjänstefel eller felaktig förvaltning vid en byrå där personen tidigare tjänstgjort, när denna person ansöker om tjänst vid en annan byrå.
14.
–
respektera en tidsfrist vid utnämningen av ledamöter till uttagningskommittéer,
–
utarbeta intervjufrågor och innehåll i skriftliga prov i förväg,
–
bedöma skriftliga prov anonymt,
–
förbereda modellsvar för intervjufrågor och skriftliga prov,
–
protokollföra alla rekryteringsbeslut,
–
använda ett elektroniskt rekryteringsverktyg för att underlätta rekryterings- och urvalsprocessen,
och betonar behovet av att konsekvent genomföra denna policy och visa att den ger resultat.
Genomförande av rekryteringsplaner
15.
16.
17.
Parlamentet uppmanar kommissionen att redogöra för om det finns bestämmelser om relevanta arbetsuppgifter och skyldigheter för tjänstemän i enlighet med artikel 16 i Tjänsteföreskrifterna för tjänstemännen i Europeiska Unionen EGT L 56, 4.3.1968, s.
1.
(så kallade tidsfrister vid byte av arbetsplats) vid alla byråerna och hur de tillämpas.
Tillfällig personal
18.
Intressekonflikter
19.
20.
Europaparlamentet uppmanar kommissionen att ge parlamentet en utförlig översikt över de kriterier som tillämpas för att se till att den rekryterade personalen är oberoende, i synnerhet när det gäller potentiella intressekonflikter, och att tillämpa avskräckande påföljder i de fall regelbrott upptäcks.
21.
Europaparlamentet uppmanar revisionsrätten att göra en heltäckande analys av byråernas sätt att hantera situationer där det kan finnas risk för intressekonflikter.
III.
GEMENSAMMA UTMANINGAR NÄR DET GÄLLER INTERNKONTROLLSYSTEM
22.
Sammanfattningar av internrevisionsrapporter
23.
Europaparlamentet uppmanar direktörerna för respektive byrå att till fullo fullgöra sin skyldighet att i sina rapporter med sammanfattningar av rapporterna från internrevisionstjänsten till den myndighet som ska bevilja ansvarsfrihet inkludera följande:
–
antal och typ av internrevisioner som utförts av internrevisionstjänsten,
–
alla rekommendationer (även sådana som byrån eventuellt skulle kunna avvisa) coh
–
alla åtgärder som vidtagits med anledning av dessa rekommendationer.
Parlamentet välkomnar i detta sammanhang Frontex initiativ att främja en enhetlig struktur för alla byråer för dessa sammanfattningar till myndigheten som ska bevilja ansvarsfrihet.
24.
Internrevisionstjänstens roll
25.
Parlamentet betonar särskilt att interrevisionstjänsten utfärdar oberoende yttranden om kvaliteten på förvaltnings- och kontrollsystemen och lämnar rekommendationer om förbättringar av villkoren för genomförandet av verksamheterna och främjandet av sund ekonomisk förvaltning från byråernas sida.
26.
Europaparlamentet uppmanar därför byråernas styrelser att vederbörligen beakta rekommendationerna från internrevisionstjänsten för att snabbt avhjälpa de upptäckta bristerna.
27.
28.
Europaparlamentet rekommenderar starkt att revisionsrätten i sina årsrapporter om byråerna gör en hänvisning till internrevisionstjänstens slutsatser samt presenterar en utvärdering av hur byråerna efterkommit internrevisionstjänstens rekommendationer.
29.
Internrevisionsfunktionens roll
30.
Europaparlamentet uppmanar eftertryckligen byråerna att inrätta en internrevisionsfunktion som ska ge direktörerna stöd och råd om förvaltningen av den interna kontrollen och utföra riskbedömningar samt interna revisioner.
31.
32.
Europaparlamentet välkomnar och uppmuntrar dessutom till att internrevisionstjänsten fungerar som ordförande för byråernas nätverk Audinet, som möts två eller tre gånger per år för att samordna internrevisionsfunktionens arbete och utbyta erfarenheter om uppläggning, metoder och bästa praxis för revisioner.
Pilotrevision för etiska frågor
33.
IV.
REVISIONSFÖRKLARING OCH ÅRLIG VERKSAMHETSRAPPORT
Revisionsförklaring
34.
Europaparlamentet uppmuntrar byråerna att offentliggöra sina direktörers revisionsförklaringar på sina webbplatser och att bifoga dem som bilagor till de årliga verksamhetsrapporterna för att bekräfta att informationen i dessa årliga verksamhetsrapporter ger en sann och rättvisande bild, om ej annat anges i reservationer i samband med särskilda inkomst- och utgiftsområden.
35.
Europaparlamentet understryker att byrådirektörerna är skyldiga att ange eventuella reservationer i sina revisionsförklaringar om revisionsrätten eller kommissionens internrevisionstjänst konstaterat allvarliga problem (dvs. kritiska revisionsrekommendationer om underliggande brister och i de fall då väsentlighetströskeln har överskridits).
Årliga verksamhetsrapporter
36.
37.
Europaparlamentet gratulerar även Europeiska centrumet för förebyggande och kontroll av sjukdomar och återigen Europeiska miljöbyrån till att i sina årliga verksamhetsrapporter ha använt lättlästa tabeller eller diagram som sammanfattar de viktigaste resultaten som uppnåtts.
38.
Europaparlamentet uppmanar revisionsrätten att inkludera en översiktlig utvärdering av respektive årlig verksamhetsrapport i sina särskilda årsrapporter om byråerna på samma sätt som redan sker i årsrapporten om kommissionen, där revisionsrätten granskar de årliga verksamhetsrapporterna från kommissionens olika generaldirektorat.
V.
BYRÅERNAS LEDNING OCH FÖRVALTNING
Byråernas styrelser
39.
40.
Europaparlamentet uppmanar dessutom byråernas direktörer att vidta åtgärder för att förstärka sina styrelsers roll genom att ta upp strategiska frågor och prioriteringar till diskussion i tillräckligt god tid för att strategiska beslut ska kunna fattas.
41.
Parlamentet uppmanar byråernas styrelser att uppnå största möjliga konvergens mellan planering av uppgifter och resurser (både ekonomiska och mänskliga) genom förbättring av sin verksamhetsbaserade budgetering och förvaltning.
Kommissionens roll
42.
43.
Disciplinära förfaranden
44.
VI.
VERKSAMHETSRESULTAT
45.
46.
Europaparlamentet konstaterar att resultat och effektivitet inte mäts på ett enhetligt sätt och uppmanar den interinstitutionella arbetsgruppen för byråerna att ta itu med detta problem.
47.
Flerårigt arbetsprogram
48.
Årligt arbetsprogram
49.
50.
Feedbackförfaranden
51.
52.
Parlamentet anser att detta är ett värdefullt verktyg som även andra byråer bör använda för att hantera sina utmaningar.
53.
Europaparlamentet anser dessutom att det är ytterst viktigt att byråerna vidareutvecklar sina system för resultatövervakning för att se till att resultaten av deras verksamhet följs upp och uppmuntrar byråerna att hänvisa till dessa i sina årliga verksamhetsplaner.
54.
Europaparlamentet uppmuntrar dessutom byråerna att regelbundet rapportera om de centrala resultatindikatorerna.
Tabell som bifogas till revisionsrättens rapport
55.
Europaparlamentet gratulerar Europeiska centrumet för kontroll av narkotika och narkotikamissbruk, Översättningscentrum för Europeiska unionens organ samt Europeiska myndigheten för livsmedelssäkerhet till att i en tabell som bifogats till revisionsrättens särskilda rapport för 2009 ha gjort en jämförelse mellan de verksamheter som genomfördes under 2008 och 2009 för att göra det möjligt för den myndighet som beviljar ansvarsfrihet att lättare bedöma deras resultat från år till år.
VII.
ÖVERVÄGANDEN OM BYRÅERNA: EN GEMENSAM STRATEGI
56.
57.
Europaparlamentet påminner om att den interinstitutionella arbetsgruppen för byråerna genom sitt gemensamma uttalande i mars 2009 inledde en ’dialog om tillsynsmyndigheter för att göra en lägesbedömning, särskilt vad gäller dessa myndigheters samstämmighet, effektivitet och ansvar samt insynen i deras arbete’ samt att arbetsgruppen skulle ’behandla en rad viktiga frågor som de deltagande institutionerna föreslagit, inklusive tillsynsmyndigheternas roll och ställning i EU:s institutionella system, inrättandet av, strukturer för och driften av dessa myndigheter samt frågor som rör finansiering, budget, övervakning och förvaltning’.
58.
Europaparlamentet påminner om att man i sin resolution av den 5 maj 2010 om ansvarsfrihet för 2008 uppmanade den interinstitutionella arbetsgruppen att ’överväga möjligheten att närmare knyta samman eller till och med slå samman vissa byråer’ samt konstaterade att ’de små byråerna [...] brottas med allvarliga effektivitetsbrister’.
59.
Europaparlamentet anser att man bör införa ett moratorium mot inrättande av ytterligare byråer, åtminstone tills man funnit en tillfredsställande lösning på de frågor som framfördes i det gemensamma uttalandet från den interinstitutionella arbetsgruppen för byråerna samt i resolutionen av den 5 maj 2010.
60.
Europaparlamentet anser att man när dessa frågor är lösta bör iaktta största försiktighet när det gäller att inrätta ytterligare byråer och försäkra sig om att dessa verkligen behövs och ger bästa valuta för pengarna för att nå ett överenskommet politiskt mål.
61.
Europaparlamentet framhåller åter vikten av att överväga om vissa byråer kan slås samman, så att dessa kan dela på omkostnader och andra kostnader.
62.
Europaparlamentet uppmanar den interinstitutionella arbetsgruppen för byråerna att överväga om vissa av de mindre byråer som inte lämpar sig för en regelrätt sammanslagning i stället kan grupperas i samma stad och om möjligt i samma byggnad, så att de kan dra nytta av gemensamma centrala resurser och minimera bördan av omkostnader och andra kostnader.
63.
Europaparlamentet välkomnar revisionsrättens planer på att hösten 2011 offentliggöra en särskild rapport om kostnadsriktmärkning för unionens byråer.
64.
65.
Europaparlamentet erinrar om att unionens budget ska bygga på solid ekonomisk förvaltning, vilket kräver att utgifterna är relevanta, effektiva och ändamålsenliga samt att onödiga utgifter åtgärdas på lämpligt sätt.
66.
Europaparlamentet uppmanar därför kommissionen att göra en utvärdering av alla unionens byråer i syfte att upptäcka förekomst av överlappande verksamheter, och i de fall överlappningar konstateras undersöka möjligheten att slå samman de berörda byråerna samt lämna en rapport om detta till parlamentet senast den 31 december 2011.
VIII.
ALLMÄNNA ÖVERVÄGANDEN OM ÖKNINGEN AV ANTALET INRÄTTADE GEMENSAMMA FÖRETAG
67.
68.
Europaparlamentet välkomnar dock det faktum att internrevisionstjänsten har för avsikt att utöva denna funktion som internrevisor för de gemensamma företagen från och med budgetåret 2011.
69.
Europaparlamentet anser att de gemensamma företagen, med hänsyn till omfattningen av deras budget och deras komplexa uppgifter, bör inrätta en revisionskommitté som rapporterar direkt till styrelsen.
o
o o
70.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till de byråer som omfattas av detta förfarande för beviljande av ansvarsfrihet samt till rådet, kommissionen och revisionsrätten.
P7_TA-PROV(2011)0227
Den årliga rapporten från rådet till Europaparlamentet om de viktigaste aspekterna och de grundläggande vägvalen när det gäller den gemensamma utrikes- och säkerhetspolitiken (Gusp) 2009, som läggs fram inför Europaparlamentet i enlighet med del II, avsnitt G, punkt 43 i det interinstitutionella avtalet av den 17 maj 2006
A7-0168/2011
Europaparlamentets resolution av den 11 maj 2011 om rådets årliga rapport till Europaparlamentet om de viktigaste aspekterna och de grundläggande vägvalen när det gäller den gemensamma utrikes- och säkerhetspolitiken (Gusp) – 2009, som läggs fram för parlamentet i enlighet med del II punkt G.43 i det interinstitutionella avtalet av den 17 maj 2006 ( 2010/2124(INI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av rådets årliga rapport till Europaparlamentet om de viktigaste aspekterna och de grundläggande vägvalen när det gäller den gemensamma utrikes- och säkerhetspolitiken (Gusp) – 2009, som läggs fram för parlamentet i enlighet med del II punkt G.43 i det interinstitutionella avtalet av den 17 maj 2006 EUT C 139, 14.6.2006, s.
1.
,
–
med beaktande av det ovannämnda interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning,
–
med beaktande av sina resolutioner av den 19 februari 2009 EUT C 76 E, 25.3.2010, s.
54.
och den 10 mars 2010 EUT C 349 E, 22.12.2010, s.
51.
om rådets årliga rapport om Gusp 2007 respektive 2008,
–
med beaktande av sin resolution av den 8 juli 2010 om den europeiska avdelningen för yttre åtgärder Antagna texter, P7_TA(2010)0280 .
,
–
med beaktande av sin resolution av den 11 november 2010 om stärkandet av OSSE: en roll för EU Antagna texter, P7_TA(2010)0399 .
,
–
med beaktande av förklaringen av vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik om politisk ansvarighet Ibid., bilaga II.
,
–
med beaktande av den höga representantens uttalande vid Europaparlamentets plenarsammanträde den 8 juli 2010 om hur den centrala förvaltningen av den europeiska avdelningen för yttre åtgärder ska organiseras i stort Antagna texter, P7_TA(2010)0280 , bilagan.
,
–
med beaktande av slutsatserna från Europeiska rådets möte den 16 september 2010 om EU:s yttre förbindelser,
–
–
med beaktande av betänkandet från utskottet för utrikesfrågor och yttrandet från budgetutskottet ( A7-0168/2011 ), och av följande skäl:
A.
EU bör utveckla sina utrikespolitiska mål ytterligare och främja sina värderingar och intressen i världen med det övergripande målet att bidra till fred, säkerhet, solidaritet, konfliktförebyggande, främjande av demokrati, skydd för de mänskliga rättigheterna, jämställdhet mellan kvinnor och män, respekt för internationell rätt, stöd för internationella institutioner, effektiv multilateralism och ömsesidig respekt mellan folken, hållbar utveckling, fri och rättvis handel samt utrotning av fattigdomen.
B.
Genomförandet av Lissabonfördraget tillför en ny dimension till EU:s yttre åtgärder och kommer att bidra till att göra unionens utrikespolitik och – i vidare mening EU:s yttre åtgärder – enhetligare, konsekventare och effektivare.
C.
Lissabonfördraget ger EU:s utrikespolitik en ny dynamik, särskilt genom att förse unionen med institutionella och operativa verktyg som kan göra det möjligt för den att spela en internationell roll som är förenlig med dess framträdande ekonomiska ställning och dess ambitioner samt att organisera sig för att bli en effektiv global aktör som kan ta medansvar för den globala säkerheten och leda arbetet för att ta fram gemensamma svar på gemensamma utmaningar.
D.
E.
Världsordningen genomgår för närvarande en stor omvandling, och det har uppkommit nya utmaningar och nya maktstrukturer som innebär att EU måste samarbeta mer aktivt med nuvarande och blivande makter och icke-statliga aktörer och med bilaterala och multilaterala partner och institutioner för att främja effektiva lösningar på problem som är gemensamma för medborgare i EU och i hela världen och som kan påverka den globala säkerheten.
F.
G.
Rådets årliga rapport om Gusp 2009
1.
2.
3.
Europaparlamentet anser att den årliga rapporten om Gusp bör grunda sig på den nya institutionella ram som skapats genom Lissabonfördraget och tjäna som ett instrument för utökad interinstitutionell dialog, där man framför allt diskuterar genomförandet av EU:s utrikespolitiska strategi, utvärderar hur effektiv den är och anger vilken väg man bör slå in på i framtiden.
Genomförandet av Lissabonfördraget
4.
Vice ordföranden/den höga representanten uppmanas att använda sina befogenheter fullt ut för att initiera och genomföra den gemensamma utrikes- och säkerhetspolitiken och se till att den följs och att parlamentets berörda organ blir fullt delaktiga i detta arbete.
5.
6.
7.
8.
9.
10.
11.
12.
13.
14.
15.
16.
Europaparlamentet understryker att en grundlig analys behöver genomföras om de långsiktiga finansiella behoven för Gusp i samband med de kommande diskussionerna om den fleråriga budgetramen 2014–2020.
17.
Vice ordföranden/den höga representanten förväntas lämna all relevant information om förhandlingarna under hela förfarandet, däribland förhandlingsdirektiv och utkast till förhandlingstexter.
18.
Tematiska huvudfrågor för Gusp
19.
20.
Europaparlamentet uppmanar vice ordföranden/den höga representanten, rådet och medlemsstaterna att motverka obalansen mellan Europeiska utrikestjänstens civila respektive militära planeringskapacitet och att öka personalen på områdena rättsliga frågor, civil förvaltning, tull och medling för att se till att GSFP-uppdragen har adekvat och tillräcklig expertis.
21.
22.
Europaparlamentet anser att det är en strategisk prioritering för EU att stärka internationella partnerskap för krishantering och fördjupa dialogen med andra viktiga aktörer för krishantering – som FN, Nato, Afrikanska unionen (AU), OSSE och tredjeländer som Förenta staterna, Turkiet, Norge och Kanada – och att samordna åtgärder, utbyta information och förena resurser för fredsbevarande och fredsbyggande, däribland samarbete om krishantering och särskilt sjöfartssäkerhet, samt kampen mot terrorism i enlighet med internationell rätt.
23.
24.
25.
26.
27.
28.
29.
Med tanke på att klimatförändringarna har blivit en viktig del av de internationella förbindelserna upprepar Europaparlamentet att EU måste stärka sitt ledarskap inom den globala klimatpolitiken och även inleda en dialog med andra huvudaktörer såsom tillväxtmakterna (Kina, Brasilien, Indien), Ryssland, Förenta staterna och utvecklingsländerna.
30.
31.
32.
Geografiska huvudprioriteringar för Gusp
Multilateral diplomati, internationella organisationer
33.
34.
Frankrike och Storbritannien uppmanas att, i egenskap av ständiga medlemmar i FN:s säkerhetsråd och i enlighet med artikel 34.2 i EU-fördraget, alltid begära att vice ordföranden/den höga representanten bjuds in för att representera EU när EU har tagit ställning i en fråga som finns på säkerhetsrådets dagordning.
EU bör vara representerat som union i de multilaterala finansiella organen, särskilt Internationella valutafonden och Världsbanken, utan att detta påverkar medlemsstaternas representation.
35.
36.
37.
38.
De transatlantiska förbindelserna
39.
40.
Västra Balkan
41.
42.
43.
44.
45.
46.
Det östliga partnerskapet
47.
48.
Europaparlamentet hoppas att den reform av den europeiska grannskapspolitiken som kommissionen har inlett kommer att leda till en ny strategisk vision och en differentierad strategi inom samma politik när det gäller intresseområdena, i enlighet med unionens olika intressen, utmaningar och regionala hot.
49.
50.
51.
52.
53.
Europaparlamentet understryker vikten av att EU spelar en mer aktiv roll i att lösa de låsta konflikterna i Transnistrien och Sydkaukasien.
54.
Europaparlamentet välkomnar och stöder de moldaviska myndigheternas engagemang för att stärka förbindelserna med Europeiska unionen när det gäller arbetet med att ingå associeringsavtalet, utveckla en dialog om liberalisering av viseringsbestämmelserna och inleda förhandlingar om ett frihandelsavtal.
Europeiska unionens strategi för Svarta havet
55.
Europaparlamentet uppmanar kommissionen att påskynda genomförandet av projekten inom Svartahavssynergin och att låta denna fråga stå kvar på Europeiska utrikestjänstens dagordning.
56.
Europaparlamentet understryker Svartahavsområdets betydelse inom det östliga partnerskapet och anser att Europeiska unionen måste visa ett större engagemang i detta sammanhang.
Centralasien
57.
Ryssland
58.
59.
60.
Turkiet
61.
Parlamentet välkomnar uttalandet från rådet av den 14 december 2010 där man efterlyste ett ökat samarbete i säkerhets- och utrikespolitiska frågor av gemensamt intresse.
Turkiets allt aktivare utrikespolitik innebär nya utmaningar och möjligheter för Gusp.
Vice ordföranden/den höga representanten uppmanas att inbegripa Turkiet i en institutionaliserad dialog om viktiga strategiska frågor, till exempel energipolitik, stabilitet i västra Balkan och Kaukasien, Irans kärnenergiprogram eller det demokratiska uppvaknande som är på gång i Mellanöstern.
På så sätt kan man se till att målen blir enhetligare och ge ny dynamik åt de bilaterala förbindelserna.
Parlamentet understryker emellertid att en sådan dialog inte får ersätta Turkiets anslutningsprocess, utan måste komplettera och stärka den.
62.
Parlamentet varnar för att det kan uppstå allvarliga problem på lång sikt om förhållandet mellan EU och Turkiet inte stabiliseras och EU och Nato även fortsättningsvis hindras från att uppnå målet om närmare samarbete.
Mellanöstern och Medelhavsområdet
63.
64.
65.
66.
67.
Europaparlamentet erinrar om sin roll i EU:s budgetförfarande och framhåller vikten av att UfM:s demokratiska legitimitet garanteras, att beslut fattas på ett öppet sätt och att Europaparlamentet, UfM:s parlamentariska församling och de nationella parlamenten blir delaktiga i beslutsprocessen.
68.
69.
70.
71.
72.
Asien
73.
74.
75.
76.
77.
78.
79.
80.
Afrika
81.
82.
Europaparlamentet uttrycket sitt stöd för beslutet att ta fram en övergripande EU-strategi för Afrikas horn, genom att bidra till återuppbyggnad av statliga institutioner i Somalia och förena mänsklig säkerhet med utveckling, rättsstatsprincipen, respekt för de mänskliga rättigheterna och kvinnors rättigheter och därvid inbegripa alla EU-instrument för att skapa långsiktiga lösningar.
83.
84.
85.
86.
87.
Latinamerika
88.
89.
o
o o
90.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik, rådet, kommissionen, EU-medlemsstaternas regeringar och parlament, FN:s generalsekreterare, Natos generalsekreterare, talmannen i Natos parlamentariska församling, OSSE:s tjänstgörande ordförande, talmannen i OSSE:s parlamentariska församling, ordföranden för Europarådets ministerkommitté och talmannen i Europarådets parlamentariska församling.
P7_TA-PROV(2011)0256
EU:s sjunde ramprogram för forskning, teknisk utveckling och demostration
A7-0160/2011
Europaparlamentets resolution av den 8 juni 2011 om den preliminära utvärderingen av Europeiska unionens sjunde ramprogram för verksamhet inom området forskning, teknisk utveckling och demonstration ( 2011/2043(INI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av fördraget om Europeiska unionen (EU-fördraget) och fördraget om Europeiska unionens funktionssätt (EUF-fördraget), i synnerhet artiklarna om forskning,
–
med beaktande av Europaparlamentets och rådets beslut nr 1982/2006/EG av den 18 december 2006 om Europeiska gemenskapens (efter Lissabonfördragets ikraftträdande Europeiska unionens) sjunde ramprogram för verksamhet inom området forskning, teknisk utveckling och demonstration (2007–2013) EUT L 412, 30.12.2006, s.
1.
,
–
med beaktande av framför allt artikel 7 i nämnda beslut avseende övervakning, utvärdering och översyn av sjunde ramprogrammet,
–
–
med beaktande av kommissionens meddelande av den 9 februari 2011 med titeln ”Meddelande från kommissionen till Europaparlamentet, rådet, Europeiska ekonomiska och sociala kommittén och Regionkommittén – Svar på rapporten från expertgruppen för preliminär utvärdering av sjunde ramprogrammet för forskning, teknisk utveckling och demonstration och rapporten från expertgruppen för preliminär utvärdering av finansieringsinstrumentet för riskdelning” ( KOM(2011)0052 ),
–
med beaktande av slutsatserna från den preliminära utvärderingen av sjunde ramprogrammet för forskning, inbegripet finansieringsmekanismen för delade risker från rådets (konkurrenskraft) (inre marknaden, industri, forskning och rymdfrågor) 3074:e möte den 9 mars 2011,
–
med beaktande av expertgruppens slutrapport ”Interim Evaluation of the Seventh Framework Programme” av den 12 november 2010,
–
med beaktande av sin resolution av den 11 november 2010 om förenklat genomförande av ramprogrammen för forskning Antagna texter, P7_TA(2010)0401 .
,
–
med beaktande av expertgruppens rapport ”Evaluation of the Sixth Framework Programmes for Research and Technological Development 2002–2006” från februari 2009,
–
med beaktande av expertgruppens rapport ”Towards a world class Frontier research Organisation – Review of the European Research Council's Structures and Mechanisms” av den 23 juli 2009,
–
med beaktande av den oberoende expertgruppens rapport ”Mid-Term Evaluation of the Risk-Sharing Financial Facility (RSFF)” av den 31 juli 2010,
–
med beaktande av expertgruppens rapport ”First Interim Evaluation of the Innovative Medicines Initiative Joint Undertaking” av den 20 december 2010,
–
med beaktande av expertgruppens rapport ”First Interim Evaluation of the ARTEMIS and ENIAC Joint Technology Initiatives” av den 30 juli 2010,
–
med beaktande av den oberoende expertgruppens rapport ”Interim Evaluation of the Ambient Assisted Living Joint Programme” från december 2010,
–
med beaktande av Regionkommitténs yttrande som antogs vid plenarsessionen den 27–28 januari 2011 om förenklat genomförande av ramprogrammen för forskning,
–
med beaktande av Europaparlamentets resolution av den 20 maj 2010 om hur synergieffekterna av medel öronmärkta för forskning och innovation enligt förordning (EG) nr 1080/2006 avseende Europeiska utvecklingsfonden och sjunde ramprogrammet för forskning och utveckling har utnyttjats i städer och regioner såväl som i medlemsstaterna och unionen Antagna texter, P7_TA(2010)0189 .
,
–
med beaktande av Europeiska revisionsrättens särskilda rapport nr 9/2007 av den 22 november 2007 med titeln ”Utvärderingen av EU:s ramprogram för forskning, teknisk utveckling och demonstration (FoTU) – skulle kommissionens tillvägagångssätt kunna förbättras?”,
–
med beaktande av Europeiska revisionsrättens särskilda rapport nr 8/2009 med titeln ”Expertnätverk och integrerade projekt i gemenskapens forskningspolitik – uppnåddes målen?”,
–
med beaktande av Europeiska revisionsrättens särskilda rapport nr 2/2010 med titeln ”Har stödsystemen för förberedande studier och uppbyggnad av ny infrastruktur inom det sjätte ramprogrammet för forskning varit ändamålsenliga?”,
–
med beaktande av yttrandet från Europeiska ekonomiska och sociala kommittén av den 15 september 2010 över kommissionens meddelande till Europaparlamentet, rådet, Europeiska ekonomiska och sociala kommittén och Regionkommittén om förenklat genomförande av ramprogrammen för forskning,
–
med beaktande av artikel 48 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för industrifrågor, forskning och energi och yttrandet från budgetutskottet ( A7-0160/2011 ), och av följande skäl:
A.
Europeiska gemenskapens sjunde ramprogram för verksamhet inom området forskning, teknisk utveckling och demonstration är världens största instrument för stöd till forskning och det viktigaste verktyget i Europeiska unionens forskningspolitik.
B.
C.
I Lissabonfördraget införs fullbordandet av det europeiska området för forskningsverksamhet som ett särskilt medel i EU:s politik.
D.
I Europa 2020-strategin görs forskning och innovation till en central del av en intelligent och hållbar tillväxt för alla.
E.
Forskning är det som omvandlar ekonomisk styrka till kunskap, medan innovation omvänt omvandlar kunskap till ekonomisk styrka.
F.
G.
Investeringar i FoU är det bästa långsiktiga svaret på dagens ekonomiska och finansiella kris, eftersom de ger EU möjlighet att bli ett konkurrenskraftigt kunskapssamhälle i världsklass.
H.
I.
Det är också uppenbart att det utöver de investerade beloppen även behövs en bättre samordning och samfinansiering mellan unionen, medlemsstaterna och regionerna, med full respekt för medlemsstaternas specifika egenskaper och etiska villkor.
J.
Endast tämligen små offentliga investeringar i FoU är föremål för europeiskt samarbete.
K.
Förbindelserna mellan den akademiska världen, forskningen och industrin måste förbättras för att forskningsresultat bättre ska kunna omvandlas till produkter och tjänster som genererar ekonomisk tillväxt och fördelar för samhället i stort.
L.
M.
N.
Åren 2011–2013 är kritiska år, och vi kommer särskilt att behöva uppmärksamma faktorer som konkurrenskraft och social sammanhållning, där forskning och innovation är avgörande inslag.
O.
En komplicerad administrativ förvaltning, omfattande pappersexercis, byråkrati, bristande insyn, ineffektivitet och omotiverade förseningar utgör fortfarande stora hinder för sjunde ramprogrammet och avskräcker forskare, industri och små och stora företag från att delta i programmet.
En av de största prioriteringarna i programmet bör därför vara att ta ett stort steg mot förenkling.
P.
Målet på 40 procent kvinnliga forskare i sjunde ramprogrammet är ambitiöst och riktigt.
1.
Europaparlamentet välkomnar den höga kvaliteten på expertgruppens rapporter om den preliminära utvärderingen av sjunde ramprogrammet samt finansieringsmekanismen med delad risk, som avser insatsernas kvalitet, genomförande och noterade resultat, trots det allmänna mandat som gruppen tilldelades.
Parlamentet påpekar dock att man i utvärderingen inte beaktar medlemsstaternas och EU:s åtgärder i deras helhet.
2.
3.
Europaparlamentet uppmanar kommissionen att särskilt följa upp expertgruppens tio specifika rekommendationer.
4.
Europaparlamentet betonar att slutsatserna från den preliminära översynen är relativa, eftersom huvuddelen av anslagen inom sjunde ramprogrammet ännu inte har tilldelats.
Sjunde ramprogrammets resultat
5.
Europaparlamentet anser att Europa visserligen fortfarande ligger efter Förenta staterna och håller på att tappa försprånget till tillväxtländerna, men att de resultat som uppnåtts i sjunde ramprogrammet tycks påvisa ett europeiskt mervärde när det gäller FoU.
Parlamentet uppmanar kommissionen att öka ansträngningarna för att kommunicera de framgångsrika resultaten till medlemsstaterna, forskarsamfundet och de europeiska medborgarna.
6.
7.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att förstärka kommunikationsarbetet om sjunde ramprogrammet (bland annat genom att använda ny teknik som smarta forskningsinformationstjänster) och att underlätta tillgången till information om deltagande, tillkännage kommande forskningsutmaningar och sprida forskningsrön.
Parlamentet stöder kommissionens initiativ att främja öppen tillgång till resultat från offentligt finansierad forskning, om detta är lämpligt och möjligt med hänsyn till immateriella rättigheter.
8.
9.
10.
11.
12.
13.
14.
15.
Europaparlamentet stöder inom ramen för programdelen ”Människor” de Marie Curie-åtgärder som är så värdefulla för forskares karriärer, säkerställer individuell forskning ”nerifrån och upp” inom många olika ämnen, hindrar kompetensflykt och gör en forskarkarriär mer lockande för unga lovande forskare både från EU och från tredjeländer.
16.
17.
18.
19.
Europaparlamentet uppmanar kommissionen att ge parlamentet tydlig och detaljerad information om hur de gemensamma teknikinitiativen fungerar och för varje enskilt fall lämna uppgifter om juridisk status, vilka personer som ingår i rådet och vilken verksamhet som har bedrivits.
20.
21.
22.
Dessutom måste kommissionens samordnande roll stärkas och medlemsstaterna bör respektera sina ekonomiska åtaganden.
23.
24.
Europaparlamentet betonar betydelsen av Gemensamma forskningscentrets direkta insatser och dess bidrag till en hållbar utveckling, konkurrenskraft, säkerhet och kärnkraftssäkerhet.
25.
26.
27.
28.
29.
Europaparlamentet anser att förfarandena för konkurrerande ansökningar för övriga partner bör bygga på grundförutsättningen att de inblandade företagen och forskarna har de mest ingående kunskaperna om projektet och vilken typ av partner som behövs, och att kommissionen inte ska tvinga dem att följa utvärderingsexperternas rankningslistor utan i stället utvärdera en skriftlig motivering av konsortiets val.
30.
Europaparlamentet välkomnar sjunde ramprogrammets resultat till förmån för små och medelstora företag, både när det gäller stödåtgärderna för små och medelstora företag i programdelen ”Kapacitet”, programmet ”Eurostars” och det mål på 15 procent som fastställts i programdelen ”Samarbete”.
31.
32.
Europaparlamentet noterar med oro vissa medlemsstaters relativt låga deltagande i sjunde ramprogrammet, vilket inte bidrar till den territoriella sammanhållningen eller till en balanserad utveckling i EU.
Parlamentet anser att en bättre samordning, enhetlighet och synergi mellan sjunde ramprogrammet och struktur- och sammanhållningsfonderna samt ett bättre utnyttjande av programdelen ”Människor” skulle kunna förbättra de underrepresenterade medlemsstaternas deltagande.
33.
Europaparlamentet välkomnar de stadiga men blygsamma framstegen mot ett jämnare deltagande av både män och kvinnor i ramprogrammet, eftersom mångfald är viktigt för kreativitet och innovation.
34.
Europaparlamentet anser att man på regional nivå bör erkänna den särskilda roll som intresseorganisationer (t.ex. handelskamrarna, nätverket Enterprise Europe Network och regionala innovationsbyråer) har som länk mellan lokala, innovativa små och medelstora företag och kommissionen.
35.
36.
Finansiering
37.
38.
39.
Europaparlamentet betonar den avgörande roll som forskningsinfrastrukturen spelar för kunskapstriangeln och understryker att utvecklingen och finansieringen av denna infrastruktur (på grundval av Esfris lista tillhandahållande av laboratorieutrustning och instrument samt underhåll av dessa) bör främjas genom bättre samordning och samfinansiering mellan sjunde ramprogrammet, Europeiska investeringsbankens instrument, strukturfonderna samt nationell och regional politik.
Parlamentet anser att man bör undvika förekomsten av flera forskningsinfrastrukturer i olika medlemsstater samt gynna en öppen och kompetensbaserad tillgång till forskningsinfrastruktur.
Parlamentet efterlyser insatser för att öka finansieringen av forskningsinfrastruktur inom sjunde ramprogrammet, i synnerhet där de största möjligheterna till ett europeiskt mervärde finns.
40.
41.
Europaparlamentet uppmanar EU och dess medlemsstater att respektera sina ekonomiska åtaganden, inklusive åtagandena om de insatser som följer av artiklarna 185 och 187, inom ramen för internationella forskningsavtal.
42.
Mot bakgrund av målet att tre procent av BNP ska investeras i forskning och teknisk utveckling senast 2020 och med hänsyn till att forskning och innovation är den enda säkra vägen till ekonomisk återhämtning i EU, uppmanar Europaparlamentet kommissionen att överväga möjligheten att fastställa en mellanliggande, bindande lägstanivå för investeringarna i forskning och teknisk utveckling på cirka en procent av BNP senast 2015.
Innovationsfunktionen
43.
Parlamentet uppmanar kommissionen att innan sjunde ramprogrammet löper ut börja finansiera demonstrations- och pilotprojekt samt koncepttest och att överväga ett finansieringssystem som belönar framgångsrika projekt och ser till att de förs in på marknaden, som ett komplement till dagens förskottsfinansiering.
I detta avseende anser parlamentet också att det behövs nära samordning mellan sjunde ramprogrammet, ramprogrammet för konkurrenskraft och innovation och strukturfonderna.
44.
45.
46.
47.
Uppföljningen av förenklingsåtgärder
48.
Europaparlamentet är bekymrat över den alltför stora administrativa börda som är förknippad med sjunde ramprogrammet.
49.
Europaparlamentet upprepar hur viktigt det är att utan dröjsmål införa förenklingsåtgärder för förfarandena, administrationen och finansieringen i den nuvarande förvaltningen av sjunde ramprogrammet, såsom de åtgärder som togs upp i parlamentets resolution av den 11 november 2010.
50.
Europaparlamentet kräver åtgärder för att minska handläggningstiden i syfte att öka antalet anslag som beviljas inom mindre än åtta månader med en viss procentenhet under 2011, och inom mindre än sex månader under den återstående programperioden.
51.
Europaparlamentet välkomnar rekommendationerna om att minska handläggningstiden och kräver en utvärdering av redan befintliga instrument innan nya upprättas inom ramen för sjunde ramprogrammet.
52.
Europaparlamentet föreslår att kommissionen hjälper de offentliga organen att förbättra sina förvaltningssystem genom att göra utvärderingar utan ekonomiska konsekvenser för att uppmuntra dessa organ att vidta en rad åtgärder som förbättrar deras projektförvaltning och genomföra dem inom en tidsfrist som är kortare än ett år.
Finansieringsinstrumentet för riskdelning
53.
Europaparlamentet anser att finansieringsinstrumentet för riskdelning har haft en avgörande kvalitativ och kvantitativ hävstångseffekt för att öka investeringarna i forskning, utveckling och innovation under krisen då banksektorn inte längre kunde fylla den funktionen, med en slutgiltig utlåning under de första åren på 8 miljarder euro som genererat mer än 20 miljarder euro i investeringar.
54.
55.
56.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att undersöka publiciteten kring tillgången till lån från finansieringsinstrumentet för riskdelning på medlemsstatsnivå och se till att potentiella deltagare får den information och hjälp de behöver för att få tillgång till lån från instrumentet, i synnerhet i de medlemsstater vars valuta inte är euro.
57.
Parlamentet betonar vikten av att se till att dessa finansieringsinstrument är utformade på ett sätt som passar små och medelstora företag.
Övergripande slutsats och framtida inriktning
58.
Parlamentet anser framför allt att sjunde ramprogrammets mål ska anpassas till EU:s strategier för resurseffektivitet, råvaror och den digitala agendan.
59.
60.
61.
Europaparlamentet betonar att det är viktigt att ta hänsyn till bedömningen av de resultat som uppnåtts på vart och ett av de områden som politiskt har prioriterats för finansiering, och till hur effektiva de varit, med målet att förbättra utvärderingen av framtida program.
o
o o
62.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet och kommissionen samt till medlemsstaterna.
P7_TA-PROV(2011)0330
Kvinnor och företagsledarskap
A7-0210/2011
Europaparlamentets resolution av den 6 juli 2011 om kvinnor och företagsledarskap ( 2010/2115(INI) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av den fjärde internationella kvinnokonferensen som hölls i Peking i september 1995, den förklaring och den handlingsplan som antogs i Peking samt de slutdokument som blev resultatet och som antogs vid FN:s särskilda sessioner Peking +5, Peking +10 och Peking +15 om ytterligare åtgärder och initiativ för att genomföra Pekingförklaringen och handlingsplanen, vilka antogs den 9 juni 2000, den 11 mars 2005 respektive den 12 mars 2010,
–
med beaktande av FN:s konvention från 1979 om avskaffande av all slags diskriminering av kvinnor,
–
med beaktande av den allmänna förklaringen om de mänskliga rättigheterna från 1948,
–
med beaktande av Europeiska unionens stadga om de grundläggande rättigheterna, särskilt artiklarna 1, 2, 3, 4, 5, 21 och 23,
–
med beaktande av artikel 2 i fördraget om Europeiska unionen, där värden som är gemensamma för medlemsstaterna betonas såsom mångfald, icke-diskriminering, tolerans, rättvisa, solidaritet och principen om jämställdhet mellan kvinnor och män,
–
med beaktande av artikel 19 i fördraget om Europeiska unionens funktionssätt, enligt vilken diskriminering på grund av kön ska bekämpas,
–
med beaktande av kommissionens rapport om utvecklingen av jämställdheten mellan kvinnor och män 2011,
–
–
med beaktande av kommissionens meddelande av den 21 september 2010, ”Strategi för jämställdhet 2010–2015” ( KOM(2010)0491 ),
–
med beaktande av kommissionens grönbok av den 6 juni 2010 om företagsstyrning i finansiella institut och om ersättningspolicy ( KOM(2010)0284 ),
–
med beaktade av kommissionens meddelande av den 5 mars 2010, ”Ett förstärkt engagemang för jämställdhet – Kvinnostadga” ( KOM(2010)0078 ),
–
med beaktande av den europeiska pakten för jämställdhet som antogs av Europeiska rådet i mars 2006, och den nya europeiska pakten för jämställdhet mellan kvinnor och män som antogs av rådet den 7 mars 2011,
–
med beaktande av rådets rekommendation 96/694/EG om en balanserad fördelning mellan kvinnor och män i beslutsprocessen,
–
med beaktande av det årliga mötet för Världsekonomiskt forum i Davos den 26-29 januari 2011 och programmet ”Women Leaders and Gender Parity”,
–
med beaktande av sin resolution av den 11 maj 2011 om bolagsstyrning i finansinstitut Antagna texter, P7_TA(2011)0223 .
,
–
med beaktande av sin resolution av den 8 mars 2011 om jämställdhet mellan kvinnor och män i Europeiska unionen – 2010 Antagna texter, P7_TA(2011)0085 .
,
–
med beaktande av sina resolutioner av den 15 juni 1995 om FN:s fjärde internationella kvinnokonferens i Peking: Jämställdhet, utveckling och fred EGT C 166, 3.7.1995, s.
92.
, av den 10 mars 2005 om uppföljningen av handlingsprogrammet från FN:s fjärde internationella kvinnokonferens (Peking + 10) EUT C 320E, 15.12.2005, s.
247.
och av den 25 februari 2010 om Peking + 15 – FN:s handlingsplan för jämställdhet EUT C 348E, 21.12.2010, s.
11.
,
–
med beaktande av artikel 48 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män ( A7-0210/2011 ), och av följande skäl:
A.
B.
Ett av EU:s viktigaste mål borde vara att undanröja de hinder och den ojämlikhet mellan könen som kvarstår och som motverkar kvinnors framsteg i karriären, så att det blir möjligt för kompetenta och kvalificerade kvinnor att få tillträde till befattningar som de i dag har svårt att nå.
C.
Jämställdhet i arbetet bör främja att ingen åtskillnad görs mellan män och kvinnor på arbetsmarknaden generellt och i fråga om befordringar till ledande befattningar på alla nivåer, för att uppnå en social rättvisa och utnyttja kvinnors kompetens fullt ut och därmed stärka ekonomin genom att kvinnor garanteras samma möjlighet att utvecklas som män.
D.
Kvinnors representation hindras även av en kombination av faktorer såsom kvardröjande könsdiskriminering, stereotypa beteenden som lever kvar i förtagen och begränsade möjligheter att få en mentor för en eventuell framtida chefskarriär.
E.
F.
G.
Därför är det viktigt att införa metoder som fallstudier och utbyte av god praxis på området samt positiv särbehandling för att uppnå ett optimalt utnyttjande av kvinnlig arbetskraft på alla nivåer i företagens verksamhet.
H.
I.
J.
K.
L.
M.
Kommissionen har meddelat att den ska lägga fram lagstiftningsåtgärder som ska se till att de börsnoterade företagen vidtar effektiva åtgärder för att uppnå en jämn fördelning mellan kvinnor och män i styrelserna, och i de fall självregleringen inte fungerar, se till att detta sker inom de följande 12 månaderna.
1.
Europaparlamentet välkomnar de åtgärder som kommissionen aviserade den 1 mars 2011, särskilt kommissionens avsikt att lägga fram förslag till EU-lagstiftning 2012 om företagen inte genom frivilliga åtgärder klarar av att uppnå målen om 30 procent kvinnor i företagsstyrelserna senast 2015 och 40 procent senast 2020.
2.
Europaparlamentet uppmanar med kraft företagen att uppnå den kritiska tröskeln 30 procent kvinnor bland ledamöterna i styrande organ senast 2015 och 40 procent 2020.
3.
Europaparlamentet konstaterar en klar förbättring av kvinnornas representation i Norge efter antagandet av en lag 2003 som föreskriver att minst 40 procent av vardera kön ska vara representerat i styrelserna för börsnoterade företag med fler än 500 anställda, med effektiva sanktioner vid överträdelser.
4.
Europaparlamentet betonar att företagen måste respektera lika möjligheter och likabehandling av kvinnor och män i arbetslivet och att de i detta syfte bör vidta åtgärder för att förhindra all diskriminering.
5.
6.
7.
Europaparlamentet framhåller att rekryteringen till poster i företagens styrande organ måste bygga på den kompetens som personerna tillägnat sig i form av färdigheter, kvalifikationer och erfarenhet, och att principerna om öppenhet, objektivitet, delaktighet, effektivitet, icke-diskriminering och jämlikhet måste iakttas i företagens rekryteringspolicy.
8.
Europaparlamentet anser att man bör överväga att införa effektiva regler för att förhindra att personer upptar flera poster i styrelserna för att ställa dessa poster till kvinnornas förfogande, men även för att sträva efter effektivitet och opartiskhet bland styrelsemedlemmarna i medelstora och stora företag.
9.
Europaparlamentet understryker att de offentliga, börsnoterade företagen bör föregå med gott exempel och vara de första som tillämpar en jämn könsfördelning i ledningen och på ledande poster på alla nivåer.
10.
Europaparlamentet uppmanar medlemsstaterna och kommissionen att vidta nya politiska åtgärder för att öka andelen kvinnor i företagsledningarna, särskilt genom att
a)
inleda en dialog som skulle kunna äga rum årligen och som inte begränsar sig till frågan om kvoter, med styrelserna för stora företag och med arbetsmarknadens parter om vilka metoder som kan användas för att öka antalet kvinnor,
b)
stödja initiativ för att utvärdera och främja jämställdheten mellan kvinnor och män i rekryteringskommittéer och på områden som löneskillnader, yrkesklassificering, utbildning och karriärutveckling,
c)
främja de europeiska företagens sociala ansvar genom insatser för att garantera kvinnorna ledaransvar och familjevänliga tjänster,
d)
stödja åtgärder som uppmuntrar unga kvinnor att i högre grad välja naturvetenskapliga och tekniska studier, vilket också FN:s ekonomiska och sociala råd har krävt,
e)
införa specifika åtgärder och arrangemang för att erbjuda tjänster av hög kvalitet och till rimliga priser, t.ex. när det gäller omsorg av barn, äldre och andra omsorgsbehövande personer, skatteincitament för företagen eller annan ersättning för att göra det möjligt för de anställda i företagen att kombinera familje- och yrkesliv,
f)
utveckla enskilda kvinnors kompetens i företagen för att förbereda dem på ett effektivt sätt för utövandet av ledande funktioner genom särskild och fortlöpande utbildning samt andra stödåtgärder, såsom riktat mentorskap och nätverksstrukturer för att effektivt förbereda dem för ledarskap på alla nivåer,
g)
utveckla utbildningen om jämlikhet och icke-diskriminering,
h)
främja exakta och kvantifierbara åtaganden från företagens sida,
i)
uppmuntra alla berörda parter att utarbeta initiativ för att ändra sättet att se på kvinnor och kvinnor och kvinnors självuppfattning när det gäller arbete, så att kvinnor får möjlighet att ta ledningsansvar på företagets operativa sida och inte bara på den funktionella sidan; enligt parlamentet bör sådana initiativ syfta till att dels uppmuntra flickor och unga kvinnor att föreställa sig bredare karriärmöjligheter med stöd av lärare, familj och olika förebilder, dels förmedla kvinnligt ledarskap på ett positivt sätt i de europeiska medierna,
j)
fastställa sätt att öka andelen kvinnor från särskilt underrepresenterade grupper, såsom kvinnor med invandrarbakgrund eller etnisk minoritetsbakgrund.
11.
12.
Europaparlamentet anser i synnerhet att företag som är skyldiga att lägga fram icke förenklade resultaträkningar borde uppnå en balanserad representation av kvinnor och män i ledningen inom en rimlig tidsperiod.
13.
Europaparlamentet uppmanar företagen att anta och tillämpa företagsstyrningskoder för att främja jämställdhet mellan könen i styrelser, använda sig av grupptryck för att påverka organisationer inifrån och införa principen följ-eller-förklara, som innebär att företagen måste förklara varför det inte finns åtminstone en kvinna i styrelsen.
14.
a)
hantera problem med tillgång till ansvarsfull barnomsorg till överkomligt pris i närmiljön,
b)
15.
Europaparlamentet uppmuntrar företagsledarna att uppmärksamma sin personal på kvinnors och mäns karriärutveckling och personligen engagera sig i kvinnliga chefers uppföljnings- och karriärstödprogram på det egna företaget.
16.
Europaparlamentet uppmanar kommissionen att
a)
snarast möjligt lägga fram en aktuell lägesbeskrivning om andelen kvinnor i alla typer av företag i EU samt om de åtgärder av både tvingande och inte tvingande karaktär som näringslivet har vidtagit och de bestämmelser som nyligen antagits i de olika medlemsstaterna för att öka andelen kvinnor,
b)
mot bakgrund av slutsatserna i lägesbeskrivningen och om företagens och medlemsstaternas frivilliga åtgärder är otillräckliga, föreslå införande av kvoter senast 2012 för att öka kvinnornas andel i företagens styrande organ till 30 procent senast 2015 och till 40 procent senast 2020 med beaktande av medlemsstaternas befogenheter samt deras ekonomiska, strukturella (storleken på företagen), rättsliga och regionala särdrag.
17.
Europaparlamentet uppmanar kommissionen att upprätta en färdplan för att nå de fastställda specifika och mätbara målen för att nå fram till en balanserad representation i företagen, oavsett deras storlek och att utarbeta en särskild vägledning för små och medelstora företag.
18.
19.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen och medlemsstaternas regeringar.
P7_TA-PROV(2011)0335
Förberedelser inför valet till ryska statsduman i december 2011
B7-0396 , 0448 , 0450 , 0451 och 0452/2011
Europaparlamentets resolution av den 7 juli 2011 om förberedelserna inför valet till ryska statsduman i december 2011
Europaparlamentet utfärdar denna resolution
–
med beaktande av partnerskaps- och samarbetsavtalet mellan Europeiska unionen och Ryska federationen som trädde i kraft 1997 och som har förlängts i väntan på att ersättas av ett nytt avtal,
–
med beaktande av de pågående förhandlingarna om ett nytt avtal som ska skapa en ny heltäckande ram för förbindelserna mellan EU och Ryssland, och av partnerskapet för modernisering som lanserades 2010,
–
med beaktande av sina tidigare betänkanden och resolutioner om Ryssland och förbindelserna mellan EU och Ryssland, särskilt resolutionen av den 9 juni 2011 om toppmötet mellan EU och Ryssland Antagna texter, P7_TA(2011)0268 .
, resolutionen av den 17 februari 2011 om rättsstatsprincipen i Ryssland Antagna texter, P7_TA(2011)0066 .
, resolutionen av den 17 juni 2010 om toppmötet mellan EU och Ryssland Antagna texter, P7_TA(2010)0234 .
, resolutionen av den 12 november 2009 inför toppmötet mellan EU och Ryssland i Stockholm den 18 november 2009 EUT C 271E, 7.10.2010, s.
2.
, resolutionen av den 17 september 2009 om morden på människorättsaktivister i Ryssland EUT C 224E, 19.8.2010, s.
27.
och resolutionen av den 17 september 2009 om de externa aspekterna av en tryggad energiförsörjning EUT C 224E, 19.8.2010, s.
23.
,
–
med beaktande av samråden om mänskliga rättigheter mellan EU och Ryssland, i synnerhet det senaste mötet den 4 maj 2011,
–
med beaktande av det ryska justitieministeriets beslut av den 22 juni 2011 om att avslå ansökan om att registrera Folkets frihetsparti (Parnas) och med beaktande av tidigare, liknande beslut som innebär att dessa partier inte kan delta i valet,
–
med beaktande av det uttalande om partiregistrering i Ryssland som Catherine Ashton, vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik, gjorde den 22 juni 2011,
–
med beaktande av Rysslands skyldighet, till följd av dess medlemskap i Europarådet och landets undertecknande av Europakonventionen om skydd för de mänskliga rättigheterna och de grundläggande friheterna, att upprätthålla demokratins principer,
–
med beaktande av resultatet av det toppmöte mellan EU och Ryssland som hölls i Nizjnij Novgorod den 9–10 juni 2011,
–
A.
Den politiska mångfalden är en hörnsten i demokratin och det moderna samhället, och en källa till politisk legitimitet.
B.
Den 12 april 2011 kritiserade Europadomstolen det tungrodda förfarandet för registrering av politiska partier i Ryssland, vilket inte är förenligt med den europeiska konventionen om skydd för de mänskliga rättigheterna och de grundläggande friheterna.
C.
Observatörer från kontoret för demokratiska institutioner och mänskliga rättigheter (ODIHR) besökte Ryssland under parlamentsvalet 2003 och föreslog att ett normalt OSSE-uppdrag skulle inledas sex veckor innan valet och bestå av 60 långtidsstationerade observatörer samt 400 observatörer med korta uppdrag.
D.
1.
Europaparlamentet är fortfarande övertygat om att Ryssland är en av EU:s viktigaste partner för strategiskt samarbete, med vilken unionen delar inte bara ekonomiska och handelsrelaterade intressen, utan även målet att föra ett nära samarbete såväl i det gemensamma grannskapet som på den internationella arenan.
2.
Europaparlamentet upprepar de åsikter parlamentet framförde i sin resolution av den 9 juni 2011 om toppmötet mellan EU och Ryssland i Nizjnij Novgorod.
3.
Europaparlamentet beklagar djupt de ryska myndigheternas beslut att avslå Folkets frihetspartis (Parnas) ansökan om registrering inför valet till statsduman i december 2011, och uppmanar de ryska myndigheterna att garantera fria och rättvisa val samt dra tillbaka alla beslut och bestämmelser som strider mot denna princip.
4.
Europaparlamentet upprepar sin oro över de svårigheter som de politiska partierna möter vad gäller registreringen inför valet, och som effektivt begränsar den politiska konkurrensen i Ryssland, minskar väljarnas valmöjligheter och visar att det fortfarande finns verkliga hinder för politisk mångfald i landet.
5.
6.
7.
8.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik, kommissionen, medlemsstaternas regeringar och parlament, OSSE, Europarådet samt Ryska federationens president, regering och parlament.
P7_TA-PROV(2011)0394
Eritrea: fallet Dawit Isaak
B7-0505 , 0507 , 0509 , 0510 , 0511 och 0512/2011
Europaparlamentets resolution av den 15 september 2011 om Eritrea: fallet Dawit Isaak
Europaparlamentet utfärdar denna resolution
–
med beaktande av den allmänna förklaringen om de mänskliga rättigheterna,
–
–
med beaktande av Afrikanska stadgan om mänskliga rättigheter och folkens rättigheter, i vilken Eritrea är part, i synnerhet artiklarna 6, 7 och 9,
–
med beaktande av artikel 9 i partnerskapsavtalet AVS–EU, i dess ändrade lydelse från 2005 (Cotonouavtalet), som Eritrea har undertecknat,
–
med beaktande av uttalandet från rådets ordförandeskap av den 22 september 2008 om politiska fångar i Eritrea samt senare uttalanden från rådet och kommissionen om Eritrea och om människorättssituationens utveckling sedan dess,
–
med beaktande av sina tidigare resolutioner om Eritrea, i synnerhet resolutionerna om de mänskliga rättigheterna och fallet Dawit Isaak,
–
A.
Det är djupt oroväckande att notera den försämrade människorättssituationen i Eritrea och de eritreanska myndigheternas uppenbara ovilja att samarbeta trots att EU och internationella människorättsorganisationer vid upprepade tillfällen vädjat om detta.
B.
C.
Rättsstatens principer får aldrig äventyras.
D.
Tusentals eritreaner, bland dem tidigare högt uppsatta medlemmar av det styrande partiet, har fängslats utan åtal, utan rättvis rättegång och utan möjlighet att träffa sina advokater eller anhöriga sedan de kritiserat president Isaias Afewerki offentligt 2001.
E.
F.
G.
I ett rättsligt yttrande som lades fram för Europaparlamentets talman i september 2010 framhålls att EU har en juridisk och moralisk skyldighet att skydda sina medborgare i enlighet med Europeiska konventionen om de mänskliga rättigheterna och i enlighet med EU-domstolens rättspraxis.
H.
Det är chockerande att Eritreas regering konsekvent vägrar att lämna ut någon information om fångarnas situation, exempelvis var de hålls fångna och om de ens är kvar i livet.
I.
Enligt rapporter från tidigare fångvaktare har mer än hälften av de tjänstemän och journalister som greps 2001 avlidit.
J.
EU är en viktig partner till Eritrea genom sitt utvecklingsstöd och bistånd till landet.
1.
Europaparlamentet noterar med stor oro den alltjämt undermåliga människorättssituationen i Eritrea, framför allt bristen på yttrandefrihet och den fortsatta förekomsten av politiska fångar, som frihetsberövats i strid med rättsstatens principer och Eritreas konstitution.
2.
3.
Europaparlamentet uppmanar de eritreanska myndigheterna att omedelbart frige Dawit Isaak och tidigare högt uppsatta tjänstemän i enlighet med den allmänna förklaringen om de mänskliga rättigheterna.
4.
Europaparlamentet uppmanar de eritreanska myndigheterna att häva förbudet mot landets oberoende press och att omedelbart frige de oberoende journalister och alla andra som har fängslats enbart för att de utövat sin rätt att yttra sig fritt.
5.
6.
Europaparlamentet uppmanar vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik att öka EU:s och dess medlemsstaters ansträngningar för att få Dawit Isaak fri.
7.
8.
Europaparlamentet vädjar till Afrikanska unionen, som är en partner till EU och som uttryckligen engagerar sig för universella värden som demokrati och mänskliga rättigheter, att intensifiera sina insatser med anledning av den beklagliga situationen i Eritrea och att arbeta tillsammans med EU för att se till att Dawit Isaak och andra politiska fångar släpps fria.
9.
Europaparlamentet följer med intresse den rättsliga processen till följd av att europeiska advokater i juli 2011 överklagade fallet Dawit Isaak till Eritreas högsta domstol under åberopande av skyddet mot godtyckliga frihetsberövanden (habeas corpus).
10.
Europaparlamentet upprepar sin begäran att det ska anordnas en nationell eritreansk konferens som för samman de olika politiska partiledarna och företrädarna för det civila samhället i syfte att komma med en lösning på den nuvarande krisen och föra landet i riktning mot demokrati, politisk pluralism och hållbar utveckling.
11.
Europaparlamentet framhåller med starkast möjliga eftertryck allvaret och den brådskande naturen i de frågor som behandlas ovan.
12.
Europaparlamentet uttrycker sitt uppriktiga stöd till och deltagande med de anhöriga till dessa politiska fångar.
13.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, vice ordföranden för kommissionen/unionens höga representant för utrikes frågor och säkerhetspolitik, medlemsstaternas parlament och regeringar, Eritreas parlament och regering, Panafrikanska parlamentet, Comesa, Igad, ordförandena för den gemensamma parlamentariska AVS–EU-församlingen samt Afrikanska unionen.
P7_TA-PROV(2011)0440
Genomförande av artikel 10 i FN:s protokoll om skjutvapen och införande av exporttillstånd samt import- och transiteringsåtgärder för skjutvapen, delar till skjutvapen och ammunition ***I
A7-0157/2011
Europaparlamentets lagstiftningsresolution av den 13 oktober 2011 om förslaget till Europaparlamentets och rådets förordning om genomförande av artikel 10 i FN:s protokoll om skjutvapen och om införande av exporttillstånd samt import- och transiteringsåtgärder för skjutvapen, delar till skjutvapen och ammunition ( KOM(2010)0273 – C7-0138/2010 – 2010/0147(COD) )
(Ordinarie lagstiftningsförfarande: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2010)0273 ),
–
–
–
–
med beaktande av artikel 55 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för internationell handel och yttrandet från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor ( A7-0157/2011 ).
1.
Europaparlamentet antar nedanstående ståndpunkt vid första behandlingen.
2.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om den har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
3.
Europaparlamentet uppdrar åt talmannen att översända parlamentets ståndpunkt till rådet, kommissionen och de nationella parlamenten.
P7_TC1-COD(2010)0147
Europaparlamentets ståndpunkt fastställd vid första behandlingen den 13 oktober 2011 inför antagandet av Europaparlamentets och rådets förordning (EU) nr .../2011 om genomförande av artikel 10 i FN:s protokoll om skjutvapen och om införande av exporttillstånd samt import- och transiteringsåtgärder för skjutvapen, delar till skjutvapen och ammunition
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om Europeiska unionens funktionssätt, särskilt artikel 207,
med beaktande av Europeiska kommissionens förslag,
efter översändande av utkastet till lagstiftningsakt till de nationella parlamenten,
, och
av följande skäl: (1)
I enlighet med rådets beslut 2001/748/EEG av den 16 oktober 2001 EUT L 280, 24.10.2001, s.
5.
13).
vägnar av protokollet mot olaglig tillverkning av och handel med eldvapen, delar till eldvapen och ammunition, bifogat till Förenta nationernas konvention mot gränsöverskridande organiserad brottslighet undertecknade kommissionen på gemenskapens vägnar nämnda protokoll (nedan kallat FN:s protokoll om skjutvapen eller protokollet) den 16 januari 2002.
(2)
(3)
För att göra det lättare att spåra skjutvapen och effektivt bekämpa olaglig handel med skjutvapen, delar och väsentliga delar till skjutvapen och ammunition är det nödvändigt att förbättra informationsutbytet mellan medlemsstaterna
, i synnerhet genom ett bättre utnyttjande av befintliga kommunikationskanaler
.
(4)
Behandlingen av personuppgifter ska genomföras i enlighet med bestämmelserna i Europaparlamentets och rådets direktiv 95/46/EG av den 24 oktober 1995 om skydd för enskilda personer med avseende på behandling av personuppgifter och om det fria flödet av sådana uppgifter EGT L 281, 23.11.1995, s.
31.
och Europaparlamentets och rådets förordning (EG) nr 45/2001 av den 18 december 2000 om skydd för enskilda då gemenskapsinstitutionerna och gemenskapsorganen behandlar personuppgifter och om den fria rörligheten för sådana uppgifter EGT L 8, 12.1.2001, s.
1.
.
(5)
5.
51.
om kontroll av förvärv och innehav av vapen.
(6)
Enligt FN:s protokoll om skjutvapen ska parterna införa eller förbättra sina administrativa förfaranden eller system för att utöva effektiv kontroll över tillverkningen, märkningen, importen och exporten av skjutvapen.
(7)
(8)
Denna förordning bör inte tillämpas på skjutvapen, delar och väsentliga delar till skjutvapen eller ammunition som är särskilt avsedda för militära ändamål.
Kraven i artikel 10 i FN:s protokoll om skjutvapen bör anpassas så att förenklade förfaranden införs för skjutvapen för civilt bruk.
På motsvarande sätt bör det sörjas för vissa lättnader när det gäller tillstånd för flera transporter, transiteringsåtgärder och temporär export för lagliga ändamål.
(9)
1.
eller på direktiv 91/477/EEC.
(10)
I direktiv 91/477/EEG behandlas överföringar av skjutvapen för civilt bruk inom Europeiska unionens territorium, medan denna förordning är inriktad på åtgärder rörande
export
till eller genom tredjeländer.
(11)
Skjutvapen, delar och väsentliga delar till skjutvapen och ammunition som importeras från tredjeländer omfattas av unionens lagstiftning och särskilt av kraven i direktiv 91/477/EEG.
(12)
Enhetligheten bör säkerställas med tanke på gällande bestämmelser om registerföring i unionens lagstiftning.
(13)
För att säkerställa en korrekt tillämpning av denna förordning bör varje medlemsstat vidta åtgärder som ger de behöriga myndigheterna nödvändiga befogenheter.
(14)
I syfte att
upprätthålla förteckningen över skjutvapen, delar och väsentliga delar till skjutvapen och ammunition för vilka tillstånd krävs enligt denna förordning
, bör befogenheten att anta akter i enlighet med artikel 290 i fördraget om Europeiska unionens funktionssätt delegeras till kommissionen med avseende på att anpassa bilaga I till denna förordning till
bilaga I till rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan EGT L 256, 7.9.1987, s.
1.
och till bilaga I till direktiv 91/477/EEG.
Kommissionen bör, då den förbereder och utarbetar delegerade akter, se till att relevanta handlingar översänds samtidigt till Europaparlamentet och rådet och att detta sker så snabbt som möjligt och på lämpligt sätt.
(15)
Unionen har antagit en samling tullbestämmelser som återfinns i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen EGT L 302, 19.10.1992, s.
1
och dess tillämpningsföreskrifter enligt kommissionens förordning (EEG) nr 2454/93 EGT L 253, 11.10.1993, s.
1.
.
Hänsyn bör också tas till Europaparlamentets och rådets förordning (EG) nr 450/2008 av den 23 april 2008 om fastställande av en tullkodex för gemenskapen (Moderniserad tullkodex) EUT L 145, 4.6.2008, s.
1.
, vars bestämmelser ska tillämpas i olika faser enligt artikel 188 i kodexen.
Ingenting i denna förordning inskränker eventuella bemyndiganden som har beviljats i kraft av och i enlighet med gemenskapens tullkodex och dess tillämpningsföreskrifter.
(16)
Dessa sanktioner bör vara effektiva, proportionella och avskräckande.
(17)
Denna förordning påverkar inte tillämpningen av unionens ordning för kontroll av export, överföring, förmedling och transitering av produkter med dubbla användningsområden som fastställts i rådets förordning (EG) nr 428/2009 av den 5 maj 2009 EUT L 134, 29.5.2009, s.1.
(18)
Denna förordning är i linje med de relevanta aspekter som förts fram om skjutvapen, delar och väsentliga delar till skjutvapen och ammunition för militär användning, säkerhetsstrategier, olaglig handel med handeldvapen och lätta vapen och export av militär teknik, däribland rådets gemensamma ståndpunkt 2008/944/Gusp av den 8 december 2008 om fastställande av gemensamma regler för kontrollen av export av militär teknik och krigsmateriel
EUT L 335, 13.12.2008, s.
99.
.
(19)
Kommissionen och medlemsstaterna bör underrätta varandra om de åtgärder som vidtas enligt denna förordning och om andra relevant uppgifter med anknytning till denna förordning som de förfogar över.
(20)
Denna förordning hindrar inte medlemsstaterna från att tillämpa sina konstitutionella bestämmelser om allmänhetens tillgång till officiella handlingar, med beaktande av Europaparlamentets och rådets förordning (EG) nr 1049/2001 av den 30 maj 2001 om allmänhetens tillgång till Europaparlamentets, rådets och kommissionens handlingar
EGT L 145, 31.5.2001, s.
43.
.
HÄRIGENOM FÖRESKRIVS FÖLJANDE:
KAPITEL I
SYFTE, DEFINITIONER OCH RÄCKVIDD Artikel 1
I denna förordning fastställs regler för exporttillstånd samt import- och transiteringsåtgärder för skjutvapen, delar och väsentliga delar till skjutvapen och ammunition, i syfte att genomföra artikel 10 i Förenta Nationernas protokoll mot olaglig tillverkning av och handel med eldvapen, delar till eldvapen och ammunition, bifogat Förenta nationernas konvention mot gränsöverskridande organiserad brottslighet (FN:s protokoll om skjutvapen).
Artikel 2
I denna förordning gäller följande definitioner:
1.
”Skjutvapen”: varje bärbart vapen med pipa som avfyrar, är avsett att avfyra, eller kan omvandlas till att avfyra ett skott, en kula eller en projektil med hjälp av ett antändbart drivämne
enligt bilaga I
.
Ett vapen anses kunna omvandlas till att avfyra ett skott, en kula eller en projektil med hjälp av ett explosivt ämne om
–
det liknar ett skjutvapen, och
–
det på grund av sin konstruktion eller sina materialegenskaper kan omvandlas på detta sätt.
2.
”Delar och väsentliga delar”: varje komponent eller ersättningskomponent
enligt bilaga I
som har utformats särskilt för ett skjutvapen och som är nödvändig för dess funktion, inbegripet pipa, stomme eller låda, glidskena eller cylinder, slutstycke samt varje anordning som formgivits eller anpassats för att dämpa det ljud som uppkommer då ett skjutvapen avfyras.
4.
”Ammunition”: alla patroner eller delar av patroner, inklusive patronhylsor, tändladdningar, drivladdningar, kulor och projektiler som används i skjutvapen
enligt bilaga I
, förutsatt att dessa delar själva omfattas av krav på tillstånd i den berörda medlemsstaten.
5.
”Skjutvapen som har gjorts obrukbara”: föremål som på annat sätt motsvarar definitionen skjutvapen som har gjorts definitivt obrukbara genom åtgärder som medför att skjutvapnets samtliga väsentliga delar gjorts definitivt oanvändbara och omöjliga att avlägsna, ersätta eller ändra med tanke på eventuell återanvändning.
Medlemsstaterna ska låta en behörig myndighet kontrollera dessa åtgärder för att göra skjutvapen obrukbara.
Medlemsstaterna ska föreskriva att det i samband med denna kontroll utfärdas ett intyg eller en annan handling av vilken det framgår att skjutvapnet är obrukbart eller att vapnet förses med en väl synlig märkning i detta syfte.
6.
”Export”:
a)
ett exportförfarande enligt artikel 161 i förordning (EEG) nr 2913/92,
b)
återexport enligt artikel 182 i förordning (EEG) nr 2913/92, med undantag av varor som
7.
”Person”: en fysisk eller juridisk person eller en sammanslutning av personer som tillerkänns rättskapacitet utan att vara juridiska personer, om det är möjligt enligt gällande lagstiftning.
8.
”Exportör”: varje ▌person
som är etablerad i unionen och som upprättar eller
på vars vägnar en exportdeklaration upprättas, dvs. den person som vid tidpunkten för deklarationens godkännande har ett avtal med mottagaren i tredje land och som har befogenhet att besluta om att föra ut varan ur unionens tullområde.
Om inget exportavtal har ingåtts eller om kontraktsinnehavaren inte agerar för egen räkning ska den person som har befogenhet att besluta om att föra ut varan ur unionens tullområde anses vara exportör.
När förfoganderätten över skjutvapen, delar och väsentliga delar till skjutvapen eller ammunition innehas av en person som är etablerad utanför unionen enligt det avtal på vilket exporten grundas, ska den avtalsslutande part som är etablerad i unionen anses vara exportör.
9.
”Gemenskapens tullområde”: de områden som avses i artikel 3 i förordning (EEG) nr 2913/92.
10.
”Exportdeklaration”: den handling genom vilken en person i föreskriven form och på föreskrivet sätt begär att få hänföra skjutvapen, delar och väsentliga delar till skjutvapen och ammunition till ett exportförfarande.
11.
”Temporär export”: utförsel från unionens tullområde av skjutvapen avsedda för återimport
inom en period som inte överstiger 24 månader.
12.
”Omlastning”: transitering där varorna fysiskt lastas av införseltransportmedlet och därefter lastas om
för återexport
, i allmänhet på ett annat transportmedel.
13.
”Transitering”: transport av varor från unionens tullområde, genom ett eller flera tredjeländers territorium med slutdestination i ett annat tredjeland.
14.
”Exporttillstånd”:
a)
ett enda
licens som ges en viss exportör för
en transport av ett eller flera skjutvapen, delar och väsentliga delar till skjutvapen och ammunition till en bestämd slutlig
mottagare eller mottagare i ett tredjeland
b)
exporttillstånd för flera transporter eller licens för flera licenser som ges en viss exportör för flera transporter av ett eller flera skjutvapen, delar och väsentliga delar till skjutvapen och ammunition till en bestämd slutlig mottagare eller mottagare i ett tredjeland, och/eller
c)
ett globalt tillstånd eller en global licens som ges en viss exportör för flera transporter av ett eller flera skjutvapen, delar och väsentliga delar till skjutvapen och ammunition till flera bestämda slutliga mottagare eller mottagare i ett eller flera tredjeländer.
▌
15.
a)
den berörda medlemsstaten inte tillåter det i enlighet med bestämmelserna i denna förordning,
b)
och 4.2
i direktiv 91/477/EEG, eller
c)
de importerade skjutvapnen inte vid tiden för införseln försetts med åtminstone en enkel märkning, varigenom det första importlandet inom Europeiska unionen kan identifieras, eller, om skjutvapnet saknar en sådan märkning, en unik märkning genom vilken de importerade skjutvapnen kan identifieras.
16.
”Spårning”: en systematisk utredning av hur skjutvapen och i förekommande fall delar och väsentliga delar till skjutvapen och ammunition går från tillverkare till köpare, i syfte att hjälpa medlemsstaternas behöriga myndigheter att upptäcka, utreda och analysera olaglig tillverkning och olaglig handel.
Artikel 3
1.
Denna förordning ska inte tillämpas på följande:
(a)
Bilaterala statliga transaktioner eller statliga överföringar.
(b)
Skjutvapen och delar och väsentliga delar till skjutvapen och ammunition, särskilt utformade för militär användning, och under alla omständigheter, helautomatiska skjutvapen.
(c)
(d)
Samlare och organ som ägnar sig åt de kulturella och historiska aspekterna hos skjutvapen, delar och väsentliga delar till skjutvapen och ammunition och som erkänts som sådana
i denna förordning
av den medlemsstat på vars territorium de är etablerade, förutsatt att de har sörjt för spårningsåtgärder.
(e)
Skjutvapen som har gjorts obrukbara.
(f)
▌
2.
KAPITEL II
EXPORTTILLSTÅND, FÖRFARANDEN OCH KONTROLLER
samt import- och transiteringsåtgärder
Artikel 4
Ett exporttillstånd
som har upprättats i enlighet med det formulär som anges i bilaga II
och ska utfärdas skriftligt eller på elektronisk väg
.
Om export av skjutvapen, delar och väsentliga delar till skjutvapen och ammunition kräver ett exporttillstånd i enlighet med denna förordning och också omfattas av krav på exporttillstånd i enlighet med rådets gemensamma ståndpunkt 2008/944/Gusp, kan medlemsstaterna tillämpa ett enda förfarande för att fullgöra sina skyldigheter enligt denna förordning och rådets gemensamma ståndpunkt.
Om skjutvapnen, delarna och de väsentliga delarna till skjutvapnen kommer att befinna sig i en eller flera medlemsstater andra än den där ansökan har lämnats in, ska detta anges i ansökan.
De behöriga myndigheterna i den medlemsstat där ansökan om tillstånd har lämnats in ska omedelbart samråda med de behöriga myndigheterna i den eller de berörda medlemsstaterna och förse dem med relevant information.
Den eller de medlemsstater som konsulteras ska inom 10 arbetsdagar framföra eventuella invändningar mot beviljandet av ett sådant tillstånd, vilka ska vara bindande för den medlemsstat där ansökan har lämnats in.
Artikel 5
Kommissionen ska
ges befogenhet att anta delegerade akter enligt artikel 6 med avseende på ändring av
bilaga I på grundval av ändringarna av bilaga I till förordning (EEG) nr 2658/87
och på grundval av bilaga I till direktiv 91/477/EEG
.
Artikel 6
1.
Befogenheten att anta delegerade akter ges till kommissionen med förbehåll för de villkor som anges i denna artikel.
2.
Befogenheten att anta delegerade akter som avses i artikel 5 ska ges till kommissionen på obestämd tid.
3.
Den delegering av befogenhet som avses i artikel 5 får när som helst återkallas av Europaparlamentet eller rådet.
Ett beslut om återkallelse innebär att delegeringen av den befogenhet som anges i beslutet upphör att gälla.
Beslutet får verkan dagen efter det att det har offentliggjorts i Europeiska unionens officiella tidning, eller vid ett senare i beslutet angivet datum.
Det påverkar inte giltigheten av delegerade akter som redan har trätt i kraft.
4.
Så snart kommissionen antar en delegerad akt ska den samtidigt delge Europaparlamentet och rådet denna.
5.
En delegerad akt som antas enligt artikel 5 ska träda i kraft endast om varken Europaparlamentet eller rådet har gjort invändningar mot den delegerade akten inom en period av två månader från den dag då akten delgavs Europaparlamentet och rådet, eller om både Europaparlamentet och rådet, före utgången av den perioden, har underrättat kommissionen om att de inte kommer att invända.
Denna period ska förlängas med två månader på Europaparlamentets eller rådets initiativ.
Artikel 7
1.
Innan en medlemsstat utfärdar ett exporttillstånd ▌ för skjutvapen, delar
och väsentliga delar
till skjutvapen, och ammunition ska den berörda medlemsstaten kontrollera att
(a)
det importerande tredjelandet har
gett sitt tillstånd till
importen, och
(b)
eventuella tredjeländer som är transitländer före transporten skriftligen har meddelat att de inte har några invändningar mot transiteringen.
Denna bestämmelse gäller inte för
–
transporter luft- eller sjövägen och transporter via hamnar eller flygplatser i tredjeländer, förutsatt att omlastning eller byte av transportmedel inte äger rum,
–
temporär export för kontrollerbara lagliga ändamål, vilket inbegriper jakt, tävlingsskytte, bedömning, utställningar utan försäljning och reparation.
2.
Medlemsstaterna får besluta
att om inga invändningar mot transiteringen inkommit inom 20 arbetsdagar från den dag då exportören ingivit sin skriftliga ansökan om godkännande av transiteringen det berörda tredjelandet som är transitland ska anses inte ha några invändningar mot transiteringen ▌.
3.
Exportören ska tillhandahålla den berörda myndighet i medlemsstaten som är ansvarig för utfärdandet av exporttillståndet ▌ de nödvändiga handlingar som visar att det importerande tredjelandet har gett sitt tillstånd till importen och att det tredjeland som är transitland inte haft några invändningar mot transiteringen ▌.
4.
Medlemsstaterna ska handlägga ansökningar om exporttillstånd ▌ inom en tidsrymd som fastställs i nationell lagstiftning eller praxis, men som ▌ inte får vara längre än
60 arbetsdagar från det datum då alla de uppgifter som krävs har lämnats till de behöriga myndigheterna
.
Under exceptionella omständigheter och av vederbörligen motiverade skäl kan denna tidsrymd förlängas till
5.
Giltighetstiden för ett exporttillstånd
får inte överstiga giltighetstiden för importtillståndet
.
inte vara kortare än
nio månader
.
6.
Medlemsstaterna får besluta att använda elektroniska dokument för handläggningen av ansökningarna om tillstånd.
Artikel 8
1.
För spårningsändamål ska exporttillståndet
och importlicensen
eller importtillståndet
som utfärdats av det importerande tredjelandet
och de åtföljande handlingarna innehålla uppgifter om bland annat följande:
(a)
Utfärdandedag och sista giltighetsdag för tillstånden.
(b)
Plats för utfärdande av tillstånden.
(c)
Exportland.
(d)
Importland.
(e)
I förekommande fall, tredjeländer eller länder som är transitländer.
(f)
Mottagare.
(g)
Slutlig mottagare, om denne är känd vid tidpunkten för avsändandet.
(h)
, delarna
2.
De uppgifter som det hänvisas till i punkt 1 ska, om de ingår i
importlicensen eller
importtillståndet, före transporten lämnas av exportören till de tredjeländer som är transitländer.
Artikel 9
1.
▌Förenklade förfaranden ▌ för temporär export
eller återexport
av skjutvapen
(a)
Inget exporttillstånd ska krävas för
(i)
temporär export som utförs av jägare eller tävlingsskyttar som en del av deras medförda personliga tillhörigheter, under en resa till ett tredjeland, förutsatt att de inför behöriga myndigheter styrker skälen för resan, lämpligen genom uppvisande av en inbjudan eller ett annat bevis på sin jakt- eller tävlingsskytteutövning i det tredjeland som är destinationsland, av
–
ett eller flera skjutvapen,
–
väsentliga delar, om detta anges, samt delar till skjutvapnen,
–
tillhörande ammunition, begränsat till högst 800 skott för jägare och högst 1200 skott för tävlingsskyttar,
(ii)
återexport som utförs av jägare eller tävlingsskyttar som en del av deras medförda personliga tillhörigheter efter tillfällig införsel för jakt- eller tävlingsskytteutövning, förutsatt att skjutvapnen fortfarande tillhör en person som är etablerad utanför unionens tullområde och att de återexporteras till denna person.
(b)
en annan medlemsstat än
den medlemsstat där de är bosatta, ▌visa upp
för behöriga myndigheter
det europeiska skjutvapenpasset enligt artiklarna 1 och 12 i direktiv 91/477/EEG ▌.
Vid lufttransport ska det europeiska skjutvapenpasset visas upp för de behöriga myndigheterna i samband med att de relevanta varorna lämnas över till lufttrafikföretaget för transport ut ur unionens tullområde.
Jägare och tävlingsskyttar får, när de lämnar unionens tullområde via
.
(c)
De behöriga myndigheterna i en medlemsstat ska, för en period som inte överstiger 10 arbetsdagar, avbryta förfarandet för export från eller, vid behov, på annat sätt förhindra att skjutvapen, delar eller väsentliga delar till skjutvapen, eller ammunition lämnar unionens tullområde via den medlemsstaten, om de har anledning att misstänka att de skäl som anförs av jägare eller tävlingsskyttar inte är förenliga med de relevanta aspekter och förpliktelser som fastställs i artikel 10.
Under exceptionella omständigheter och av vederbörligen motiverade skäl kan den tid tidsrymd som anges i detta led förlängas till 30 dagar.
2.
Medlemsstaterna ska i enlighet med sin gällande nationella lagstiftning införa förenklade förfaranden för
(a)
återexport av skjutvapen efter temporär införsel för bedömning eller utställning utan försäljning, eller i enlighet med förfarandet för aktiv förädling för reparation, förutsatt att skjutvapnen fortfarande tillhör en person som är etablerad utanför unionens tullområde och att de återexporteras till denna person,
(b)
återexport av skjutvapen, delar och väsentliga delar till skjutvapen, och ammunition i tillfällig förvaring från den tidpunkt då de förs in i unionens tullområde fram till utförseln,
(c)
temporär export av skjutvapen för bedömning och reparation samt utställning utan försäljning, förutsatt att exportören styrker sitt lagliga innehav av dessa skjutvapen och exporterar dem i enlighet med förfarandet för passiv förädling eller tullförfarandet för temporär export.
Artikel 10
1.
Vid beslut om beviljande av exporttillstånd ▌ enligt denna förordning ska medlemsstaterna vid behov beakta alla relevanta aspekter, inbegripet
(a)
▌
(b)
nationella utrikes- och säkerhetspolitiska aspekter, inbegripet de som täcks av rådets gemensamma ståndpunkt 2008/944/GUSP,
(c)
aspekter rörande den avsedda slutanvändningen, mottagaren
, den bestämda slutliga mottagaren
och risken för omdirigering.
2.
När medlemsstaterna bedömer en ansökan om exporttillstånd ▌ska de utöver kriterierna i punkt 1 även beakta huruvida exportören tillämpar proportionella och tillräckliga åtgärder och förfaranden i syfte att se till att bestämmelserna och målen i denna förordning och de krav och villkor som gäller för tillståndet iakttas.
När beslut fattas om huruvida ett exporttillstånd i enlighet med denna förordning ska beviljas, ska medlemsstaterna respektera sina förpliktelser med hänsyn till de sanktioner som införts genom beslut som antagits av rådet eller ett beslut av Organisationen för säkerhet och samarbete i Europa (OSSE) eller genom en bindande resolution av Förenta nationernas säkerhetsråd, särskilt rörande vapenembargon.
Artikel 11
1.
Medlemsstaterna ska
(a)
(b)
upphäva, tillfälligt upphäva, ändra eller återkalla ett exporttillstånd om villkoren för beviljande
inte uppfylldes eller
inte längre är uppfyllda.
Denna punkt hindrar inte tillämpningen av strängare regler enligt nationell lagstiftning.
2.
Om de behöriga myndigheterna i en medlemsstat tillfälligt har upphävt ett exporttillstånd ska deras slutliga bedömning meddelas medlemsstaterna när perioden för det tillfälliga upphävandet löper ut.
3.
Innan de behöriga myndigheterna i en medlemsstat ▌beviljar ett exporttillstånd
i enlighet med denna förordning
ska de
beakta
Om den behöriga myndigheten i medlemsstaten efter dessa samråd beslutar att bevilja ett tillstånd, ska den meddela de behöriga myndigheterna i de övriga medlemsstaterna och lämna alla relevanta uppgifter för att förklara beslutet.
4.
Artikel 12
Denna artikel ska inte tillämpas på ▌export ▌enligt artikel 9.
Artikel 13
1.
Medlemsstaterna
ska vid misstanke
begära att det importerande tredjelandet bekräftar mottagandet av transporten av skjutvapen, delar eller väsentliga delar till skjutvapen eller ammunition.
2.
Medlemsstaterna ska på begäran underrätta det exporterande tredjelandet om mottagandet inom unionens tullområde av transporten av skjutvapen, delar eller väsentliga delar till skjutvapen eller ammunition.
En sådan bekräftelse ska i princip ske genom uppvisande av de relevanta tullhandlingarna för import.
Det första stycket ska tillämpas endast om det anmodande exporterande tredjelandet var en part i FN:s protokoll om skjutvapen redan vid tidpunkten för exporten till unionen.
3.
Medlemsstaterna ska följa bestämmelserna i punkterna 1 och 2 i enlighet med deras gällande nationella lagstiftning eller praxis.
Särskilt när det gäller export ▌får medlemsstatens behöriga myndighet besluta att antingen vända sig till exportören eller ta kontakt direkt med det importerande tredjelandet.
Artikel 14
Kontroll och validering kan i förekommande fall säkerställas via diplomatiska kanaler.
Artikel 15
För att säkerställa en korrekt tillämpning av denna förordning ska varje medlemsstat vidta nödvändiga och proportionella åtgärder för att göra det möjligt för dess behöriga myndigheter att
(a)
(b)
fastställa att exportkontrollåtgärderna tillämpas korrekt, vilket särskilt får inbegripa rätt till tillträde till lokaler som tillhör personer som berörs av en exporttransaktion.
Artikel 16
KAPITEL III
Artikel 17
1.
Vid fullgörandet av
tullformaliteterna
för export av skjutvapen, delar och väsentliga delar till skjutvapen och ammunition vid
exporttullkontoret
ska exportören framlägga bevis för att nödvändigt exporttillstånd har erhållits.
2.
Exportören får anmodas att av varje dokument som framläggs som bevis tillhandahålla en översättning till ett officiellt språk i den medlemsstat där exportdeklarationen uppvisas.
3.
Medlemsstaterna
ska
även, utan att det påverkar befogenheter som de tilldelats i enlighet med förordning (EEG) nr 2913/92, för en period som inte överstiger 10
dagar
avbryta förfarandet för export från
sina territorier
eller, vid behov, på annat sätt förhindra att skjutvapen, delar eller väsentliga delar till skjutvapen eller ammunition som omfattas av ett giltigt exporttillstånd lämnar
unionens tullområde
▌via
deras
territorium, om
de
har anledning att misstänka att
(a)
relevanta uppgifter inte beaktades när tillståndet beviljades, eller
(b)
omständigheterna har ändrats väsentligt sedan tillståndet beviljades.
Under exceptionella omständigheter och av vederbörligen styrkta skäl kan denna tidsrymd förlängas till 30 dagar.
4.
Artikel 18
1.
Medlemsstaterna får besluta att tullformaliteterna för export av skjutvapen, delar och väsentliga delar till skjutvapen eller ammunition endast kan fullgöras vid tullkontor som bemyndigats för detta ändamål.
2.
KAPITEL IV
ADMINISTRATIVT SAMARBETE Artikel 19
1.
vidta alla lämpliga åtgärder för att upprätta ett direkt samarbete och informationsutbyte mellan de behöriga myndigheterna, i syfte att öka effektiviteten av de åtgärder som fastställs i denna förordning.
Denna information får omfatta
(a)
uppgifter om exportörer vars ansökan om tillstånd har avslagits eller exportörer som omfattas av beslut av medlemsstaterna i enlighet med artikel 11,
(b)
uppgifter om mottagare eller andra aktörer som deltar i misstänkt verksamhet och, om sådana uppgifter är tillgängliga, om transportvägar.
2.
1.
KAPITEL V
ALLMÄNNA BESTÄMMELSER OCH SLUTBESTÄMMELSER Artikel 20
1.
En samordningsgrupp för frågor rörande export av skjutvapen, med en företrädare för kommissionen som ordförande, ska inrättas.
Varje medlemsstat skall utse en företrädare till denna.
Samordningsgruppen ska undersöka varje fråga som avser tillämpningen av denna förordning som kan tas upp antingen av ordföranden eller av en företrädare för en medlemsstat.
Den ska vara bunden av reglerna om sekretesskydd i förordning (EG) nr 515/97.
2.
Artikel 21
1.
Varje medlemsstat ska informera kommissionen om de lagar och andra författningar som antas för genomförandet av denna förordning, inbegripet de åtgärder som avses i artikel 16.
2.
Senast när denna förordning träder i kraft ska varje medlemsstat
informera de
På grundval av de uppgifter som lämnas av medlemsstaterna ska kommissionen offentliggöra och årligen uppdatera en förteckning över dessa myndigheter i C-serien av Europeiska unionens officiella tidning.
3.
ska kommissionen se över tillämpningen av den här förordningen och lägga fram en rapport till Europaparlamentet och rådet om tillämpningen, vilken kan innehålla ändringsförslag.
Medlemsstaterna ska förse kommissionen med alla relevanta uppgifter som den behöver för att utarbeta denna rapport
.
Artikel 22
Denna förordning träder i kraft den tjugonde dagen efter den dag då denna förordning offentliggörs i
EUT: Vänligen för in datumet 18 månader efter det att denna förordning har offentliggjorts.
har trätt i kraft i Europeiska unionen,
.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Utfärdad i
På Europaparlamentets vägnar På rådets vägnar
Ordförande Ordförande
BILAGA I
Bygger på kombinerade nomenklaturen för varor enligt rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan.
Förteckning över skjutvapen, delar och väsentliga delar till skjutvapen och ammunition såsom avses i artiklarna 2.1 och 4.1:
▌
Varuslag
KN-nummer
Där ”ex” anges före KN-numret skall tillämpningen av förmånssystemet bestämmas såväl av KN-numret som av den motsvarande varubeskrivningen.
1
Halvautomatiska eller repeterande korta vapen
ex 9302 00 00
2
Korta vapen med enkelskott med centralantändning.
ex 9302 00 00
3
Korta vapen med enkelskott med kantantändning, vars totala längd är mindre än 28 cm.
ex 9302 00 00
4
Halvautomatiska långa skjutvapen, vars magasin och patronläge tillsammans kan innehålla mer än tre skott.
ex 9303 20 10
ex 9303 20 95
ex 9303 30 00
ex 9303 90 00
5
Halvautomatiska långa skjutvapen, vars magasin och patronläge tillsammans inte kan innehålla mer än tre skott och där laddningsmekanismen kan tas bort eller det inte är uteslutet att vapnet med hjälp av vanliga verktyg kan omändras på sådant sätt att magasin och patronläge tillsammans kan innehålla mer än tre skott.
ex 9303 20 10
ex 9303 20 95
ex 9303 30 00
ex 9303 90 00
6
Repeterande och halvautomatiska långa skjutvapen med slätborrade lopp som inte överstiger 60 cm i längd.
ex 9303 20 10
ex 9303 20 95
7
Halvautomatiska skjutvapen för civilt bruk som liknar vapen med automatisk mekanism.
ex 9302 00 00
ex 9303 20 10
ex 9303 20 95
ex 9303 30 00
ex 9303 90 00
8
Repeterande långa skjutvapen andra än de som står upptagna i punkt 6.
ex 9303 20 95
ex 9303 30 00
ex 9303 90 00
9
Långa skjutvapen med räfflade lopp för enkelskott.
ex 9303 30 00
ex 9303 90 00
10
Halvautomatiska långa skjutvapen som inte omfattas av punkterna 4–7.
ex 9303 90 00
11
Korta vapen med enkelskott med kantantändning, vars totala längd inte är mindre än 28 cm.
ex 9302 00 00
12
Enkelskotts långa skjutvapen med slätborrade lopp.
9303 10 00
ex 9303 20 10
ex 9303 20 95
13
Delar som har utformats särskilt för ett skjutvapen och som är nödvändig för dess funktion, inbegripet pipa, stomme eller låda, glidskena eller cylinder, slutstycke samt varje anordning som formgivits eller anpassats för att dämpa det ljud som uppkommer då ett skjutvapen avfyras.
Varje väsentlig del av sådana skjutvapen: slutstycket, patronläget och pipan till ett skjutvapen tillhör som separata delar samma kategori som det skjutvapen de är eller är tänkta att vara monterade på.
ex 9305 10 00
ex 9305 21 00
ex 9305 29 00
ex 9305 99 00
14
Ammunition: alla patroner eller delar av patroner, inklusive patronhylsor, tändladdningar, drivladdningar, kulor och projektiler som används i skjutvapen, förutsatt att dessa delar själva omfattas av krav på tillstånd i den berörda medlemsstaten.
ex 3601 00 00
ex 3603 00 90
ex 9306 21 00
ex 9306 29 00
ex 9306 30 10
ex 9306 30 90
ex 9306 90 90
15
Samlingar och samlarobjekt av historiskt intresse
Antikviteter med en ålder av över 100 år
ex 9705 00 00
ex 9706 00 00
I denna bilaga gäller följande definitioner:
(a)
korta vapen: ett skjutvapen med en pipa som inte överstiger 30 cm eller vars totala längd inte överstiger 60 cm.
(b)
långa vapen: alla skjutvapen som inte är korta vapen.
(c)
automatvapen: ett skjutvapen som laddar om automatiskt varje gång ett skott avfyras och som kan avfyra mer än ett skott med ett tryck på avtryckaren.
(d)
halvautomatiskt skjutvapen: ett skjutvapen som laddar om automatiskt varje gång ett skott avfyras och som bara kan avfyra ett skott med ett tryck på avtryckaren.
(e)
repeterande skjutvapen: ett skjutvapen som efter att ett skott har avfyrats är avsett att laddas om från ett magasin eller cylinder med hjälp av ett manuellt tillvägagångssätt.
(f)
skjutvapen för enkelskott: ett skjutvapen utan magasin som laddas för varje skott genom att man manuellt sätter in ett skott i patronläget eller i ett laddningsutrymme där pipan bryts.
Bilaga II
(förlaga till formulär för exporttillstånd)
(som det hänvisas till i artikel 4 i denna förordning)
När medlemsstaterna beviljar exporttillstånd ska de se till att det på formuläret framgår vilken typ av tillstånd som avses.
Detta exporttillstånd gäller till sista giltighetsdag i alla Europeiska unionens medlemsstater.
EUROPEISKA UNIONEN
EXPORT AV SKJUTVAPEN (förordning (EG) nr…/20…
* EUT: Vänligen för in referensnumret på denna förordning.
)
Typ av tillstånd
1
1.
Exportör
(EORI-nummer i förekommande fall)
nr
2.
Tillståndets identifikationsnummer
Fylls i av utfärdande myndighet.
3.
Sista giltighetsdag
Där ”ex” anges före KN-numret skall tillämpningen av förmånssystemet bestämmas såväl av KN-numret som av den motsvarande varubeskrivningen.
TILLSTÅND
4.
Uppgifter om kontaktställe
5.
Mottagare (EORI-nummer i förekommande fall)
6.
Utfärdande myndighet
7.
Ombud/representant
(om annan än exportören) (EORI-nummer i förekommande fall)
nr
8.
Exportland
Kod (
Se förordning (EG) nr°1172/95 (EGT L 118, 25.5.1995, s.
10) i dess gällande lydelse.
)
9.
Importland och antal importtillstånd
Kod (
1
)
10.
Slutlig mottagare (om denne är känd vid tidpunkten för avsändandet) (EORI-nummer i förekommande fall)
11.
Tredjeländer som är transitländer (i förekommande fall)
Kod (
1
)
12.
Medlemsstat där varorna kommer att hänföras till exportförfarande
Kod (
1
)
13.
Se förordning (EG) nr 1172/95 (EGT L 118, 25.5.1995, s.
10) i dess gällande lydelse.
)
14.
Varukod enligt Harmoniserade systemet eller Kombinerade nomenklaturen (i förekommande fall med 8 siffror)
13.a Märkning
15.
Valuta och värde
16.
Varumängd
19.
Exportförfarande
17.
Slutanvändning (i förekommande fall)
18.
Kontraktsdatum (i förekommande fall)
20.
Ytterligare upplysningar som krävs enligt nationell lagstiftning (anges på formuläret)
Fält för eventuell förtryckt information
från medlemsstaterna
Fylls i av utfärdande myndighet
Underskrift
Utfärdande myndighet
Stämpel
Fält för eventuell förtryckt information
från medlemsstaterna
Ort och datum
EUROPEISKA UNIONEN
1a
Ett separat formulär ska fyllas i för varje mottagare.
1.
Exportör
2.
Identifikationsnummer
9.
Importland och antal importtillstånd
TILLSTÅND
5.
Mottagare
13.1.
Beskrivning av produkterna
14.
Varukod (i förekommande fall med 8 siffror)
13.a Märkning
15.
Valuta och värde
16.
Varumängd
13.1.
Beskrivning av produkterna
14.
Varukod (i förekommande fall med 8 siffror)
13.a Märkning
15.
Valuta och värde
16.
Varumängd
13.
3.
Beskrivning av produkterna
14.
Varukod (i förekommande fall med 8 siffror)
13.a Märkning
15.
Valuta och värde
16.
Varumängd
13.
4.
Beskrivning av produkterna
14.
Varukod (i förekommande fall med 8 siffror)
13.a Märkning
15.
Valuta och värde
16.
Varumängd
13.
5.
Beskrivning av produkterna
14.
Varukod (i förekommande fall med 8 siffror)
13.a Märkning
15.
Valuta och värde
16.
Varumängd
13.
6.
Beskrivning av produkterna
14.
Varukod (i förekommande fall med 8 siffror)
13.a Märkning
15.
Valuta och värde
16.
Varumängd
13.
7.
Beskrivning av produkterna
14.
Varukod (i förekommande fall med 8 siffror)
13.a Märkning
15.
Valuta och värde
16.
Varumängd
Anmärkning: Ett separat formulär ska fyllas i för varje mottagare, i linje med 1a.
I kolumn 22 ska i fält 1 anges den återstående kvantiteten och i fält 2 den mängd som dras av vid detta tillfälle.
21.
Nettomängd/-värde (nettovikt eller annan specificerad enhet)
24.
Tulldokument (typ och nummer) eller utdrag (nr) och datum för avdraget
25.
Medlemsstat, namn och underskrift, avdragande myndighets stämpel
22.
Med siffror
23.
Avdragen mängd/avdraget värde med bokstäver
1
2
1
2
1
2
1
2
1
2
1
2
P7_TA-PROV(2011)0452
Motorer som släpps ut på marknaden enligt flexibilitetssystemet ***I
A7-0080/2011
Europaparlamentets lagstiftningsresolution av den 25 oktober 2011 om förslaget till Europaparlamentets och rådets direktiv om ändring av direktiv 97/68/EG vad gäller bestämmelser om motorer som släpps ut på marknaden enligt flexibilitetssystemet ( KOM(2010)0362 – C7-0171/2010 – 2010/0195(COD) )
(Ordinarie lagstiftningsförfarande: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2010)0362 ),
–
–
–
med beaktande av yttrandet från Europeiska ekonomiska och sociala kommittén av den 16 september 2010 EUT C 48, 15.2.2011, s.
134.
,
–
–
med beaktande av artikel 55 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för miljö, folkhälsa och livsmedelssäkerhet och yttrandet från utskottet för transport och turism ( A7-0080/2011 ).
1.
Europaparlamentet antar nedanstående ståndpunkt vid första behandlingen.
2.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om den har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
3.
Europaparlamentet uppdrar åt talmannen att översända parlamentets ståndpunkt till rådet, kommissionen och de nationella parlamenten.
P7_TC1-COD(2010)0195
Europaparlamentets ståndpunkt fastställd vid den första behandlingen av den 25 oktober 2011 inför antagandet av Europaparlamentets och rådets direktiv 2011/.../EU om ändring av direktiv 97/68/EG vad gäller bestämmelserna om motorer som släpps ut på marknaden enligt flexibilitetssystemet
(Text av betydelse för EES)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av fördraget om Europeiska unionens funktionssätt, särskilt artikel 114,
med beaktande av Europeiska kommissionens förslag,
efter översändande av utkastet till lagstiftningsakt till de nationella parlamenten,
med beaktande av Ekonomiska och sociala kommitténs yttrande EUT C 48, 15.2.2011, s.
134.
,
i enlighet med det ordinarie lagstiftningsförfarandet Europaparlamentets ståndpunkt av den 25 oktober 2011 (ännu ej offentliggjord i EUT) och rådets beslut av den …
, och
av följande skäl: (1)
Europaparlamentets och rådets direktiv 97/68/EG av den 16 december 1997 om tillnärmning av medlemsstaternas lagstiftning om åtgärder mot utsläpp av gas- och partikelformiga föroreningar från förbränningsmotorer som skall monteras i mobila maskiner som inte är avsedda att användas för transporter på väg EGT L 59, 27.2.1998, s.
1.
reglerar avgasutsläpp
och fastställer utsläppsgränser för luftföroreningar
från motorer monterade i maskiner som inte är avsedda att användas på väg
samt bidrar till skyddet av människors hälsa och miljön
.
(2)
Översynen av direktiv 97/68/EG förbereds för närvarande av kommissionen i enlighet med kraven i artikel 2 i Europaparlamentets och rådets direktiv 2004/26/EG av den 21 april 2004 om ändring av direktiv 97/68/EG
EUT L 146, 30.4.2004, s.
1.
.
För att säkerställa att direktivet efter översynen följer unionens normer för god luftkvalitet och mot bakgrund av erfarenheten, vetenskapliga rön och tillgänglig teknik bör kommissionen i samband med den kommande översynen av direktiv 97/68/EG, om inte annat följer av konsekvensbedömningen, överväga
–
att införa ett nytt utsläppssteg – steg V – som, under förutsättning att det är tekniskt möjligt, bör grundas på kraven för Euro 6-normerna för tunga nyttofordon,
–
att införa nya krav på minskning av partiklar, det vill säga en gräns för antalet partiklar vilken, om det är tekniskt möjligt, ska gälla för alla kategorier av motorer med kompressionständning i syfte att säkerställa en effektiv minskning av ultrafina partiklar,
–
att inta en helhetssyn på främjandet av utsläppsminskande föreskrifter och eftermontering av efterbehandlingssystem i de befintliga maskiner som inte är avsedda att användas på väg, på grundval av de diskussioner som just nu pågår under överinseende av FN:s ekonomiska kommission för Europa beträffande harmoniserade krav på eftermontering av utsläppsbegränsande anordningar ; detta förhållningssätt bör stödja medlemsstaterna i deras arbete för att förbättra luftkvaliteten och främja arbetstagarskyddet,
–
att införa en metod för regelbunden testning av mobila maskiner och fordon som inte är avsedda att användas på väg, särskilt för att fastställa om deras utsläppsprestanda faktiskt motsvarar de värden som angetts vid registreringen,
–
möjligheten att under vissa omständigheter tillåta utbytesmotorer som inte uppfyller kraven i steg III A för rälsbussar och lokomotiv,
–
möjligheten att harmonisera de specifika utsläppsnormerna för järnvägsfordon med relevanta internationella normer i syfte att säkerställa tillgången till överkomligt prissatta motorer som följer de fastställda utsläppsgränserna.
(3)
Övergången till steg III B kräver en drastisk teknikändring som innebär avsevärda kostnader för omkonstruktion av motorerna och framtagning av avancerade tekniska lösningar.
Den rådande globala finansiella och ekonomiska krisen eller eventuella ekonomiska konjunkturfluktuationer bör dock inte medföra sänkta miljönormer.
Denna översyn av direktiv 97/68/EG bör därför anses utgöra ett undantag.
Dessutom är investeringar i miljövänlig teknik viktiga för främjande av framtida tillväxt, sysselsättning och hälsoskydd.
(4)
I direktiv 97/68/EG föreskrivs ett flexibilitetssystem, så att utrustningstillverkarna under tiden mellan två utsläppssteg kan köpa in ett begränsat antal motorer som inte uppfyller de utsläppsgränser som gäller under den perioden men som är godkända enligt kraven i det närmast föregående steget av utsläppsgränser.
(5)
(6)
Under steg III B bör det maximala antal motorer som används för andra tillämpningar än framdrivning av rälsbussar
,
lokomotiv och
kvantitet
utrustning med motorer i den kategorin som utrustningstillverkaren
Alternativet att ett fast
antal motorer får släppas ut på marknaden enligt flexibilitetssystemet bör
.
Detta fasta antal motorer bör också granskas och det bör inte överskrida värdena i avsnitt 1.2.2 i bilaga XIII till direktiv 97/68/EG.
(7)
Reglerna för flexibilitetssystemet bör anpassas för att utöka systemets tillämpning till motorer för framdrivning av lokomotiv
under en strikt begränsad tidsperiod
.
(8)
Att förbättra luftkvaliteten är ett viktigt mål för unionen, som eftersträvas genom Europaparlamentets och rådets direktiv 2008/50/EG av den 21 maj 2008 om luftkvalitet och renare luft i Europa
EUT L 152, 11.6.2008, s.
1.
.
Att utsläppen åtgärdas vid källan har stor betydelse för uppnåendet av detta mål, inklusive en minskning av utsläppen från sektorn för mobila maskiner som inte är avsedda att användas på väg.
(9)
Företag som arbetar med maskiner som omfattas av detta direktiv bör kunna utnyttja europeiska ekonomiska stödprogram eller relevanta stödprogram i medlemsstaterna.
Dessa stödprogram bör syfta till att främja ett tidigt införande av högsta möjliga utsläppsnormer.
(10)
I direktiv 97/68/EG stadgas det om ett undantag för utbytesmotorer, vilket inte gäller för rälsbussar och lokomotiv.
Med tanke på vikt- och storleksrestriktioner är det dock nödvändigt att införa ett begränsat undantag även för utbytesmotorer för rälsbussar och lokomotiv.
(11)
De åtgärder som anges i detta direktiv återspeglar tillfälliga svårigheter som tillverkningsindustrin drabbats av
.
(12)
Med hänsyn till den speciella infrastrukturen i Förenade kungarikets järnvägsnät, som medför andra strukturella mått och därmed även vikt- och storleksrestriktioner och som därför behöver en längre period för anpassningar till nya utsläppsgränser, är det lämpligt att medge ökad flexibilitet för denna specifika marknad när det gäller motorer för användning i lokomotiv.
13)
Direktiv 97/68/EG bör därför ändras i enlighet med detta.
Direktiv 97/68/EG ska ändras på följande sätt:
1.
Förbränningsmotorer med kompressionständning som är avsedda att användas för andra ändamål än framdrivning av
rälsbussar och
fartyg i inlandssjöfart får släppas ut på marknaden inom ramen för ett flexibilitetssystem i enlighet med förfarandet i bilaga XIII och förfarandet i punkterna 1–5.
2.
Artikel 10 ska ändras på följande sätt:
a)
I punkt 1a ska andra stycket utgå.
b)
Följande punkter ska införas:
1b.
a)
utbytesmotorer som överensstämmer med gränserna enligt steg III A och som ersätter motorer för rälsbussar och lokomotiv som
i)
inte uppfyller normerna enligt steg III A, eller
ii)
uppfyller normerna enligt steg III A men inte normerna enligt steg III B,
b)
utbytesmotorer som inte överensstämmer med gränserna enligt steg III A och som ersätter motorer för rälsbussar som saknar körkontroll och inte är självgående, om dessa utbytesmotorer uppfyller normer som inte är lägre än de normer som uppfylls av de motorer som är monterade i befintliga rälsbussar av samma typ.
Tillstånd enligt denna punkt får beviljas enbart i fall då godkännandemyndigheten i medlemsstaten är säker på att användningen i rälsbussen eller lokomotivet i fråga av en utbytesmotor som uppfyller kraven enligt det senast tillämpbara utsläppssteget kommer att medföra betydande tekniska svårigheter.
1c.
Motorer som omfattas av punkt 1a eller 1b ska märkas med texten ’UTBYTESMOTOR’ och den unika hänvisningen till det aktuella undantaget.
1d.
Kommissionen ska bedöma de negativa miljöeffekterna av punkt 1b och eventuella tekniska svårigheter beträffande efterlevnaden av bestämmelserna i den punkten.
Mot bakgrund av denna bedömning ska kommissionen senast den 31 december 2016 lägga fram en rapport till Europaparlamentet och rådet med en översyn av punkt 1b, i lämpliga fall åtföljd av ett lagstiftningsförslag som inbegriper ett slutdatum för tillämpningen av den punkten.
c)
Punkt 7 ska ersättas med följande: 7.
Medlemsstaterna ska tillåta att motorer enligt de definitioner som ingår i punkterna A i, A ii och A v i avsnitt 1 i bilaga I släpps ut på marknaden i enlighet med det flexibilitetssystem som definierats i enlighet med föreskrifterna som anges i bilaga XIII.
▌
3.
Bilaga XIII ska ändras i enlighet med bilagan till det här direktivet.
Artikel 2 Införlivande
1.
Medlemsstaterna ska senast den ... * EUT: Vänligen för in datumet: Tolv månader efter offentliggörandet av detta direktiv.
anta och offentliggöra de lagar och andra författningar som är nödvändiga för att följa detta direktiv.
De ska genast överlämna texten till dessa bestämmelser till kommissionen.
När en medlemsstat antar dessa bestämmelser ska de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs.
Närmare föreskrifter om hur hänvisningen ska göras ska varje medlemsstat själv utfärda.
2.
Medlemsstaterna ska till kommissionen överlämna texten till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 3 Ikraftträdande
Detta direktiv träder i kraft den tjugonde dagen efter det att det har offentliggjorts i
Europeiska unionens officiella tidning
.
Artikel 4 Adressater
Detta direktiv riktar sig till medlemsstaterna.
Utfärdat i
På Europaparlamentets vägnar På rådets vägnar
Ordförande Ordförande
BILAGA
Avsnitt 1 i bilaga XIII ska ersättas med följande: 1.
UTRUSTNINGSTILLVERKARENS ÅTGÄRDER
1.1
Med undantag för steg III B ska en utrustningstillverkare som vill utnyttja flexibilitetssystemet
, med undantag för motorer för framdrivning av rälsbussar och lokomotiv,
.
får inte överskrida de tak
som beskrivs i avsnitten 1.1.1 och 1.1.2.
1.1.1
årliga
släpper ut på marknaden
(beräknat som ett medelvärde av de senaste fem årens försäljning på unionsmarknaden).
ska
1.1.2
Som alternativ till avsnitt 1.1.1 och med undantag för motorer för framdrivning av rälsbussar och lokomotiv får utrustningstillverkaren söka tillstånd för sina
motortillverkare
att släppa ut ett fast antal motorer på marknaden
vilka är avsedda att användas enbart av utrustningstillverkaren
.
Antalet motorer i varje motorkategori får inte överskrida följande tak:
Motorkategori
P (kW)
Antal motorer
19 ≤ P < 37
200
37 ≤ P < 75
150
75 ≤ P < 130
100
130 ≤ P ≤ 560
50
1.2
Med undantag för motorer för framdrivning av rälsbussar och lokomotiv ska, under steg III B
men inte längre än tre år efter det att detta steg har börjat tillämpas
motortillverkare att släppa ut motorer på marknaden vilka är avsedda att användas enbart av utrustningstillverkaren
.
1.2.1
Antalet motorer som släpps ut på marknaden enligt flexibilitetssystemet får för varje motorkategori inte överskrida
37,5 %
årliga
släpper ut på marknaden
(beräknat som medelvärdet av de senaste fem årens försäljning på unionsmarknaden).
ska
1.2.2
Som alternativ till avsnitt 1.2.1 får utrustningstillverkaren söka tillstånd för sina
motortillverkare
att släppa ut ett fast antal motorer på marknaden
vilka är avsedda att användas enbart av utrustningstillverkaren
.
Antalet motorer i varje motorkategori får inte överskrida följande tak:
Motorkategori
P (kW)
Antal motorer
37 ≤ P < 56
200
56 ≤ P < 75
175
75 ≤ P < 130
250
130 ≤ P ≤ 560
125
▌
1.4
När det gäller motorer för framdrivning av lokomotiv får en utrustningstillverkare under steg III B,
men inte längre än tre år efter det att detta steg har börjat tillämpas,
söka tillstånd för sina
motortillverkare
att släppa ut högst
16 motorer
på marknaden
vilka är avsedda att användas enbart av utrustningstillverkaren
Lokomotiv ska anses uppfylla detta krav endast om de har ett säkerhetscertifikat för drift i Förenade kungarikets nät, eller om ett sådant certifikat kan utfärdas för dem.
Ett sådant tillstånd ska beviljas endast när det finns tekniska skäl till att utsläppsgränserna för steg III B inte kan uppfyllas.
1.5
Utrustningstillverkaren ska i sin ansökan till godkännandemyndigheten lämna följande upplysningar:
a)
Ett prov på den märkning som ska anbringas på varje mobil maskin som inte är avsedd att användas på väg i vilken en motor som släppts ut på marknaden enligt flexibilitetssystemet är avsedd att installeras.
Märkningen ska innehålla följande text: ’MASKIN nr … (maskinens löpnummer) AV … (totalt antal maskiner i respektive effektkategori) MED MOTOR nr … TYPGODKÄND (dir.
97/68/EG) MED nr …’.
b)
Ett prov på den tilläggsmärkning som ska anbringas på motorn med den text som avses i avsnitt 2.2.
1.6
Utrustningstillverkaren ska förse godkännandemyndigheten med alla nödvändiga upplysningar om tillämpningen av flexibilitetssystemet som godkännandemyndigheten kan begära för att kunna fatta ett beslut.
1.7
Utrustningstillverkaren ska förse alla godkännandemyndigheter i medlemsstaterna som begär det med alla upplysningar som godkännandemyndigheten begär för att bekräfta att en motor som påstås vara utsläppt eller som är märkt som utsläppt på marknaden enligt flexibilitetssystemet verkligen är det.
P7_TA-PROV(2011)0473
Det hot mot folkhälsan som antimikrobiell resistens utgör
B7-0538/2011
Europaparlamentets resolution av den 27 oktober 2011 om det hot mot folkhälsan som antimikrobiell resistens utgör
Europaparlamentet utfärdar denna resolution
–
med beaktande av sin resolution av den 12 maj 2011 om antibiotikaresistens, som främst tar upp djurhälsa,
–
med beaktande av det vetenskapliga yttrandet från Europeiska myndigheten för livsmedelssäkerhet (Efsa) från augusti 2011 med titeln ”on the public health risks of bacterial strains producing extended-spectrum β-lactamases and/or AmpC β-lactamases in food and food-producing animals”,
–
med beaktande av kommissionens arbetsdokument av den 18 november 2009 om antimikrobiell resistens (SANCO/6876/2009r6),
–
med beaktande av den gemensamma tekniska rapporten från september 2009 från Europeiska centrumet för förebyggande och kontroll av sjukdomar (ECDC) och från Europeiska läkemedelsmyndigheten (EMA) om ”The bacterial challenge: time to react – A call to narrow the gap between multidrug-resistant bacteria in the EU and the development of new antibacterial agents”,
–
med beaktande av rådets rekommendation av den 15 november 2001 om återhållsam användning av antimikrobiella medel inom humanmedicin (2002/77/EG) och av Europaparlamentets resolution av den 23 oktober 2001 om förslaget till denna rådsrekommendation ( KOM(2001)0333 – C5-0411/2001 – 2001/2164(COS) ),
–
med beaktande av kommissionens meddelande av den 20 juni 2001 om en gemenskapsstrategi mot antibiotikaresistens ( KOM(2001)0333 ),
–
A.
Antimikrobiella medel kan förstöra eller hindra tillväxt av bakterier, virus och andra mikroorganismer (antibiotika är mikrobiella medel som endast verkar mot bakterier) och har därför spelat en viktig roll för att förbättra folkhälsan genom att minska antalet dödsfall orsakade av sjukdomar och infektioner som förut inte kunde botas eller var dödliga.
B.
Användningen av dessa medel har lett till att vissa mikroorganismer som förut var känsliga för dessa antimikrobiella medel har utvecklat så kallad antimikrobiell resistens.
C.
Denna naturliga process har accelererats genom överdriven och okontrollerad användning av de antimikrobiella medlen, vilket sätter de uppnådda medicinska framstegen på spel.
D.
E.
F.
Antimikrobiell resistens är en viktig, till stor del olöst fråga, och har blivit ett hot mot folkhälsan i Europa och i hela världen, som leder till längre, mer komplicerade behandlingar, minskad livskvalitet, högre dödlighet (varje år dör 25 000 patienter i EU av en infektion som orsakats av resistenta mikroorganismer), extra sjukvårdskostnader och produktivitetsförluster som uppgår till minst 1,5 miljarder euro årligen.
G.
H.
I.
Olämplig och irrationell användning av antimikrobiella läkemedel skapar gynnsamma villkor för att resistenta mikroorganismer ska dyka upp, spridas och bestå.
J.
Antimikrobiell resistens hos människor beror ofta på olämpliga doser av antibiotika, felaktig behandling och på att patogener konstant exponeras för antimikrobiella medel på sjukhus.
K.
God hygien i form av effektiv tvättning och torkning av händerna kan minska behovet av antibiotika och antimikrobiella medel.
L.
M.
God djurhållningspraxis minimerar behovet av antibiotika.
N.
Åtgärder mot resistens mot antimikrobiella medel i humanläkemedel kan därför inte diskuteras isolerat från åtgärder för att bekämpa resistens mot antimikrobiella medel inom veterinärläkemedel, djurfoder och växtodling.
O.
Epruma European Platform for the Responsible Use of Medicines in Animals.
P.
Antimikrobiell resistens är en företeelse som helt klart har gränsöverskridande konsekvenser och man kan inte utesluta effekter inom andra områden, som högst sannolikt inte skulle vara hanterbara med nuvarande resurser och kunskaper och kan leda till oförutsedda medicinska, sociala och ekonomiska bakslag.
1.
Europaparlamentet är bekymrat över att antimikrobiell resistens, trots de åtgärder som vidtas på europeisk och internationell nivå, utgör ett allt större hot mot folkhälsan i Europa och i hela världen.
2.
Europaparlamentet efterlyser ytterligare upptrappning av kampen mot resistens mot antimikrobiella medel i läkemedel, och att man i följande prioritetsordning ska fokusera på:
–
Återhållsam användning av antimikrobiella medel både när det gäller människor och djur, och att man därvid säkerställer att de endast används när de verkligen behövs för själva sjukdomsbehandlingen och att doseringen, doseringsintervallet och behandlingstiden stämmer.
–
Övervakning och kontroll av antimikrobiell resistens.
–
Behovet av forskning om och utveckling av nya antimikrobiella medel och alternativ.
–
Kopplingar till åtgärder för att bekämpa resistens mot antimikrobiella medel i veterinärläkemedel, djurfoder och växtodling.
3.
Europaparlamentet uppmanar kommissionen att utan dröjsmål föreslå en lagstiftningsram för åtgärder mot antimikrobiell resistens genom att främja initiativ för ansvarsfull användning och stödja spridningen av och information om dessa.
Återhållsam användning av antimikrobiella medel
4.
Europaparlamentet bekräftar än en gång att det behövs brådskande åtgärder för att undvika, eller till och med vända, den ytterligare ökningen av resistenta mikroorganismer, genom att minska onödig och oriktig användning av antimikrobiella medel.
5.
Europaparlamentet understryker att det huvudsakliga målet är att bevara antimikrobiella medel som ett effektivt verktyg för att bekämpa sjukdomar, både hos djur och hos människor, samtidigt som användningen av antimikrobiella medel begränsas till det absolut nödvändiga.
6.
Europaparlamentet konstaterar att det i en rapport om genomförandet av rådets rekommendation Kommissionens arbetsdokument, tillhörande dokument till Andra rapporten från Kommissionen till Rådet på grundval av medlemsstaternas rapporter om genomförandet av Rådets rekommendation (2002/77/EG) om återhållsam användning av antimikrobiella medel inom humanmedicin.
från 2001 och i en Eurobarometer-undersökning från 2010 fastställdes en rad brister och luckor i stödet till återhållsam användning av mikrobiella medel.
7.
Europaparlamentet konstaterar att det fortsätter att finnas skillnader inom unionen när det gäller graden av tillgång till information om antimikrobiell resistens och effekterna på medborgarnas konsumtionsmönster, särskilt med avseende på genomförandet av lagstiftning om obligatorisk receptbeläggning av antibiotika, eftersom procentandelen antibiotika som sålts receptfritt 2008 visat sig variera avsevärt mellan medlemsstaterna.
8.
Europaparlamentet påpekar att när det gäller denna företeelse är Europa inte starkare än den svagaste länken, och därför bör länder med höga nivåer av antimikrobiell resistens ägnas särskild uppmärksamhet.
9.
10.
Europaparlamentet är medvetet om att det förekommer många missuppfattningar om antibiotika och deras effekter och att 53 procent av européerna fortfarande tror att antibiotika dödar virus och 47 procent tror att de hjälper mot förkylningar och influensa, enligt en undersökning som kommissionen låtit utföra (Eurobarometerundersökningen ”Special Eurobarometer 338 on Antimicrobial Resistance” från april 2010).
11.
Europaparlamentet framhäver att patienters brist på efterlevnad när det gäller recept, t.ex. att strunta i att fullfölja behandlingen eller att inte följa rekommendationer för dosering, bidrar stort till antimikrobiell resistens.
12.
Europaparlamentet uppmanar kommissionen att utreda frågan om oriktig användning och försäljning av antimikrobiella medel med eller utan recept längs hela kedjan – från läkaren och farmaceuten till patienten – och att undersöka samtliga inblandade aktörers beteende och genomföra en bred strategi på lång sikt om hur medvetna alla dessa aktörer är.
13.
Europaparlamentet understryker att inom ramen för återhållsam användning av antimikrobiella medel bör de berörda aktörerna uppmärksamma bättre användning av sådana antibiotika som för närvarande finns tillgängliga, genom att noga granska dosering, behandlingstid och läkemedelskombinationer.
14.
Europaparlamentet uppmanar kommissionen och medlemsstaterna att främja god tvättning och torkning av händerna – särskilt på sjukhus – för att förebygga spridning av infektioner och minska behovet av antibiotika.
15.
Europaparlamentet ser därför positivt på den årliga europeiska antibiotikadagen som infaller den 18 november, vars syfte är att öka kunskaperna om det hot mot folkhälsan som antimikrobiell resistens utgör och uppmana till en mer ansvarstagande användning av antibiotika, genom att vidta ett flertal åtgärder i medlemsstaterna.
Övervakning och kontroll av antimikrobiell resistens
16.
17.
18.
Europaparlamentet understryker vikten av diagnostik i kampen mot antimikrobiell resistens och uppmanar till större investeringar på detta område samt en effektivare och bättre användning av gängse diagnostiska verktyg.
19.
Europaparlamentet uppmanar kommissionen, Europeiska centrumet för förebyggande och kontroll av sjukdomar (ECDC) och andra berörda EU-organ att utan dröjsmål föreslå ett harmoniserat och integrerat system för övervakning av antimikrobiell resistens (Antimicrobial Resistance Surveillance System) och antimikrobiell användning i Europa, som inbegriper tidig varning för nya mekanismer för resistens och nya resistenta stammar.
Behovet av forskning om och utveckling av nya antimikrobiella medel och alternativ
20.
Europaparlamentet erkänner att den växande klyftan mellan frekvensen infektioner orsakade av resistenta mikroorganismer och nedgången inom forskning och utveckling av nya antimikrobiella medel nu hotar att kasta folkhälsosektorn tillbaks till tiden före antibiotika.
21.
Europaparlamentet anser att nedgången inom forskning och utveckling orsakats av att marknadsmekanismerna slutat fungera och uppmanar kommissionen att, genom lagstiftning och andra typer av åtgärder, lägga fram förslag om att inrätta eller förbättra incitament för läkemedelsbranschen att trappa upp investeringar i forskning och utveckling av nya antimikrobiella medel och av eventuella alternativ.
22.
Europaparlamentet upprepar att det behövs mer forskning om nya antimikrobiella medel liksom om eventuella alternativ inom EU:s ramprogram för forskning och uppmuntrar till gemensam forskning på EU-nivå som kan leda till effektivitetsökning.
23.
Europaparlamentet påpekar att avsaknaden av snabb diagnostik har bidragit till både överanvändning av antibiotika och ökade utvecklingskostnader.
24.
Europaparlamentet erkänner behovet av att främja kompletterande åtgärder, såsom användningen av effektiva vacciner för att förebygga infektioner, i enlighet med rådets slutsatser av den 1 december 2009 om innovativa incitament till effektiva antibiotika.
Helhetssyn
25.
Europaparlamentet uppmanar kommissionen att se till att åtgärder avseende antimikrobiell resistens och folkhälsa ingår i en helhetssyn på antimikrobiell resistens, och är medvetet om kopplingarna till åtgärder för att bekämpa resistens mot antimikrobiella medel i veterinärläkemedel, djurfoder och växtodling, särskilt med tanke på risken för korsöverföring.
26.
Europaparlamentet uppmanar kommissionen att ta itu med bristen på information om användningen av antibiotika inom veterinärläkemedel över hela EU genom att samla in jämförbara artspecifika uppgifter av hög kvalitet för varje medlemsstat.
27.
Europaparlamentet välkomnar ansträngningarna att anpassa och förbättra den lagstadgade bedömningen av nya antibiotika.
28.
Europaparlamentet uppmanar kommissionen att fortsätta stödja EARRS och Esvac i fråga om uppgiftsinsamling om användningen av antibiotika som en grund för framtida åtgärder för att säkerställa ansvarsfull användning.
29.
Europaparlamentet uppmanar kommissionen att lägga fram lagstiftningsförslag om att avveckla användning av antibiotika som profylax inom djuruppfödning.
30.
Europaparlamentet betonar att sektorerna för djurproduktion och intensiv fiskodling bör inrikta sig på att förebygga sjukdomar genom god hygien, bra anläggningar att hålla djuren i och god djurhållning samt strikta biosäkerhetsåtgärder, snarare än att använda antibiotika profylaktiskt.
31.
32.
33.
34.
Europaparlamentet anser att användning av antibiotika av typen ”sista utvägen”, som riktar sig mot problematiska patogener hos människor, bör tillåtas inom jordbruket endast på licens i kombination med övervakning av resistens, företrädesvis utifrån en bedömning från fall till fall.
Internationellt samarbete
35.
36.
Europaparlamentet uppmanar kommissionen att se till att tillräckliga ekonomiska och mänskliga resurser finns tillgängliga för att genomföra de aktuella strategierna.
o
o o
37.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet och kommissionen.
P7_TA-PROV(2011)0586
Utvidgning av bestämmelserna i partnerskaps- och samarbetsavtalet EG/Uzbekistan till att omfatta bilateral handel med textilprodukter
A7-0427/2011
Europaparlamentets resolution av den 15 december 2011 om förslaget till rådets beslut om ingående av ett protokoll till avtalet om partnerskap och samarbete som upprättar ett partnerskap mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Republiken Uzbekistan, å andra sidan, vilket utvidgar bestämmelserna i partnerskaps- och samarbetsavtalet till att omfatta bilateral handel med textilprodukter, med hänsyn till att det bilaterala avtalet om handel med textilprodukter löper ut (16384/2010 – C7-0097/2011 – 2010/0323(NLE))
Europaparlamentet utfärdar denna resolution,
–
med beaktande av förslaget till rådets beslut (16384/2010),
–
–
med beaktande av sina tidigare resolutioner av den 15 november 2007 EUT C 282 E, 6.11.2008, s.
478.
, av den 26 oktober 2006 EUT C 313 E, 20.12.2006, s.
466.
om Uzbekistan, av den 12 mars 1999 om partnerskaps- och samarbetsavtalet mellan EU och Uzbekistan EGT C 175 E, 21.06.1999, s.
432.
, av den 8 juni 2011 om den yttre dimensionen av socialpolitiken, främjande av arbetsnormerna och de sociala normerna och de europeiska företagens sociala ansvar Antagna texter, P7-TA(2011) 0260.
och av den 25 november 2010 om mänskliga rättigheter samt sociala normer och miljönormer i internationella handelsavtal Antagna texter, P7-TA(2010) 0434.
,
–
med beaktande av avtalet mellan Europeiska ekonomiska gemenskaperna och Uzbekistan om handel med textilprodukter EGT L 123, 17.5.1994, s.
745.
och rådets beslut 2000/804/EG av den 4 december 2000 om ingående av avtal om handel med textilprodukter med vissa tredje länder (däribland Uzbekistan) EGT L 326, 22.12.2000, s.
63.
,
–
med beaktande av avtalet om partnerskap och samarbete som upprättar ett partnerskap mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Republiken Uzbekistan, å andra sidan EGT L 229, 31.8.1999, s.
–
med beaktande av rådets slutsatser om Uzbekistan, exempelvis av den 25 oktober 2010 http://www.consilium.europa.eu/uedocs/cms_data/docs/pressdata/EN/foraff/117329.pdf
, av den 27 oktober 2009 http://www.consilium.europa.eu/uedocs/cms_data/docs/pressdata/en/gena/110783.pdf
, av den 16 december 2008 http://ec.europa.eu/sport/information-center/doc/timeline/european_council_12-12-2008_conclusions_en.pdf
, av den 27 oktober 2008 http://www.consilium.europa.eu/uedocs/cms_data/docs/pressdata/en/gena/110783.pdf
, av den 13 oktober 2008 http://www.consilium.europa.eu/uedocs/cmsUpload/103295.pdf
och av den 29 april 2008 http://www.eu2008.si/si/News_and_Documents/Council_Conclusions/April/0428_GAERC4.pdf
, i vilka frågor som rör mänskliga rättigheter, demokratisering och rättsstatliga principer i in Uzbekistan togs upp,
–
med beaktande av de avslutande iakttagelserna av FN:s kommitté för mänskliga rättigheter (2005 Kontoret för FN:s högkommissarie för mänskliga rättigheter, konventionsförkortning: CCPR.
26/04/2005.
)), http://www.unhchr.ch/tbs/doc.nsf/(Symbol)/CCPR.CO.83.UZB.En?Opendocument
Avslutande iakttagelser av kommittén för mänskliga rättigheter, Uzbekistan
, www2.ohchr.org/english/bodies/hrc/docs/co/Uzbekistan98_AUV.doc)
), de avslutande iakttagelserna av FN:s kommitté för ekonomiska, sociala och kulturella rättigheter (2006) http://www.unhchr.ch/tbs/doc.nsf/%28Symbol%29/E.C.12.UZB.CO.1.En?Opendocument
, de avslutande iakttagelserna av kommittén för avskaffande av diskriminering av kvinnor (2010) Förenta nationerna, konvention om avskaffande av alla former av diskriminering av kvinnor, CEDAW/C/UZB/CO/4, Distr.: General 5 februari 2010.
Avslutande iakttagelser av kommittén om avskaffande av diskriminering av kvinnor, Uzbekistan,
(http://www2.ohchr.org/english/bodies/cedaw/docs/co/CEDAW-C-UZB-CO-4.pdf)
, de avslutande iakttagelserna av FN:s kommitté för barnets rättigheter (2006) Kontoret för FN:s högkommissarie för mänskliga rättigheter, kommittén för barnets rättigheter,
avslutande iakttagelser: Uzbekistan.
02/06/2006.
(CRC/C/UZB/CO/2.
), (http://www.unhchr.ch/tbs/doc.nsf/(Symbol)/CRC.C.UZB.CO.2.En?Opendocument)
, rapporten från arbetsgruppen för allmän regelbunden översyn av Uzbekistan (2009) http://lib.ohchr.org/HRBodies/UPR/Documents/Session3/UZ/A_HRC_10_82_Add1_Uzbekistan_E.pdf
), rapporten från ILO:s expertkommitté för tillämpning av konventioner och rekommendationer avseende konventionen om de värsta formerna av barnarbete (2010 Internationella arbetskonferensen, 99:e sammanträdet, 2010, Rapport från expertkommittén för tillämpning av konventioner och rekommendationer, (http://www.ilo.org/wcmsp5/groups/public/@ed_norm/@relconf/documents/meetingdocument/wcms_123424.pdf)
och 2011 Internationella arbetskonferensen, 100:e sammanträdet, 2011, Rapport från expertkommittén för tillämpning av konventioner och rekommendationer (ILC.
100/III/1A), (http://www.ilo.org/wcmsp5/groups/public/@ed_norm/@relconf/documents/meetingdocument/wcms_151556.pdf)
) samt rapporten från ILO:s expertkommitté för tillämpning av konventioner och rekommendationer avseende konventionen om avskaffande av tvångsarbete (2010 http://www.ilo.org/wcmsp5/groups/public/@ed_norm/@relconf/documents/meetingdocument/wcms_123424.pdf
och 2011 http://www.ilo.org/wcmsp5/groups/public/@ed_norm/@relconf/documents/meetingdocument/wcms_151556.pdf
), som alla uttrycker oro över den fortsatta användningen av barnarbete i Uzbekistan,
–
med beaktande av kommissionens meddelande ”Anständigt arbete för alla – EU:s bidrag till agendan för anständigt arbete i världen” ( KOM(2006)0249 ),
–
med beaktande av kommissionens meddelande ”En särskild plats för barnen i EU:s yttre åtgärder” ( KOM(2008)0055 ) samt Europeiska kommissionens arbetsdokument om bekämpning av barnarbete ( SEK(2010)0037 ),
–
med beaktande av rådets slutsatser om barnarbete av den 14 juni 2010 och dess ”uppmaning till kommissionen att studera och före 2011 års utgång rapportera om de värsta formerna av barnarbete och handel, med hänsyn till internationell erfarenhet och yttrandena från behöriga internationella organisationer” Europeiska unionens råd, rådets slutsatser om barnarbete, 3023:a sammanträdet i rådet (urtrikesfrågor), Luxemburg den 14 juni 2010, (http://www.consilium.europa.eu/uedocs/cms_data/docs/pressdata/EN/foraff/115180.pdf)
,
–
, vilka ratificerades av Uzbekistan 2009 respektive 2008 och som följdes av antagandet av en nationell handlingsplan i Uzbekistan,
–
med beaktande av artikel 15 i rådets förordning (EG) nr 732/2008 av den 22 juli 2008 om tillämpning av Allmänna preferenssystemet under perioden 1 januari 2009 – 31 december 2011 EUT L 211, 6.8.2008 s.
1.
samt artikel 19 i förslaget till Europaparlamentets och rådets förordning om tillämpning av ett system med allmänna tullpreferenser ( KOM(2011)0241 ),
–
med beaktande av uppmaningar av olika icke-statliga organisationer Business Social Compliance Initiative, C.W.F Children Worldwide Fashion, Anti-Slavery International, Uzbek-German Forum for Human Rights and Ethical Trading Initiative.
och av fackföreningar ITUC-ETUC.
om utredningar avseende de allmänna preferenserna för Uzbekistan,
–
med beaktande av det vägledande DCI-programmet för Centralasien 2011–2013 Europeiska kommissionen, generaldirektoratet för yttre förbindelser, direktoratet för Östeuropa, södra Kaukasus, centralasiatiska republiker, vägledande DCI-program 2011–2013, s.
54, (http://www.eeas.europa.eu/central_asia/docs/2010_ca_mtr_en.pdf)
,
–
–
med beaktande av interimsbetänkandet från utskottet för internationell handel och yttrandet från utskottet för utrikesfrågor ( A7-0427/2011 ), och av följande skäl:
a.
Textilprodukter är undantagna från partnerskaps- och samarbetsavtalet och reglerades i stället genom ett bilateralt avtal som upphörde att gälla 2005, vilket skapar en rättsosäkerhet för EU:s exportörer, eftersom Uzbekistan (som inte är medlem i WTO) har friheten att höja sina importtullar, medan EU behandlar alla länder i världen som mest gynnad nation (i fråga om tullar).
b.
Syftet med detta protokoll är att inkludera textilprodukter i partnerskaps- och samarbetsavtalet, vilket kommer att leda till att båda parterna beviljar varandra status som mest gynnad nation, vilket gör att det oklara rättsläget upphör för EU:s textilexportörer.
c.
EU har tidigare avhjälpt detta oklara rättsläge för EU:s textilexportörer genom ändringar av partnerskaps- och samarbetsavtal med olika länder (exempelvis Azerbajdzjan 2007 och Kazakstan 2008).
d.
I artikel 2 i avtalet om partnerskap och samarbete med Uzbekistan fastställs att ”respekten för demokratin, den internationella rättens principer och de mänskliga rättigheterna, såsom de definieras särskilt i Förenta nationernas stadga, Helsingforsslutakten och Parisstadgan för ett nytt Europa samt för de marknadsekonomiska principerna, inbegripet dem som uppställs i handlingarna från ESK-konferensen i Bonn, ligger till grund för parternas inrikes- och utrikespolitik och utgör väsentliga beståndsdelar i partnerskapet och i detta avtal”.
e.
Rådet uppgav den 25 oktober 2010 att det ”fortfarande är allvarligt bekymrat över den övergripande situationen när det gäller mänskliga rättigheter, demokratisering och rättsstatliga principer i Uzbekistan”.
f.
Den uzbekistanska regeringen tar viktiga steg för att uppnå demokrati.
g.
Den uzbekistanska regeringen handlar i strid med slutsatserna från ministermötet mellan Europeiska unionen och Centralasien i Tasjkent den 7 april 2011, där parterna erinrade om att utveckling av ett starkt civilsamhälle utgör en integrerad del av demokratiutvecklingen.
h.
Uzbekistan ärvde och behöll ett i stort sett oreformerat statligt drivet jordbrukssystem, medan andra länder i samma region, exempelvis Kazakstan och i mindre utsträckning Tadzjikistan, moderniserar sitt jordbruk och åtgärdar många av problemen What has changed?
En verklig reform och mekanisering av jordbruket skulle göra det möjligt att betydligt minska mängden tvångsarbete för barn och slöseriet med vatten samt göra jordbruket mer lönsamt.
i.
Uzbekistanska jordbrukare kan officiellt vara fria aktörer, men de arrenderar sin mark, köper sitt gödningsmedel och är skyldiga att uppfylla kvoter, allt från regeringen, medan regeringen köper sin bomull till fasta priser och tjänar betydande summor på försäljning av bomull till det mycket högre världsmarknadspriset.
j.
Rådets ordförandeskap erinrade i EU:s uttalande vid ILO i juni 2011 om ”de väldokumenterade påståendena och den breda enigheten bland Förenta nationernas organ, Unicef, representantorganisationerna för arbetsgivare och arbetstagare och ickestatliga organisationer, och uppgav att trots de juridiska åtagandena av Uzbekistans regering om att utrota tvångsarbete för barn tvingas i praktiken uppskattningsvis mellan 0,5 och 1,5 miljoner barn i skolåldern år efter år att delta i det farliga arbetet i bomullsskörden i upp till tre månader varje år”.
k.
Skolorna är stängda under skördeperioden på hösten, vilket hämmar utbildningen.
l.
Barn, deras lärare och föräldrar riskerar att straffas om de inte lyder.
m.
Uzbekistans regering har uppgett att ”det är tradition att äldre barn hjälper till i familjeföretagen” och att ”påståendena om utbrett tvångsarbete i jordbruket saknar grund” ILO-rapport 2011 från expertkommittén för tillämpning av konventioner och rekommendationer, s.
429, (http://www.ilo.org/wcmsp5/groups/public/@ed_norm/@relconf/documents/meetingdocument/wcms_151556.pdf)
.
n.
Oberoende internationella observatörer har samlat in bevis för att tvångsarbete, särskilt tvångsarbete för barn, är systematisk och organiserad praxis, och innebär press på lärare och familjer samt polisens och säkerhetsstyrkornas medverkan.
o.
Den uzbekistanska regeringen har hittills vägrat att ge tillträde för oberoende övervakningsuppdrag för att få fram fakta och informera om längden på höstens skördeperiod, arbetshälsovillkoren för skolelever, hur gamla de är och vilka eventuella bestraffningar de hotas av om de inte lyder.
p.
Enligt kommissionen står EU:s textil- och klädexport till Uzbekistan för 0,05 procent av EU:s textil- och klädexport.
q.
EU är en av de viktigaste importörerna av bomull från Uzbekistan, och denna import beräknas ha uppgått till mellan 6 Källa: Europeiska kommissionen GD Handel och
och 23 http://unctad.org/infocomm/anglais/cotton/market.htm
procent av den uzbekistanska bomullsexporten de senaste tio åren.
r.
s.
Rättvis och öppen internationell handel kräver konkurrens på lika villkor och de ekonomiska faktorer som avgör priset på produkter som exporteras till EU bör inte snedvridas av seder som strider mot de grundläggande principerna om mänskliga rättigheter och barnets rättigheter.
t.
Många textilförsäljare, däribland europeiska, har beslutat att de inte längre ska köpa bomull från Uzbekistan och att de kommer att underrätta alla sina leverantörer om detta åtagande Internationellt forum om arbetsrätt, http://www.laborrights.org/stop-child-forced-labor/cotton-campaign/company-response-to-forced-child-labor-in-uzbek-cotton)
.
u.
Rådet uppgav i sina slutsatser om barnarbete av den 14 juni 2010 att det är fullt medvetet om EU:s roll och ansvar i kampen för att få barnarbete att upphöra.
v.
Kommissionens ordförande José Manuel Barroso har uppmanat den uzbekistanske presidenten, Islam Karimov, att tillåta ett ILO-övervakningsuppdrag i landet för att ta upp frågan om barnarbetsseder som eventuellt kvarstår Uttalande av Europeiska kommissionens ordförande José Manuel Barroso efter hans möte med Uzbekistans president Islam Karimov, (http://europa.eu/rapid/pressReleasesAction.do?reference=MEMO/11/40&type=HTML)
.
w.
EU:s stöd till Uzbekistan inom ramen för EU:s strategi för Centralasien har hittills inte uppmärksammat jordbruksreformer i högre grad.
x.
Kommissionen insisterar också kraftigt på att ILO:s övervakningsuppdrag ska vara det enda relevanta övervakningsorganet i samband med undersökningar av ett tillfälligt återtagande av referenser till det allmänna preferenssystemet, och kommissionens förslag att avskaffa detta krav inom ramen för översynen av förordningen om det allmänna preferenssystemet välkomnas.
y.
1.
Europaparlamentet begär att rådet och kommissionen ska ta följande rekommendationer i beaktande:
i)
Fördöm kraftfullt användningen av tvångsarbete för barn i Uzbekistan.
ii)
Ge starkt stöd åt ILO:s krav på Uzbekistans regering att acceptera ett observatörsuppdrag med tre parter på hög nivå, vilket skulle ha full rörelsefrihet och snabbt tillträde till alla platser och relevanta parter, däribland på bomullsfälten, för att bedöma ILO-konventionens genomförande.
iii)
Förklara vikten av utländska observatörer för att övervaka utvecklingen av tvångsarbetssituationen i Uzbekistan och andra länder i regionen.
iv)
Uppmana enträget Uzbekistans president Islam Karimov att tillåta en övervakningsdelegation från ILO att besöka landet för att undersöka frågan om tvångsarbete för barn.
v)
Uppmana Uzbekistans regering att ta emot en övervakningsdelegation från ILO och se till att användningen av tvångsarbete för barn och annat tvångsarbete verkligen är på väg att upphöra på nationell, regional och lokal nivå.
vi)
Påminn de uzbekistanska myndigheterna om att trots att principerna om respekt för mänskliga rättigheter ingår i Republiken Uzbekistans författning, och att Uzbekistan har undertecknat och ratificerat de flesta FN-konventioner avseende mänskliga rättigheter, medborgerliga och politiska rättigheter och barnets rättigheter, återstår fortfarande den faktiska tillämpningen av denna formella uppsättning rättsakter.
vii)
viii)
ix)
Kommissionen bör undersöka och, om så är lämpligt, lägga fram ett lagstiftningsförslag för Europaparlamentet om en effektiv spårbarhetsmekanism för de varor som framställs genom tvångsarbete för barn.
x)
Stöd parlamentets krav på bomullshandlare och återförsäljare av bomull att avstå från att köpa bomull från Uzbekistan som framställts genom tvångsarbete för barn och att underrätta konsumenter och alla leverantörer om detta åtagande.
xi)
xii)
Förklara hur viktiga förbindelserna mellan unionen och Uzbekistan är, grundade på partnerskaps- och samarbetsavtalet och dess demokratiska principer och människorättsprinciper, och påminn om unionens löften om ytterligare och fördjupade bilaterala förbindelser, vilka inbegriper handel liksom alla områden med koppling till demokratiska principer, respekt för humanitära och grundläggande rättigheter samt rättsstatsprincipen.
xiii)
Bidra aktivt till förbättringen av de sociala, ekonomiska och mänskliga rättigheterna för befolkningen i Uzbekistan genom att främja ett tillvägagångssätt som utgår från gräsrotsnivå och genom att stödja civilsamhällets organisationer och medierna för att åstadkomma en hållbar demokratiseringsprocess.
xiv)
Förse regelbundet parlamentet med betydande information om situationen i Uzbekistan, i synnerhet när det gäller avskaffandet av tvångsarbete för barn.
2.
Sammanfattningsvis konstaterar Europaparlamentet att man inte kommer att ge sitt godkännande förrän ILO-observatörer getts tillstånd av de uzbekistanska myndigheterna att göra en noggrann granskning utan att hindras, och har bekräftat att konkreta reformer har genomförts och gett påtagliga resultat på ett sådant sätt att praxis med tvångsarbete för barn och annat tvångsarbete i praktiken är på väg att avskaffas på nationell, regional och lokal nivå.
3.
Europaparlamentet uppdrar åt talmannen att begära ytterligare diskussioner med kommissionen och rådet.
4.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet och kommissionen samt Uzbekistans regering och parlament.
P7_TA-PROV(2012)0003
En gemenskapskodex om viseringar ***I
A7-0441/2011
Europaparlamentets lagstiftningsresolution av den 19 januari 2012 om förslaget till Europaparlamentets och rådets förordning om ändring av förordning (EG) nr 810/2009 av den 13 juli 2009 om införande av en gemenskapskodex om viseringar (viseringskodex) ( KOM(2011)0516 – C7-0226/2011 – 2011/0223(COD) )
(Ordinarie lagstiftningsförfarande: första behandlingen)
Europaparlamentet utfärdar denna resolution
–
med beaktande av kommissionens förslag till Europaparlamentet och rådet ( KOM(2011)0516 ),
–
–
–
–
med beaktande av artikel 55 i arbetsordningen,
–
med beaktande av betänkandet från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor ( A7-0441/2011 ).
1.
Europaparlamentet antar nedanstående ståndpunkt vid första behandlingen.
2.
Europaparlamentet uppmanar kommissionen att lägga fram en ny text för parlamentet om den har för avsikt att väsentligt ändra sitt förslag eller ersätta det med ett nytt.
3.
Europaparlamentet uppdrar åt talmannen att översända parlamentets ståndpunkt till rådet, kommissionen och de nationella parlamenten.
P7_TC1-COD(2011)0223
Europaparlamentets ståndpunkt fastställd vid första behandlingen den 19 januari 2012 inför antagandet av Europaparlamentets och rådets förordning (EU) nr .../2012 om ändring av förordning (EG) nr 810/2009 om införande av en gemenskapskodex om viseringar (viseringskodex)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
efter översändande av utkastet till lagstiftningsakt till de nationella parlamenten,
i enlighet med det ordinarie lagstiftningsförfarandet Europaparlamentets ståndpunkt av den 19 januari 2012.
, och
av följande skäl: (1)
Det är nödvändigt att förtydliga reglerna om transitering genom det internationella transitområdet på flygplatser för att säkerställa rättssäkerhet och öppenhet.
(2)
1.
, som innehar en giltig visering som utfärdats av en medlemsstat, Kanada, Japan eller Förenta staterna, eller som innehar ett giltigt uppehållstillstånd som utfärdats av en medlemsstat, Andorra, Kanada, Japan, San Marino eller Förenta staterna är undantagna från kravet på visering för flygplatstransitering.
(3)
I fråga om personer som innehar en giltig visering bör undantaget gälla när de reser till det utfärdande landet eller till ett annat tredjeland, och när de återvänder från det utfärdande landet efter att ha använt viseringen.
(4)
Eftersom målet för denna förordning, nämligen att förtydliga reglerna om transitering genom det internationella transitområdet på flygplatser, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna och det därför bättre kan uppnås på unionsnivå, kan unionen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget om Europeiska unionen.
I enlighet med proportionalitetsprincipen i samma artikel går denna förordning inte utöver vad som är nödvändigt för att uppnå detta mål.
(5)
36.
31.
.
(6)
52.
1.
.
(7)
21.
19.
.
(8)
(9)
43.
.
(10)
Irland deltar därför inte i antagandet av denna förordning, som inte är bindande för eller tillämplig på Irland.
(11)
i 2003 års anslutningsakt.
(12)
i 2005 års anslutningsakt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
b)
c)
Artikel 2
Europeiska unionens officiella tidning
.
Denna förordning är till alla delar bindande och direkt tillämplig i medlemsstaterna i enlighet med fördragen.
Utfärdad i
På Europaparlamentets vägnar På rådets vägnar
Ordförande Ordförande
P7_TA-PROV(2012)0042
Utdelning av livsmedel till de sämst ställda i unionen ***II
A7-0032/2012
Europaparlamentets lagstiftningsresolution av den 15 februari 2012 om rådets ståndpunkt vid första behandlingen inför antagandet av Europaparlamentets och rådets förordning om ändring av rådets förordningar (EG) nr 1290/2005 och (EG) nr 1234/2007 vad gäller utdelning av livsmedel till de sämst ställda i unionen (18733/1/2011 – C7-0022/2012 – 2008/0183(COD) )
(Ordinarie lagstiftningsförfarande: andra behandlingen)
–
med beaktande av rådets ståndpunkt vid första behandlingen (18733/1/2011 – C7-0022/2012 ),
–
med beaktande av de motiverande yttranden från det danska folketinget, Sveriges riksdag och Förenade kungarikets överhus som lagts fram i enlighet med protokoll (nr 2) om tillämpning av subsidiaritets- och proportionalitetsprinciperna, och enligt vilka utkastet till lagstiftningsakt inte är förenligt med subsidiaritetsprincipen,
–
med beaktande av yttrandena från Europeiska ekonomiska och sociala kommittén av den 20 januari 2011 EUT C 84, 17.3.2011, s.
49.
och den 8 december 2011 Ännu ej offentliggjorda i EUT.
,
–
med beaktande av yttrandet från Regionkommittén av den 27 januari 2011 EUT C 104, 2.4.2011, s.
44.
,
–
med beaktande av sin ståndpunkt av den 26 mars 2009 EUT C 117 E, 6.5.2010, s.
258.
,
–
,
–
med beaktande av de ändrade förslagen från kommissionen ( COM(2010)0486 ) och COM(2011)0634 ),
–
–
med beaktande av artikel 72 i arbetsordningen,
–
med beaktande av andrabehandlingsrekommendationen från utskottet för jordbruk och landsbygdens utveckling ( A7-0032/2012 ).
1.
Europaparlamentet godkänner rådets ståndpunkt vid första behandlingen.
2.
Europaparlamentet konstaterar att rättsakten är antagen i enlighet med rådets ståndpunkt.
3.
4.
5.
Europaparlamentet uppdrar åt talmannen att översända parlamentets ståndpunkt till rådet, kommissionen och de nationella parlamenten.
P7_TA-PROV(2012)0046
Möjligheten att införa stabilitetsobligationer
B7-0016/2012
Europaparlamentets resolution av den 15 februari 2012 om möjligheten att införa stabilitetsobligationer ( 2011/2959(RSP) )
Europaparlamentet utfärdar denna resolution
–
med beaktande av Europaparlamentets och rådets förordning (EU) nr 1173/2011 av den 16 november 2011 om effektiv övervakning av de offentliga finanserna i euroområdet EUT L 306, 23.11.2011, s.
1.
, som är en del av den så kallade ”six-pack”,
–
med beaktande av kommissionens grönbok av den 23 november 2011 om möjligheten att införa stabilitetsobligationer,
–
med beaktande av presentationen av den 23 november 2011 av kommissionens vice ordförande Olli Rehn i utskottet för ekonomi och valutafrågor och av diskussionerna av den 29 november 2011 med det tyska rådet av ekonomiska experter om en europeisk skuldinlösenfond,
–
med beaktande av Europeiska rådets ordförande Herman Van Rompuys interimsrapport av den 6 december 2011: Mot en starkare ekonomisk union,
–
A.
Parlamentet har begärt att kommissionen ska lägga fram en rapport om möjligheten att införa eurovärdepapper.
B.
Situationen i euroområdet är unik, eftersom länderna i euroområdet har samma valuta men saknar en gemensam skattepolitik och en gemensam obligationsmarknad.
C.
Emissionen av obligationer med solidariskt ansvar skulle kräva en djupare integrationsprocess.
1.
Europaparlamentet är mycket oroat över de fortsatta spänningarna på euroområdets statsobligationsmarknader, vilket återspeglats i större spreadar, hög volatilitet och sårbarhet för spekulativa attacker under de två senaste åren.
2.
Europaparlamentet anser att euroområdet, som ger ut världens andra internationella valuta, är medansvarig för det internationella valutasystemets stabilitet.
3.
Europaparlamentet understryker att det ligger i euroområdets och medlemsstaternas långsiktiga intresse att utnyttja alla fördelar med att ge ut euron, som har förutsättning att bli en internationell reservvaluta.
4.
5.
Europaparlamentet anser också att euroområdet och medlemsstaterna bär ansvaret för att en valuta som används av mer än 330 miljoner människor och många företag och investerare är stabil på lång sikt, något som indirekt påverkar resten av världen.
6.
7.
8.
Europaparlamentet tar del av kommissionens bedömning, som utgör en del av kommissionens grönbok om möjligheten att införa stabilitetsobligationer, att stabilitetsobligationer skulle underlätta penningpolitiken i euroområdet och även effektivisera statsobligationsmarknaden och det finansiella systemet i hela euroområdet.
9.
10.
Europaparlamentet anser att de mål som ligger till grund för besluten i Europeiska rådet av den 8–9 december 2011 om att ytterligare stärka de offentliga finansernas hållbarhet också bidrar till att skapa nödvändiga villkor för ett eventuellt införande av stabilitetsobligationer.
11.
–
Effektiva marknadsincitament för att minska skulderna.
–
Kriterier för inträde och utträde, överenskommelser om villkor och löptid, omfördelning av finansieringsfördelar för de nuvarande AAA-länderna.
–
Ett system för differentiering av räntesatser mellan medlemsstater med olika kreditbetyg.
–
Budgetdisciplin och ökad konkurrenskraft.
–
Procykliska effekter och effekter av skulddeflation.
–
Tillräcklig attraktionskraft för marknadsinvesterare, samtidigt som man är försiktig med eller undviker alltför högt ställda säkerheter eller en omfördelning av riskerna mellan länderna.
–
Förmånsrätt för stabilitetsobligationer i förhållande till nationella obligationer om medlemsstaten inte kan betala sin skuld.
–
Kriterier för tilldelning av lån till medlemsstater och kapaciteten att hantera skulden.
–
Mätbara och genomförbara skuldprogram.
–
Formaliteterna för en bindande färdplan, i likhet med Maastrichtkriterierna för införandet av den gemensamma valutan.
–
Samverkan mellan EFSF och ESM för medlemsstater som har likviditetsproblem.
–
Lämpliga rättsliga krav, inklusive ändringar av fördrag och konstitutioner.
12.
13.
Europaparlamentet påpekar att denna resolution är ett preliminärt svar på kommissionens grönbok och kommer att följas upp av en mer omfattande resolution i form av ett initiativbetänkande.
14.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen och Europeiska centralbanken.
P7_TA-PROV(2012)0062
Framtiden för det europeiska jordövervakningsprogrammet (GMES)
B7-0063/2012
Europaparlamentets resolution av den 16 februari 2012 om framtiden för det europeiska jordövervakningsprogrammet (GMES) ( 2012/2509(RSP) )
–
med beaktande av kommissionens meddelande av den 30 november 2011 om det europeiska jordövervakningsprogrammet (GMES) och dess operationer (från 2014 och framöver) ( COM(2011)0831 ),
–
med beaktande av kommissionens meddelande av den 29 juni 2011 om en budget för Europa 2020 ( COM(2011)0500 ),
–
med beaktande av sin resolution av den 19 januari 2012 om en rymdstrategi för Europeiska unionen i allmänhetens tjänst Antagna texter, P7_TA(2012)0013 .
,
–
med beaktande av rådets slutsatser av den 31 maj 2011 om en rymdstrategi för Europeiska unionen i allmänhetens tjänst,
–
med beaktande av den muntliga frågan av den 13 februari 2012 till kommissionen om framtiden för det europeiska jordövervakningsprogrammet ( O-000025/2012 – B7–0037/2012 ),
–
A.
B.
GMES är politiskt, strategiskt och tekniskt mycket betydelsefullt för Europa och ger god valuta för pengarna sett till de ekonomiska, sociala och tekniska fördelarna.
C.
GMES har utformats som ett unionsprogram under EU:s förvaltning och ansvar, med finansiering från EU:s budget på sammanlagt cirka 3,2 miljarder fram till 2013.
D.
E.
1.
Europaparlamentet beklagar att kommissionen den 30 november 2011 endast offentliggjorde ett meddelande och inte presenterade något lagstiftningsförslag om GMES, med tanke på att nuvarande förordning (EU) nr 911/2010 endast omfattar de inledande operationerna och kommer att löpa ut i slutet av 2013.
2.
3.
Europaparlamentet ser inte en finansiering av GMES utanför den fleråriga budgetramen – med den finansiering och de styrstrukturer som kommissionen föreslår i sitt meddelande – som ett gångbart alternativ.
4.
Europaparlamentet påpekar att en osäkerhet kring GMES-programmets framtid och finansiering är förödande för utvecklingen och introduktionen på marknaden av GMES-tjänster och -tillämpningar, som är tänkta att generera ekonomisk tillväxt och välfärd för EU:s medborgare.
5.
Europaparlament uppmanar därför kommissionen att snabbt lägga fram ett lagstiftningsförslag om en långsiktig styrning, stöd och drift av GMES-programmet, finansierat genom den fleråriga budgetramen, för att programmet ska kunna införas och drivas korrekt samt nå sitt mål som är att vara i full drift från 2014.
6.
Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen samt medlemsstaternas regeringar och parlament.
