10.
Finansiella instrumentet för miljön (LIFE+) (omröstning)
6.
Begränsning av utsläppande på marknaden och användning av perfluoroktansulfonat (omröstning)
8.
Befrielse från mervärdesskatt och punktskatt på varor som införs av resande från tredjeländer (omröstning)
1.
Tjänster på den inre marknaden (omröstning)
Omröstningen är härmed avslutad.
Avslutande av sammanträdet
(Sammanträdet avslutades kl. 23.30.)
5.
Övergångsbestämmelser i fråga om språkordningen (omröstning)
Öppnande av sammanträdet
(Sammanträdet öppnades kl. 9.05.)
Undertecknande av rättsakter som antagits genom medbeslutandeförfarandet: se protokollet
Omröstning
3.
Olagligt fiske (omröstning)
8.
Reformering av den gemensamma organisationen av marknaden för vin (omröstning)
Avtalstexter översända av rådet: se protokollet
Förbud mot produkter som härrör från säl i Europeiska unionen (debatt)
Inkomna dokument: se protokollet
Debatter om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer (debatt)
Avtalstexter översända av rådet: se protokollet
13.
Flerårig plan för torskbestånden i Östersjön och det fiske som utnyttjar de bestånden (omröstning)
- Betänkande: Chmielewski
Inkomna dokument: se protokollet
Öppnande av sammanträdet
(Sammanträdet öppnades kl. 9.05.)
2.
Samordnade åtgärder för att förebygga och begränsa föroreningar (kodifierad version) (omröstning)
- Betänkande: Wallis
9.
Läget i förhandlingarna om rambeslutet om kampen mot rasism och främlingsfientlighet (omröstning)
- Betänkande: Roure
19.
Bulgariens och Rumäniens anslutning till konventionen av den 29 maj 2000 (omröstning)
- Betänkande: Genowefa Grabowska
6.
Uttjänta fordon (kommissionens genomförandebefogenheter) (omröstning)
- Betänkande: Florenz
14.
Demokratisk övervakning inom ramen för instrumentet för samarbete och utveckling (omröstning)
- Resolutionsförslag
Uttalande av talmannen
Avslutande av sammanträdet
(Sammanträdet avslutades kl. 21.45.)
Rättelser till avgivna röster och röstavsikter: se protokollet
(Sammanträdet avbröts kl. 12.25 och återupptogs kl. 15.00.)
Avtalstexter översända av rådet: se protokollet
Föredragningslista för nästa sammanträde: se protokollet
2.
Bulgariens och Rumäniens anslutning till konventionen om tillämplig lag för avtalsförpliktelser, öppnad för undertecknande i Rom den 19 juni 1980 (omröstning)
- Betänkande: Cristian Dumitrescu
Avtalstexter översända av rådet: se protokollet
Fastställande av en ram för markskydd - Temainriktad strategi för markskydd (debatt)
Nästa punkt är den gemensamma debatten om
ett betänkande av Cristina Gutiérrez-Cortines för utskottet för miljö, folkhälsa och livsmedelssäkerhet om förslaget till direktiv för Europaparlamentet och rådet om inrättande av rambestämmelser för markskydd och om ändring av direktiv 2004/35/EG - C6-0307/2006 -, samt
ett betänkande av Vittorio Prodi för utskottet för miljö, folkhälsa och livsmedelssäkerhet om en temainriktad strategi för markskydd.
(DE) Fru talman! Jag skulle inte ha begärt ordet igen om kommissionsledamot Franco Frattini inte försökt spela offer i sina avslutande kommentarer.
Herr kommissionsledamot! Ni måste inse det faktum att ni befinner er i ett europeiskt forum där ni har en specifik skyldighet att vara mycket noga med vad ni säger; och det ni uttalade i intervjun i Il Messaggero var fel i sak.
Ingen myndighet i Europa har rätt att gå in i ett läger och fråga någon: ”Vad gör du för din försörjning?” och deportera vederbörande om han/hon inte svara omedelbart.
Det är fullständigt och totalt fel, men det är just det ni sa i intervjun med Il Messaggero, så bli inte förnärmad när man påpekar det för er.
Den här debatten är avslutad.
Jag beklagar men det är omöjligt.
Jag trodde ni ville lägga till en punkt till dagordningen.
Debatten är avslutad.
Låt oss gå vidare. ...
Jag motsätter mig denna intervention.
Vi kan inte gå vidare i den här frågan, jag trodde att Martin Schulz ville lägga till en punkt till dagordningen.
Fru talman! Låt mig först tacka Europaparlamentet och särskilt föredragandena Cristina Gutiérrez-Cortines och Vittorio Prodi, utskottet för miljö, folkhälsa och livsmedelssäkerhet och övriga utskott för deras bidrag under den första behandlingen.
Kommissionens förslag om on en temainriktad strategi för markskydd härrör från arbete som påbörjades 1998 på initiativ av det tyska miljöministeriet.
Som resultat av långa överläggningar med intresserade parter och med medlemsstaterna har marken erkänts som en värdefull naturresurs och markförstöringen i Europa håller på att bli problematisk.
Kommissionen har därefter samarbetat med de berörda parterna, framför allt med parlamentet och rådet, för att frågor om markskydd ska förstås bättre och samförstånd uppnås inom detta område.
Parlamentets resolution om meddelandet om markskydd från 2002 innehöll viktiga rekommendationer till kommissionen om den inriktning som behövs för att säkerställa lämpligt markskydd i Europa.
Med slutsatserna från Mallorca 2002 gav rådet en uppmaning till kommissionen att föreslå en heltäckande, långtgående strategi beträffande markskydd. Uppmaningen omfattade generella principer, lämpliga kvantitativa och kvalitativa mål och tidtabeller för bedömning och utvärdering av de planerade åtgärderna.
Låt mig övergå till några mer specifika frågor.
Det är mycket tillfredsställande att nedbrytning av marken har erkänts som ett allvarligt problem som måste övervinnas.
Med tanke på det nuvarande parlamentets stora oro för exempelvis ökenspridning är det angeläget att vi här i Europa öppet deklarerar vårt engagemang för att ta itu med orsakerna till problemet, såväl i Europa som i den övriga världen.
Klimatförändringar och olämpliga markförvaltningsåtgärder äventyrar markens tillstånd.
Att bestämma graden av förstöring och att därefter utveckla metoder för att se till att marken används på ett hållbart sätt, är en direkt tillämpning av den kunskapsbaserade strategi som parlamentet med rätta värderar högt.
På detta sätt skapas garantier för att åtgärderna ska bli mer riktade och för att resurserna ska användas mer effektivt för att tjäna våra syften.
Företagen har rätt att förvänta sig en konsekvent tillämpning av gemenskapslagstiftningen i de olika medlemsstaterna.
I den miljökonsekvensbedömning som utarbetats av kommissionen har man kommit fram till att det inom EU sannolikt finns 3,5 miljoner platser som är kontaminerade.
En andel av dessa, kanske 15 procent, har definitivt blivit kontaminerade.
Det är därför av största vikt att företagen kan lita på att vi inför samma metoder för klassificering av kontaminerade platser, för att kunna planera investeringar.
Vi måste komma ihåg att det finns en direkt relation mellan klimatförändringar och mark.
Enligt en forskningsartikel som nyligen publicerats i den vederhäftiga internationella vetenskapliga tidskriften Nature, har marken bara inom Storbritannien under de senaste 25 åren, varje år frisatt 13 miljoner ton koldioxid till atmosfären - lika mycket som skulle avges varje år av ytterligare 5 miljoner bilar.
Det är också värt att notera att markens förmåga att absorbera kol och omvandla det till nyttig humus ännu inte blivit fullständigt exploaterad.
Låt mig mot bakgrund av detta sammanfatta de grundläggande syftena med de åtgärder som kommissionen föreslagit.
För det första måste vi utveckla en mycket flexibel, men konsekvent och övergripande europeisk markpolitik.
Genom att skapa en ram för hållbar markanvändning och genom åtgärder som utförs vid källan kommer denna politik att förhindra ytterligare förstöring av marken, vars viktiga och livsnödvändiga sociala, miljömässiga och ekonomiska funktioner kommer att bevaras.
För det andra måste vi samla nödvändig information om marktillståndet i Europa så att vi kan fatta politiska beslut som grundar sig på kunskap och koncentrera våra insatser till platser där den svåraste markförstöringen konstaterats.
För det tredje bör förstörd mark där så är möjligt återställas, baserat på en analys av markens tillstånd och utföras av medlemsstaterna.
Syftet med återställandet bör vara att åstadkomma en markkvalitet som stämmer med åtminstone den nuvarande och den avsedda markanvändningen.
För det fjärde bör vi anta ett minimum av gemensamma regler för EU som helhet för att bland medlemsstaterna säkerställa en konsekvent strategi när det gäller markskyddsfrågor.
Dessa gemensamma regler ska hjälpa oss att åstadkomma öppenhet och att undvika snedvridning av den inre marknaden.
Syftet med strategin och direktivet är att lansera en långsiktig politik beträffande markskydd inom EU, så att alla medlemsstater redan inom några år ska ha gjort betydande framsteg inom området.
Jag vill ta upp vissa nyckelaspekter i ramdirektivet om markskydd.
För det första måste det dokument som produceras efter medbeslutandeprocessen vara entydigt och ge rättslig klarhet för intresserade parter som påverkas av lagstiftningen.
Vi får inte införa ändringar som ger kryphål i lagstiftningen och som på ett onödigt sätt begränsar direktivets omfång.
För det andra innehåller förslaget redan en hög grad av subsidiaritet och flexibilitet.
Jag inser att vissa ändringar redan föreslagits för att ytterligare öka graden av subsidiaritet.
Man måste emellertid vara övertygad om att ändringarna inte skapar problem när direktivet ska tillämpas av samtliga medlemsstater.
Detta gäller särskilt ändringsförslag som rör åtgärdsprogram inom de prioritetsområden som specificerats i direktivet.
För det tredje, för att uppnå en hög grad av miljöskydd måste vi komma överens om en konsekvent strategi för identifiering av kontaminerad mark, som ska följas av samtliga medlemsstater.
Den föreslagna strykningen av bilaga II skulle hindra oss från att nå vårt syfte.
Låt mig avslutningsvis säga att kommissionen från och med nu kommer att följa utvecklingen när kommissionens förslag diskuteras i rådet och i Europaparlamentet.
Därefter kommer kommissionen att ta ställning.
föredragande. - (ES) Fru talman! Innan vi diskuterar det förslag som vi ska rösta om i dag, vill jag tacka alla föredraganden från alla politiska grupper och jag vill särskilt tacka María Sornosa från socialdemokratiska gruppen i Europaparlamentet och vår vän Vittorio Prodi, som verkligen har arbetat tätt tillsammans med oss och som berikat direktivet, liksom De gröna/Europeiska fria alliansen och många andra ledamöter.
Det dokument vi ska rösta om i morgon innehåller många ändringar som härrör från ett avtal och därför har det berikats genom bidrag från andra politiska partier.
Det är ett dokument som till stora delar är enhälligt, något som är oväntat i en miljöpolitik som kan sägas leda till en ny EU-strategi och bana nya vägar.
Dokumentet är ytterst innovativt eftersom det svarar mot ett nytt sätt att gripa sig an direktiv.
Vi stod inför problemet att av 27 länder hade bara nio en lagstiftning om markskydd. Detta är en fråga vi måste ta itu med på nytt i framtiden.
EU har utvecklats asymmetriskt och det finns många länder som ligger på en hög nivå när det gäller markpolitik medan andra knappt har kommit i gång.
Hur ska vi komma fram till en samförståndspolitik, en gemensam politik, när skillnaderna är så stora?
Detta är den utmaning som vi har ställts inför.
Vad har vi för lösning?
Vi gick till fördraget och såg att vid definition av direktivbegreppet konstateras i artikel 249 att direktiv är gemensamma mål, men att deras genomförande och tillämpning kan överlämnas till medlemsstaterna, och det var vad vi gjorde.
Artiklarna 1 och 2 har skärpts fram till artikel 6 för att tydliggöra de gemensamma målen.
Vi har med andra ord angett målet.
Vi vet vilket mål vi måste nå och vi måste inse att hållbarhet är en process som måste ha tydliga mål, men det kan inte gå lika snabbt för alla länder att komma dit.
Vi begär inte att de som ännu inte har kommit i gång ska hålla jämna steg med de andra.
Därför vill vi att genomförandet ska lämnas i medlemsstaternas händer, med maximal respekt för subsidiaritet, för att de länder som redan kommit en bit på väg inte ska behöva upprepa sina officiella arrangemang.
De länder som har ett tydligt markskydd ska inte behöva göra om det hela.
I flexibilitetspolitiken ingår också att varje land, med tanke på att klimat och förhållanden är olika i olika länder, måste komma överens med sina medborgare om att genomföra den här politiken.
I till exempel artikel 8 garanterar vi därför att jordbrukarna ska kunna upprätta avtal om markskydd med sina medlemsstater och att de som redan har gjort det inte ska behöva göra om lagstiftningen.
Det betyder att vi samtidigt måste se till att det finns en tydlig politik för kontaminerad mark och att i detta avseende se till att medborgarnas hälsa går före allt annat, parallellt med målen att skydda hälsa och öppenhet när det gäller information till medborgarna; det är klart.
Varför anser jag att det är viktigt att det finns ett direktiv, trots alla kritiker som inte tycker så?
Mina damer och herrar! Det behövs eftersom vi ska bygga Europa på våra starka sidor och vi måste följa de länder som utfört saker på ett lyckat sätt.
Om vi inte lagstiftar hamnar vi i ovisshet och osäkerhet; och ovisshet och osäkerhet undergräver både marknad och hälsa.
Låt oss bygga Europa på dess starka sidor, inte på de svaga.
Detta är den väg vi måste välja.
Dessutom garanteras subsidiaritet och vi har redan sagt att ingen ska behöva gå igenom sina officiella arrangemang eller sin lagstiftning en gång till.
Medlemsstaterna får ansvaret för genomförandet och frihet betyder ansvar.
I ett EU med 27 medlemsstater måste vi lära oss att miljöpolitiska åtgärder inte kommer till stånd om de ska införas genom rättsväsendet.
Vi kan inte bara förlita oss på åklagare och domstolar för att de ska tillämpas.
Vi måste förlita oss på en gemensam politik och på tilltro till medlemsstaternas trovärdighet och kapacitet att komma i gång och genomföra de bästa politiska åtgärderna.
Det är därför som vi i stort har studerat god praxis.
En annan sak som är innovativ med det här direktivet är att det för första gången tar itu med klimatförändringar som rör mark, och tar upp sådana frågor som lämplig behandling av mark som översvämmas och bekämpning av ökenspridning och erosion.
Det finns en sak till som vi måste beakta: Europa och dess landsbygd är resultatet av människans arbete, den har producerats av bönder som fungerat som landsbygdens trädgårdsmästare.
Vi måste räkna med att det framtida Europa kommer att byggas av dess medborgare och därför säger jag igen att vi måste sätta upp gemensamma mål, men hjälpa medborgarna att ta den väg som också säkerställer hälsa och ger överblickbarhet.
Jag tackar för ordet, och tackar de politiska partierna ännu en gång.
föredragande. - (IT) Fru talman, herr kommissionsledamot, mina damer och herrar! Jag tackar er och jag vill också rikta ett tack till föredraganden Cristina Gutiérrez-Cortines.
Vi fick en rejäl uppgift att samarbeta om och jag hoppas vi har lyckats förbättra texten.
Det direktiv som diskuteras i dag syftar till att skydda Europas mark från sådana företeelser som ökenspridning, erosion och försaltning som i allt högre grad sammankopplas med klimatförändringar och specifik markförstöring.
Trots alla föreskrifter som gäller användning och frisättning av föroreningar till miljön har det paradoxalt nog inte funnits något direktiv som inför bestämmelser om åtaganden för att identifiera och certifiera mark som varit svårt förorenad innan den åtgärdades.
Detta verkar dock bekymra vissa personer i parlamentet och även andra som är kritiska till något de kallar för ”angrepp på subsidiariteten” och ”EU-institutionernas kvävande närvaro”, och som använder åtgärder som ramdirektivet för mark till att oroa grupper av jordbrukare eller företag och som talar om orättvisa lagar, orättvisa bestämmelser och nya administrativa och/eller ekonomiska bördor.
Vad är det vi talar om?
Vi talar om samma direktiv som ger medlemsstaterna en tidsperiod på cirka 25 år för att identifiera alla områden inom det nationella territoriet som kan anses allvarligt förorenade och således riskabla att använda för flera ändamål, såväl allmänna som privata, och alla områden som riskerar att omvandlas till öken, utsättas för erosion, saltbildning och förlust av kompaktering.
Vi talar om riktlinjer för att organisera en plan för systematisk förbättring, där så krävs, i vårt gemensamma intresse.
Vi talar om att skydda människors hälsa samtidigt som vi skyddar miljön.
Vi talar om ett ramdirektiv som respekterar medlemsstaternas autonomi och som inte innebär några betungande bestämmelser.
Jag frågar er alltså - varför denna motvilja i vissa medlemsstater och i parlamentet - de vanliga misstänkta - mot att acceptera en lista med åtgärder och platser som måste utredas noga av de nationella myndigheterna?
Vad kan de ha att dölja?
Varför så mycket motvilja när deras företrädare i rådet redan har accepterat den bindande verkan när det gäller undersökning av alla platser som föreslagits av kommissionen i bilaga II, och öppenhetsprincipen som måste råda vid markrelaterade transaktioner?
Det finns också ett mervärde med en EU-strategi för markkontroll som ska ge medlemsstaterna bättre möjlighet till kunskap om marken i de egna länderna.
I alla händelser kommer rapporteringen till kommissionen att ske praktiskt taget automatiskt eftersom rapporterna kommer att baseras på satellitbesiktningar.
Det är kanske inte allmänt känt att kommissionen redan genomfört ett liknande projekt som lett fram till den europeiska markatlasen. Det är ett bra exempel på vad vi kan åstadkomma om vi arbetar tillsammans.
Men det finns ytterligare ett argument för en gemenskapsbaserad strategi mot markförstöring, och det är klimatförändringarna, som är den utmaning som hela Europa står inför.
Den utmaningen kommer att innebära extrema väderförhållanden: mer nederbörd, längre torkperioder, mindre snömängder och höjning av havsnivån.
Det betyder att vi måste sköta om marken, för att kämpa mot dessa utmaningar, öka vattenretentionstiderna över hela territoriet för att förhindra översvämningar och gynna absorption av grundvatten, i synnerhet längs kusterna, och förhindra saltvattensinfiltration, som kan inträffa på grund av höjda havsnivåer.
Skogsskötsel för att begränsa risken för skogsbrand, eftersom längre torkperioder kommer att innebära större risk för ökenspridning i händelse av brand.
Den här typen av markskötsel kommer för övrigt att gynna användning av förnybara energikällor, till exempel vattenkraft och biomassa.
Slutligen bör vi komma ihåg markens roll när det gäller att balansera växthusgaser.
Under onsdagens omröstning vill jag be er betänka att vi mer än något annat behöver en strategi och ett direktiv som kan garantera att kommande generationer kan bruka och glädjas åt den mark som vi för tillfället har i vår vård, och betänka att alla medlemsstater står inför samma hot och samma miljörisker.
Marken är en resurs som det är ont om i Europa, och vi måste maximera dess tillgänglighet.
föredragande för yttrandet från utskottet för industrifrågor, forskning och energi. - (ES) Tack, fru talman, och tack också till kommissionsledamot Stavros Dimas för det fasta stödet till detta direktiv!
Vi välkomnar kommissionens förslag eftersom det syftar till att skydda marken och bevara dess förmåga att kontinuerligt utföra sina miljömässiga, ekonomiska och sociala funktioner och sina odlingsfunktioner, som givetvis alla är väsentliga för människors verksamhet.
Som kommissionsledamot Stavros Dimas så riktigt framfört, föreslås i direktivet flexibla regler som har ambitiösa mål och som inte är alltför normativa till sitt innehåll.
Inom ett gemensamt ramverk, en minsta gemensam nämnare, ska medlemsstaterna definiera sin egen interventionsnivå, vilket möjliggör en mer effektiv användning av administrativ kapacitet på nationell nivå.
Trots det mycket starka motståndet mot detta direktiv från vissa sektorer är det uppenbart att mark är en livsnödvändig resurs som väsentligen är icke-förnybar, och som drabbas av ökande miljömässigt tryck till följd av människors verksamhet.
Enligt de betänkanden som diskuterats här har man beräknat att markförstöringens kostnader uppgår till cirka 40 000 miljoner euro varje år, en kostnad som bärs av samhället i form av skador på infrastrukturen, ökade sjukvårdskostnader och många andra faktorer.
Det här direktivet är givetvis baserat på principer om försiktighet och förebyggande åtgärder och på principen att miljöskador ska rättas till vid källan och att förorenaren betalar.
Lagstiftningen kommer att mildra markförstöringens gränsöverskridande verkan, vilket också är ett faktum, och hjälpa till att säkerställa lika villkor inom den inre marknaden.
Jag vill betona denna aspekt eftersom de olika åligganden som ekonomiska aktörer kan införa i linje med skiljaktiga nationella markskyddslagstiftningar, skulle kunna snedvrida konkurrensen.
Avslutningsvis är markskyddsdirektivet ett steg framåt som möjliggör konkurrens med större insyn och som skyddar områden av gemensamt intresse, till exempel vatten, livsmedelssäkerhet och människors hälsa.
föredragande för yttrandet från utskottet för jordbruk och landsbygdens utveckling. - (EN) Fru talman! Jag skulle föredra att detta direktiv aldrig lagts fram.
Jag stöder att det förkastas - inte för att jag inte vill ha markskydd, eftersom det ligger i vårt intresse att ha det, utan därför att jag undrar om ett direktiv verkligen är rätt väg att gå.
Kommissionsledamoten Dimas sa själv att för tillfället är det endast nio medlemsstater som har en gällande lagstiftning för markskydd.
Jag anser att det ankommer på de övriga 18 medlemsstaterna att genomföra en lagstiftning för markskydd istället för att vi ska behöva lägga fram ytterligare ett direktiv.
Vi har redan ett grundvattendirektiv och ett nitratdirektiv.
När det gäller jordbruket har vi en omfattande lagstiftning avseende tvärvillkor om mark och markkompaktering.
Jag vet att föredraganden gör sitt bästa för att betona jordbruket i detta förslag, men jag är snarare rädd för att det kommer att innebära ännu mer byråkrati och ännu fler svårigheter för våra jordbrukare.
Kommissionsledamoten konstaterade också att det finns 300 olika marktyper i Europeiska unionen.
Det är väldigt svårt att ha ett generellt direktiv som ska omfatta samtliga markvarianters behov.
Det räcker med att man tittar på jordbruket under det gångna året, där det i vissa medlemsstater har varit torka medan det i andra har varit mycket vått på grund av kraftiga skyfall.
Om man i år gräver upp potatisen i flera av medlemsstaterna i norr där det har regnat mycket, kommer det självklart att orsaka kompaktering.
Det är nödvändigt för att kunna få tag i grödan.
Det kan rättas till nästa år genom att man alvplöjer och reparerar skador på marken.
Det krävs flexibilitet.
Jag anser att idén att lägga fram ännu ett direktiv som skapar ännu fler lagar för våra jordbrukare och vår industri är fel väg att gå.
för PPE-DE-gruppen. - (DE) Fru talman, mina damer och herrar! Direktivet om markskydd och ramdirektivet om markskydd hör, tillsammans med den temainriktade strategin för markskydd, till de viktigaste frågorna under denna sammanträdesperiod på samma sätt som de gjort under de senaste veckorna och månaderna i utskotten.
I regel behandlas en strategi - i det här fallet om markskydd - före respektive direktiv, och det av goda skäl.
Fördelen med att gå fram stegvis är att olika intressen diskuteras öppet i god tid, så att de synpunkter som kommer fram kan beaktas när direktivet utformas.
När det gäller den kraftiga kritik som riktats mot kommissionens förslag till direktiv om markskydd skulle en diskussion om frågan i förväg utan tvekan ha varit nyttig, inte minst för att dämpa känslorna på olika håll.
Till skillnad från hur ramdirektiv i regel brukar vara utformade innehåller kommissionens förslag - och jag håller med om det - många fyrkantiga, detaljerade bestämmelser som tvingar medlemsstaterna att utföra undersökningar och skicka in rapporter, vilket skulle medföra en stor administrativ belastning.
Detta är oacceptabelt.
De nya medlemsstaterna har redan nationell lagstiftning om markskydd som fungerar bra.
För dem skulle kommissionens förslag i vissa fall kräva att deras system läggs om helt, vilket skulle medföra en dubblering av regelverket och ytterligare byråkratiska bördor.
Därför ställer sig som sagt många medlemsstater skeptiska till direktivet.
Under de senaste månaderna har jag emellertid arbetat intensivt med att göra om kommissionens förslag, skriva om det.
Det handlade i grunden om att ge medlemsstaterna mer handlingsutrymme, samtidigt som vi bevarar målsättningen att stoppa den ökande markförsämringen på europeisk nivå.
Jag hoppas verkligen att vi i slutändan, tillsammans med vår vän Cristina Gutiérrez-Cortines, lyckades nå ett vettigt resultat, inte minst med tanke på hur viktig den övergripande frågan om markskydd är, ett resultat som kan bli en global modell, inte bara en europeisk.
Låt mig därför än en gång uttrycka mitt varma tack till föredraganden för att ha erbjudit en lösning som gjorde det möjligt att nå en kompromiss.
för PSE-gruppen. - (ES) Fru talman, herr kommissionsledamot, mina damer och herrar! Inom ramen för gemenskapsrätten har viktiga naturresurser (vatten, luft, arter, livsmiljön för växter och djur) sina egna specifika lagar, medan marken som resurs inte har det.
Det är dags att råda bot på denna obalans och därför vill jag tacka kommissionen för dess förslag, och också tacka föredraganden Cristina Gutiérrez-Cortines för det arbete hon har utfört.
Som många av oss redan har påpekat är marken en icke förnybar och därför begränsad naturresurs som utför många viktiga ekologiska och ekonomiska funktioner. Den utgör grunden för praktiskt taget all mänsklig verksamhet.
Det råder inget tvivel om att det europeiska institutionella rättssystemet kan komma att stimulera till en förbättring av den lagstiftning som just nu utarbetas i många länder genom att erbjuda ett sammanhängande ramverk som stöds av europeiska regler och helst också av europeiska resurser.
När det gäller markens stationära natur, som många verkar utnyttja som ett argument för att motivera valet av nationell eller subsidiär behandling snarare än en europeisk politik, så innehåller Europeiska kommissionens meddelande tillräckliga argument för behovet av en strategi på EU-nivå. Några av mina kolleger, till exempel Joan Calabuig Rull, har också nämnt detta.
Det finns några länder som inte är så pigga på att standardisera markskyddet på europeisk nivå, och därför anser vi att både strategin och direktivet har fått rätt fokus, eftersom direktivet är ett flexibelt rättsligt instrument, ambitiöst och inte överdrivet preskriptivt.
Det innebär att varje medlemsstat kan anpassa det efter sina egna behov och den egna sociala och ekonomiska situationen, eftersom en ram har fastslagits och långsiktiga mål har bestämts.
Jag tror med andra ord att metoden att föreslå ett direktiv som bygger på prevention, som ökar medborgarnas medvetenhet, ger information, identifierar prioriterade eftersatta områden och inventerar förorenade markområden, i kombination med program för nationella åtgärder och återställningsstrategier, är en konsekvent, effektiv och flexibel strategi för att hantera problemet markförstöring i Europa, samtidigt som man respekterar mångfalden av nationella förhållanden och alternativ.
Jag ber därför kammaren att först av allt med ett rungande ”nej!” avvisa det totala förkastandet av förslaget från vissa sektorer och stödja kompromissändringsförslagen som vi nådde fram till efter långvariga förhandlingar.
Detta är kanske inte det direktiv som alla önskade sig, men just på grund av att vi alla på något sätt är emot detta direktiv kan det kanske bli användbart i framtiden.
för ALDE-gruppen. - (DE) Fru talman! För det första skulle jag också vilja framföra mitt uppriktiga tack till föredraganden Cristina Gutiérrez-Cortines, som under de senaste månaderna har lagt ner stor energi på att medla mellan dem som stöder och dem som motsätter sig ett direktiv och som i slutändan lyckades lägga grunden till en fungerande kompromiss.
Trots det hyser jag, vilket jag alltid har gjort, samma åsikt som de ledamöter i parlamentet som vill avvisa kommissionens förslag.
Naturligtvis är det så att marken utgör själva grunden för vår existens.
Utan en frisk mark finns det inget jordbruk, ingen naturlig cykel av näringsämnen och, på lång sikt, inget liv.
Vi är skyldiga att om möjligt skydda våra marker från skadliga effekter och hålla dem i gott skick.
Men detta direktiv är inte rätt sätt att göra det på.
Jag tror inte frågan här är om vi vill skydda våra marker bättre eller inte.
På europeiska nivå är frågan snarare, som jag ser det: ligger detta inom vår behörighet eller inte?
Jag tror inte det gör det.
Många medlemsstater har naturligtvis infört sin egen fungerande lagstiftning om markskydd, med mer omsorg om och bättre lösningar för lokala problem än vad som skulle vara möjligt med en centraliserad reglering från Bryssel.
Därför skulle jag vilja be parlamentet stödja de ändringsförslag som skyddar medlemsstaternas handlingsutrymme.
Bortsett från detta är vi på väg att skapa en mängd ny byråkrati och nya kostnader för administrativa organ och verksamheter.
Det finns ändringsförslag som skulle utnyttja etablerandet av en industriell verksamhet till att kräva detaljerade undersökningar och rapporter.
Låt mig snabbt ge er bara ett exempel, nämligen när man ska bygga en industrigasanläggning.
Sådana anläggningar separerar luft, som är en blandning av olika gaser, i dess komponenter. Och det skadar inte marken på något sätt.
Jag tycker inte vi ska oroa oss för sådana saker, utan bara sådant där det finns en berättigad oro för att det skulle kunna förorena marken.
Jag tror det är hög tid att vi avstår från att utarbeta och offentliggöra markstatusrapporter.
De innebär ett intrång i den fria avtalsrätten.
Försäljningen av mark omfattas av civilrätten, av goda skäl, och så bör det förbli.
Mina damer och herrar, jag hoppas att vi i slutändan ska komma fram till ett direktiv som verkligen garanterar markskyddet och som inte i första hand ökar de administrativa bördorna.
Fru talman! Det finns ett ordspråk som är välkänt i många länder: ”Bättre sent än aldrig”.
Vi har kommit sent till markskyddet, efter decennier av ödeläggelse som märks tydligast i industriområdena, men det är bra att vi har insett att marken ger oss näring och att vi inte får förstöra den.
Vi får inte behandla den som en vara och bedriva en politik som innebär att den bästa affären är att köpa jordbruksmark och sedan använda den till annat än jordbruksproduktion.
Den här politiken har redan slagit tillbaka.
Det är bra att vi äntligen kan se det och börjar skydda marken, vår försörjning.
Får jag påminna om den tanke som kommer till uttryck i yttrandet från utskottet för jordbruk och landsbygdens utveckling, nämligen att ett villkor för ett effektivt markskydd är att marken bevaras och utvecklas genom jordbruket.
Mark som vårdas av bönder förblir fruktbar, men när den berövas den omvårdnaden förvandlas den till en öken.
Som företrädare för gruppen nationernas Europa stöder jag betänkandena från Cristina Gutiérrez-Cortines och Vittorio Prodi.
för Verts/ALE-gruppen. - (DE) Fru talman! Vi säger klart ”ja” till ett gemensamt markskydd för EU.
Vi har fått höra att marken är vår viktigaste icke förnybara resurs.
Markförstöringen kostar EU över 38 miljarder euro varje år.
I Tyskland är bara 2 procent av marken fortfarande orörd.
Tolv procent av marken i EU har drabbats av erosion.
Markförstörelsen respekterar inga nationsgränser.
Därför håller vi på att rycka undan mattan för oss själva genom vårt sätt att utnyttja marken.
EU-förslaget var bra. Det gick i rätt riktning och vi hade gärna förbättrat det.
Jag vet att föredraganden kämpade för det, men dessvärre såg utskottet för miljö, folkhälsa och livsmedelssäkerhet till att förslaget blev urvattnat och att ett stort antal punkter förstördes efter påtryckningar från konservativa grupper med anknytning till jordbruket.
Jag kan inte förstå varför vi i utskottet för miljö har gått med på att bibehålla sekretessen för mark som innehåller ärvda föroreningar.
Jag hoppas att vi ska kunna rätta till detta i morgon.
Det strider mot öppenheten och även mot Århuskonventionen.
Vi vet också att klimatförändringar och mark av god kvalitet går hand i hand, att marken är en viktig koldioxidkälla och att den hela tiden förlorar sin förmåga att binda koldioxid.
På grund av den urvattning som skedde i utskottet för miljö är jag rädd att ett ambitiöst markskyddsdirektiv dessvärre blir omöjligt.
Men vi behöver verkligen ett effektivt markskydd med en gemensam tidsram och gemensamma kriterier.
Vi behöver helt enkelt effektiva mål för att kunna sätta stopp för markförsämringen i Europeiska unionen.
Vi får inte ge upp försöken att skapa något som är rättsligt bindande på grund av denna så kallade kompromiss.
Endast rättsligt bindande åtgärder kommer att göra det möjligt för oss att utarbeta och genomföra en ambitiös markstrategi.
för GUE/NGL-gruppen. - (IT) Fru talman, mina damer och herrar! Vi har här ett mycket viktigt och positivt direktiv.
Jag vill tacka kommissionsledamoten Stavros Dimas, som har hanterat frågan.
Jag är medlem av en grupp som ofta kritiserar direktiv och kommissionen, men det är inte aktuellt i det här fallet.
Detta direktiv kommer att innebära enorma framsteg för EU, både vad gäller politikens kvalitet och dess effektivitet.
Tack vare ramdirektiven om naturelementen kommer marken att betraktas som en viktig del av biosfären, en grundförutsättning för den miljö- och klimatmässiga balansen och inte bara som en plattform för byggnader.
Marken lever, den absorberar koldioxid, den producerar biomassa. Den måste skyddas.
Den måste till och med förbättras, för den europeiska marken är särskild förorenad.
Europa inser detta. Vi genomförde en lång och svår diskussion i utskottet, och jag vill tacka Cristina Gutiérrez-Cortines för hennes stora engagemang i frågan.
Men det finns en risk för att Europaparlamentet ska lägga sig i kommissionens text.
Jag hoppas verkligen att det inte blir så. Jag föredrar alltid när parlamentet ligger före kommissionen.
Vissa har till och med rekommenderat att direktivet ska avvisas, men det skulle vara ett allvarligt misstag.
Europa måste blicka framåt.
Marken under våra fötter är mark som vi alla delar. Den är en del av vår planet.
Det är den enda mark vi har och vi måste ta hand om den.
för IND/DEM-gruppen. - (EN) Fru talman! Jag kan se en viss logik i en EU-lagstiftning som reglerar vatten- och luftkvaliteten.
Vi delar resurserna med andra medlemsstater och resten av världen.
Men jag anser att logiken haltar när det gäller markskyddet.
Mark är en resurs med begränsad rörlighet och uppgiften att upprätta rimliga skyddsnormer bör tillfalla varje enskild medlemsstat och dess lokala myndigheter.
Innan Europeiska unionen tar över för mycket av markkontrollen bör vi stanna upp ett ögonblick och rannsaka oss själva.
I Irland har en del av problemen i politiken om markförstöring kommit uppifrån-och-ned från Europeiska unionen.
Till exempel EU:s sockerreform, som tog bort betan från växelbruket för vete.
Införandet av betan gav marken egenskaper som gjorde den lämpligare för spannmål.
Även EU:s skogsstöd under åren har lett till olämpliga granodlingar som under sin tillväxt har gjort marken surare och i vissa fall pressat samman marken vid skörd så mycket att den blivit ofruktsam, medan den i andra fall har fått marken att lossna från kullarna och spolas ner i floder och sjöar.
Markvariationen är enorm, men mark ska alltid leva och förnyas.
EU bör förbjuda markförstöring men lämna markvård och markförvaltning till experterna på varje särskild typ i varje område.
(SK) Innan vi går in på texten i det föreslagna ramdirektivet om markskydd bör vi fundera på om EU-lagstiftning på detta område verkligen behövs.
Vi bör beakta yttrandet från utskottet för rättsliga frågor. I det yttrandet avvisades klart behovet av lagstiftning om markskydd på EU-nivå, eftersom marken inte har några gränsöverskridande egenskaper.
Därför är detta en rent regional fråga. Trots att andra utskott i sina respektive yttranden i allt väsentligt var för EU-lagstiftning på detta område, är vissa grupperingar något tveksamma.
Ändringsförslaget till artikel 5 i yttrandet från utskottet för jordbruk och landsbygdens utveckling anger till exempel klart att markförsämringen har lokala eller regionala orsaker och effekter och att det därför är viktigt att vidta nationella, till skillnad från europeiska, åtgärder.
Detta verkar strida mot resten av texten, som helt klart stöder ramdirektivet.
Samma formuleringar hittar man i ändringsförslaget till artikel 2 från utskottet för miljö, folkhälsa och livsmedelssäkerhet.
Å andra sidan är det viktigt att inse att förstöring av marken som icke förnybar resurs får betydande konsekvenser för andra aspekter där det redan finns lagstiftning, såsom vattenkvalitet, livsmedelssäkerhet, klimatförändring etc. Även om båda sidor delvis hade rätt när det gällde behovet av ett ramdirektiv, så tror jag beslutet att anta eller förkasta det europeiska ramdirektivet blir ett politiskt beslut.
Jag vill gärna kommentera förändringen av betänkandets karaktär från negativ till positiv.
Ett exempel är att termen ”riskområde” ersatts av ”prioriterat område”.
Jag anser att vi bör använda starka ord när det gäller områden där markförstöringen måste stoppas snabbt. Markområden i riskzonen ska betecknas med en negativ term för att understryka att läget är allvarligt.
(CS) Fru talman, herr kommissionsledamot! Jag vill först av allt tacka föredragandena för deras arbete med förslaget.
Dessvärre måste jag emellertid ställa mig bakom den ståndpunkt som redovisats av utskottet för rättsliga frågor som uppmanar det ansvariga utskottet att föreslå att kommissionens förslag avvisas.
De skäl som anges av utskottet är giltiga och de förblir giltiga trots de omfattande ändringar som gjorts av förslaget under de senaste månaderna.
Marken har verkligen inga gränsöverskridande effekter och bör därför förbli en fråga för medlemsstaterna.
Trots de positiva ändringarna strider därför detta förslag fortfarande mot subsidiaritetsprincipen. När det gäller proportionaliteten skulle antagandet av ett sådant lagförslag kunna ses som ett slöseri med resurser.
Vi får dessutom inte glömma att det finns många olika typer av mark inom EU, mark som används på många olika sätt.
Det är sant att direktivet har blivit vad som skulle kunna beskrivas som ett flexibelt ramdirektiv.
Som resultat av vår nya filosofi är direktivet dessutom bindande vad gäller resultaten, medan det överlåter besluten om form och metod till medlemsstaterna. Det är mycket positivt att den befintliga lagstiftningen i medlemsstaterna som täcker direktivets mål inte behöver revideras.
Därför är vi på allvar på väg mot principerna subsidiaritet och proportionalitet.
En positiv sidoeffekt av denna lagstiftning skulle vara det tryck som medlemsstater med otillräcklig markskyddslagstiftning utsätts för för närvarande, men jag är inte säker på att detta är det bästa sättet att utöva sådana påtryckningar.
Efter att ha vägt alla fördelar och nackdelar mot varandra har jag kommit fram till att det inte är nödvändigt att anta det föreslagna direktivet.
Medlemsstaterna kan skydda sin mark på egen hand.
Avslutningsvis vill jag upprepa den franska filosofens ord att om en lag inte är absolut nödvändig, så bör den inte skrivas.
(DE) Fru talman! Jag ansluter mig till de ledamöter som anser att markskydd absolut är en uppgift för Europeiska unionen, och att Europaparlamentet därför bör anta detta ramdirektiv.
Uppriktigt sagt förstår jag inte heller kommentarerna om att olika marktyper i våra medlemsstater inte skulle ha beaktats.
Jag tänker läsa igenom direktivet igen och försöka se vad de andra ledamöterna menar, för jag hittade inga av dessa stelbenta åtgärder och förslag.
Låt mig också nämna jordbrukets roll, för som jag ser det är kompromissändringsförslaget från de olika parterna mycket viktigt.
Enligt det ska medlemsstaterna när de använder mark i jordbrukssyfte uppmuntra grödor och beskogning som kan få positiv effekt på organiska ämnen och markens fruktbarhet för att förhindra jordskred och ökenomvandling.
På samma sätt bör man också stödja jordbruksmetoder som förebygger kompaktering och erosion.
Vi vet att jordbruket ofta kan skapa problem för markens kvalitet, och jag anser att ett sådant förtydligande är absolut avgörande.
Jag tror inte tanken att ”stödja jordbruket till varje pris” räcker för att skydda marken på regional, nationell eller till och med europeisk nivå.
- (PL) Fru talman! Ett ramdirektiv om markskydd kommer enligt min mening att bli ett instrument som främjar produktionen av livsmedel och tillräcklig tillgång på rent vatten för kommande generationer av EU-medborgare.
Marken har också flera andra viktiga uppgifter: den är ett underlag för mänskliga aktiviteter, tillsammans med städer och infrastruktur, och också för natur och värdefulla landskap.
Markskydd är avgörande om vi ska kunna bevara vårt naturarv och våra råmaterial.
Mot bakgrund av detta blir ett flexibelt ramdirektiv som erkänner subsidiaritetsprincipen ett instrument som uppmuntrar medlemsstaterna att skydda sin mark.
Ett direktiv längs de riktlinjerna blir bindande för medlemsstaterna när det gäller de resultat som ska uppnås på området markskydd, men det låter medlemsstaterna välja de former och metoder som ska tillämpas för att uppnå ett sådant skydd.
Direktivets förslag att medlemsstaterna ska göra upp förteckningar över förorenade områden, bland annat på regional nivå, som ska offentliggöras och uppdateras vart femte år, är värt att notera.
Detta är viktig information för att skydda EU-medborgarnas liv och hälsa.
(FR) Fru talman! Jag vill också först av allt tacka våra föredragande och berömma Cristina Gutiérrez-Cortines för det svåra arbete hon har utfört för att kunna nå resultatet att skydda vår mark.
Till skillnad från mina kolleger i parlamentet anser jag att en mer restriktiv lagstiftningsstrategi hade gett ett bättre skydd.
Jag tycker också det är synd att de av våra kolleger vilkas länder har strängare regler än vad som föreslås här, fortfarande försöker urvattna betänkandet med ändringsförslag som jag starkt rekommenderar att ni förkastar i morgon.
Våra aktiviteter inom jordbruk och transporter har drastiskt förändrat kvaliteten på vår mark.
Men den marken utgör själva grunden för vår biologiska mångfald och våra livsmedel.
Den filtrerar och lagrar organiska ämnen och mineraler och hjälper oss också att få tillgång till vatten.
Den spelar en viktig roll i kampen mot klimatförändringen.
När vi nu ställs inför ett ökat behov av livsmedels- och energiproduktion är det dessutom viktigt att vi skyddar och återställer kvaliteten på vår mark och förhindrar ökenomvandling.
Utan lagstiftning på EU-nivå kan vi inte hoppas på att uppnå resultat.
(NL) Fru talman! Jag talar som företrädare för min kollega Johannes Blokland.
Den här diskussionen har återigen visat att den föreslagna markpolitiken är mycket kontroversiell.
När det nu finns två förslag - strategin och direktivet - så verkar det som om en ny gren på miljöpolitiken har introducerats.
Jag säger ”verkar”, eftersom inget kunde ligga längre från sanningen.
Hållbar förvaltning av markanvändningen intar redan en framträdande plats i 33 olika europeiska direktiv, till exempel ramdirektivet om vatten.
Varför ska vi då lägga fram förslag på överlappande lagstiftning som innebär ännu fler bördor, framför allt för medlemsstater som redan har en väl fungerande markpolitik?
Jag kommer att stödja Vittorio Prodis tematiska strategi.
Jag anser att de medlemsstater som fortfarande inte har utvecklat en markpolitik måste göra detta på grundval av den strategin.
Ramdirektivet är däremot oproportionerligt och strider dessutom enligt min mening mot subsidiaritetsprincipen.
Till skillnad från luft och vatten har marken ingen gränsöverskridande dimension, och politiken tillämpas ofta regionalt eller lokalt.
Detta är också skälet till att jag - dvs. Johannes Blokland - har undertecknat ändringsförslaget som förkastar kommissionens förslag.
(EN) Fru talman! Vi känner alla till att ett otillåtet beslagtagande av någon annans egendom är stöld.
Jag tycker det verkar som om detta markdirektiv innebär en omotiverad maktstöld från Bryssels sida och förorsakar onödig extra byråkrati.
Som tidigare nämnts i denna debatt skiljer sig mark från luft och vatten genom att inte färdas från stat till stat.
Den har ingen gränsöverskridande dimension.
Därför bör mark vara och förbli en fråga för varje enskild medlemsstat.
IPPC-direktivet, skyldigheter avseende tvärvillkor, direktivet om deponering av avfall och nitratdirektivet ger oss redan mer än vad som egentligen behövs av EU-inblandning.
Därför behövs det inga ursäkter för en uppmaning att förkasta detta makthungriga förslag.
Men om Europeiska unionen typiskt nog beslutar att blanda sig i denna nationella fråga skulle ett förslag kunna vara att införa en betalning till jordbrukarna som motprestation för en markförvaltning och jordbrukspraxis som främjar kolbindning.
(FR) Fru talman! Min första tanke när jag såg detta förslag till direktiv var att avvisa texten.
Jag tror inte heller att ett ramdirektiv egentligen var en lämplig lösning.
Varför ska vi utarbeta en ny text om markskydd när vi redan har ett helt batteri av förordningar om mark, avfall, bekämpningsmedel och naturskydd?
Inom ramen för en bättre lagstiftning slog det mig att det inte får verka som om vi ska gå igenom Europeiska kommissionens grottekvarn igen.
Jag försökte tänka mig in i hur borgmästarna i våra städer skulle reagera när de ställs inför ytterligare en text att analysera.
Men verkligheten är denna: människans aktiviteter har inte respekterat marken.
Vi har utarmat marken genom intensiv produktion.
Dessutom har vi klimatförändringen och ökenomvandlingen.
Vår stadsplanepolitik har mineraliserat och utarmat marken. Våra medborgare blir nu förvånade när de drabbas av katastrofala översvämningar på grund av att marken inte längre kan absorbera regnvattnet.
Vem av oss har inte sett de öppna såren i landskapet som orsakas av dagbrott som förser oss med värdefulla råvaror?
Utarmad, uttorkad, förstörd, förorenad och skadad - det är vad som har hänt med denna mark som tidigare generationer talade om med vördnad. Marken var allt för dem: deras arbete, deras mat, deras liv och för många också deras egendom.
Det som en gång var Moder jord betraktas nu med misstänksamhet.
Vad blir konsekvenserna för miljö och hälsa av denna försämring, denna förorening?
Cristina Gutiérrez-Cortines har gjort ett fantastiskt jobb för att försöka hitta en acceptabel strategi, för att försöka sammanföra dem som inte ville ha detta direktiv och de som ville ha det.
Hon har lyssnat på parlamentet.
Hon har hittat balanserade ståndpunkter som respekterar behovet av subsidiaritet i valet av metoder, för det finns enorma skillnader mellan medlemsstaterna.
Sluttexten har utvecklats en hel del.
Den undviker att öka bördorna på grund av administrativa kostnader genom att uppmuntra oss att rätta till de misstag vi gjort i det förgångna, våra strategier inom jordbruk, näringsliv och stadsplanering som inte respekterar marken.
Detta betänkande, som helt gjorts om av Cristina Gutiérrez-Cortines, är bra.
Det finns en sådan mångfald av olika marktyper i Europeiska unionen att subsidiaritetsgarantin är av avgörande betydelse, samtidigt som man garanterar skydd och ett hållbart utnyttjande av marken.
(HU) Vårt övergripande mål är att garantera en sund miljö för våra medborgare och det finns strikta EU-bestämmelser som reglerar de flesta aspekter av vår miljö.
Marken är den enda komponenten i miljön som vi hittills inte har kunnat reglera, så för närvarande finns det inget EU-instrument för att stoppa föroreningen av marken och devalveringen av dess kvalitet, även om detta leder till skador för tiotals miljoner euro för oss alla.
Enligt den nuvarande lagstiftningen är vi enbart tvungna att ingripa mot föroreningar av marken när föroreningen hamnar i andra delar av miljön, grundvatten, sötvatten, jordbruksprodukter, eller när det är för sent att göra något i praktikern.
Jag välkomnar detta nya direktiv och hoppas det antas av Europeiska unionen. Det gläder mig att ett kompromisspaket har tagits fram som är ännu mer acceptabelt ur miljöskyddssynpunkt.
Det är också viktigt ur ungerskt perspektiv att lagstiftningen, på det sätt som många av oss har föreslagit, också omfattar åtgärder mot försurning av marken.
Detta är ett allvarligt hot mot vår jordbruksproduktion, så det måste även av den anledningen bekämpas med hjälp av EU-instrument.
En registrering av förorenade områden kommer att uppmuntra till åtgärder, så vi kan förhindra en förorening av vattenresurser för dricksvatten, och naturligtvis att växter förorenas.
Markreglering ligger därför i böndernas intresse.
Jag hoppas därför att vissa parlamentsledamöter från högern, inklusive, vilket är förvånande, vissa ungerska ledamöter, inte ska lyckas förhindra att det utarbetas ett direktiv som skyddar det ungerska jordbrukets och miljöns intressen.
I direktivets anda kommer återställningen av de förorenade eller markförstörda områden som upptäcks att bli en uppgift för unionen, en uppgift som vi måste avsätta resurser till i kommande gemenskapsbudgetar.
(EN) Fru talman! Detta förslag till direktiv om markskydd har stora trovärdighetsproblem.
För det första varierar markens innehåll och kvalitet i olika delar av en medlemsstat enormt.
Hur mycket större markvariationer är det då inte i 27 olika medlemsstater med högst varierande klimat?
Det är absurt att ens föreslå att Europeiska unionen skulle införa ett direktiv som skulle gälla för all mark från Medelhavet till Skandinavien.
När det gäller våra redan hårt ansatta jordbrukare, har många av dem skrivit till mitt valkretskontor för att starkt ifrågasätta behovet av ett direktiv för markskydd.
De har mycket riktigt påpekat att de har ett bestående intresse av att skydda marken, eftersom den är deras levebröd.
De menar också att det skulle lägga ännu en tung börda på deras axlar på grund av att gällande nationell lagstiftning inte erkänns tillräckligt.
Det andra stora trovärdighetsproblemet beror på EU:s kortfristiga öppna gränspolitik, som har uppmuntrat till massinvandring från Östeuropa till mitt land.
Även grönområden är hotade.
Att begrava omfattande arealer under massiv betong räknar inte jag som det bästa sättet att skydda marken.
(NL) Fru talman, herr kommissionsledamot! Jag stöder den markstrategi som utarbetats i Prodibetänkandet, men jag motsätter mig markdirektivet.
Mitt motstånd mot direktivet grundas entydigt på subsidiaritets- och proportionalitetsprincipen.
Jag har därför lagt fram ett ändringsförslag som förkastar direktivet, men också ett ändringsförslag som väljer ett annat instrument, nämligen öppen samordning.
Målen kan nås fullt ut med den metoden.
Trots allt står det väldigt klart att detta handlar om stimulans, kunskapsdelning och övervakning.
Allt är möjligt, inklusive finansiellt stöd från unionen.
Risken för dubbleringar kvarstår. Men än en gång: de prioriterade områdena har valts ut och till och med havsbotten har dragits in i diskussionen.
Medborgarna i mitt land, Nederländerna, förstår inte motiven för att införa onödig lagstiftning från ovan, från EU-nivå.
Det finns som sagt redan över 30 direktiv som gäller markens kvalitet, antingen direkt eller indirekt.
Vad är det för mening med central lagstiftning om det också går att tillämpa en decentraliserad strategi?
Men trots allt uppskattar jag Cristina Gutiérrez-Cortines försök att styra reglerna mer i riktning mot subsidiaritet.
Slutligen har jag lagt fram många fler förslag, med 40 namnteckningar, ändringsförslag som syftar till att ytterligare lyfta fram kvalitet och markskydd och reagera på de nya utmaningarna, bland annat klimatförändringen.
Ingen lagstiftning bör emellertid införas på EU-nivå.
Jag vädjar till mina kolleger i parlamentet att stödja mina ändringsförslag i det syftet.
(NL) Fru talman! Ett hjärtligt tack till Cristina Gutiérrez-Cortines, men jag måste säga att dessvärre håller vi inte med henne.
Det finns många platser i Europa med förorenad mark eller andra markproblem såsom erosion.
De problemen måste lösas så snabbt som möjligt, Jag antar att alla håller med om detta.
Kommissionen föreslår att vi ska lösa markproblemen på EU-nivå, och så vitt jag kan se är det här problemet ligger.
Trots allt är markproblemen ofta lokala och det är bara i enskilda fall som de verkligen får gränsöverskridande effekter.
Ett europeiska samarbete är önskvärt när det gäller markproblem med gränsöverskridande effekter, och i det sammanhanget är solidaritet och samarbete viktiga.
När det gäller lokala och nationella markproblem är emellertid en europeisk politik totalt överflödig.
Många medlemsstater har redan en bra nationell politik för att lösa och förebygga markproblem.
Deras politik erbjuder ett skydd som är minst lika bra som det som nu ligger på bordet.
Markdirektivet bör ta hänsyn till de medlemsstaterna. De bör undantas från europeiska skyldigheter.
(HU) Tack, herr talman!
För det första vill jag gratulera Cristina Gutiérrez-Cortines till att ha lagt ned så mycket tid och energi på att utarbeta ett utkast som faktiskt har lyckats ta sig ända till diskussion och omröstning i kammaren trots det motstånd som märks i parlamentet.
I dag, när extrema väderförhållanden orsakade av klimatförändring och civilisation medför en ökad belastning på marken och därför på hela den levande världen, är den här lagstiftningen särskilt viktig.
För min del anser jag direktivet vara ett av de viktigaste dokumenten om jordbrukets betydelse, och ett erkännande av de människor som arbetar för att bibehålla, skydda och förbättra marken.
Utan dem skulle vi inte bara sakna livsmedel. Miljön omkring oss skulle också drabbas av allvarliga skador.
Ett hållbart jordbruk som bedrivs med kunskaper är en av huvudpelarna i miljöskyddet.
Men en av de viktigaste förutsättningarna för detta är information.
Information om i vilket skick marken befinner sig, tillgänglig för allmänheten, skulle bli ett av resultaten av den nya lagstiftningen och något som äntligen skulle skydda människor och jordbrukare i stället för förorenare.
I mitt hemland Ungern är bilden redan splittrad: å ena sidan finns det mark av utmärkt kvalitet och ett starkt skydd i lagstiftningen.
Att rensa upp det kommer att ta minst fyrtio år till och kosta fyra miljarder euro. Just nu håller vi på att åtgärda detta med unionens pengar, men vi skulle vilja att processen gick ännu snabbare i framtiden, och där skulle denna lagstiftning bli till god hjälp.
Mina damer och herrar! Genom att anta direktivet om markskydd håller vi dessutom på att slutföra en process även i teologisk mening.
Vi har redan reglerat alla element som skapade världen, luft, vatten, eld, dvs. energi, och deras betydelse skyddas grundligt och på lämpligt sätt av unionen. Därför har nu turen kommit till det fjärde elementet, marken, och cirkeln sluts.
Tack så mycket!
(NL) Herr talman, herr sekreterare! Jag vill börja med att framföra mina uppriktiga gratulationer till vår föredragande Cristina Gutiérrez-Cortines och tacka henne för hennes enorma ansträngningar att försöka nå en balans mellan dem som stöder och dem som motsätter sig detta direktiv om en fråga som trots allt är väldigt komplicerad.
Personligen är jag fast övertygad om att ett europeiskt direktiv om markskydd är en nödvändighet, av olika skäl.
Jag hoppas att det fortfarande ska finns en chans att övertyga Mairead McGuinness.
Vissa ledamöter avvisar ramdirektivet, eftersom deras land redan har vittgående lagstiftning om markskydd.
Min region, Flandern, har också bedrivit en progressiv markpolitik under flera år.
Ett system med obligatoriska markcertifikat i samband med fastighetsöverlåtelser, något som fortfarande är otänkbart i många medlemsstater, har till exempel funnits på plats under lång tid.
Jag skulle vilja få dessa medlemmar att resonera på ett annat sätt.
Ett flexibelt direktiv erbjuder inte bara en ram för de medlemsstater som ännu inte har en markpolitik, utan det kan dessutom helt klart förhindra att man undergräver konkurrenspositionen för de länder och regioner som redan gör vad de kan.
Därför är det mycket viktigt att samtliga medlemsstater vidtar de åtgärder som anges i betänkandet.
Det finns helt klart gränsöverskridande effekter på många håll: erosion i Flandern skulle till exempel kunna ge slam i Nederländerna och tvärtom.
Direktivet ger också ett sammanhängande ramverk för befintlig lagstiftning om markskydd.
Jag skulle kunna redovisa fler skäl, men eftersom min tid är begränsad tänker jag avsluta med att säga att betänkandet som diskuteras i dag uppfyller alla de krav som nämnts ovan mycket bättre än kommissionens ursprungliga förslag.
Jag har också själv lagt fram många ändringsförslag och är mycket nöjd med resultatet.
Förslaget ger medlemsstaterna tillräckligt utrymme, skapar inga ytterligare administrativa bördor eller dubbleringar och det innebär också ett erkännande av de regionala myndigheternas roll.
Jag hoppas därför på ett starkt stöd från mina kolleger i morgondagens omröstning.
(EN) Herr talman! Jag vill börja med att gratulera Cristina Gutiérrez-Cortines.
Hon har gjort ett alldeles fantastiskt arbete med ett betänkande som varken behövs eller önskas av majoriteten av oss. Dessutom anser jag att det ger denna kammare och kommissionen dåligt rykte.
Ni tar fram lagstiftning som är helt och hållet onödig.
Vad ni istället borde göra är att tillämpa den lagstiftning som vi redan har.
Kommissionen misslyckas vanligtvis totalt med att tillämpa befintlig lagstiftning.
Jag kan nämna flera fall, men jag vill inte uppehålla mig vid detta nu.
Om jag exempelvis skulle vända mig till er kollega kommissionsledamot Markos Kyprianou: vi har precis haft ännu ett utbrott av mul- och klövsjuka i Storbritannien, vi har bluetongue och i dag meddelades att vi har fågelinfluensa.
Han lovade att han skulle stoppa allt detta.
Han skulle göra allt för att stoppa detta.
Jag trodde honom.
Jag tror på kommissionen när den säger en sak, och ändå tillämpar den inte den lagstiftning som redan finns för att undvika att dessa virus kommer in.
Jag uppmanar kammaren att fullständigt förkasta denna lagstiftning.
Jag anser att Cristina Gutiérrez-Cortines har gjort ett helt fantastiskt jobb och jag kommer att stödja henne fullt ut om denna kammare beslutar att inte förkasta betänkandet, men jag vill kort nämna något som Karin Scheele och Dorette Corbey sa om erosion.
Jag håller fullständigt med dem.
Erosion är ett stort problem, men inte nödvändigtvis i Europeiska unionen.
Den är ett problem vid skogsskövling och det är något som vi kan göra någonting åt.
Jag håller fullständigt med Jim Allister.
Jag anser att kommissionen sviker oss.
Den misslyckas med att tillämpa gällande förordningar.
Avslutningsvis vill jag bara säga att som jordbrukare kan jag konstatera att marken är mitt liv.
Jag kommer att skydda den så gott jag kan.
Skapa därför inte mer lagstiftning.
Tillåt mig fortsätta att skydda marken som ger oss föda och som försörjer de människor som bor på landsbygden.
(DE) Herr talman, herr kommissionsledamot, mina damer och herrar! Det kommissionen säger, nämligen att marken är den viktigaste basen för en långsiktig, hållbar produktion av livsmedel, foder och biomassa, är sant.
Det är också sant att vi inte kan vara nöjda med markförhållandena i Europeiska unionen. Men att därav dra slutsatsen att vi behöver ett direktiv på europeisk nivå är att ge sig av i fel riktning.
Varför?
Vi tar inte hänsyn till att det redan finns ett antal förordningar i Europeiska unionen som gäller marken och som vi skulle kunna utnyttja effektivt.
Exempel på sådana direktiv är till exempel livsmiljödirektivet, direktivet om integrerad miljöförebyggande verksamhet och kontroll, ramdirektivet om vatten, grundvattendirektivet och reglerna om tvärvillkor.
Genom dem har vi möjligheter att ekonomiskt påverka förbättringen av situationen i enskilda länder.
Allt detta är åtgärder som redan existerar. Om vi lägger till markskyddsdirektivet så kommer det att leda till en dubblering av reglerna, parallell lagstiftning, vilket faktiskt bara skapar mer byråkrati.
Vi säjer att vi vill minska byråkratin med 25 procent till 2010, men resultat av detta blir raka motsatsen!
Det kommer att leda till en ökning med 25 procent.
I fördraget lovade vi att reglera lokalt allt som bäst kunde regleras på den nivån, och det är det vi måste göra, och vi måste skynda på processen.
Påståendet att försämringen av marken skulle leda till klimatförändring är emellertid oacceptabelt.
Forskarna är helt överens om att denna försämring är ett resultat av klimatförändringen, och inte orsaken.
Föredraganden har sannerligen lagt ner mycket arbete på detta, men när vi ser att de regler som finns i andra direktiv är prioriterade, så är det oacceptabelt.
Vi har inga direktiv som är högt prioriterade och sedan sådana som är lågt prioriterade.
Om vi verkligen vill uppnå resultat måste vi hålla oss till metoden med öppen samordning och föra över expertis från ett land till nästa.
Det är rätt strategi och kommer säkert att ge resultat.
Detta direktiv kommer i stället enbart att skapa mer byråkrati och förvirrad lagstiftning.
(DE) Herr talman! Var finns mervärdet?
Hur motiverar man europeiska regler om markskydd?
Kommissionens argument om gränsöverskridande effekter är ganska artificiella, åtminstone ur ekologisk synpunkt.
Jag kan inte heller acceptera argumentet att den inre marknaden snedvrids av att det finns olika nationella lagar om markskydd.
Om kommissionen verkligen menade det, så skulle den inte lägga fram ett förslag på ramdirektiv som ger medlemsstaterna största möjliga självbestämmande när det gäller att definiera målen för markskyddet.
Det skulle öka skillnaderna i markskyddslagstiftning mer än det skulle jämna ut dem.
Avslöjar denna strategi att kommissionen är osäker på hur den ska gå vidare i samband med subsidiaritet när det gäller marklagstiftningen på vissa platser?
Men borde vi inte i första hand utnyttja verktyget öppen samordning i ett sådant fall, när vi alla vill se ett bättre markskydd, men de nationella lagarna skiljer sig åt?
Det anser jag.
I ramdirektivet tar kommissionen ett andra steg före det första.
Länder som saknar lagstiftning går miste om möjligheten att lära från länder med mycket goda markskyddsrutiner.
Vi kommer också att få se mer byråkrati, framför allt i de länder som redan har en tuff lagstiftning.
Varför ska de behöva undersöka hela landet och ange riskområden, trots att de redan har en föredömlig lagstiftning?
Vi behöver inte den här byråkratin, och vi behöver inte heller det guldkantade markskyddssystem som Europa nu tänker kräva av oss.
Avslutningsvis en kommentar till argumentet att parlamentet självt bad om det här direktivet för flera år sedan.
Ja, så var det för fem år sen och ännu tidigare.
Men sedan dess har vi skaffat oss erfarenheter av livsmiljödirektivet, direktivet om integrerat förebyggande och kontroll av föroreningar, ramdirektivet om vatten och många andra.
Dessutom ställs vi till svars lokalt, till skillnad från kommissionen.
Därför håller vi inte fast vid några fem- eller tioårsplaner när företag och lokala myndigheter på marken talar om för oss att det skulle bli för mycket av det goda.
Jag inser att föredraganden har lagt mer mycket arbete på att göra direktivet mindre tvingande, men byråkrati undviker man bäst vid källan.
Vi har fortfarande en chans att göra det genom att förkasta direktivet.
Jag hoppas att detta skickar en stark signal till rådet om att det inte kan förvänta sig att medlemsstaterna ska acceptera denna våg av byråkrati.
skriftlig. - (DE) Mot bakgrund av överenskommelsen om reformfördraget måste Europaparlamentet, och med det hela EU, stödja och stärka den bekräftelse på en anda av samhörighet med medborgarna och skydd av subsidiariteten som inleds i och med dessa initiativ.
Förslaget om ett ramdirektiv om markskydd lever inte upp till den målsättningen.
Den byråkrati som krävs i samband med direktivet står inte alls i proportion till direktivets faktiska nytta, och det finns inga möjligheter att motivera det inför Europas medborgare.
Tvärtom strider det mot Europeiska rådets beslut att minska byråkratin i EU med 25 procent till 2012.
Marken är i första hand en lokal resurs.
Ett effektivt markskydd måste därför genomföras på den lämpligaste nivån - på regional eller lokal nivå.
Enbart på de nivåerna kan det mycket breda urvalet av olika markegenskaper hanteras konsekvent.
Trots de omfattande förbättringar som gjorts av föredraganden avvisar jag förslaget, eftersom det innebär ett intrång i subsidiaritetsprincipen.
Vissa medlemsstater har redan mycket goda förordningar, som till och med skulle kunna försvagas genom detta direktiv.
Vid behov skulle den öppna samordningsmetoden kunna erbjuda en lösning.
- (PL) Markförstöringen är ett faktum.
En faktor som orsakar den är ... den gemensamma jordbrukspolitiken.
Självförsörjning av livsmedel har uppnåtts till priset av ett intensivare jordbruk och en utarmning av marken.
Den ökande ekonomiska avkastningen leder till att de små och medelstora jordbruken försvinner. Den övervägande majoriteten av dem var miljövänligare än de stora, vinstorienterade jordbruksföretagen.
Detta är sista chansen att bromsa trenden att överge jordbruken och återgå till en rationell och balanserad jordbruksmodell som skyddar marken.
Den nuvarande fördelningen av jordbruksbidrag är emellertid oförenlig med denna modell.
Bidragen går framför allt till jordbrukskoncerner och stora intensivjordbruk. 1,39 procent av bidragsmottagarna får nästan 30 procent av bidragen!
Den gemensamma jordbrukspolitiken måste ändras.
Huvudsyftet borde vara att producera sunda livsmedel, inte ökad konkurrenskraft.
Bra mark borde vara ett huvudinslag i denna nya politik.
Därför stöder jag alla åtgärder som syftar till att skydda marken och återställa dess fruktbarhet.
Låt oss inte konkurrera med produkter från monokulturer och intensiv djuruppfödning.
Låt oss säga NEJ till billigt kött, fullpackat med hormoner.
Låt oss inte konkurrera med frukt som har lågt näringsvärde, med billiga viner av låg kvalitet eller med genmanipulerade livsmedel, vilkas konsekvenser vi fortfarande vet mycket litet om.
Den europeiska jordbruksmodellen borde verkligen skilja ut oss från övriga världen och vara en förebild för den.
2.
Europeiska unionen och humanitärt bistånd (omröstning)
- Betänkande: Cornillet
(PL) Herr talman! Jag vill uppmärksamma er på att vi, efter diskussionen om kompromissversionen av denna resolution, hade exakt 16 minuter på oss att lägga fram ändringsförslag och se över resultatet av vårt arbete.
Jag anser att detta undergräver rätten för varje parlamentsledamot och varje politisk grupp här i parlamentet att fritt kunna påverka våra resolutionstexter, även genom att lägga fram ändringsförslag.
Jag vill be om att vi inte låter detta upprepas i framtiden.
- Före omröstningen om ändringsförslag 1:
för PSE-gruppen. - (EN) Herr talman! Vi talar om låsta konflikter.
Vi nämner två konflikter - Abchazien och Sydossetien - men jag skulle, för min grupps räkning, vilja lägga till frasen ”såsom Transnistrien” efter ”låst konflikt” så att Transnistrien också nämns i skäl O.
för PSE-gruppen. - (EN) Herr talman! Hannes Swoboda har redan informerat er om vårt ändringsförslag, som handlar om Transnistrien.
(Det muntliga ändringsförslaget beaktades.)
5.
Det europeiska intresset - För framgång i en globaliserad värld (omröstning)
- Gemensamt resolutionsförslag
- Före omröstningen om rubriken ovanför punkt 1:
för ALDE-gruppen. - (EN) Jag vill föreslå att rubriken i den första delen ändras till ”Lissabonstrategins externa dimension”.
Det vill säga att ändra ”extern politik” till ”Lissabonstrategins externa dimension”.
(Det muntliga ändringsförslaget antogs.)
- Före omröstningen om punkt 5:
- (DE) Herr talman! På grund av att ett muntligt ändringsförslag till punkt 5 har dragits tillbaka vill gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater rösta nej, tvärt emot vad som står i dess listor.
- Före omröstningen om punkt 14:
- (DE) Herr talman! Det finns ledamöter som har problem med mittpartiet, den del av texten som börjar med ”påpekar att” och slutar med ”inhemsk efterfrågan”.
Tillsammans med Daniel Caspary från gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater, föreslår jag därför att vi lägger till orden ”i vissa medlemsstater” efter ”den europeiska ekonomin”, och jag hoppas att detta kommer att lösa problemen med mittpartiet.
Jag tror att detta också kan vara till hjälp för gruppen Alliansen liberaler och demokrater för Europa.
(Det muntliga ändringsförslaget antogs.)
- Före omröstningen om punkt 30:
- (DE) Herr talman! Det finns inget att invända mot att texten senareläggs, men jag skulle ändå vilja att vi hade en omröstning om den.
Om parlamentet röstar för texten hör den hemma någon annanstans, men det skulle kunna inträffa att texten inte får något stöd, vilket är anledningen till att jag ber om en omröstning om den ursprungliga texten.
Det har inte framförts någon yrkan på en delad omröstning.
- Efter den slutliga omröstningen:
Herr talman. Nu har parlamentet röstat för att de integrerade riktlinjerna ska uppdateras och förändras.
Det handlar till exempel om den sociala dimensionen.
Hittills har kommissionen inte velat lyssna på det.
Jag skulle vilja höra herr Špidlas kommentarer till det beslut som parlamentet nu har tagit och om han inom kommissionen kommer att driva frågan om uppdaterade och förändrade integrerade riktlinjer.
ledamot av kommissionen. - (CS) Det beslut som parlamentet har fattat har en viss tyngd, och kommissionen måste ta hänsyn till detta vid utarbetandet av ytterligare handlingar. Av denna anledning väger parlamentets omröstning naturligtvis tungt och frågan om de integrerade riktlinjerna var grundläggande i den debatt vi hade i parlamentet.
Vi utgår från att ”viss tyngd” betyder ”stor tyngd” och rekommenderar att kommissionen antar vår bedömning.
Situationen i Georgien (ingivna resolutionsförslag): se protokollet
11.
Samordning av vissa bestämmelser om sändningsverksamhet för television (omröstning)
- Betänkande: Ruth Hieronymi
23.
Utnämning av en ledamot av revisionsrätten (Henri Grethen) (omröstning)
- Betänkande: Inés Ayala Sender
27.
Proklamation av samförståndet kring det humanitära biståndet (omröstning)
- Förslag till resolution
Bortfallna skriftliga förklaringar: se protokollet
17.
En papperslös förvaltning för tull och handel (omröstning)
- Betänkande: Christopher Heaton-Harris
1.
Kommissionens arbets- och lagstiftningsprogram för 2008 (omröstning)
- Resolutionsförslag
3.
Stabiliserings- och associeringsavtal mellan EG och Montenegro (omröstning)
- Rekommendation: Marcello Vernola
Avbrytande av sessionen
Jag förklarar Europaparlamentets session avbruten.
(Sammanträdet avslutades kl. 16.20.)
Skattemässig behandling av förluster i gränsöverskridande situationer (debatt)
Nästa punkt är betänkandet av Piia-Noora Kauppi, för utskottet för ekonomi och valutafrågor (ECON), beträffande skattemässig behandling av förluster i gränsöverskridande situationer.
föredragande. - (EN) Herr talman! Jag vill börja med att förtydliga vad mitt betänkande, som vi debatterar idag, handlar om.
Betänkandet handlar till synes om skattepolitik, men den verkliga frågan är den om en fungerande inre marknad i EU.
Den globala ekonomin utvecklas på ett sätt som lägger ett allt större tryck på EU att upprätthålla sin konkurrenskraft, något som har understrukits och bekräftats i olika sammanhang, särskilt i Lissabonfördraget och dess reviderade versioner.
Vi måste ta oss an utmaningen aktivt och jag tror att ett fullt funktionellt gemensamt handelssystem är första prioritet om vi vill uppnå målet.
Förutom fri rörlighet för varor, människor och tjänster, kräver detta också lika villkor för europeiska företag så att de kan göra affärer varsomhelst i EU, som om det vore ett enda land, en inre marknad - en riktig inre marknad - där beslut fattas på grundval av äkta ekonomiska fördelar, inte en snedvriden marknad skapad av byråkratiska bestämmelser.
Om denna frihet hindras leder det inte bara till suboptimala ekonomiska val, utan hindrar också europeiska företag från att växa.
Det är tråkigt att det fortfarande finns sådana hinder, eftersom en EU-omfattande inre marknad är ett måste för att europeiska företag ska kunna växa, och en förutsättning för att vi ska kunna skapa fler europeiska världsledande företag.
Gränsöverskridande konsolidering av förluster - ämnet för mitt betänkande - är ett steg på väg mot en sådan fungerande inre marknad. För tillfället är skattereglerna för en koncern som arbetar i en enskild medlemsstat i det avseendet mycket mer fördelaktiga än för en gränsöverskridande koncern.
I en enskild medlemsstat kan ett företag vanligtvis dra av förluster som orsakats av dess filialer och dotterbolag genom beskattning av moderbolaget. I fråga om filialer och dotterbolag i andra medlemsstater, varierar den nationella lagstiftningen markant.
I de flesta fall, om konsolidering av förluster för skattesyften är möjligt inom samma koncern, beviljas detta icke desto mindre med märkbara och varierande fördröjningar.
Denna diskrepans får svåra konsekvenser för den inre marknadens funktion.
Den stör investeringsbeslut och skapar ett hinder för inträde på vissa marknader, samtidigt som den orättvist gynnar de stora marknaderna där förluster kan tacklas lättare.
Det hämmar i synnerhet de små och medelstora företagens förmåga att expandera, eftersom de ofta får förluster när företaget bildas som inte omedelbart kan absorberas - även tidsfaktorn är mycket relevant för små och medelstora företag.
Lagstiftningen är olika i medlemsstaterna, vilket leder till ökade kostnader för överensstämmelse, något som är dyrt för de små och medelstora företag och som kan hanteras av de större företagen genom skattestyrning.
Till sist är fördröjd förlustutjämning dyr och nedtyngande för alla europeiska företag.
Det innebär en betydande kostnad när kapital som rättsligen kan återkrävas är uppbundet, ofta i flera år, eftersom den aktuella nationella lagstiftningen om förlustutjämning inte tillåter konsolidering utan fördröjning.
I betänkandet föreslås en lösning genom att man verkar för möjligheten att dra av förluster samma räkenskapsår, vilket skulle flytta den orimliga tidsåtgången bort från företaget till den offentliga sektorn.
Det skulle också skapa mer jämlika konkurrensvillkor samtidigt som det sänkte företagens kostnader för överensstämmelse.
Det skulle också innebära att skatteområdet är ett område där det är mycket kvar att göra för att få ut mesta möjliga av den inre marknaden.
Detta innebär inte harmonisering av skattesatser, utan snarare att skattekonkurrens är ett sundhetstecken i den europeiska ekonomin.
Det innebär dock en lagstiftning för att främja gränsöverskridande affärsverksamhet och upprätta lika villkor där investeringar baseras på sunda ekonomiska fördelar.
Jag välkomnar därför kommissionens verksamhet på det här området: att främja åtgärder för gränsöverskridande förlustutjämning.
Jag skulle vilja att parlamentet stöder den här lagstiftningen, som behövs omedelbart, och jag är tacksam för det stöd som vi har fått under processen.
Parlamentets åsikt i frågan kommer också i rätt tid, eftersom EG-domstolen har efterlyst politisk vägledning i fallet.
Jag vill också uppmana kommissionen att fortsätta med CCCTB som en mer långsiktig lösning, en punkt i betänkandet som jag hoppas att kammaren stöder.
CCCTB är dock ett långsiktigt projekt vars förverkligande ligger långt in i framtiden.
Under tiden finns det ett trängande behov av gränsöverskridande lagar, lättnader och konsolidation av förluster som en övergångsåtgärd mot några av de allvarliga problem som återfinns i den inre marknadens funktion.
ledamot av kommissionen. - (EN) Herr talman! För några veckor sedan diskuterade vi som ni säkert minns hur beskattning och tullpolitik bidrog till Lissabonstrategin för tillväxt, sysselsättning och konkurrenskraft.
Gränsöverskridande förlustutjämning är ett nyckelelement för att kunna upprätta en konkurrenskraftig inre marknad utan hinder och på så sätt bidra till tillväxt och sysselsättning.
Låt mig förklara vikten av att tillåta gränsöverskridande förlustutjämning för den inre marknaden.
Föreställ er ett litet eller medelstort företag som driver en lönsam affärsverksamhet på hemmaplan.
När det väl planerar att utöka verksamheten till andra medlemsstater, till den inre marknaden, kommer det inte bara att stöta på problem angående extra kostnader för regelefterlevnad. Därför kan detta företag i många fall inte avräkna några förluster i ett inledningsskede mot vinster som det skulle kunna generera i sin egen medlemsstat.
Att icke inhemska förluster resulterar i dubbel beskattning avskräcker många små och medelstora företag från att investera i andra medlemsstater.
Med det nya initiativet om gränsöverskridande förlustutjämning kan stora företag - men även små och medelstora företag - lättare utöka sin verksamhet utomlands och till fullo dra nytta av den inre marknaden.
Initiativet om gränsöverskridande förlustutjämning utgör en riktad lösning på kort till medellång sikt och utgör en tillfällig åtgärd.
Men observera att detta initiativ i framtiden kan utgöra ett komplement till en gemensam konsoliderad bolagsskattebas (CCCTB), särskilt för företag som inte omfattas av CCCTB.
Initiativet om gränsöverskridande förlustutjämning är mer begränsat än den konsolidering av skatteunderlaget som CCCTB innebär, eftersom detta innebär automatisk och omfattande utjämning av alla vinster och förluster inom en företagsgrupp.
Jag uppskattar det starka stöd för kommissionens initiativ om gränsöverskridande förlustutjämning som uttrycks i Piia-Noora Kauppis betänkande, för samordningsmetoden och naturligtvis också för vårt arbete med CCCTB.
Jag är liksom ni övertygad om att vi bör fortsätta med att montera ner skattehinder på den inre marknaden.
PPE-DE-gruppen - (HU) Tack, herr talman!
Jag vill tacka kommissionsledamoten och fru Kauppi för betänkandet.
De har tagit upp ett viktigt problem som väcker starka och motsatta reaktioner.
Två kommentarer.
Å ena sidan anser jag att det ur den inre marknadens synpunkt är viktigt att det inte finns någon risk för att ett moderbolag och ett dotterbolag ska missgynnas bara av den orsaken att de har verksamhet i två olika medlemsstater, jämfört med företag som har verksamhet i bara en medlemsstat.
Jag yrkar därför på att dubbelbeskattningen ska upphöra, som kommissionsledamoten framfört, kanske genom elektroniskt samarbete.
Med tiden skulle vi kunna uppmuntra effektiv verksamhet över gränserna hos de ekonomiska aktörerna och utnyttja avräknings- och undantagsmetoder.
Samtidigt anser jag att vi måste bli betänksamma när ett dotterbolag går med vinst medan moderbolaget går med förlust.
I till exempel de nya medlemsstaterna är detta ännu mer intressant ur vår synvinkel.
Min andra synpunkt som gäller inkassering av dubbel beskattning har att göra med den gemensamma konsoliderade bolagsskattebasen (CCCTB).
Vi måste förstås diskutera det, men jag har vissa betänkligheter.
Jag är ingen förkämpe för suverän beskattningsrätt men jag har ingen riktigt klar uppfattning om vilken effekt som CCCTB kan få.
Jag fruktar också att det kommer att bli en mängd politiska påtryckningar för att få fram en minsta nivå, precis som med momsen eller inkomstskatten.
Detta bevisas av de förslag som framförts av socialist- och kommunistgrupperna, och kanske också av representanterna på vänsterkanten, även om jag tror att Maastrichtkriterierna satt stopp för det.
Det jag oroar mig över är att jag inte vet vilken effekt det här kan ha på de nya kapitalsvaga östeuropeiska medlemsländerna, mot bakgrund av kapitalflödet inom den inre marknaden.
Var kommer administrationen att ligga?
Kommer vi att kunna behålla individuella skattelättnader för att väga upp en situation med ofördelaktiga infrastrukturer?
Jag kommer därför inte att ta upp dessa frågor men jag vill än en gång tacka kommissionsledamoten och föredraganden.
Tack, herr talman!
PSE-gruppen. - (IT) Herr talman, herr kommissionsledamot, mina damer och herrar! Det resolutionsförslag som vi ska rösta om i morgon är symptomatiskt för behovet av en skattepolitik på EU-nivå.
Detta betyder inte att den nationella skattepolitiken ska försvagas eller kontrolleras - ingen betvivlar de enskilda medlemsstaternas kompetens inom detta område.
Men det betyder att den ska ges en ram och samordnas, i synnerhet när beslut om sammanslagning och omlokalisering, som fattats av företag inom och utanför Europa, överskrider nationella gränser, vilket är fallet i fråga om företagsförluster i gränsöverskridande situationer.
Helt klart är inte bara nationella föreskrifter utan också bilaterala överenskommelser otillräckliga, mot bakgrund av att det i vår tidsålder med globaliserade finansmarknader och globaliserad produktion inträffar en mängd fenomen som överskrider de enskilda ländernas gränser.
Förslagets innehåll är ett resultat av att vi är överens på många punkter och jag tänker här nämna de viktigaste. Jag vill också passa på att tacka föredraganden för hennes osvikliga samarbetsvilja.
EU:s tjugosju olika skattesystem hindrar den inre marknaden från att fungera smidigt och är ett hinder för all affärsverksamhet, i synnerhet småskalig affärsverksamhet, såsom kommissionsledamoten Kovács påpekat.
Det första påståendet i texten är självklart, det uttrycker djup oro över de negativa konsekvenser som medlemsstaternas olika system vid behandling av förluster i gränsöverskridande situationer kan ha för den inre marknaden.
Den föreslagna lösningen är fortfarande en temporär övergångslösning eftersom den enda perfekta lösningen är en gemensam konsoliderad bolagsskattebas (CCCTB).
Därför stöder vi kommissionens meddelande som ett betydelsefullt steg mot att ta itu med situationen, och uppmanar samtidigt till lämplig samordning mellan medlemsstaterna när det gäller tidsplanering och lösningar - jag citerar en del av den fjärde punkten.
Det är viktigt att minnas att det finns gemensamma europeiska institutioner som till exempel Europabolaget och Europeisk kooperativ förening, liksom EU-förfaranden när det gäller grupper av gemenskapsföretag.
Vi måste bygga vidare på det, eftersom det inte bara ger oss möjlighet att knyta industriella kontakter och således påverka sysselsättningen, utan också ger oss möjlighet att bekräfta bildandet av stabila grupper av gemenskapsföretag.
Den fråga som vi trots allt vill stödja är utveckling och införande av ett produktionssystem tillsammans med EU, och inte med enskilda medlemsstater, ett produktionssystem som inte ger efter för falska lockrop och som med taktiska beslut etablerar sig i andra länder där det finns skatteförmåner, och på så sätt jämnar ut kostnader och förluster som det faller sig.
Produktionssystemet måste kunna förlita sig på lika behandling och undvika olika slags bokföring beroende på om det kontrollerande företaget har sin bas i något visst land eller verkar i flera länder.
Ett sådant resultat kan inte uppnås utan lämpliga regler och enhetliga villkor.
Att erkänna att lönsam skattekonkurrens skulle undergräva innehållet i detta förslag är inte detsamma som att höja den ideologiska fanan i opposition mot förslaget.
för ALDE-gruppen. - Herr talman! Ett tack till vår kollega Piia-Noora Kauppi för ett bra betänkande.
På ett balanserat sätt redogör hon för de problem och svårigheter som uppstår på den inre marknaden när vi har 27 olika skattesystem.
Globaliseringen, som har nämnts, har ju ytterligare ökat kraven på en gemensam syn inom EU på skattefrågor, så att konkurrenshinder kan undvikas.
Olika regler och byråkrati gör också att företagen förlorar i ekonomisk styrka och att vi förlorar jobb inom EU.
Vi behöver tydligare regler och ett synsätt som gynnar företagande, såsom Kauppi föreslår.
Kanske också vissa av oss behöver ta bort en del skygglappar.
Skatter är som bekant ett mycket känsligt ämne.
Det känsliga ordet heter skattekonkurrens och självständighet för nationerna att bestämma skattesatser.
Det långsiktiga målet för kommissionen är en konsoliderad företagsskattebas.
Då detta inte går att uppnå bör riktade åtgärder eftersträvas inom de områden som gynnar effektiviteten på den inre marknaden.
Betänkandet redovisar olika handlingsmöjligheter och visar på att enskilda länder har valt olika vägar, vilket är bra men inte tillräckligt. Det är principiellt rimligt att företag kan kvitta förluster inom ett bolag eller mellan bolag i ett konsortium även över gränser.
För att underlätta en sådan ordning behövs en gemensam syn på vad som ska beskattas, dvs. en konsoliderad bolagsskattebas.
Vi inom ALDE-gruppen tycker att detta är en riktig väg.
Införandet av CCCTB förhindrar i sig inte skattekonkurrens, snarare tvärtom.
Basen blir gemensam och överskådligheten bättre.
Denna nyordning kommer att förbättra möjligheterna särskilt för små och medelstora företag att kvitta sina förluster.
Oroade finansministrar - det finns ju många sådana - kan känna sig lugna.
Er makt att beskatta kvarstår.
I fråga om ändringsförslag 1 vill vi från vår grupp ha en delad omröstning där den första delen, som handlar om punktskatter, kan behandlas separat.
För övrigt kan vi tänka oss att lägga ned rösterna i omröstningen om Donata Gottardis ändringsförslag till skälen E och F för att möjliggöra en bred samsyn och ett brett stöd här i kammaren för detta utmärkta betänkande.
UEN-gruppen. - (PL) Herr talman! Föredraganden har gjort ett mycket bra arbete, men det här är ett kontroversiellt betänkande.
Vi kommer att rösta emot och jag ska nu förklara varför.
Det här är ett försök att skapa enhetliga skattesystem inom unionen, och att påtvinga medlemsstaterna skattelösningar.
Det innebär också att man vill gynna gränsöverskridande företag, framför små och medelstora företag. Detta skulle i sin tur leda till att många nationella företag skulle etablera filialer och dotterbolag i andra länder, inte för att det är ekonomiskt försvarbart, utan för att utnyttja bestämmelser som tillämpas på gränsöverskridande företag.
Jag skulle vilja peka på att gränsöverskridande företag under många år har kunnat dra fördel av den bristande kompetensen och korruptionen hos tjänstemän i postkommunistiska länder, där man tillgripit skattefiffel och bokföringsfiffel för att deklarera förluster och undgå skatt.
Unionen har sett mellan fingrarna med detta.
De nya bestämmelserna innebär att den här hanteringen kan fortsätta på laglig grund.
Det som förvånar mig särskilt är att följderna förmodligen blir negativa för länderna i den gamla unionen, eftersom deras skatter kommer att minska.
Jag anser att man först måste lösa problemet med skatte- och bokföringsfiffel hos gränsöverskridande bolag inom unionen och förbättra skatteinstrumentet, i synnerhet i de nya medlemsstaterna.
Det skulle bidra till att man förebygger och upptäcker skatteförseelser.
GUE/NGL-gruppen. - (DE) Herr talman, mina damer och herrar! Vi kan vara någorlunda överens om en sak: den situation som nu råder inom EU, där vi har 27 olika skattesystem som tillämpas parallellt, inom en enda marknad med fullständigt fri rörlighet för kapital, är alldeles ohållbar.
Den kommer att göra slut på sammanhållningen.
Skattekonkurrens innebär skattedumpning för de rika och mäktiga men ökar skattebördan på normalinkomsttagare och konsumenter.
Det är knappast förvånande att en sådan situation är särskilt tilltalande för fastighetsägare och storföretag.
Vad som verkligen är förvånande och alarmerande är emellertid att man i parlamentet fortfarande talar sig varm för en sådan verklighet, trots att ledamöterna i stället borde företräda de mångas intressen och inte bara elitens.
Trots alla nyanser och nyanserade bedömningar är fru Kauppis betänkande bara tomma ord.
Detta gäller både den ståndpunkt som intagits när det gäller skattekonkurrensens påstådda positiva konsekvenser och det sätt på vilket betänkandet behandlar ämnet för denna debatt, nämligen den skattemässiga behandlingen av förluster i gränsöverskridande situationer.
Det är en offentlig hemlighet att företag regelbundet utnyttjar förlustutjämning vid gränsöverskridande situationer, för att undgå skatt genom att flytta vinsterna till lågskatteområden och lågskatteländer.
Det här brukar gå mycket bra, som framgår av tillgänglig statistik: sådan faktisk förlustutjämning har i själva verket inneburit att den skatt som betalas på de multinationella företagens vinster sjunkit kontinuerligt under de senaste 20 åren.
Utslagen i EG-domstolen har bara tjänat till att underlätta sådana skattearrangemang och har därför kraftigt inkräktat på medlemsstaternas beskattningsrätt.
Allt detta underblåser dumpning av bolagsbeskattningen.
De som stöder denna utveckling vill tydligen se ett Europa där omätliga rikedomar kan ackumuleras på toppen, samtidigt som armodet ökar nere på botten och den tidigare medelklassen måste klara sig på inkomster som i realiteten faller.
Vi vill ha ett annat Europa och vi vill ha en skattepolitik som är rättvis rakt igenom samhällsskikten. Vår grupp kommer därför att förkasta betänkandet.
för IND/DEM-gruppen. - (EN) Herr talman! Föredraganden hävdar att detta initiativ kommer att uppmuntra små och medelstora företag att utöka sin gränsöverskridande affärsverksamhet.
Men jag blir inte förvånad om det har fått ett massivt stöd av de stora multinationella företagen, eftersom det är de som tjänar mest på det. I mitt land, Storbritannien, är den stora majoriteten av företag små och står för ca 70 procent av sysselsättningen.
Endast en liten del av dessa är intresserade av affärer i utlandet.
Men min huvudsakliga invändning är att det innebär mer inblandning av EU i skattefrågor.
Att döma av EU:s tidigare inblandning när det gäller mervärdesskatt, kommer det att innebära en oändlig rad av lagändringar.
Vi har haft åtta direktiv om moms hittills, och det är fortfarande en enda röra som kan utnyttjas till bedrägeri.
Företag fungerar bäst när det finns enkla, lättförståeliga regler, som Olle Schmidt precis sa. EU vet hur man gör en enda sak, och gör den perfekt.
Och det är att komplicera saker.
Så, tvärtemot andra ledamöter anser jag att det vore en mycket bättre plan att uppmuntra skattekonkurrens.
Då kan de nationer som har de lättaste och enklaste skatterna attrahera flest företag.
(PT) Herr talman! De olika medlemsstaternas olika behandling av förluster snedvrider konkurrensen inom den inre marknaden, den är orättvis och uppmuntrar en dålig skattetillämpning.
Vi välkomnar därför kommissionens initiativ att föreslå en lägsta nivå för harmonisering av dessa regler och hoppas att rådet godkänner förslaget.
Det här är ett område där regleringen måste bli bättre, i synnerhet för att undanröja den rådande osäkerheten, som lett till upprepade hänvändelser till EG-domstolen och till ökad osäkerhet om ekonomiska förhållanden till men för aktiebolag liksom för mindre och medelstora företag.
Det är ett absolut krav att de olika skattereglerna ska vara förenliga med en effektivt fungerande inre marknaden.
Kvaliteten i det betänkande som utarbetats av Piia-Noora Kauppi innebär att vi kan uppnå bred samstämmighet mellan de politiska huvudgrupperna om grundprinciperna.
En del mindre väsentliga sidor av betänkandet i dess första version, kan emellertid bli till hinder för en sådan överenskommelse.
Enligt socialistgruppen är denna process inte förenlig med ett öppet försvar för skattekonkurrens.
Skattekonkurrens gynnar konstlad förflyttning av bolag, kapital och människor.
Sådana omflyttningar leder ofta till tecken på sociala, miljömässiga och produktionsrelaterade misslyckanden.
Inom vissa ekonomier orsakar skattekonkurrensen dessutom allvarliga problem för den makroekonomiska balansen med varierande följdverkningar, i synnerhet när det gäller kvaliteten och kvantiteten hos den allmänna egendom som medborgarna i dessa länder har tillgång till.
Socialistgruppen i Europaparlamentet anser att i ett ämne av så stor strategisk vikt skulle det vara mycket lämpligt om parlamentet kunde lägga fram en ståndpunkt med brett stöd inför kommissionen och rådet . Inom detta initiativområde har EU fortfarande lång väg kvar, i synnerhet när det gäller att skapa en gemensam konsoliderad bolagsskattebas (CCCTB).
Vi måste skapa politiska villkor för det fortsatta arbetet.
En enighet om detta betänkande finns inom räckhåll.
Vi hoppas att kompromissviljan hos de största politiska grupperna gör att vi kan upprätthålla den enighet som uppnåtts om dess huvudbudskap och att vi får ett brett godkännande när vi kommer till slutomröstningen.
Sekundära aspekter som inte innebär oöverstigliga politiska skiljaktligheter får inte hindra oss från ett godkännande.
I denna process välkomnar vi det aktiva engagemanget från flera medlemmar i PPE-DE-gruppen, i synnerhet från gruppens föredragande, liksom deras kompromissvilja och öppenhet som gjort att vi kan nå enighet om de grundläggande punkterna i detta betänkande.
Tack för ordet.
(LT) Jag skulle vilja rikta er uppmärksamhet på något som vi kan tala mycket om, nämligen alla tillkortakommanden inom den inre marknaden, och betona att utvecklingen av den inre marknaden skulle ge många fördelar.
Detta dokument är viktigt genom att det gynnar en förbättrad arbetsproduktivitet hos företag med verksamhet inom den inre marknaden.
Det finns ytterligare en aspekt.
Jag representerar ett land där den övervägande delen företag tillhör europiska multinationella bolag. De är alltså inte nationella.
Därför är det ibland mycket svårt för oss att styra vår ekonomi i makroekonomisk bemärkelse eftersom bolagsstrategier inte tar hänsyn till målen för den nationella ekonomin, som t.ex. skattebalansen.
Vi behöver finna en lämplig kompromiss mellan fördelarna med en utveckling av den inre marknaden och makroekonomisk stabilitet.
Jag vill ännu en gång rikta kommissionsledamotens uppmärksamhet mot behovet att samordna politiska och ekonomiska frågor och med herr Almunia.
(PL) Herr talman! När jag nu tar ordet i denna debatt beträffande tvister som rör skattemässig behandling av förluster i gränsöverskridande situationer, vill jag betona följande frågor.
För det första ligger direkt beskattning, t.ex. bolagsbeskattning, inte inom kommissionens behörighetsområde.
Rent principiellt borde kommissionen därför inte befatta sig med det.
För det andra är jag förvånad över att betänkandet innehåller uttalanden som ogillar den minskning av bolagsskattesatser som införts i vissa medlemsstater, i synnerhet de nya medlemsstaterna.
För det tredje oroar jag mig över kommissionens krav på att påskynda arbetet med att införa en konsoliderad bolagsskattebas inom EU.
En sådan skatt, skatteskala och fastställande av skattebas är några av de mycket få instrument som fortfarande finns kvar inom ramen för medlemsstaternas befogenheter och som kan användas för att påskynda den ekonomiska utvecklingen i mindre utvecklade länder.
För det fjärde visar ett närmare studium av kommissionens förslag till en konsoliderad skattebas att syftet är att alla medlemsstater ska utvecklas i en takt som innebär en höjning av BNP på högst 2 procent per år.
Hur ska i så fall de nya medlemsstaterna, som ligger 20 eller 30 år efter EU:s mer utvecklade medlemsstater, kunna komma i kapp?
(EL) Herr talman, herr kommissionsledamot! Frågan om beskattning och möjligheten för företagsgrupper med gränsöverskridande verksamhet inom EU att överföra förluster, kan inte hanteras blott och bart under förutsättning att man vill underlätta företagens gränsöverskridande verksamhet.
Detta ändamål är givetvis av betydelse för att den inre marknaden ska fungera smidigt, men när det handlar om beskattning av en affärsrörelse, såsom anges i Piia-Noora Kauppis betänkande, bör detta betraktas i ett vidare sammanhang, nämligen större harmonisering av beskattningen inom EU.
Om vi nu antar att skattekonkurrens inte existerar på lika villkor och att det inte finns något krav på minimiavtal när det gäller en gemensam, enhetlig skattebas för företag, så att man kan fastställa enhetliga, öppna regler för att bedöma denna skattebas, måste vi gå fram mycket försiktigt när det gäller bestämmelser som rör möjlighet till skattelättnader för förluster i gränsöverskridande situationer.
I annat fall riskerar vi att snedvrida medlemsstatens beskattnings- och intäktssystem, liksom själva funktionen för den inre marknaden och konkurrensen mellan olika verksamheter.
(EN) Herr talman! Med den här nya formen av debatt kunde jag förstås använda min minut till att fråga kommissionsledamoten hur läget är angående CCCTB i rådet, eftersom vi vet att en del finansministrar inte är särskilt nöjda.
Skulle ni vilja berätta om hur debatten förs i rådet och vad de 27 medlemsstaterna föreslår idag?
ledamot av kommissionen. - (EN) Herr talman! Jag har följt debatten med stort intresse och den har bekräftat min övertygelse att införandet av gränsöverskridande förlustutjämning utgör en viktig del i att fördjupa den inre marknaden.
Jag delar Piia-Noora Kauppis åsikter om att det på ytan handlar om skatter, men att det egentligen handlar om att få den inre marknaden att fungera korrekt.
Jag är särskilt tacksam för att ni stöder och underlättar de små och medelstora företagens ekonomiska gränsöverskridande verksamhet, något som ligger mig mycket varmt om hjärtat.
Jag vill tacka föredraganden, Piia-Noora Kauppi för det mycket uppmuntrande betänkandet, samt utskottet för ekonomi och valutafrågor och utskottet för rättsliga frågor. Kommissionen kan hålla med om de flesta slutsatser.
Parlamentets stöd välkomnas som en faktor som kan ha en positiv verkan på de väntade diskussionerna i rådet.
Som antyds i betänkandet kan jag försäkra er om att vi fortsätter arbeta på CCCTB och samordningen av medlemmarnas direkta skattesystem.
CCCTB ligger mig också varmt om hjärtat och skälet är att jag är övertygad om att det gynnar de små och medelstora företagen mer än vad det gynnar de multinationella företagen.
Jag förstår dock oron, och för att svara på frågan i slutet av debatten, kan jag säga att det ligger på rådets bord, men inte som ett konkret förslag. Just nu existerar det som ett koncept och vad gäller konceptet har två tredjedelar av medlemsstaterna uttryckt sitt stöd och färre än en tredjedel har uttryckt tvekan eller missnöje.
Det vore alltför tidigt för en diskussion, särskilt en diskussion som skulle påverka den aktuella debatten om gränsöverskridande förlustutjämning, eftersom det för tillfället inte finns något konkret lagstiftningsförslag. I kommissionens lagstiftningsprogram finns dock en punkt som säger att vi ska lägga fram ett konkret, lagstiftningsförslag om CCCTB under andra halvåret, med den konsekvensbedömning som krävs.
Då kan vi diskutera om oron är befogad eller inte.
Om det dessutom inte föreligger en enhällig överenskommelse, något som jag för tillfället tror vara fallet, kan vi falla tillbaka på förstärkt samarbete som en lösning.
Ingen enskild medlemsstat kommer alltså att tvingas acceptera CCCTB eller använda sig av det.
Även i de länder som väljer CCCTB kommer inga företag att tvingas använda det, eftersom det inte är någon mening med att tvinga företag som inte opererar på den inre marknaden - som inte bedriver verksamhet på den inre marknaden - att använda den här allmänna skattebasen.
De kan fortsätta att använda sina inhemska, nationella skattebas.
Jag delar er slutsats att, för att främja följdriktig utveckling och en fungerande inre marknad, måste man ta itu med de hinder som beror på olika regler för bolagsskatter i medlemsstaterna, helst genom gemensamma metoder och samordnade åtgärder.
Med hänsyn till förlustutjämningen, visar ert betänkande på flera specifika områden som vi behöver arbeta med, bland annat frågan om de små och medelstora företagens specifika behov, hur koncerner ska definieras och omfattningen av automatiskt informationsutbyte.
Mina tjänsteavdelningar kommer att studera dessa förslag och kommentarer och, där det är möjligt, belysa frågorna.
Frågan om de små och medelstora företagen ingår redan som en viktig del i vice talmannen Günther Verheugens arbete.
En annan fråga, definitionen av företagskoncerner, är en väsentlig del i arbetet med CCCTB.
Jag kan också försäkra er om att era rekommendationer för gränsöverskridande förlustutjämning inom företag och företagskoncerner till viss del kommer att styra vårt arbete de kommande månaderna.
I ert betänkande nämns skatteflykt ett flertal gånger.
Det kan påpekas att kommissionen i december förra året antog ett meddelande om hur åtgärder mot missbruk ska tillämpas inom området direkta skatter.
Kommissionen delar de farhågor om skatteflykt som ert betänkande uttrycker.
Medlemsstaterna måste kunna förhindra att deras skatteunderlag urholkas på grund av missbruk och aggressiv skatteplanering.
Samtidigt är det viktigt att se till att man inte inskränker friheterna i fördraget.
Med detta initiativ vill kommissionen främja ytterligare diskussioner med andra institutioner om hur nationella åtgärder mot skattemissbruk kan uppfylla de kraven.
Era observationer om riskerna med skatteflykt kommer att tas i beaktande.
Slutligen gäller det ändringsförslagen i betänkandet. Kommissionen avråder från ändringsförslagen 1, 2, 3, 4, 5 och 6, men kan stödja ändringsförslagen 7 och 8, som ligger i linje med andan i meddelandet.
föredragande. - (EN) Herr talman! Jag ska fatta mig kort.
Det gläder mig förstås att de flesta grupper kommer att bifalla betänkandet vid omröstningen i morgon.
Min grupp har föreslagit att ledamöterna ska lägga ner sin röst angående ändringsförslagen 7 och 8.
Jag anser att det ligger i linje med kommissionens rekommendationer och att 7 och 8 förmodligen kommer att antas, vilket innebär att vi har en stor majoritet som stöder förslaget imorgon.
Jag skulle också vilja påminna en aning om det förflutna: hur svårt det var att tala om dessa frågor innan vi accepterade de första direktiven om bolagsbeskattning - ett direktiv om moder- och dotterbolag och ett direktiv om räntor och royalties på 1990-talet.
Men de finns nu, efter ingående diskussioner, och jag menar fortfarande att vi kan lösa alla praktiska frågor, som åtgärder mot missbruk, att vi kan förbättra direktivet om moder- och dotterbolag och att vi kan förbättra resultaten från forumet för internprissättning, och att sådana initiativ i allra högsta grad behövs.
Men till syvende och sist behöver vi en mycket bred lösning och CCCTB.
För tillfället är detta det bästa alternativet och vi måste ta allvarligt på det.
Jag hoppas att det kommer att ske under innevarande mandatperiod, före valet 2009.
Någonting måste göras före valet 2009 och vi har inte råd att vänta på medlemsstaternas ratificeringar och folkomröstningar.
Vi måste agera nu, innan tiden är slut för det här parlamentet.
Diskussionen avslutas.
Omröstning äger rum imorgon.
2. (
- Före omröstningen:
Inkomna dokument: se protokollet
Fullständigt genomförande av gemenskapens inre marknad för posttjänster (debatt)
Nästa punkt är andrabehandlingsrekommendationen från utskottet för transport och turism om fullständigt genomförande av gemenskapens inre marknad för posttjänster (13593/6/2007 - C6-0410/2007 - (föredragande: Markus Ferber).
Den tog sin början 1992, då EU-kommissionen offentliggjorde sin vitbok om utvecklingen av posttjänster, som följdes av antagandet av det första postdirektivet 1997 och översynen av detta direktiv 2002. Nu, vid början av 2008, efter över 15 år, hoppas jag att vi är redo att tillsammans anta ett rationellt regelverk som ska hjälpa oss att förlika konsumenternas intressen, intressena hos de företag som hittills haft monopol på tillhandahållandet av posttjänster, intressena hos konkurrenterna som vill ge sig in på den här lukrativa marknaden, och intressena hos de anställda inom postsektorn.
Vi i Europaparlamentet har arbetat mycket hårt för att uppnå de här målen under de gångna månaderna.
Herr talman, jag måste påpeka att klockan går för fort - jag har inte talat i tre och en halv minut än!
Jag tycker att vi har lyckats här i Europaparlamentet med att uppnå en acceptabel kompromiss mellan alla dessa olika intressen.
Jag vill tacka alla som har hjälpt till att uppnå detta - mina kolleger i Europaparlamentet, och i synnerhet Brian Simpson. Våra ansträngningar på området för posttjänster lade grunden för en 14-årig vänskap.
Vi har följt den här viktiga frågan tillsammans här sedan 1994.
Jag vill även tacka kommissionen, som har spelat en mycket konstruktiv roll, både med sina förslag och vid förhandlingsbordet.
Jag måste nog faktiskt rikta ett särskilt tack inte till det nuvarande slovenska ordförandeskapet, utan till det portugisiska ordförandeskapet för rådet, som lyckades formulera en gemensam ståndpunkt 1 oktober förra året.
Det som jag är särskilt stolt över, och som vi i Europaparlamentet alla kan vara stolta över, är att rådet i sin gemensamma ståndpunkt tagit till sig resultaten från våra överläggningar grupperna emellan, och införlivat mer än 95 procent av dem i grunderna för den gemensamma ståndpunkten.
Det är en stor framgång för Europaparlamentet, och visar att parlamentet kan lösa så komplexa frågor som avreglering av marknaden för posttjänster, vilket ytterligare berättigar de större befogenheter som anförtrotts till parlamentet genom reformfördraget.
Under diskussionerna i utskotten före den andra behandlingen försökte vi identifiera områden som vi kunde förbättra i den gemensamma ståndpunkten.
Vi gjorde det inte lätt för oss, för varje kompromiss har oundvikligen en eller annan aspekt där det kan finnas utrymme för förbättringar.
Men i december konstaterade vi i utskottet för transport och turism genom ett överväldigande godkännande i en omröstning att alla de punkter som parlamentet ansåg som viktiga faktiskt hade beaktats, och att vi inte kunde förbättra något mer.
Att ändra något skulle ha varit ett steg tillbaka.
Därför kan jag som föredragande nu säga att rekommendationen som gjorts av en stor majoritet av det ledande utskottet är att den gemensamma ståndpunkten antas utan ändringar, och det skulle glädja mig om det inträffade i morgon.
Vi skulle också föregå med gott exempel genom att avsluta den komplicerade frågan om liberaliseringen av posttjänsterna, som har sysselsatt parlamentet i 15 år, utan att en enda gång ha behövt tillgripa förlikningsförfarandet.
Låt mig bara påminna parlamentet om att vi alltid har lyckats nå en överenskommelse vid den andra behandlingen.
Att göra det igen skulle bli pricken över i vid slutet på en lång lagstiftningsprocess.
Jag ber därför om ert stöd och upprepar mitt tack till alla som har samarbetat mycket konstruktivt i den här processen.
rådets ordförande. - (SL) Jag är mycket hedrad över att vara här vid ert plenarsammanträde i dag.
Kommissionens förslag till direktiv om fullständigt genomförande av gemenskapens inre marknad för posttjänster har varit ett av de mest krävande lagstiftningsförslagen för medlagstiftarna under de senaste 15 månaderna.
När kommissionen lade fram förslaget i oktober 2006, förväntade sig alla ändlösa meningsskiljaktigheter och livliga debatter inom våra institutioner om framtiden för en av de äldsta och mest traditionsbundna offentliga tjänsterna i Europa.
Att diskutera det här ämnet var en extremt krävande uppgift för det tyska ordförandeskapet och särskilt för det portugisiska ordförandeskapet under 2007.
Från första början av debatterna fastslog våra institutioner en gemensam målsättning om att undvika populism och demagogi och fokusera på de viktigaste faktorerna, inklusive sociala aspekter för anställda inom postsektorn och permanent finansiering av en samhällsomfattande tjänst.
Som vi vet hotas postsektorn av strukturella förändringar och måste anpassas till nya ekonomiska och sociala omständigheter.
Slutfasen av den fullständiga reformen av den inre marknaden för posttjänster innebär en unik tillväxtmöjlighet för alla berörda entreprenörer.
När allt kommer omkring förväntar sig allmänheten att vi ska bevara och förbättra posttjänsternas kvalitet och effektivitet, så att användarna ska vinna på förändringen, oavsett var de bor.
Öppnandet av marknaden för posttjänster har hittills varit en framgångssaga.
Nya aktörer har kommit in på marknaden och nya möjligheter har utnyttjats, inte enbart av de nya aktörerna utan också av de etablerade.
Nya tjänster för användarna har utvecklats.
Det är uppenbart att fullständig liberalisering av posttjänsterna är en nödvändig förutsättning för att ge nytt liv åt den här sektorn och trygga dess existens vid sidan av nya former av konkurrens och alternativa tjänster.
Våra två institutioners tillvägagångssätt är ytterligare bevis på de grundläggande principerna om att bevara pålitliga tjänster av hög kvalitet och till ett överkomligt pris för alla användare, och att inte tillåta diskriminerande hinder för nya aktörer på marknaden.
Samtidigt inser både Europaparlamentet och rådet att villkoren för vissa marknader för posttjänster inom EU skiljer sig från de övriga.
När rådet uttryckte sin gemensamma ståndpunkt antog man därför beslutet att sätta slutet av 2010 som det gemensamma slutdatumet för liberaliseringen.
Vissa medlemsstater har dock blivit beviljade en övergångsperiod fram till slutet av 2012 för att införa de nya reglerna.
I likhet med den grundläggande principen för alla tidigare direktiv om posttjänster tillåter subsidiaritetsprincipen att medlemsstaterna avpassar de gemensamma reglerna till särskilda nationella omständigheter och ser till att det finns en fristående tillsynsmyndighet som övervakar marknaden för posttjänster.
Låt mig avsluta det här korta anförandet med att gratulera Markus Ferber och föredragandena från alla de inblandade politiska grupperna, dvs. skuggföredragandena, till deras bidrag till våra givande och konstruktiva diskussioner.
Jag vill påminna er om att även om vi inte alltid instämde helt i deras särskilda påpekanden, tog rådet ändå med ett antal lämpliga ändringar i sin gemensamma ståndpunkt i november 2007 och visade därigenom prov på sin politiska beslutsamhet, öppenhet och konstruktiva flexibilitet.
Jag vill särskilt framhäva kommissionens fina arbete under hela den gemensamma beslutsprocessen och dess ansträngningar för att effektivt stödja och vägleda medlemsstaterna i alla frågor om genomförandet av det nya direktivet.
I morgon kommer ni att få det slutliga beslutet och återigen bekräfta vår överenskommelse enligt rådets gemensamma ståndpunkt och rekommendationen från utskottet för transport och turism den 9 december förra året.
Vi är säkra på att ha hittat den rätta balansen mellan de olika målsättningarna och att öppet och lyhört ha behandlat de politiska utmaningarna utan att sätta rättssäkerheten för entreprenörer och konsumenter inom postsektorn i fara.
Ännu en gång tack för ert samarbete och för texten, som jag säkert tror kommer att antas, och tack för er uppmärksamhet.
ledamot av kommissionen. - (EN) Fru talman! I morgon väntas Europaparlamentet fatta ett historiskt beslut som markerar slutet på en process som inleddes för drygt femton år sedan.
Det tredje direktivet om posttjänster slutför på ett bra sätt den väl förberedda och gradvisa processen mot ett fullständigt genomförande av den inre marknaden för posttjänster.
Vad som idag syns vara en självklar och uppenbar lösning var långt ifrån oomstridd när diskussionen startade.
Den 18 oktober 2006 lade kommissionen fram sina förslag.
De följdes av intensiva och konstruktiva förhandlingar inom institutionerna.
Till sist var det Europaparlamentet som med sitt betänkande vid första behandlingen den 11 juli 2007 beredde väg för de kompromissförslag som ni idag har framför er.
Många här i kammaren har aktivt medverkat till detta viktiga resultat, och på min kollega, kommissionsledamot Charlie McCreevys vägnar vill jag särskilt berömma föredraganden, Markus Ferber, och hans kolleger och skuggföredragande från andra politiska grupper som har varit med och utformat kompromissförslaget.
Detsamma gäller det finska, tyska, portugisiska och, sist men inte minst, det slovenska ordförandeskapet.
Några kommentarer om innehållet: den text som vi nu ska besluta om är balanserad.
De olika politiska gruppernas och medlemsstaternas intressen beaktas.
Enligt kommissionens förslag skulle liberaliseringen av marknaden ske tidigare och slutdatumet i det befintliga direktivet om posttjänster fastställdes.
Två extra år är en väsentlig tidsperiod.
Det kommer att ge alla aktörer tid att slutföra sina förberedelser.
Det bör emellertid inte leda till att vi slår oss till ro.
Det viktiga för postsektorn, dess kunder, operatörer och anställda är att vi får ett slutligt och ovillkorligt datum då den fullständiga liberaliseringen av marknaden ska vara genomförd.
Genom den gemensamma ståndpunkten får vi rättvisa villkor och åläggs att undanröja marknadshinder.
Ett begränsat antal ändringsförslag har lagts fram inför morgondagens omröstning.
I de flesta fall rör det sig om ändringsförslag som avvisades redan av utskottet för transport och turism i december.
Som min kollega Charlie McCreevy konstaterade den gången tillför dessa ändringsförslag inget mervärde för den inre marknaden, för användarna av posttjänster, eller för de anställda vid posten.
Tiden är inne att fullborda postreformen.
Sammanfattningsvis är den text ni har förelagts balanserad, bra i sak, och om ni ser till de viktigaste bestämmelserna håller ni säkert med mig om att den ligger i linje med vår målsättning, som är en verklig liberalisering av marknaden, inte som ett självändamål, utan som ett verktyg för att uppfylla det övergripande målet om en högeffektiv och långsiktigt hållbar postsektor av hög kvalitet, som är anpassad till 2000-talets behov.
för PPE-DE-gruppen. - (DE) Fru talman! Under de senaste åren har vi alla, inklusive jag själv, upprepade gånger beklagat att de flesta platserna i rådets bänk har stått tomma även vid mycket viktiga lagstiftningsprojekt.
Vi borde därför tydligt uttrycka vår glädje över att det slovenska ordförandeskapet finns representerat på hög nivå vid den här viktiga lagstiftningsdebatten, och över att Slovenien redan anammar andan av Lissabonfördraget, som Slovenien förstås just har ratificerat.
Den inre marknaden för posttjänster har länge varit på väg.
Vi är mycket glada över att om allt går väl kommer vårt nuvarande utkast att bidra till att föra processen till en lyckad avslutning.
Det första förslaget från kommissionen var i princip sammanhängande och godtagbart, men för oss i Europaparlamentet var den grundläggande principen i många fall alltför allmänt tillämpad, och vi kände att viktiga detaljer förblev olösta.
På gruppen för Europeiska folkpartiet och Europademokraters vägnar framför jag varma gratulationer till vår föredragande, Markus Ferber. Det var bra att vårt utskott under hans ledning kunde fatta beslut med mycket stor majoritet om att lägga till flera viktiga punkter till kommissionens förslag vid första behandlingen, och tolka och vidareutveckla bestämmelserna.
I synnerhet på den finansiella sidan har vi lagt till ett extra alternativ - ett viktigt alternativ, eftersom det ser till att en nyckelfråga inte förbises.
Vi förstärkte de sociala bestämmelserna, särskilt i frågor som arbetsvillkor, arbetstider och semesterrättigheter.
Framför allt införde vi en tillfällig ömsesidighetsklausul för att se till att direktivet inte ger upphov till lättförtjänsta vinster för ett fåtal kvarvarande monopolinnehavare genom att de expanderar sin verksamhet in på avreglerade marknader.
I gengäld godtog vi att direktivet ska träda i kraft två år senare.
Vi anser att förslaget i stort var väl avvägt, och vi känner oss bekräftade genom rådets agerande, som i mycket hög grad stödde Europaparlamentets ståndpunkt.
Vi borde anta den ståndpunkten i morgon och liksom rådet, kommissionen och föredraganden vara nöjda över resultatet.
för PSE-gruppen. - (EN) Fru talman! På PSE-gruppens vägnar vill jag tacka Markus Ferber för hans betänkande och stora arbetsinsats som varat i flera år.
PSE-gruppen godtar att en stor del av parlamentets ståndpunkt vid den första behandlingen har godkänts av rådet. Härigenom kommer samhällsomfattande tjänster att garanteras, liksom finansieringen av de tjänsterna, och man erkänner att det måste finnas en social trygghet, samtidigt som genomförandet skjuts upp två år fram till slutet av 2010 för alla gamla medlemsstater och fram till 2012 för de nya.
Enligt min åsikt är detta en bra kompromiss.
Det finns fortfarande de som vill utkämpa antiliberaliseringsstriden.
Men den striden förlorade vi för femton år sedan när parlamentet gick med på att liberalisera sektorn för posttjänster - den gången mot min vilja.
En del av oss ledamöter har i femton års tid förhalat det fullständiga genomförandet, men till sist kommer det en tid då vi måste se verkligheten i vitögat.
Även om jag personligen skulle vilja ha en andra behandling utan ändringsförslag, anser min grupp att det är rätt att klargöra hur de samhällsomfattande tjänsterna ska finansieras och skydda de tjänster som erbjuds synskadade och blinda.
Vi stöder därför ändringsförslagen 1, 2, 6, 18 och 19.
Vi måste se till att posttjänsterna kan konkurrera, inte nödvändigtvis med varandra, men med annan teknik.
Men vi behöver rättvisa konkurrensvillkor och jag hoppas, med de reservationer jag har nämnt, att vi ska kunna avsluta vårt arbete i denna fråga på grundval av vår ståndpunkt i första behandlingen och återvända till den viktigaste frågan, som är att erbjuda medborgarna pålitliga och regelbundna posttjänster till överkomliga priser, och erkänna att alla brevbärare i hela unionen utför ett viktigt arbete.
Till sist: när Markus Ferber och jag började arbeta med den här frågan var ingen av oss gråhåriga.
Och titta på oss nu!
för ALDE-gruppen. - (IT) Fru talman! Mina damer och herrar!
Liksom alla mina kolleger vill jag gratulera föredraganden, Markus Ferber, till hans arbete. Det här arbetet påbörjades för länge sedan och under arbetets gång har vi haft betydande stunder av samförstånd och en del stunder av konstruktiv diskussion.
För min och min grupps del har det aldrig funnits något motstånd på principiell eller ideologisk nivå mot idén om liberalisering, som vi alla instämmer med och stöder, samtidigt som vi förstås försöker att se till att samhällsomfattande tjänster garanteras.
I det nuvarande förslaget till direktiv, som antogs av parlamentet vid den första behandlingen och sedan behandlades på nytt av rådet, kan vi se att en sådan garanti finns med, även om vissa av villkoren kunde ha gjorts mer precisa, specifika och detaljerade.
Vi vill inte framstå som om vi inte kan se skogen för alla träd, men å andra sidan vill vi inte heller ignorera att ibland kan detaljer vara avgörande.
Av det skälet skulle vi ha föredragit att vissa frågor hade behandlats mer i detalj. Detta gäller områdena för tillstånd, konkurrens, avgifter mellan operatören som tillhandahåller den samhällsomfattande tjänsten och andra individuella tjänster, samt rättigheter och skyldigheter kring nätverksåtkomst.
Vi skulle ha föredragit det, men majoriteten av åsikterna från parlamentet, som också fanns representerade i utskottet, var nog att det var onödigt att göra garantierna mer precisa, och man föredrog i stället att inte riskera att komplicera överenskommelsen.
Sammanfattningsvis är det så här vi ställer oss till förslaget nu. Angående ändringsförslagen om villkoren för blinda och synskadade vill vi tydligt säga att om dessa och enbart dessa ändringsförslag skulle tvinga fram en förlikning, skulle vi inte stödja det.
Om däremot andra ändringsförslag skulle antas ska vi också rösta för det.
Annars skulle vi rösta emot alla ändringsförslag som lagts fram.
Tack, fru talman, herr kommissionsledamot, herrar och fruar rådsmedlemmar.
Först av allt vill jag tacka Markus Ferber för hans arbete med att försöka uppnå en kompromiss mellan parlamentet och rådet på ett så politiskt känsligt område som posttjänster.
Jag vill betona att de objektiva svårigheterna med att liberalisera samhällsomfattande tjänster, framför allt för de nya medlemsstaterna, bemöttes i direktivet med en adekvat extra tidsfrist på två år då man kan behålla de här tjänsterna.
Samtidigt har en solid rättslig ram upprättats för att garantera samhällsomfattande tjänster.
Jag anser därför att bollen ligger hos medlemsstaternas myndigheter.
Trots de svårigheter som mött postföretag i vissa medlemsstater, däribland i mitt land Lettland, tror jag att en liberalisering av marknaden kommer att lösa den till synes hopplösa situationen med föråldrade tillhandahållare av posttjänster.
Vid omröstningen i morgon uppmanar jag er att inte stödja de tidigare nämnda förslagen, eftersom medlemsstaterna måste använda sina befogenheter till att även gynna de synskadade.
Tack.
för Verts/ALE-gruppen. - (DE) Fru talman! Tyvärr hindrar de faktiska omständigheterna mig från att delta i firandet.
Faktum nummer ett: vem kommer att vinna på det här?
Konsumenter som bor i storstäder och som älskar att få reklam i brevlådan - de kommer att vinna på det.
Likaså företag som specialiserar sig på massutskick och reklamkampanjer via post.
De som är blinda eller synskadade har däremot ingenting att vinna på det här förslaget.
Jag ber er därför att stödja vårt ändringsförslag i den frågan.
Inte heller de anställda i postsektorn har något att vinna - de kommer att få arbeta för låg lön och under enorm press, som bara kan öka under de planerade villkoren.
En annan grupp som inte kommer att vinna på liberaliseringen är de som är bosatta i glesbygdsområden och kommer att bli beroende av privata posttjänster, för vi kommer att få se en smygande nedvittring av servicenivåerna ner till det minsta möjliga och tillåtna.
Framför allt kommer inte skattebetalarna att vinna något på detta, eftersom de åter måste finansiera den samhällsomfattande tjänst som tidigare finansierades internt, eftersom den i själva verket subventionerades av inkomster från massutskick och privatpost.
Av de här anledningarna kommer jag att rösta mot direktivet.
Jag anser att det är missriktat.
Konkurrens är nog bra, men man måste se till att den sker på lika villkor.
Det har inte gjorts i det här fallet.
för GUE/NGL-gruppen. - (NL) Fru talman! Posttjänster är en arbetsintensiv offentlig tjänst.
Under artonhundratalets andra hälft beslutade staterna i Europa att de behövde ha monopol på posttjänster, eftersom den privata sektorn inte klarade av att sköta dem.
Det har alltid funnits privata företag som försökt ta sig runt den här situationen.
De erbjöd billigare tjänster, men selektivt - de valde ut de livligaste delarna av postutdelningstjänsten och erbjöd sämre arbetsvillkor och anställningsvillkor.
Sedan 1990-talet har en politisk majoritet försökt att skapa allt större utrymme för sådana företag, och det föreslagna beslutet ger dem nästan helt fria händer.
Min grupp befarar att detta kommer att leda till sämre utdelningstjänster för konsumenterna, försämrade villkor för arbetstagarna och merkostnader för medlemsstaterna för att underhålla och återupprätta sina samhällsomfattande posttjänster.
Till och med nu, när de tre största grupperna har kommit överens om en kompromiss om tidsgränser och kompletterande åtgärder, ser min grupp det här valet som ett steg tillbaka.
Utöver åtgärder för att förbättra vissa detaljer, som striktare garantier för blinda kunder och för de anställda, föreslår vi därför att denna liberalisering bör avslås.
Detta skulle också ligga i linje med vad som nyligen hände i Leipzig, där väljarna sa nej till försäljning av offentliga företag.
för IND/DEM-gruppen. - (EN) Fru talman! Jag noterar uttrycket ”ett bestämt och oåterkalleligt datum”.
En sak som EU-fadern Jean Monnet avskydde med demokrati var att ingenting är oåterkalleligt.
Ingen demokratisk regering kan binda sina efterträdare vid något oåterkalleligt.
Det finns ett demokratiskt underskott i EU, eftersom den allt hårdare sammanknutna unionen utformades som något oåterkalleligt.
Inga demokratiska öppningar.
Folk får bara rösta för att stödja vad EU-eliten har bestämt.
Det är som en enkelriktad gata.
De franska och nederländska folken röstade nej till denna oåterkalleliga union.
Att man inte beaktar deras åsikt utan återvänder till samma ratade konstitution bevisar min tes.
Ni drar inte lärdom av historien.
Sovjetunionen föll.
Hitlers tusenåriga rike varade i tolv år.
Genom att inte låta folket rösta kommer ni att få detta intoleranta EU-välde på fall lika säkert som dag följer på natt.
(HU) Fru talman! I slutet av 2012 kommer posttjänstområdet att vara fullständigt liberaliserat, och vi kommer att ha förverkligat den gemensamma marknaden också inom det området.
Eftersom ett öppnande av marknaden kommer att påverka marknaderna i de olika medlemsstaterna på olika sätt, har vi genom lagstiftningen åstadkommit en stegvis liberalisering av marknaden.
Vi har också uppnått en situation där de berörda postkontoren kan behålla och förfoga över sin vinst fram till dispensperiodens slut, vilket jag personligen betraktar som ett resultat.
Efter lång tid har vi lyckats skapa en EU-förordning som är sådan att alla befinner sig i en konkurrenssituation.
Ett särskilt tack till föredraganden för detta.
Efter liberaliseringen av marknaden är förordningen inte till nackdel utan innebär nya framtidsutsikter för de konkurrerande företagen.
Men det är bara en halv seger om vi inte också tar nästa steg.
Vilka är då dessa steg?
För det första, måste de postkontor som nu har dispens inom de närmaste åren fokusera på att motsvara de krav som konkurrensen inom EU ställer, det vill säga, de måste ta vara på de tidsfördelar som de fått.
För det andra, måste vi genom statliga förordningar och program se till att den samhällsomfattande tjänsten ligger kvar på en jämförbar nivå även om postkontoren bantas med konkurrenskraft som motto.
Vi får inte glömma att serviceansvar är och förblir ett statligt åtagande.
Förordningen har utformats så att EU-medborgare ska ha tillgång till posttjänster till lämpligt pris och med lämplig kvalitet, var de än bor, också på mycket små orter.
Tack för uppmärksamheten.
(FR) Fru talman! Jag anser att den fråga som vi ska rösta om i morgon är en historisk fråga, eftersom posten har varit i allmänhetens tjänst från allra första början, ända från monarkins dagar.
Distributionen av brevförsändelser var strategisk och utvecklades också till en samhällsomfattande och snabb service.
Vi har just avslutat den offentliga styrningen av posttjänsterna, eller kommer att göra det i morgon, och ska ersätta den med en i stort sett avreglerad postmarknad.
Det som föreslås i direktivet är först och främst en fantastisk marknad för advokater och jurister, eftersom liberaliseringen inte innebär harmonisering.
Varje medlemsstat kan besluta om sin egen finansieringsmetod och det finns fyra olika metoder.
I direktivet föreslås också något fullständigt paradoxalt: att den samhällsomfattande tjänsten ska kompenseras genom statligt stöd, precis som man i vissa länder finansierat sådant som inte var ekonomiskt livskraftigt genom överföring av medel från lönsamma sektorer.
Jag tycker att vi gör ett misstag.
Det kommer att visa sig med tiden, men vissa tecken märks redan i dag.
I Storbritannien har man investerat över 880 miljoner euro inom posttjänstområdet.
I Spanien har man just tillkännagett att landsbygden inte längre kommer att få direkta posttjänster på grund av konkurrenstrycket.
I Tyskland har man problem med att minimilönerna inte är i linje med marknaden för posttjänster.
Jag har en känsla av att vi gynnar företagen, vi låter dem skumma grädden av de bästa marknadsandelarna men vi ser inte till allmänhetens intresse eller till EU:s internationella konkurrenskraft inom posttjänstområdet.
(NL) Fru talman! Jag stöder den kompromiss som Markus Ferber kommit fram till och som tillstyrkts av rådet, eftersom jag är för en öppen marknad inom posttjänstområdet.
Jag tror att direktivet ger medlemsstaterna tillräckligt vida ramar för att liberalisera sina marknader på lämpligt sätt, och att det finns olika typer av tjänsteleverantörer som kan konkurrera om kunderna förutsatt att de levererar med given kvalitet.
Avsikten är inte att medlemsstaterna ska utnyttja ramarna för att hindra marknaderna från att liberaliseras, även om det finns viss risk för det.
Det skulle vara lätt att tillämpa direktivet så att nya företag ställs inför så stränga krav att inga nya aktörer vill besvära sig med brevförsändelser.
Om medlemsstaterna tillämpar direktivet på det sättet kommer vi att ha antagit ett stycke lagstiftning, utan att i praktiken ha ändrat någonting för postkunderna.
Jag anser att vi ska godkänna texten, men jag vill be kommissionen se till att syftet med att skapa en liberaliserad posttjänstmarknad inte kringgås av medlemsstaterna genom olika åtgärder.
Jag ser till exempel att man nyss har vidtagit åtgärder som faktiskt på nytt avliberaliserat postmarknaden i föredragandens hemland Tyskland.
(GA) Herr talman! Posttjänsterna på Irland är av central betydelse för livet på landsbygden, i synnerhet för landsbygds- och glesbygdsbor med långt till närmaste granne.
Jag välkomnar bestämmelsen om samhällsomfattande tjänster - det är av vitalt intresse för folket på Irland, liksom i övriga medlemsstater.
Jag gratulerar föredraganden till att han hållit fast vid den principen.
För att gagna kunderna borde vi ta in det i våra dokumentutkast. I det sammanhanget vill jag också säga att jag glad över den nya finansiella tjänst som Irish Post Office nu etablerar på Irland.
Det visar att företag som utför posttjänster kan anpassa sig till nya marknadskrav samtidigt som de fortsätter att leverera samhällsomfattande postservice.
Jag välkomnar också domstolens senaste förordnande om att företag som levererar posttjänster har rätt att sluta avtal om att sköta utbetalning av socialbidrag.
(PT) Rådet har samtyckt till full liberalisering av EU-marknaden inom posttjänstområdet från den 31 december 2010 under Portugals ordförandeskap. Liberaliseringen innebär att man ska tillämpa konkurrensregler på något som av många uppfattas som ett allmännyttigt organ, för att skapa en inre marknad inom posttjänstområdet. ”Det är utmärkt!”, skulle Portugals premiärminister säga.
Beslutet är emellertid ett hårt slag för de samhällsomfattande posttjänsterna, särskilt genom att man avskaffar monopoliserade områden och startar en process för att avveckla dem för att sedan överlämna dem till vinningslystna multinationella företag. Beslutet innebär att man på det allmännas bekostnad äventyrar nationella rättigheter och sparkar ut dem som arbetar inom postsektorn.
Om det funnits några tvivel beträffande den verkliga betydelsen av uttrycket ”regler för tjänster i allmänhetens intresse” i fördragsutkastet, kommer det här direktivet att skingra dem: fortsatt avveckling och nedbrytning av allmännyttiga tjänster, hinder mot att äga och ombesörja dessa tjänster via demokratiskt förvaltade och styrda offentliga bolag.
Vårt förslag är därför att direktivet förkastas.
Fru talman! Posten är en av de mest uppskattade samhällstjänsterna bland medborgarna, gammal som ung.
Detta gör att utformningen av beslutet är särskilt angeläget.
Vid tidigare behandlingar av direktivet har jag uttryckt oro för att glesbygdens behov inte skulle tillgodoses.
Det har inte varit klart att samma service skulle garanteras till alla.
Under en frågestund med kommissionär McCreevy har jag lovats att ingen förändring av förpliktelserna i den allmänna servicen skulle ske.
I dag kan vi se en kompromiss som lämnar garantier för att vi i glesbygden kommer att få vår post hämtad och lämnad fem dagar i veckan precis som alla andra.
Jag kommer att stödja kompromissen av postdirektivet i morgon.
Förhoppningsvis kommer detta att leda till att alla får bättre service, lägre pris och ett effektivare postsystem när vi avreglerar den inre marknaden på ytterligare ett område.
(NL) Fru talman! Jag vill rikta ett varmt tack till föredraganden Markus Ferber för hans arbete.
Han har lyckats ena parlamentet i den här besvärliga frågan vid första behandlingen, även om både han och jag kände att vi borde ha kommit lite längre.
Det var förstås vårt eniga ställningstagande som vägledde rådet, och jag ansluter mig helhjärtat till den gemensamma ståndpunkten.
Medlemmar i socialistgrupperna och de gröna grupperna har tyvärr börjat tveka och inser inte de stora möjligheter som direktivet erbjuder när det gäller nya verksamheter och arbetstillfällen.
Jag är helt och fullt övertygad om det och jag stöder mig på exempel från flera medlemsstater.
Allt hänger nu på om kommissionen håller fast vid direktivet så att det inte stannar vid en pappersprodukt.
Om direktivet införs kommer det helt säkert att uppnå sitt syfte och öppna marknaderna.
Konsumenterna får bättre service, och det blir inte som i Tyskland, där nya aktörer, och inte bara nya aktörer utan också nya företag, nya tjänster och nya arbetstillfällen, slås ut från marknaden under förevändning av socialt skydd.
Jag är förstås glad över det gensvar jag fick från kommissionen i går.
Om jag förstått det rätt ska kommissionen titta närmare på situationen i Tyskland.
Jag uppmanar er att göra det mycket snart eftersom de nya aktörerna på den tyska marknaden har det besvärligt, och det skulle vara hemskt om situationen inte reds upp; det får så att säga en prejudicerande verkan.
Det finns risk för att Frankrike och andra länder följer efter och till slut kommer vi inte att ha uppnått någonting alls.
Kommissionen har ett mycket stort ansvar i den här frågan.
Jag hoppas att ni använder alla lagliga möjligheter som står till buds och dessutom utövar politiskt tryck för att direktivet ska tillämpas på den europeiska postmarknaden.
(PL) Fru talman! Det är ett kontroversiellt beslut att låta privata aktörer utföra posttjänster.
Tiden kommer att utvisa om det är till konsumenternas fördel.
I vissa nya medlemsstater med lägre utvecklingsnivå har institutioner som försvarar konkurrens- och konsumentintressen har ganska svag förankring i det allmänna medvetandet.
Det finns risk för att balansen mellan kapitalets och konsumenternas intressen rubbas.
Därför är det bra att fastställa datumet till 2012.
Samtidigt föreslår jag att vi analyserar hur postmarknaden fungerar i de länder som redan antagit de nya reglerna, för att identifiera och förebygga oegentligheter i de övriga länderna, och att vi gör det före 2012.
Jag funderar också på om en aktör som utför allmännyttiga tjänster bör få ersättning av myndigheterna och inte bara kompensation - såsom föreslås av författarna till det här betänkandet.
Många års arbete på det här lagförslaget har gett Markus Ferber gråa hår.
Jag hoppas att införandet av de nya bestämmelserna inte ska ge honom ännu mer bekymmer så att han börjar tappa håret.
(DE) Fru talman! Markus Ferbers ståndpunkt är tydligen rakt motsatt mot Corien Wortmann-Kools och de övriga ledamöternas ståndpunkter.
Jag anser det är fel att privatisering och liberalisering av allmännyttiga tjänster används som standardsvar på globaliseringsfrågor.
Jag har också skäl att tro att allt fler människor tar avstånd från det förhållningssättet.
Under en omröstning i Leipzig förra helgen röstade 80 procent av de röstande mot privatisering, och har på så sätt hindrat fullmäktige från att genomföra fler privatiseringar under de närmaste tre åren.
Låt mig också säga att det direktiv som vi diskuterar i dag verkligen inte innehåller några garantier för att skydda människor - det vill säga anställda - från social dumpning.
I Tyskland har vi har sett hur företag som byggt upp sin verksamhet på rena bottenlöner är motståndare till att införa minimilöner inom posttjänstområdet.
Jag är också allvarligt bekymrad över vilka följder det kan få om offentliga institutioner tecknar avtal med sådana företag.
(PL) Fru talman! Vi har arbetat med att liberalisera postsektorn i mer än 15 år.
Inom EU som helhet är den värderad till mer än 90 miljarder euro per år. Vi står nu inför omröstning och att skriva in den här lagstiftningen i unionens historia och jag vill gratulera föredraganden till ett utmärkt arbete.
I sin nuvarande version är till projektet till stora delar en kompromiss där vi tycks ha uppnått följande huvudsyften: fullständigt genomförande av den inre marknaden inom posttjänstområdet, huvudsakligen genom att monopolet på ordinarie brevförsändelser upphör, och säkrat fortbestånd för allmännyttiga tjänster av hög kvalitet och till låg kostnad.
Den version av direktivet som nu föreligger är emellertid inte lika ambitiös som kommissionens ursprungliga förslag.
Under den pågående liberaliseringen har avsteg från liberaliseringens idé till förmån för en gradvis och ganska försiktig liberalisering av postmarknaden när det gäller brev som väger mindre än 50 gram blivit allt tydligare.
Det framgår av det kompromissdatum då direktivet ska träda ikraft, särskilt ifråga om nya medlemsstater och länder med liten befolkning, små geografiska områden och klausuler om allmännyttiga tjänster.
Det angivna datumet, 31 december 2012, för medlemsstater som blivit EU-medlemmar 2004 tycks onödigt avlägset.
Jag inser att det är en del av den kompromiss som vi förhandlat fram och godkänt, men det kan bromsa de föreslagna förändringarna.
Jag är rädd att en så lång period - mer än fyra år - innan direktivet träder ikraft, gör att förändringar som skulle ha blivit genomförda nästan genast om det varit fråga om en tvåårsperiod, kommer att tappa fart.
Slutligen vill jag stödja fru Mrs Pleštinskás begäran om att klausuler som rör blinda och personer med nedsatt synförmåga åter ska införas i förslaget.
De saknas i den nu aktuella versionen.
(NL) Fru talman! Jag vill tacka föredraganden och mina medledamöter som hjälpt oss att komma fram till ett resultat som är avsevärt bättre än kommissionens första förslag.
Jag förstår varför många av oss tycker att det kan räcka nu, men bakom de positiva inslag som lagts till direktivet finns det också flera riskfaktorer.
Vi har fortfarande inte uppnått någonting, eftersom medlemsstaterna ges ett så stort ansvar på två viktiga punkter.
Den första punkten är att det finns mängd frågetecken när det gäller hur den samhällsomfattande tjänsten ska finansieras.
Medlemsstaterna har flera alternativ, men det är inte alltid klarlagt om de fungerar i praktiken.
I många fall kommer det att leda till tvister, bland annat rättstvister.
Jag skulle därför vilja klargöra två saker: för det första att medlemsstaterna åläggs att garantera samhällsomfattande tjänster och finansiera dem, vilka omständigheterna än må vara, och för det andra att medlemsstaterna grundligt och i god tid måste förebereda sig för den nya situationen.
Den andra viktiga punkten gäller det sociala området.
Här är det viktigt att peka på att direktivet innebär att medlemsstaterna via ett licenssystem kan kräva att alla postföretag ska följa till exempel samma kollektivavtal eller andra miniminormer.
Det är en bra ide, men den är ändå bara frivillig och kommer att tillämpas olika från ett land till ett annat.
Därför tycker jag att direktivet bör skärpas något, inte för att jag är rädd för vad som kommer att hända, utan för att en fri marknad måste regleras och för att en liberalisering måste vara noga förberedd.
(EL) Fru talman! Vi är inte nöjda med varken Europeiska kommissionen, rådet eller föredraganden, eftersom ingen av dem har hänvisat till variationer inom antalet sysselsatta inom sektorn, arbetsvillkor, antal arbetstimmar eller löner.
Man har inte heller utformat några bestämmelser som rör effektiv kontroll av företagens avgiftsstrategi eller privata monopolsituationer vid pakettransport och expresspost.
I betänkandet betonar man vidare att sysselsättningen i medlemsstaterna är stabil, även om lokala variationer kan förekomma, men man har inte tagit fram några data för att bevisa det.
Underlaget ger alltså ingen möjlighet att göra en riktig utvärdering av arbetstagarnas intressen.
Jag vill slutligen betona att rådet i viss mening ratificerat parlamentets ändringsförslag och samtidigt gett oss tillfälle att ingående diskutera de sociala konsekvenserna, både för dem som är sysselsatta inom posttjänstområdet och för konsumenterna.
(DE) Fru talman! Fullbordandet av den inre marknaden för posttjänster illustrerar mer än väl sanningen i talesättet: ”Den som väntar på något gott väntar aldrig för länge”.
Till och med jag kan stödja det framlagda utkastet som är ett resultat av femton års hårda förhandlingar.
Jag råkar vara en av de som hellre hade behållit monopolet för nationell postutdelning av brevförsändelser under 50 gram.
Nu är det sista stadiet i den kontrollerade avregleringen av postmarknaden fastställt till den 1 januari 2011.
Med tanke på de luxemburgska posttjänsternas struktur samt det lagstadgade kravet att anställa volontärer från väpnade styrkor i offentlig tjänst och de påföljande kostnaderna kunde jag inte skriva under på en snabb och otillräckligt kontrollerad avreglering av marknaden för posttjänster eftersom detta kunde ha fått oacceptabla konsekvenser för postanställda och kunder.
Inför den första behandlingen bad jag därför föredraganden, Markus Ferber, att tillåta en tvåårig förlängning av tidsfristen för införlivande för små länder med relativt få invånare, så att dessa länder kan fortsätta att begränsa tillhandahållandet av vissa tjänster till leverantören av samhällsomfattande tjänster, och jag tackar herr Ferber för hans förståelse.
Jag hade diskret skrivit om överenskommelsen för att garantera att Luxemburg skulle gagnas av undantaget, men ministrarna föredrog att förebygga eventuella missförstånd genom att namnge de berörda länderna.
Detta gör oss säkra.
Det viktiga är att kravet på att tillhandahålla samhällsomfattande tjänster garanterar insamling och snabb utdelning av brev till avsedda privatpersoner och företag under alla arbetsdagar, även i avlägsna eller glesbefolkade områden.
Det kan vara nödvändigt med extern finansiering för att täcka nettokostnaderna för de samhällsomfattande tjänsterna. Denna finansiering, och således även problemet med överkomliga taxor, har också reglerats på ett tillfredsställande sätt.
Slutligen har bästa möjliga åtgärder vidtagits för att garantera varaktiga kvalificerade arbetstillfällen hos leverantörer av samhällsomfattande tjänster, samt för att garantera att man följer anställningsvillkor och sociala trygghetssystem som baseras på existerande lagbestämmelser eller kollektivavtal, i motsats till vad vänstern ville få oss att tro.
De borde läsa utkastets formuleringar.
Det är nämligen uttryckligen fastställt att förberedelserna för avregleringen av postmarknaden måste respektera sociala hänsyn.
Vad gäller förslaget om kostnadsfria posttjänster för synskadade, som lades fram av våra filantropiska missionärer, kan jag personligen inte förstå varför förmögna människor med nedsatt syn skulle få skicka sina brev gratis på skattebetalarnas bekostnad.
De som föreslår denna ändring är helt ute och cyklar, eftersom det är medlemsstaterna som ska garantera sådana arrangemang.
Subsidiarité oblige!
(HU) Tack, fru talman. Mina damer och herrar!
Den gradvisa liberaliseringen av marknaden för posttjänster är en viktig milstolpe för fullbordandet av den inre marknaden.
Detta kommer att bidra till att sätta stopp för speciella rättigheter inom posttjänsterna, och leda till att ett bestämt och oåterkalleligt datum för liberaliseringen av marknaden fastställs. På samma gång garanteras samhällsomfattande tjänster på en hållbar och hög nivå.
Liberaliseringen av marknaden kommer att stärka konkurrensen, och på så sätt kan tjänstenivån förbättras med avseende på kvalitet, pris och valmöjligheter.
Denna åtgärd kommer att främja en harmonisering av de grundläggande principerna för reglering av posttjänster och den kommer troligen att ge lägre avgifter liksom bättre och mer nyskapande tjänster. Dessutom kommer den att leda till att bättre förutsättningar för tillväxt och sysselsättning alltjämt skapas.
Förslaget till ändring av direktivet är ett resultat av en utmärkt kompromiss som respekterar de skillnader som uppstår på grund av att medlemsstaternas historia och ekonomi skiljer sig åt.
Man tar hänsyn till att det tar längre tid att förbereda liberaliseringen i vissa länder, framförallt i de östeuropeiska länderna. På samma gång tar man även med andras intressen i beräkningen.
För att förhindra snedvridning av marknadskonkurrensen kan inte de länder som ännu inte har liberaliserat sin marknad tillhandahålla tjänster i de länder där postsektorn redan är fullständigt liberaliserad före 2012. Då går tidsfristen för undantaget ut.
Jag skulle vilja tacka Markus Ferber för hans arbete, men jag vill naturligtvis också tacka Brian Simpson, vår skuggföredragande.
(PT) Jag gratulerar Markus Ferber och Brian Simpson för kvaliteten i deras betänkande, och jag tackar även alla inblandade medlemmar och parter för deras öppenhet under förhandlingsprocessen.
Liberaliseringen av marknaden för posttjänster har fortfarande långt ifrån lett fram till en konkurrenskraftig marknad där konsumenter och företag är de största vinnarna.
Därför hävdade jag att kommissionens strategi kanske inte kan garantera tillgång till samhällsomfattande tjänster i tillräckligt stor utsträckning.
Således stödde jag skuggföredraganden Brian Simpsons ståndpunkt om att man bör garantera de samhällsomfattande tjänsterna och inrätta en kompensationsfond. Jag stödde även hans ståndpunkt om att man ska liberalisera posttjänster under 50 gram 2010, eller i särskilda fall, som de nya medlemsstaterna med yttersta randområden, senast den 31 december 2012.
Jag är också nöjd med tanke på de stater som omfattades av de särskilda villkoren, även om jag måste påpeka att dessa villkor kanske inte är tillräckliga. I så fall kommer ytterligare åtgärder att krävas.
När det gäller sysselsättningen är jag glad över det tidigare införda tillägget om att en rapport måste läggas fram om den allmänna utvecklingen av sysselsättningen inom sektorn, de arbetsvillkor som tillämpas av alla operatörer i en medlemsstat och eventuella framtida åtgärder.
Jag är väldigt nöjd med den gemensamma ståndpunkt som uppnåtts, men jag stöder ändringsförslagen som lagts fram av mina kolleger Gilles Savary, Saïd El Khadraoui och Inés Ayala Sender, bland andra, och av min parlamentariska grupp. De befäster nämligen idén om att liberaliseringsprocessen måste vara genomtänkt för att jämlik allmän tillgång, utveckling och sysselsättning ska förstärkas.
På grund av alla dessa orsaker uppmanar jag er att stödja betänkandet och rådet, samt att stödja parlamentets ståndpunkt.
(EN) Fru talman! Parlamentet bör godkänna våra ändringsförslag om att återinföra obligatoriska kostnadsfria posttjänster för blinda i direktivet.
Herr Vizjak! Trots att ni säger att ni var öppen och flexibel avvisade ni helt parlamentets ändringsförslag om obligatoriska kostnadsfria posttjänster för blinda.
Vi har i kväll hört Leonard Orban säga, på kommissionsledamot Charlie McCreevys vägnar, att våra ändringsförslag inte tillför något mervärde för användarna av posttjänster.
Herr Orban! Använder inte blinda posttjänster?
Och är inte det verkliga mervärde ni talar om den faktiska merkostnad som blinda kommer att tvingas betala?
Till Markus Ferber måste jag tyvärr säga att jag tror att ni gjorde fel som accepterade en kompromiss och gav upp det krav som parlamentet godkände vid första behandlingen.
Igår underlät ni också att besvara min fråga om huruvida posttjänsterna för blinda är hotade.
Jag hoppas att ni besvarar min fråga idag.
För om det inte finns något sådant hot, vilka skäl kan ni då ha för att inte vilja ta med det i direktivet?
Om det finns ett hot visar det att vi måste ta med det i direktivet.
I Italien, Tyskland, Finland, Nederländerna, Grekland och Portugal är det postkontoret och inte regeringen som tillhandahåller dessa kostnadsfria posttjänster.
Nya och befintliga tjänsteleverantörer på en liberaliserad marknad kommer oundvikligen att försöka hålla nere kostnaderna, och då får blinda inte drabbas.
Efter liberaliseringen på Nya Zeeland upphörde posttjänsterna för blinda.
Vi får inte låta samma sak hända här.
Slutligen några ord till dem som sympatiserar med funktionshindrade personer, men som inte tycker att det här är rätt forum eller sätt att uttrycka det. Ni sa detsamma till oss om hissdirektivet och om bussdirektivet, andra exempel på inremarknadslagstiftning.
Men parlamentet sa nej, och vi insisterade på tvingande lagstiftning om tillgänglighet för funktionshindrade.
Idag måste vi återigen insistera på tvingande rättigheter för Europas blinda och synskadade.
(SK) Fru ordförande! Tack för att ni ger mig ordet.
Rådets gemensamma ståndpunkt inkluderar inte ändringsförslagen om kostnadsfria posttjänster för blinda trots att parlamentet vid första behandlingen röstade för att behålla dessa tjänster även efter liberaliseringen av den europeiska postmarknaden.
Jag hade för avsikt att rösta för ändringsförslag 3 som Eva Lichtenberger lagt fram.
I detta förslag upprepades parlamentets ståndpunkt vid första behandlingen.
Tidigare hade man enats om en kompromiss att anta direktivet om fullbordandet av gemenskapens inre marknad för posttjänster vid andra behandlingen. Efter dagens diskussion med föredraganden Markus Ferber, blev jag informerad om att godkännandet av något av ändringsförslagen skulle äventyra denna kompromiss, vilket skulle kunna betyda att man blir tvungen att ingå förlikning.
Jag inser vikten av att anta direktivet.
När det införlivats i nationell lag, kommer medlemsstaterna att kunna lösa detta problem i enlighet med principen om subsidiaritet och krav på samhällsomfattande tjänster.
Jag uppmanar därför alla medlemsstater att tillhandahålla kostnadsfria posttjänster för blinda och synskadade i enlighet med principen om subsidiaritet och kravet på samhällsomfattande tjänster.
(PL) Fru talman! Jag skulle också vilja stödja ändringsförslagen om synskadade personer.
Om EU deklarerar för alla och envar att man inte tillåter diskriminering innebär detta att tillgången till posttjänster måste vara lika för alla. För de synskadade betyder det att de får assistans i sin tillgång.
(EN) Fru talman! Det här direktivet är bara ännu ett exempel på hur oflexibel och dålig EU-lagstiftning påverkar det brittiska folket negativt.
Direktivet leder till att postkontor slår igen och till att postanställda blir arbetslösa.
Postkontoren spelar en viktig roll i samhället, i synnerhet för gamla, fattiga, personer med nedsatt rörlighet och funktionshindrade.
Detta är bara en av otaliga EU-lagar som har skadat mitt land och kommer att fortsätta göra det.
Det brittiska medborgarna är medvetna om detta och det är ett av skälen till att de inte får rösta om EU-konstitutionen.
Om konstitutionen ratificeras kan de se fram emot mycket mer av samma slag.
(EN) Fru talman! Jag anser att föredraganden i stort - om än inte helt - har uppnått en bra balans.
Genom tillhandahållandet av samhällsomfattande posttjänster garanteras konsumenterna full tillgång till posttjänster, samtidigt som medlemsstaterna flexibelt får bestämma hur de bäst och mest effektivt kan tillhandahålla de samhällsomfattande posttjänsterna.
De samhällsomfattande posttjänsterna innebär också att ett tillräckligt antal inlämningsställen måste inrättas för att fullt ut beakta användarnas behov i landsbygdsområden och glesbefolkade områden, något som jag vet kommer att välkomnas, i synnerhet i mitt hemland Irland.
Jag måste säga att jag från början hade en del reservationer när det gäller direktivets konsekvenser för de postanställda, men medlemsstaterna har fortfarande befogenhet att reglera anställningsvillkoren och kollektivavtalen inom sektorn, så detta leder inte till orättvis konkurrens.
Slutligen vill jag säga att jag stöder ändringsförslaget om obligatoriskt tillhandahållande av kostnadsfria tjänster för blinda och synskadade.
Jag är inte av samma uppfattning som Leonard Orban - eller var det kommissionsledamot Charlie McCreevy? Jag tror faktiskt att detta innebär ett mervärde, då kostnadsfria tjänster för blinda och synskadade kommer att försvinna på en fullt liberaliserad marknad, och därför är det ett mervärde om vi kan garantera dessa människor att de kostnadsfria tjänsterna finns kvar.
(SK) Fru ordförande!
Tack för att ni ger mig ordet. Först av allt skulle jag vilja tacka Markus Ferber för ett enastående betänkande.
Tack vare det kommer snart det efterlängtade direktivet att träda i kraft, vilket betyder att gemenskapens inre marknad för posttjänster kommer att vara fullständigt genomförd 1 januari 2009.
Jag är framför allt nöjd över att principen om subsidiaritet har behållits och att det konkreta implementerandet har överlåtits åt medlemsstaterna, som kommer att skapa en lagstiftning som är specifik för deras egen situation.
Jag skulle dock även vilja betona den sociala aspekten av denna lagstiftning vad gäller rättigheterna för handikappade, i synnerhet blinda eller synskadade, och deras rätt att utnyttja kostnadsfria posttjänster.
Jag uppmanar mina kolleger i parlamentet att stödja de relevanta ändringsförslag som togs upp i plenum i veckan och som antogs av parlamentet vid första behandlingen.
Dessa tjänster är adekvata och fundamentala för följande befolkningsgrupper: människor med exceptionellt låg inkomst, områden med mycket höga nivåer av arbetslöshet och människor i svåra sociala situationer, för att inte nämna de som drabbas av social uteslutning.
(EN) Fru talman! Tack för detta tillfälle att bidra till debatten.
Jag lyckönskar föredraganden till hans arbete.
Jag tror att det är allmänhetens uppfattning att denna process redan har inletts, eftersom det i många medlemsstater inte finns postservice som är likvärdig för alla regioner.
Jag är glad över att subsidiaritet ska gälla i denna fråga så att medlemsstaterna får besluta hur de bäst ska genomföra principen om en liberaliserad marknad.
Jag måste stödja min gruppordförande Richard Howitt i frågan om funktionshinder.
Tyvärr var det någon som sa att förmögna blinda kommer att gynnas.
Beklagligt nog finns det alldeles för få förmögna, blinda människor i Europa och världen.
Jag önskar att vi kunde säga att de var förmögna och berömda allihop, men så är inte fallet.
Jag menar att vi måste ta tydlig ställning i denna fråga, bara för att visa att EU visserligen handlar om fri rörlighet för kapital och tjänster, men att EU också bryr sig om dem som saknar röst och dem som inte kan se.
Rådets ordförande. - (SL) Dagens livliga debatt har visat att det finns många berättigade olika åsikter om regleringen av denna traditionella och äldsta offentliga tjänst.
Det var också riktigt att många olika åsikter och frågor uttrycktes.
Likväl måste vi poängtera att den föreslagna texten är en balanserad kompromiss mellan, å ena sidan, liberaliseringen av den inre marknaden som säkrar konkurrenskraft och det mervärde som därigenom uppstår och, å andra sidan, konsumentskydd och skydd av rättigheter för konsumenter och sårbara konsumentgrupper samt för de som bor i avlägsna områden.
I korthet är det enligt rådets uppfattning en bra kompromisstext, och jag skulle vilja uttrycka mitt stöd för denna åsikt.
Vi är också medvetna om avsikten bakom vissa ändringsförslag, men genom diskussioner i tidigare debatter framkom en slutlig kompromisslösning.
Vi anser därför att detta är en bra text, och jag hoppas att ni kommer att använda mycket politisk visdom i morgon när ni har er sista chans att stödja den.
Kommissionen. - (RO) Först av allt skulle jag vilja tacka alla deltagare i debatten och betona att denna debatt har bevisat att parlamentsledamöterna har ett stort intresse i denna fråga.
Detta intresse hör även samman med den avgörande roll som posttjänster spelar i den europeiska ekonomin och i det dagliga livet för EU-medborgarna.
Jag skulle även vilja betona att fullbordandet av denna process kommer att garantera en bestående hög kvalitet av samhällsomfattande tjänster för alla EU-medborgare och för affärsvärlden.
Huvudmålet för postreformen är att gynna alla konsumenter och användare av posttjänster, inklusive grupper med särskilda behov.
I detta sammanhang tog jag särskild hänsyn till flera medlemmars inlägg om att man även i fortsättningen ska tillhandahålla kostnadsfria tjänster för blinda och synskadade.
Kommissionen är mycket medveten om att detta är en angelägen fråga.
Vi anser att liberaliseringen av marknaden inte kommer att förändra situationen och att de internationella kraven även fortsättningsvis kommer att uppfyllas helt och hållet.
Jag skulle vilja understryka att man i den gemensamma ståndpunkten förtydligar att marknadsliberaliseringen inte kommer att förhindra tillhandahållandet av kostnadsfria tjänster för blinda och synskadade.
I enlighet med artikel 23 i direktivet måste kommissionen utarbeta en rapport om tilämpningen av direktivet, och denna rapport måste även innehålla information om ovan nämnda grupper.
Kommissionen anser att direktivet, i sin nuvarande utformning, är den bästa rättsliga ramen, och att det kommer att leda till hög kvalitet och hållbarhet hos de europeiska posttjänsterna, samtidigt som det uppfyller internationella krav.
Sammanfattningsvis anser vi att betänkandet, som det sammanställts av Markus Feber och antagits av en bred majoritet i transportutskottet, borde stödjas.
föredragande. - (DE) Fru talman, herr ordförande, herr kommissionsledamot, mina damer och herrar! Tillåt mig att bara göra några få anmärkningar.
För det första skulle jag vara glad om de medlemmar som höll passionerade anföranden för hela världen åtminstone stannade i kammaren under resten av debatten.
De gjorde mig snarare besviken och jag måste säga att jag syftar i synnerhet på ledamöter som Eva Lichtenberger.
För det andra måste jag påpeka att i det här fallet talar vi om liberalisering och inte om privatisering.
Ägandestrukturen hos de existerande posttjänsterna intresserar inte EU och nämns inte i direktivet.
För det tredje, låt mig säga att när de första posttjänsterna inrättades för 500 år sedan var det privata företag som tillhandahöll dess tjänster.
Det var inte förrän senare som regeringarna bestämde att de själva kunde göra det bättre.
Så låt oss inte snedvrida historien, tack.
För det fjärde skulle jag vilja påminna kammaren om att statliga monopol också missbrukas.
Jag är glad över att Gabriele Zimmer uppmärksammade detta problem.
Hon kommer från ett område där staten nästan helt säkert missbrukade sitt postmonopol 1990, till skada för oskyldiga människor.
Detta är en annan punkt som särskilt måste betonas i den aktuella debatten.
Låt mig göra en sak klar: vi glömde inte bort de blinda i lagstiftningen.
De är inkluderade, men på ett sätt som stämmer överens med andan i direktivet.
Genom sina bestämmelser berättar EU för medlemsstaterna att de är ansvariga för de samhällsomfattande tjänsterna och för att finansiellt se till att kravet på att tillhandahålla dessa tjänster uppfylls. De är dessutom ansvariga för att genom licensiering och tillståndsförfaranden se till att vissa tjänster, som posttjänster för blinda, kan upprätthållas på lång sikt.
Jag är kommissionsledamoten väldigt tacksam för att han har tillkännagett att kommissionen avser att ta detta i beaktande i sin rapport, i enlighet med artikel 23 i direktivet.
Vi har inte glömt någonting, vi har inte glömt de blinda.
Likväl undrar jag om blinda ska ha fri tillgång, garanterad genom EU:s lagstiftning, medan rullstolsburna inte ska ha det.
Det är också en fråga som bör övervägas.
Debatten är härmed avslutad.
Omröstningen kommer att äga rum imorgon, den 31 januari 2008.
Skriftliga förklaringar (Artikel 142)
skriftlig. - (FR) Jag välkomnar godkännandet vid andra behandlingen av rådets gemensamma ståndpunkt om ändring av 1997 års posttjänstdirektiv om fullständigt genomförande av den inre marknaden för posttjänster, och jag gratulerar min hedervärda tyska kollega Markus Ferber för det enorma arbete han har utfört.
I synnerhet är jag nöjd med att man sköt upp liberaliseringen av den allmänna marknaden till den 31 december 2010, med en tvåårig förlängning för de länder som blivit medlemmar i EU efter 2004. Jag är också nöjd med att man behållit principen om en samhällsomfattande tjänst som omfattar åtminstone en utdelning och en insamling om dagen fem dagar i veckan för alla EU-medborgare med tillräckligt många inlämningsställen på landsbygden samt i avlägsna och glesbefolkade områden.
Slutligen är jag nöjd med att man följer subsidiaritetsprincipen när det gäller sociala hänsyn - en fråga som jag hoppas att arbetsmarknadens parter kommer att arbeta med på EU-nivå.
Jag är ledsen över att bestämmelser för att skapa en europeisk regleringsmekanism inte finns med. Min sista anmärkning är att jag är angelägen att se att operatörer snart kommer överens om att införa ett EU-frimärke för försändelser som väger 50 gram, och jag har för avsikt att ta ett politiskt initiativ för detta syfte inom en snar framtid.
skriftlig. - (RO) Den gemensamma ståndpunkten tillfredsställer såväl de krav som parlamentet genom sina röster ställde inför första behandlingen som de ändringsförslag som föreslogs av utskottet för sysselsättning och sociala frågor.
Kommissionen måste emellertid alltjämt tillhandahålla tydliga undersökningar om vilka effekter liberaliseringen av posttjänsterna kommer att ha på sysselsättningen.
I sitt yttrande efterfrågade utskottet en konsekvensanalys av denna åtgärds effekter på de fem miljoner eller fler arbetstillfällen som hänger samman med eller är beroende av posttjänsterna.
Denna studie underlättas av att posttjänsterna redan har liberaliserats i åtskilliga medlemsstater, såsom Storbritannien, Sverige och Nederländerna.
Erfarenheterna i dessa länder har ännu så länge inte visat på att liberaliseringen har lett till fler arbetstillfällen inom sektorn, eller till arbeten med högre kvalitet.
Jag anser att vissa skyddsmekanismer borde tillåtas i de fall då uppkomsten av nya leverantörer av posttjänster på marknaden kommer att leda till ett stort överskott.
En av de tillgängliga mekanismerna för de drabbade företagen och medlemsstaterna skulle kunna vara Europeiska fonden för justering för globaliseringseffekter.
skriftlig. - (PL) Fru talman! Vägen till liberaliseringen av posttjänster blir längre, och detta kan man delvis beskylla parlamentet för eftersom det har förlängt kommissionens tidsfrist med två år.
De nationella delegationernas ståndpunkter speglar de olika marknadssituationerna i de 27 medlemsstaterna.
Sverige, Storbritannien och Finland, som är förgrundsgestalter för den liberaliserade marknaden, liksom Tyskland och Nederländerna, som har gått långt i den riktningen, ser alla den slutliga tidsfristen som en seger för protektionismen.
Med utgångspunkt i sin statligt kontrollerad ekonomi ser de nya medlemsstaterna inte bara det ursprungliga förslaget 2009 utan även kompromissen 2011 som ett hot för jobben i postsektorn.
I till exempel Polen har Poczta Polska 100 000 anställda, och Poczta Polska kan inte möta öppen konkurrens på medellång sikt.
Eftersom dessa länder har funnit allierade bland offentliga tjänsteföretag i Västeuropa, först och främst i Frankrikes La Poste, har de lyckats att förhandla till sig särskilda villkor som senarelägger införandet av den fria marknaden till slutet av 2012.
Således har de postanställdas gemensamma intresse vägt tyngre än intresset hos konsumenterna, som blev utsatta för hårda prövningar under julruschen i december 2007 när postmonopolets oförmåga tydligt demonstrerades.
Den långsamma utvecklingen av sektorns liberalisering på EU-marknaden, en liberalisering som började så tidigt som 1989 med det första utkastet till direktiv, visar styrkan hos de gemensamma intressen som försvarar status quo mot en utvidgning av det allmänna intresset.
skriftlig. - (EN) Än en gång ser vi ett ideologiskt motiverat förslag, denna gång om posttjänster.
Det har inte föregåtts av någon analys av sociala konsekvenser, och inget seriöst samråd med postkontor, anställda eller konsumenter.
Det finns ingen efterfrågan på att marknaden för posttjänster ska liberaliseras, ingen logik i och inga skäl till att göra det.
Folk vill inte ställas inför en rad konkurrerande postkontor som marknadsför sina produkter.
De vill inte att deras lokala postkontor ska slå igen bara för att marknaden inte är tillräckligt lönsam för de privata postföretag som kommer att översvämma marknaden och tvinga offentliga operatörer som An Post på knä.
Folk vill ha en pålitlig postservice som levererar deras post så smidigt som möjligt och låter de lokala postkontoren ligga kvar mitt i de samhällen de betjänar.
Hur ska folk kunna ta idén om ett EU som främjar ett socialt Europa på allvar när man med detta förslag slår ännu en spik i dess kista?
Det är dags att sätta stopp för den ideologiskt motiverade tvångsmarschen mot liberalisering och privatisering.
Det irländska folket har möjlighet att hejda detta genom att rösta nej till Lissabonfördraget.
Jag är för att en liberalisering av marknaden genomförs så snabbt som möjligt och jag välkomnar det direktiv som fullbordar genomförandet av den inre marknaden för posttjänster.
Nedläggningen av små postkontor i Estland har retat upp befolkningen, men det är tydligt att efterfrågan på traditionella posttjänster har avtagit i och med att ny teknik som till exempel Internet har börjat användas.
Om det finns konkurrens kan en ny affärsverksamhet för Internetbaserade tjänster växa fram, och detta måste välkomnas.
Jag förstår även medlemsstaternas behov av att få ett fastställt datum.
Det är därför viktigt att principen om ömsesidighet tillämpas när medlemsstater tillåts vägra att öppna sina marknader för tillhandahållare av posttjänster från grannstater vars tillhandahållare skyddas av lagen.
Viktigt är också att samhällsomfattande posttjänster är garanterade för alla, även för de som är bosatta i avlägset belägna områden eller på öar.
Posttjänsterna måste ha rimliga priser, hålla hög kvalitet och vara tillgängliga för alla.
Det är nödvändigt att utarbeta planer för kostnadsrelaterade samhällsomfattande posttjänster, eftersom man ser olika på konceptet i olika medlemsstater.
Jag tror att det finns skäl till att kräva att kostnadsöverväganden för alla tjänster ska vara undantagna från indikatorn för de samhällsomfattande posttjänsterna.
skriftlig. - (DE) En liberalisering av posttjänsterna kommer att ske i hela EU - inte 2009 som ursprungligen planerats, men 2011.
Ekonomiskt sett är postsektorn mycket viktig och den har även inverkan på andra ekonomiska sektorer.
Precis som på alla andra områden med ekonomisk verksamhet är det klokt med mer konkurrens vid leverans av postförsändelser.
Inte bara företagen gagnas av detta, utan även konsumenterna får stora fördelar.
Så blir dock inte fallet om de grundläggande villkoren inte stämmer.
Med andra ord måste man garantera att breven precis som tidigare kommer att levereras på ett effektivt sätt och till rimliga priser.
Man måste se till att de allmänna bestämmelserna för samhällsomfattande posttjänster är garanterade på lång sikt - och detta överallt, även i avlägset belägna områden.
Särskilt viktigt är att det finns goda arbetsvillkor och framför allt arbetstrygghet för alla som arbetar med posttjänster.
Det är också viktigt att samma villkor gäller för verksamhet hos alla tillhandahållare av posttjänster.
Det fastslogs klart och tydligt redan från början att det här inte skulle vara en tygellös liberalisering.
Vi måste skapa bra och hållbara förutsättningar för alla - postföretagen, deras anställda och naturligtvis också deras kunder.
skriftlig. - (FI) Öppnar man upp för fri konkurrens för posttjänster kommer detta oundvikligen att innebära en försämring av tjänsterna, särskilt i glest befolkade länder som Finland.
Posten bör vara en offentlig tjänst, och vi måste garantera att den har tillräckligt med kapital genom att använda de pengar som tjänas in via tjänster som är ”lätta” att förvalta, för att kunna bistå de områden som är ”svårare”.
En nation som vill bevara sin sammanhållning och gemenskapskänsla kommer inte att privatisera offentliga posttjänster.
Vi är också beroende av en offentlig tjänst för att kunna garantera integritetsskydd och det slags säkerhet som vi kräver av posten.
Privatisering skulle kunna resultera i en osund personalpolitik som skadar förtroendet för posten.
Av denna anledning röstar vår grupp emot rådets ståndpunkt om privatisering.
skriftlig. - (EN) Liberaliseringen av marknaden för posttjänster är ett viktigt område för den europeiska inre marknaden.
Medan den här diskussionen har pågått har det funnits många frågetecken kring de samhällsomfattande posttjänsterna.
Jag tror att vi kan luta oss mot erfarenheterna från en del europeiska postmarknader som redan har avreglerats.
Posttjänsterna har tryggats i dessa länder, samtidigt som kvaliteten och servicen har förbättrats genom en mer affärsmässig verksamhet.
Samtidigt möter jag när jag reser omkring i Europa dålig och långsam service i många av de länder som försöker få så många undantag som möjligt från den planerade liberaliseringen.
Dessutom ger det här betänkandet medlemsstaterna stor handlingsfrihet vid genomförandet av liberaliseringen.
Många av de källor till oro som har nämnts kan på så vis hanteras av de nationella myndigheterna.
Jag vill tacka Markus Ferber för hans envishet i hanteringen av denna mycket besvärliga process.
skriftlig. - (RO) En fullständig liberalisering av posttjänsterna i medlemsstaterna kommer inte bara ha en positiv inverkan på användarna av posttjänster och konsumenterna, vilka kommer att dra fördel av nya och innovativa tjänster och lägre postavgifter, utan även på medlemsstaternas ekonomi totalt sett.
Det direktivförslag som diskuteras är komplett i sin nuvarande form, då det för vissa medlemsstater är möjligt med en förlängning av fristen för en fullständig liberalisering av marknaden för posttjänster.
Rumänien är ett av de länder som gagnas genom de nya bestämmelser som antagits av Europaparlamentet.
De rumänska leverantörerna av samhällsomfattande tjänster är under omstrukturering enligt ett program för 2007-2010 som antagits av den rumänska regeringen, och förberedelserna för liberalisering kommer att påbörjas först därefter.
Detta tidsschema gagnar de rumänska konsumenterna, eftersom en liberalisering av marknaden efter den 1 januari 2013 innebär tjänster med förbättrad kvalitet till överkomligt pris.
Inkomna dokument: se protokollet
8. (
Kontroll av gemenskapsrättens tillämpning 2005 (debatt)
Nästa punkt är ett betänkande av Monica Frassoni, för utskottet för rättsliga frågor, om kommissionens tjugotredje årsrapport om kontroll av gemenskapsrättens tillämpning (2005).
Herr talman, mina damer och herrar! Tillämpningen av gemenskapslagstiftningen är en central del av agendan för bättre lagstiftning som lanserats av Barrosokommissionen.
Under en tid har den varit ett slags Askungen, förlorad i trenden med konsekvensanalyser och kostnadsminskning.
I dag har kommissionen börjat rätta till detta, delvis på grund av påtryckningar från parlamentet.
Detta är ett förfarande som under flera år ofta bara har varit en form av byråkratiskt malande, där en överträdelse följer en annan utan mycket väsen, men det är ändå ett helt avgörande förfarande.
Siffrorna talar sitt tydliga språk.
Hittills har omkring 2 518 överträdelseförfaranden inletts i de mest skiftande sektorer, särskilt miljön och den inre marknaden.
Utöver detta mottar parlamentet vare år hundratals, till och med tusentals, framställningar som ofta hänvisar till specifika överträdelser av gemenskapslagstiftningen, inför vilka medborgarna känner sig hjälplösa och därför vänder sig till parlamentet.
Frågan är: Vilken chans har de att få upprättelse?
Överträdelseförfarandet beskrivs i artiklarna 226 och 228 i fördraget, och därför finns det inte mycket utrymme för kreativitet.
De gällande reglerna tvingar oss till långsamma, röriga förfaranden där den effektivaste åtgärden - böter - sällan tillämpas och bara efter en mycket lång tid, till och med årtionden.
Emellertid kan faktiskt en hel del göras, och jag tackar kommissionen för att den under de senaste två åren, och i september förra året i ett särskilt meddelande, har föreslagit en rad åtgärder som analyseras och utvärderas i mitt betänkande, och om vilka jag skulle vilja komma med några kommentarer.
För det första, tillåt mig dock att komma med en anmärkning som jag anser är avgörande för denna debatt, eftersom genomdrivande av lagar kan vara en mycket politisk fråga och kan vara ett enastående verktyg för att öka gemenskapsinstitutionernas trovärdighet och synlighet.
Jag skulle vilja nämna två specifika exempel på lite annorlunda beteenden från kommissionens sida: sopkrisen i Neapel och motorvägen Via Baltica i Rospudadalen i Polen.
Sopkrisen i Neapel var en direkt konsekvens av överträdelser, som skedde år efter år, av praktiskt taget alla gemenskapsregler om avfall.
En stor mängd överträdelseförfaranden hade inletts mot Italien under åren, och domstolen hade uttalat sig mot Italien vid många tillfällen.
Men först nu, flera år senare, när situationen har blivit oacceptabel för alla och omöjlig att dölja, har kommissionen beslutat att slå näven i bordet.
Kommissionens besök följs med stort intresse, och medborgare som protesterar mot olaglig avfallshantering meddelar på tv att framställningar skickas till Europaparlamentet.
Jag undrar: skulle detta inte ha kunnat göras tidigare?
Skulle vi verkligen inte ha kunnat inta en annorlunda hållning för att förhindra denna situation?
Jo, det kunde vi ha gjort!
Detta är faktiskt vad kommissionsledamot Stavros Dimas gjorde i fallet med Rospudadalen i Polen, som riskerade att förstöras av infrastrukturen för Via Baltica.
För första gången begärde kommissionsledamoten ett beslut om suspendering från domstolen, och detta beviljades.
Detta är ett mycket viktigt prejudikat som utsänder ett mycket tydligt budskap: Kommissionen kan och måste vara bestämd och tydlig mot medlemsstater som agerar som om inget hade hänt, och den måste använda alla de verktyg som det demokratiska systemet tillåter: medierna och den allmänna opinionen.
En av de viktigaste innovationerna som kommissionen introducerar i meddelandet gäller ett ”nytt” arbetssätt.
Vi har uttryckt många tvivel om detta nya arbetssätt, som till största delen består i att skicka ut klagomål direkt tillbaka till den medlemsstat mot vilken klagomålet har riktats, för att försöka att lösa problemet.
Vi gav uttryck för dessa tvivel, och kommissionen gav oss några försäkringar som jag hoppas att vi också kommer att höra i dag, men vi kommer att hålla ett mycket vaksamt öga på frågan och hoppas verkligen att, i fråga om överträdelseförfarandena, öppenheten och möjligheten att ”peka ut” medlemsstater samt det gemensamma arbetet med parlamentet kommer att leda till framsteg.
Vid slutet av debatten kommer jag att tala igen under två minuter för att använda min talartid.
ordförande för rådet. - (SL) Tack, herr talman, mina damer och herrar!
Fru Frassoni! För rådets räkning skulle jag vilja välkomna ert betänkande om kommissionens årsrapport om kontroll av gemenskapsrättens tillämpning, och den ytterligare analys som framställs i kommissionens meddelande ”En Europeisk Union som bygger på resultat - tillämpningen av gemenskapsrätten”.
Enligt vår uppfattning är Europaparlamentets betänkande ett mycket nyttigt bidrag till vårt gemensamma mål att säkra en lämplig och korrekt tillämpning av gemenskapslagstiftningen.
För rådets räkning skulle jag vilja välkomna slutsatserna i Monica Frassonis betänkande, som enligt vår uppfattning är av central betydelse, nämligen att säkrandet av gemenskapsrättens positiva effekter på EU-medborgarnas dagliga liv främst beror på hur effektiv EU:s politik är och på tillsynen och kontrollen av medlemsstaternas metoder för att efterleva gemenskapsrätten.
Vi är positivt inställda till Europaparlamentets åtagande att stödja utbytet av bästa praxis bland medlemsstaterna.
Enligt vår uppfattning skulle sådana utbyten på ett avgörande sätt bidra till en effektivare och mer enhetlig tillämpning av gemenskapsrätten.
Jag måste förklara här att rådets ordförandeskap inte kan kommentera de flesta av de frågor och förslag som framlagts i detta värdefulla betänkande.
Som vi vet är det administrativa genomförandet av gemenskapsrätten i princip medlemsstaternas ansvar i enlighet med deras konstitutionella bestämmelser, och kommissionens ansvar. I egenskap av fördragens väktare är kommissionen ansvarig för övervakning och enhetlig tillämpning av gemenskapsrätten.
Herr talman, herr rådsordförande, mina damer och herrar! Kommissionen är tacksam för möjligheten att diskutera dessa viktiga frågor med Europaparlamentet i dag, och jag är mycket tacksam över Monica Frassonis betänkande och bidrag, som innehåller viktiga punkter.
Jag kan försäkra er, fru Frassoni, att kommissionen tar era synpunkter på största allvar.
Europeiska unionen är en gemenskap under rättsstatsprincipen och som sådan är den unik i världen.
Bara lagen kan garantera de friheter som medborgarna har rätt till, och bara lagen kan forma marknadsekonomin på ett sådant sätt att den verkar till allas fördel.
Europeiska kommissionen är fördragens väktare.
Dess roll är att se till att gemenskapsrätten genomförs överallt och att den tillämpas korrekt på alla platser.
Till och med de bästa lagar har inget värde så länge de bara finns på papper.
Varje utskott kommer därför att finna att en av dess viktigaste uppgifter är att se till att vår lagstiftning inte bara består av tomma ord.
I fördragsbrottsförfarandena och EG-domstolen har vi ett kraftfullt verktyg.
Detta vapen måste användas när det inte finns något annat sätt att avhjälpa lagöverträdelser.
Det är dock inte ett självändamål, och det skulle kunna bli ett trubbigt verktyg om det överanvänds.
Kommissionen anser inte att antalet fördragsbrottsförfaranden är ett mått på det allvar och den beslutsamhet med vilken den kontrollerar hur väl gemenskapsrätten efterlevs.
Snarare anser kommissionen att det är en fråga om att hitta lösningar på problem.
Det verkliga måttet är hur många problem med tillämpningen av gemenskapsrätten som vi har löst, och hur pass snabbt.
Vi har kritiskt sett över vårt arbetssätt och kommit fram till följande slutsatser: när problem väl har fastställts måste de hanteras snabbt och effektivt.
Medborgare och näringslivet har rätt till snabba svar.
Därför, fru Frassoni, kommer jag att återvända till kommissionen med vad ni har sagt om avfall i Kampanien, och detta ämne kommer att behöva diskuteras.
Jag håller helt med om att ett noggrant, snabbt och beslutsamt arbetssätt är helt avgörande där gemenskapsrätten uppenbarligen förbigås.
En strategi grundad på partnerskap är i princip att föredra framför en som präglas av konfrontation.
Kommissionen vill därför se mer dialog och mer öppenhet i dessa frågor.
Vi vill också göra tydliga prioriteringar: hantera de viktigaste frågorna först, och snabbt, och inte skjuta myggor med kanoner.
Vi måste också se till att nödvändiga resurser finns tillgängliga.
Tillåt mig att komma med en kommentar i denna fråga.
Om problemen hopar sig i samband med tillämpningen av gemenskapsrätten i särskilda frågor kan detta vara för att lagen i sig själv är otydlig eller motsägelsefull.
Vi bör inte från början anta att medlemsstaten har en dålig inställning.
Som en konsekvens av dessa överväganden tog vi ett antal steg, och jag skulle vilja säga från början att vi kommer att fortsätta att ta till fördragsbrottsförfaranden och inleda dem omedelbart när den nödvändiga informationen finns tillgänglig.
Emellertid föreslår vi ett nytt arbetssätt, med vilket vi hoppas få den nödvändiga informationen snabbare.
Denna metod grundar sig på att förbättra samarbetet med medlemsstaterna innan det kommer till ett stadium där officiella förfaranden inleds, utom självklart - och detta är mycket viktigt, fru Frassoni - om det från början är uppenbart att ett fördrag med all sannolikhet överträds.
I sådana fall är vårt första steg inte att tala med medlemsstaterna, utan att agera.
Det är inte en helt ny process, utan ett inledande förfarande där vi kräver ytterligare förfaranden för att nå en lösning snabbare utan att inleda fördragsbrottsförfaranden.
Alla förfrågningar och klagomål besvaras direkt och snabbt och, beroende på fakta i frågan, kan de leda till fördragsbrottsförfaranden.
Detta innebär att varje inlägg registreras och behandlas.
Om det formuleras som ett klagomål, eller kan ses som ett klagomål, behandlas det som ett klagomål, och kommissionen vidtar lämpliga åtgärder.
Vi testar för närvarande denna nya arbetsmetod i en pilotfas.
Femton medlemsstater deltar i pilotprojektet, som har utformats för att säkra att vi faktiskt gör framsteg.
Naturligtvis kommer vi att informera parlamentet om resultaten från pilotfasen och diskutera eventuella ytterligare steg med parlamentet.
I alla fall är vi redan i en position där vi kan hitta en lösning på 90 procent av alla problem som kommer till vår kännedom utan att dra ärendet inför domstol.
Emellertid delar vi er åsikt att detta bör göras snabbare.
En övergång till en beslutprocess varje månad, som inleddes i januari, borde hjälpa.
Detta säkrar snabbare, effektivare genomförande av fördragsbrottsförfaranden.
Vi strävar efter att göra hela processen så öppen för insyn som möjligt samtidigt som vi bevarar konfidentialiteten i lämplig utsträckning, vilket EG-domstolen kräver att vi gör.
Allmänheten kommer att via Internet ha tillgång till regelbundet uppdaterade sammanfattningar av alla fördragsbrottsförfaranden som för närvarande dragits inför EG-domstolen.
För att uppnå öppenhet och rättssäkerhet behöver vi också veta hur medlemsstaterna tillämpar gemenskapsrätten i sina respektive nationella sammanhang.
Därför behöver vi jämförelsetabeller - vilket begärs i betänkandet - som tydligt visar genomförandestatusen i varje medlemsstat.
Jag tror att vi alla här delar samma mål.
Vi vill ha en gemenskapsrätt som EU-medborgarna kan ha fullt förtroende för.
föredragande för yttrandet från utskottet för framställningar. - (EN) Herr talman! Under den minut som jag har för utskottet för framställningars räkning vill jag göra tre saker.
För det första skulle jag vilja tacka Monica Frassoni för hennes samarbete om denna årsrapport, men mest av allt skulle jag vilja visa hur viktigt utskottet för framställningar är i detta förfarande för övervakning och genomförande.
Jag tror att denna betydelse slutligen har erkänts av kommissionen.
Jag tackar kommissionsledamoten för detta, eftersom vi i denna fråga verkligen borde ha ett partnerskap mellan våra båda institutioner, och särskilt med deltagande av utskottet för framställningar, vilket faktiskt är våra ögon och öron som lagstiftare, tack vare våra medborgare som kommer till oss med direkta problem som de upplever.
Men för att våra medborgare ska kunna göra detta kommer jag till min andra punkt.
Herr kommissionsledamot! Ni talade om att vår rätt är en levande rätt.
För att det ska vara en levande rätt behöver den vara begriplig för våra medborgare.
Jag har fört en lång dialog med er kollega Margot Wallström om sammanfattningar för medborgarna, så att medborgarna förstår våra lagar.
Hon har vid många tillfällen lovat oss att dessa kommer att komma med varje rättsakt.
Vi väntar fortfarande på verkliga bevis för att detta ska ske.
Avslutningsvis behöver utskottet för framställningar - och detta riktar jag till mina egna kollegor - en mycket mer framträdande plats och större resurser i vårt eget parlament.
Det är inte bara ett beskäftigt utskott som lägger sig i.
Det gör ett verkligt jobb genom att anknyta till våra medborgare inom detta område.
för PPE-DE-gruppen. - (EL) Herr kommissionsledamot! Ni har helt rätt.
Rättsstatsprincipen är grunden för EU. Ni påpekade korrekt att gemenskapsrätten är rätta sättet att uppnå målen med EU-fördragen, eftersom dess typexempel är de europeiska medborgarnas intresse, som har rätt att begära att denna lag genomförs.
Lagstiftningens omfattning, bredd och komplexitet ökar hela tiden.
Vi parlamentsledamöter från Europeiska folkpartiet skulle vilja uttrycka vår belåtenhet. Genom sin tjugotredje årsrapport om kontroll av gemenskapsrättens tillämpning och även genom tillkännagivandet av resultaten i EU visar kommissionen sin önskan att vara fördragens väktare och att se till att lagstiftningen genomförs.
Ni har helt rätt i att vi vill ha jämförelsetabeller, om vilka rådet fattade ett beslut i dag.
Föredraganden samarbetade mycket med er för att upprätta Monica Frassonis betänkande, som vi hade en intressant utfrågning om i parlamentet.
Låt oss säga er att vi också vill att parlamentet ska delta i kontrollförfarandet och att vi önskar hållas underrättade om er verksamhet.
Vi vill att ni kommer till våra utskott, såsom ni kommer till utskottet för miljö, folkhälsa och konsumentfrågor.
Vi vill höra er lägesrapport.
Vi vill att ni beaktar de framställningar som vi mottar, vilket ni påpekar i ert betänkande.
Vi skulle också vilja betona att vi, när det gäller våra beslut om immunitet, skulle vilja att ni ingriper för att se till att nationella domstolar upprätthåller dessa.
Genomförandet av gemenskapsrätten låter europeiska medborgare hoppas att demokrati, lag och ordning kommer att stärkas, och att EU:s myndigheter kommer att närma sig dem.
I dag, efter resolutionen om det nya reformerade Lissabonfördraget, önskar vi alla en bättre framtid för EU.
Herr talman! Ett mål med gemenskapsrätten är att EU ska kunna genomföra olika politiska strategier.
Tillämpningen av denna lagstiftning bör vara en prioritet för alla medlemsstater som, samtidigt som de är underställda kontroll och övervakning från kommissionens sida, kommer att garantera att lagstiftningen har de önskade positiva resultaten för EU-medborgarna.
Under tidigare år har det totala antalet förfaranden som inletts av kommissionen för att hantera överträdelser av rättsliga bestämmelser stadigt ökat, för att 2005 uppgå till nära 2 700.
Trots EU:s utvidgning med 10 nya stater har det under de följande åren inte blivit någon generell ökning av antalet överträdelser.
Det finns dock en fara att denna situation kan ha uppstått på grund av en brist på registrerade klagomål, eller på grund av administrativa problem inom de institutioner som är ansvariga för att beakta överträdelser.
Betänkandet bör lovordas först och främst för att det inkluderar detaljerade undersökningar av överträdelser i samband med framställningar, samt den information som tillhandahållits om enskilda generaldirektorats villighet till ett brett samarbete i sådana frågor.
Vi bör också välkomna kommissionens omfattande meddelande ”En Europeisk Union som bygger på resultat - tillämpningen av gemenskapsrätten”.
Emellertid behöver kommissionen mer i detalj utarbeta frågorna om tillgängliga medel för att beakta överträdelser, förfarandenas längd i fall av överträdelser, den begränsade tillämpningen av artikel 228 i fördraget och utvärderingen av hur prioriteringskriterierna tillämpas.
Den föreslagna nya arbetsmetoden som införs 2008, som ett pilotprojekt som inbegriper flera medlemsstater och som syftar till att effektivisera aktuella förfaranden, förtjänar erkännande.
Men ett skede i förfarandet ger anledning till oro, nämligen att ärendet skickas till en berörd medlemsstat som framför allt är den part som är ansvarig för en oriktig tillämpning av gemenskapsrätten. Detta kan leda till en försvagning av kommissionens roll som fördragens väktare.
Skapandet av gemenskapsrätten bör möta medborgarnas problem på ett sådant sätt att det möjliggör att snabba svar kan ges på deras frågor och klagomål, vilket kommer att göra det lättare för dem att förstå och utnyttja sina rättigheter, medan man samtidigt effektivt minskar antalet förfaranden som gäller lagöverträdelser.
Låt mig slutligen varmt gratulera Monica Frassoni till ett mycket väl förberett dokument.
för ALDE-gruppen. - (EN) Herr talman! Jag skulle vilja rikta uppmärksamheten mot våra tre institutioner och betona hur viktigt det är att var och en av dessa deltar i den genomförande och övervakande rollen.
Det står helt klart att vi här tittar på kommissionens rapport.
Självklart har kommissionen det främsta ansvaret för genomförande och genomdrivande, och vi vill inte trampa den på tårna i detta avseende.
Jag anser dock att kommissionen kan räkna med att vi i framtiden kommer att hålla en mycket noggrannare uppsikt.
Vi är tacksamma över att många av de lärdomar som togs upp i vårt betänkande om Equitable Lifes fall har tagits in.
Men när vi går över i en ny period och kanske prövar några nya idéer måste vi vara mycket försiktiga.
För det första, om vi ser på rådet, återstår det fortfarande för oss att komma överens - och jag var nöjd över att höra kommissionsledamoten nämna det - om tanken på jämförelsetabeller för varje rättsakt, så att alla kan se exakt vad som sker på medlemsstatsnivå och var varje rättsakt passar in.
Pilotprojektet är en utmärkt idé.
Det är i sin ordning, så låt oss se hur det fungerar.
Men - och här är problemet - jag är lite skeptisk över att så många medlemsstater har skrivit på detta.
Jag hoppas att de inte upplever det som ett lätt val, och jag hoppas att kommissionen kommer att ta dem ur villfarelsen att detta på något sätt skulle vara fallet.
Slutligen kommer jag till vårt eget parlament.
Tydligen måste vi efter Lissabonfördraget ha en mycket större roll när det gäller övervakning.
När vi har slutbehandlat en rättsakt här kan vi inte anta att det är det sista som händer.
Våra utskott kommer att behöva anta en mycket större roll när det gäller kontroll.
En eller två genomföranderapporter görs redan - detta kommer att öka - och vi kommer att behöva axla vårt ansvar, tillsammans med de andra institutionerna.
Bara som ett postskriptum - men ett mycket viktigt sådant - måste vi också rikta uppmärksamheten mot utbildningen av vår domarkår vid våra nationella domstolar för att se till att även de vet hur de ska genomföra gemenskapsrätten.
för Verts/ALE-gruppen. - (EN) Herr talman! Jag gratulerar min gruppkollega och gruppens vice ordförande Monica Frassoni till en lägligt och väl uttänkt betänkande.
Jag instämmer helt i Diana Wallis' kommentarer.
Att stifta lagar är vår uppgift, men genomförandet av lagar ger faktiska resultat för våra folk, och ett misslyckande att genomdriva lagar får oss ärligt talat att se dumma ut.
Jag gratulerar kommissionen till ett antal åtgärder som har varit mycket positiva.
Men vi måste verkligen föra upp detta högre på vår dagordning här i parlamentet. I Skottland finns det utan tvekan ännu ett starkt intryck av att det finns en lag för ett land och en annan lag för ett annat.
Jag är mycket medveten om att inte allt detta är kommissionens fel, men vi måste alla fullgöra vår uppgift i att lösa detta om vi är ett enda EU.
Så när jag gratulerar min gruppkollega är jag glad över att höra att många av dessa punkter kommer att tas upp av kommissionsledamoten.
Jag skulle vilja komma med en kommentar till, särskilt i samband med miljölagstiftningen, där många av konflikterna uppkommer.
Många av de mycket hedervärda målen i enskilda rättsakter står i konflikt med varandra, och vi måste inse detta när vi utarbetar dem.
Det finns knapphändig vägledning för lokala myndigheters tillämpning i fråga om hur de bör hantera de ofta mycket goda målen när dessa är motstridiga.
Vi utlovades en översyn av detta i energipaketet, så om vår kommissionsledamot skulle kunna upplysa oss om denna pågående process skulle jag vara mycket tacksam.
(NL) Herr talman! Även jag vill gratulera Monica Frassoni till hennes betänkande.
Vi har nu behandlat ett antal betänkanden om genomförandet av gemenskaprätten, och en tydlig gemensam tråd löper genom dessa betänkanden.
Detta innebär ökad uppmärksamhet på genomförandet, även från Europaparlamentets sida.
Vi kan nu använda oss av genomföranderapporter.
Jag kommer själv att lägga fram en rapport om genomförandet av det åttonde direktivet om tillsyn av revisorer i juli.
Det är bra att parlamentet även tar en ordentlig titt på införlivandet av gemenskapsrätten i medlemsstaternas lagstiftning.
Jag vill inrikta mig på frågan om tillsynsmyndigheter i detta sammanhang.
Vi talar om införlivandet av lagstiftningen av myndigheterna i medlemsstaterna och om de rättsinstanser som tillämpar lagstiftningen.
Många medlemsstater har emellertid oberoende tillsynsmyndigheter som tillämpar och utarbetar lagstiftning.
I praktiken har stora skillnader uppstått mellan de olika medlemsstaterna och tillsynsmyndigheterna.
Företag från flera medlemsstater som är verksamma internationellt ställs allt oftare inför problemet med skilda krav från olika tillsynsmyndigheter i olika medlemsstater.
Detta är ytterst olämpligt och hämmar den inre marknadens fungerande.
Jag vill diskutera ytterligare en punkt.
Vi kan inte heller undvika en ytterligare granskning av de lagstiftningsinstrument som tillämpas inom EU.
Hittills har vi huvudsakligen arbetat med direktiv när det gäller harmoniseringen.
Kommissionsledamot Günter Verheugen har redan vid flera tillfällen förklarat att det inför framtiden är vettigt att utnyttja regleringsinstrumenten inom ramen för inremarknadslagstiftningen i högre grad för att undvika alla möjliga problem, som cherry picking eller gold-plating, dvs. selektiv eller överdriven tolkning, under införlivandet av direktiven.
Jag vet att man även i de nationella parlamenten, särskilt i det nederländska parlamentet, sakta men säkert börjar inse att genomförande som omfattar selektiv eller överdriven tolkning kan skada den inre marknadens fungerande och även de nationella ekonomierna.
Eftersom det förhåller sig på det viset är steget mot reglering, där det är möjligt, inte längre så stort.
(ES) Herr talman! Vi är medvetna om hur viktigt ert uppdrag att övervaka tillämpningen av gemenskapsrätten är.
Vi talar om förhållandet mellan en överstatlig institution och nationella regeringar.
De nationella regeringarna är starka organ med stor makt; de är offentliga myndigheter.
Normalt sett är kommissionen EG-rättens och medborgarnas väktare, och i många fall är kommissionen den enda garanti som medborgarna har (eftersom EG-rätten är lagstiftning) för att den kommer att tillämpas korrekt.
Målsättningen med Monica Frassonis betänkande är att förstärka det som jag skulle vilja kalla kommissionens ryggrad, för att kommissionen ska vara medveten om denna uppgift och för att den, om vi vill ha en föregående förhandlingsfas med regeringarna om de svårigheter som kan uppstå, när det verkligen gäller agerar som medborgarna förväntar sig, kraftfullt och energiskt, och tillämpar gemenskapsrätten.
Det är oroande att vi efter utvidgningen har intrycket av att kommissionen tillämpar mindre strikta kriterier för de nya medlemsstaterna än den tillämpade för de gamla.
Detta skulle inverka negativt på EU:s konsolidering och anseende i dessa medlemsstater.
Eftersom jag har följt många av kommissionens överträdelseförfaranden kan jag försäkra kommissionen om att när den ingriper känner sig medborgarna, och även de offentliga myndigheterna, styrkta av kommissionens agerande på detta område.
Med andra ord anser jag att syftet med parlamentets betänkande, det förslag som Monica Frassoni har lagt fram, och även yttrandet från Diana Wallis, är att stärka kommissionen, så att den inte känner att den står ensam och försvarslös mot regeringarna, utan vet att den har parlamentet bakom sig för att förstärka den tillsyns- och övervakningsroll som kommissionen har över tillämpningen av gemenskapsrätten.
(DA) Herr talman! EU-medborgarna är av avgörande vikt för EU:s lagstiftning.
De är inte bara offren för de överträdelser som begås, som till exempel i Neapel, utan har ofta varit nyckelaktörer i många miljöfrågor.
De vakar som vakthundar för att försäkra sig om att lagstiftningen tillämpas korrekt överallt i EU, och i många fall är medborgarna de enda som gör detta.
Därför bör EU också stödja medborgarna genom att säkra en stark ställning för dem.
När de uppmärksammar överträdelser av gemenskapsrätten bör deras klagomål behandlas seriöst och med respekt.
Jag hoppas uppriktigt att detta inte är ett försök från kommissionens sida att sätta stopp för många av dessa klagomål, eftersom det skulle vara ett dåligt agerande.
Jag vill därför tacka Monica Frassoni för att hon har uppmärksammat dessa risker.
Hennes utmärkta betänkande blir nu ett viktigt generellt steg i rätt riktning.
EU-medborgarnas ställning kommer att stärkas genom Lissabonfördraget, men om det ska bli något annat än en meningslös prydnad måste medborgarnas bidrag till EU tas på allvar.
(PL) Herr talman! Även jag vill gratulera Monica Frassoni till ett utmärkt betänkande.
Jag vill även säga att jag är mycket nöjd med att de tio nya medlemsstaternas anslutning inte har påverkat antalet registrerade överträdelser enligt den statistik som kommissionen har lagt fram om antalet förfaranden som gäller överträdelser av EU-lagstiftningen.
Statistiken ger emellertid inte hela bilden.
En av de viktigaste mekanismer som vi har för att kontrollera hur väl EU-lagstiftningen verkligen tillämpas är systemet med förhandsavgöranden, vars målsättning är att hjälpa de lokala domstolarna att tillämpa EU-lagstiftningen enhetligt i alla medlemsstater.
Det grundläggande problemet med detta förfarande är väntetiden på ett svar från EG-domstolen, som fortfarande är mycket lång (omkring 20 månader).
Det huvudsakliga skälet till väntetiden - den tid som översättningen tar - utgör cirka nio månader.
Det är oroande att vi från många nationella parlament hör krav på ett tak för budgeten, särskilt för skriftliga översättningar.
Kommissionens rekommendationer till medlemsstaterna och kandidatländerna bygger på antagandet att EU-lagstiftningen kommer att kunna införas effektivt om man anställer personal med passande kvalifikationer och anslår lämpliga resurser.
Jag håller inte helt med om den åsikten.
Antalet anställda och tillgängliga medel är inte den rätta måttstocken.
Det krävs även beslutsamhet och engagemang i arbetet för att införa EU-lagstiftningen.
För att utföra de uppgifter som medlemsstaterna och kandidatländerna ställs inför krävs tre faktorer: kunskap, kompetens och vilja.
Den första av dessa faktorer - det vill säga att besitta kunskap - är inte ett problem i dag.
Den andra faktorn - förmågan att införliva det som har åstadkommits av gemenskapen - är kopplad till frågan om att ha tillgång till lämpliga medel och kunna anställa mer personal.
För närvarande lägger kommissionen mest tonvikt vid just denna aspekt.
Den tredje faktorn - att de som har ansvar för att införa och tillämpa EG-rätten har en vilja att göra detta - är den mest underskattade.
Viljan att tillämpa EG-rätten beror i praktiken på institutionerna och hur systemet för förfaranden, incitament och begränsningar är utformat.
Om införandet av EU-lagstiftningen blir en framgång eller ett misslyckande avgörs i sista hand av varje specifik institutionell modell.
Kunskap och pengar är inte allt.
En god vilja att agera krävs också.
(DE) Herr talman! Herr vice ordförande, i ert inledningsanförande förklarade ni att kommissionen inte vill treva i blindo, utan ta reda på om något behöver göras genom att diskutera det med medlemsstaterna.
Inom kommissionen - som trots allt är en kollegial institution - är man emellertid inte alltid enig om vissa frågor.
På transportområdet anser jag att det för närvarande finns en fråga som kommer att bli alltmer problematisk för oss under de kommande åren - och förmodligen även inom kommissionen - och det är konceptet att pengarna ska riktas om till miljövänligare transportsätt genom att korssubventionera inkomster som intjänats på ett mindre miljövänligt område - vägtullar, parkeringsavgifter osv. Detta är i själva verket en subvention.
Har denna fråga diskuterats, och hur ser situationen ut?
(HU) Tack, herr talman.
Som flera talare före mig redan har nämnt kommer våra framgångar när det gäller att nå de mål som fastställs i fördragen att bero på hur effektivt medlemsstaterna tillämpar gemenskapsrätten och hur de införlivar den i den nationella lagstiftningen.
Om de misslyckas med att tillämpa eller verkställa lagstiftningen på lämpligt sätt eller inte kan uppfylla lagstiftningens målsättningar fullt ut kommer vi att få problem.
Under de senaste åren har tendensen förbättrats när det gäller efterlevnaden av lagstiftningen, och jag anser att de tio nya medlemsstaternas efterlevnad av lagstiftningen är god.
Jag hoppas att detta inte beror på att kommissionen har mer överseende med oss, med de nya medlemsstaterna, utan att det beror på att vi gör verkliga insatser för att uppfylla kriterierna och infria förväntningarna.
Att hitta fram i den byråkratiska djungeln är tyvärr fortfarande långtifrån enkelt. Vi vet hur enormt stort antalet lagstiftningsåtgärder är, och att införliva dem i den nationella och regionala lagstiftningen är ofta oerhört tidskrävande.
Att möjliggöra en förenkling av det byråkratiska språket och en allmännare tillämpning av konsekvensbedömningar är mycket viktigt, eftersom detta skulle garantera att så lite tid som möjligt tas i anspråk för klagomålsförfaranden.
Tack så mycket.
(PL) Herr talman! De enskilda medlemsstaternas genomförande av gemenskapsrätten är en av Europeiska unionens grundläggande principer.
Därför är övervakning och undanröjande av avvikelser målet för ett antal åtgärder.
Att kontrollera enskilda medlemsstater och offentliggöra resultatet av dessa kontroller skulle ge medborgarna en möjlighet att känna sig delaktiga i införlivandet av EU-lagstiftningen i medlemsstaterna.
Samtidigt förhåller det sig emellertid så att till exempel Polen fortfarande lägger på nationell mervärdesskatt, moms, trots det sjätte direktivet och domstolsutslag.
Detsamma gäller dubbelbeskattning på inkomst av tjänst.
Det finns kända fall där tullavgifter har tillämpats för fordon som köpts av polska medborgare i EU-länder, trots utslag från EG-domstolen, och förseningar av återbetalningar av felaktigt beräknade avgifter.
Särskilt underligt är det att våra medborgare kan sitta häktade i åratal utan att någon dom avkunnas.
Polens medborgare väntar otåligt på kommissionens reaktion på de exempel som jag har nämnt och att den sätter stopp för de olagliga åtgärder som begås av vår regering.
Avslutningsvis vill jag uppriktigt gratulera Monica Frassoni. Det är bara synd att detta betänkande rör en relativt avlägsen dåtid; det skulle ha varit trevligare om det hade handlat om 2007.
(DA) Herr talman! Kommittéförfarandet är en studie i hur man begränsar demokratin utan att väljarna inser det.
För det första överförs makt från väljarna och de folkvalda företrädarna till regeringstjänstemän och lobbyister bakom stängda dörrar i Bryssel.
Omröstningen underställs därefter komplicerade regler som ingen kan komma ihåg, ingen journalist kan skriva om och ingen läroboksförfattare kan förklara.
Själva kontentan av detta är helt enkelt att de icke-valda företrädarna i kommissionen kommer att besluta om inte en kvalificerad majoritet kan uppbådas mot kommissionen.
Det är lagstiftande makt som förvandlas till verkställande makt, det är öppen lagstiftning som förvandlas till hemliga dekret, det är en majoritetsdemokrati som förvandlas till en minoritetsregering.
Det är inte en absolut autokrati, men det är på väg i den riktningen med ett stänk av Mussolinis korporativa idéer.
I och med det nya interinstitutionella avtalet kan parlamentet föra tillbaka frågan på dagordningen igen, men bara om parlamentets vänster- och högerpartier är eniga och en absolut majoritet av ledamöterna röstar för detta.
Slopa blandningen av autokrati, och styr med skarpsinne och korporatism!
Inför demokrati i all lagstiftning!
Låt det bli en grundläggande princip att en majoritet av de folkvalda företrädarna står bakom varje lag, vare sig det handlar om de nationella parlamenten eller här i Europaparlamentet!
Lagstiftande av regeringstjänstemän och lobbyister borde höra till det förflutna, och ändå förankras det fast i Lissabonfördraget.
Detta är ännu ett gott skäl till att göra fördraget avhängigt av en folkomröstning.
rådets ordförande. - (SL) Jag vill i en avslutande kommentar betona på ordförandeskapets vägnar att det är medvetet om att en effektiv övervakning av gemenskapsrätten är centralt om lagstiftningen ska respekteras allmänt och om de allmänna rättsliga principer som gemenskapens fungerande grundas på ska tryggas.
I första hand är det emellertid viktigt att garantera rättslig säkerhet för EU-medborgarna.
Vi får inte glömma bort att de spelar en viktig roll i genomförandet av gemenskapsrätten.
Denna roll avspeglas även av det antal klagomål som medborgarna inger om överträdelser av EG-rätten.
Under debatten, som jag följde mycket uppmärksamt, var flera personer förvånade över att antalet överträdelser, eller åtminstone rapporterade överträdelser, inte har ökat sedan EU:s utvidgning.
Flera talare misstänkte att kommissionen inte är lika hård mot de så kallade nya medlemsstaterna.
Jag måste betona att ordförandeskapet inte har någon anledning att tro att det är på det sättet eller har några bevis som underbygger dessa tvivel.
Jag kan emellertid komma med minst en möjlig förklaring.
När det gäller de så kallade nya medlemsstaterna måste man ta hänsyn till att de blev medlemmar efter många års intensivt införlivande av gemenskapsrätten i sina rättsliga system, och sedan dess har de haft lättare att fortsätta processen i mindre skala.
Detta är bara en kommentar om misstanken att kommissionen inte behandlar alla medlemsstater lika strängt, men jag anser att det är lämpligast om kommissionsledamoten kommenterar denna fråga.
Jag vill betona att ordförandeskapet fäster stor vikt vid de gemensamma ansvarsuppgifter och målsättningar som fastställs i det interinstitutionella avtalet om bättre lagstiftning.
Slutligen vill jag uppmana alla institutioner och medlemsstater att uppfylla sina skyldigheter inom ramen för införlivandet och tillämpningen av gemenskapsrätten.
Jag har redan sagt att dagens debatt inte får bli utan konsekvenser, och jag vill betona det igen. Jag kommer att informera Franz Josef Jung om innehållet i denna debatt och parlamentets bidrag och även förslag, eftersom flera mycket viktiga förslag har framförts under debatten, som kommissionen måste ta på allvar.
Jag vill göra ytterligare en kommentar som bygger på rättsfilosofin: en gemenskap av nationer som styrs av rättstatsprincipen bygger på förtroende.
Den kan endast fungera om de deltagande staterna kan lita på varandra.
Det är skälet till att rättsliga förfaranden måste genomföras offentligt i en konstitutionell stat, och det är också skälet till att jag fullständigt instämmer i det som Diana Wallis sa.
Information är centralt i det här sammanhanget, och öppenhet är absolut nödvändigt.
Det får inte finnas några hemligheter i tillämpningen och tolkningen av lagen.
Allt måste vara öppet och offentligt.
Det är vad jag tar med mig från den här debatten, och det har jag alltid varit övertygad om personligen.
Jag håller med om det som Diana Wallis sa om den roll som utskottet för framställningar spelar.
Som hennes kund, så att säga, erkänner jag gärna att det ibland krävs en hel del arbete och ansträngningar, men medborgarna har rätt att förvänta sig att vi gör denna insats.
Genom de framställningar som vi mottar lär vi oss dessutom mycket om hur våra medborgare uppfattar vår lagstiftning och politik.
Fru Frassoni! Kommissionsledamot Margot Wallström har redan lovat att vi i framtiden kommer att införa systemet med sammanfattningar för medborgare.
Sedan dess har kommissionen även antagit ett formellt beslut om detta, så det kommer att ske, och jag är övertygad om att ni kommer att försäkra er om att vi genomför detta.
Det har beslutats, och det kommer att genomföras.
Många ledamöter har funderat över frågan om de nya medlemsstaterna och hur det kan vara så att antalet rättegångar om överträdelser av fördragen inte har ökat trots det ökade antalet medlemsstater.
Kommissionen har en mycket klar åsikt om detta, nämligen att det finns två skäl. För det första - och i det här sammanhanget känner jag mig tämligen självmedveten, eftersom jag måste påpeka att det beror på det goda arbete som den tidigare kommissionsledamoten med ansvar för utvidgningen har gjort - beror det på att de nya medlemsstaterna förberedde sitt regelverk så noggrant att de vid tidpunkten för anslutningen uppfyllde kraven mer exakt än de gamla medlemsstaterna.
Jag kan bara bekräfta detta.
Det är helt sant.
Vi skulle aldrig ha kunnat slutföra anslutningsfördragen om inte gemenskapens regelverk hade uppfyllts.
Det andra skälet är kanske lite mer praktiskt. Medborgarna i de nya medlemsstaterna måste successivt lära sig att de kan inge klagomål, och hur de gör detta.
Jag förutsätter därför att antalet klagomål kommer att öka.
Alyn Smith nämnde att lagstiftningen även måste vara lättfattlig och tillämpbar, särskilt miljölagstiftningen.
Som vi vet genomför kommissionen en översyn av all gemenskapslagstiftning som kommer att vara klar i slutet av nästa år för att ta reda på var och hur den kan förenklas.
För bara några dagar sedan lovade vi i samband med vår presentation av framstegen med projektet ”Bättre lagstiftning” att hela denna process verkligen kommer att slutföras i slutet av nästa år.
Herr Medina! Ni behöver inte oroa er för att kommissionen sopar klagomål under mattan.
Utifrån min egen erfarenhet av över åtta år som kommissionsledamot kan jag försäkra er om att jag har blivit tvungen att bromsa övernitiska kommissionsavdelningar mycket oftare än jag har behövt säga till dem att elda på med det tunga artilleriet och inleda ett fördragsöverträdelseförfarande.
Jag måste mycket oftare säga till dem, ”vänta lite, ta det lugnt och tala med dem först för att se om detta kan göras upp i godo”.
Risken för att kommissionens tjänsteavdelningar tenderar att sopa saker under matten är nästan obefintlig.
Jag är övertygad om att detta inte sker.
När det gäller Reinhard Racks fråga: beslut om överträdelser av fördraget, vare sig det är inledningen eller avslutningen eller något enskilt steg däremellan, kräver ett formellt beslut av kommissionskollegiet.
Det är så det är organiserat.
Jag kan inte här och nu besvara er specifika fråga om korssubventioner, men jag kommer att försäkra mig om att ni får ett svar före slutet av veckan.
Angående Wiesław Stefan Kucs yttranden om häktningstider före rättegång medger jag att det skulle vara en skandal om det förekom, men det faller inte inom EU:s behörighetsområde.
Europeiska domstolen för de mänskliga rättigheterna är behörig domstol för sådana ärenden.
Jag tackar för alla era förslag och den konstruktiva andan i debatten.
Jag är övertygad om att vi kommer att ha gjort ytterligare framsteg när vi diskuterar dessa frågor igen nästa år.
Herr talman, mina damer och herrar! Jag vill tacka mina ledamotskolleger, kommissionsledamoten och ordförandeskapet för att ha deltagit i denna diskussion som, vilket kommissionsledamot Günter Verheugen påpekade, inte slutar här.
Jag vill bara helt kort nämna ett par punkter.
Jag vill kommentera frågan om att fastställa prioriteringar, som kommissionsledamot Günter Verheugen talade om.
Jag anser att detta faktiskt skulle kunna vara riskabelt. Det har emellertid aldrig gjorts hittills.
Jag har alltid varit relativt skeptisk till möjligheten att verkligen fastställa prioriteringar.
Hur som helst, om ni verkligen vill gå den vägen, ta risken att vara öppna, varför inte till och med ta upp dessa prioriteringar till diskussion?
Annars skulle en misstanke kunna slå rot om att prioriteringarna har valts för att ni vill bli kvitt besvärliga överträdelser.
Det skulle inte vara bra enligt min mening.
Det andra jag vill påpeka är att trots att kommissionen förnekar att den behöver mer resurser, särskilt mänskliga resurser, för att behandla överträdelserna är det i själva verket så att jag, under nästan alla möten som jag har haft med era kolleger i kommissionen, har fått höra att de inte har tillräckligt med resurser, inte har tillräckligt med personal, för att hantera denna fråga.
Under debatten kom frågan om antalet överträdelser i de nya medlemsstaterna upp, och det som kommissionsledamoten och ordförandeskapet sa är förmodligen sant.
Vi bör emellertid också veta att det, till exempel för miljöfrågor, endast finns två, eller kanske tre tjänstemän som har hand om alla de nya medlemsstaterna, så det finns uppenbarligen ett problem med personalbrist.
Avslutningsvis har vi frågan om parlamentets roll.
Vi diskuterar internt flera olika sätt för att göra vår roll som medlagstiftare effektivare, genom att följa upp tillämpningen av de direktiv som vi antar.
Jag anser att det finns två saker som vi absolut måste göra: för det första måste vi absolut, genom ett politiskt beslut, förstärka utskottet för framställningars roll som, vilket Diana Wallis påpekade, är vårt fönster mot världen, och för det andra måste vi systematiskt hålla sammanträden om tillämpningen, vilket emellertid kräver öppet samarbete från kommissionens sida.
Om vi håller sammanträden där vi diskuterar tillämpningen av direktiv och den kommissionstjänsteman som deltar håller tyst eller berättar saker för oss som är av föga intresse - kanske för att han eller hon inte kan berätta det vi verkligen vill veta - är allt detta meningslöst.
Tack så mycket ändå, och vi kommer otvivelaktigt att återkomma till detta igen.
Debatten är härmed avslutad.
Omröstningen kommer att äga rum i morgon kl. 12.00.
Ändringsbudget nr 1/2008 - Solidaritetsfonden - Utnyttjande av EU:s solidaritetsfond (debatt)
Nästa punkt är den gemensamma debatten om
betänkandet av Kyösti Virrankoski, för budgetutskottet om förslaget till Europeiska unionens ändringsbudget nr 1/2008 för budgetåret 2008, Avsnitt III - kommissionen, och
betänkandet av Reimer Böge för budgetutskottet om förslaget till Europaparlamentets och rådets beslut om utnyttjande av EU:s solidaritetsfond i enlighet med punkt 26 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning - C6-0036/2008 -.
föredragande. - (FI) Fru talman! Europeiska unionens solidaritetsfond inrättades 2002 till följd av de katastrofala översvämningarna som drabbade Centraleuropa och som påverkade både EU:s medlemsstater och kandidatländerna.
Man kom då överens om att fonden skulle uppgå till 1 miljard euro om året.
Tanken med fonden var att den skulle underlätta för dem som hade lidit skada på grund av stora katastrofer.
Omfattningen av katastrofskadan måste vara minst 3 miljarder euro eller minst 0,6 procent av medlemsstatens BNP.
Om skadan är begränsad till ett litet område kan omfattningen vara mindre, men regionalt kan den vara relativt större.
Den skada som nu diskuteras uppkom på grund av stora översvämningar i Storbritannien i juni och juli 2007.
Skadans omfattning har uppskattats till 4,6 miljarder euro, så den är alltså berättigad till ersättning.
Kommissionen föreslår 162 miljoner euro.
Budgetutskottet rekommenderar i sin budget stöd till finansiering på det sätt som kommissionen föreslår.
Utskottet kräver dock att parlamentet godkänner utnyttjandet av stödet.
Av det skälet måste Reimer Böges betänkande om utnyttjande av EU:s solidaritetsfond antas först.
I andra hänseenden gäller den första ändringsbudgeten huvudsakligen organ och förvaltningen av Galileoprogrammet.
I budgeten har ett genomförandeorgan för Europeiska forskningsrådet inrättats.
Det har upprättats i enlighet med det budgetförfarande som har överenskommits för detta år.
I enlighet med ändringsbudgeten inrättas också ett gemensamt genomförandeorgan, genomförandeorganet för forskning (REA) för de andra programmen inom sjunde ramprogrammet för forskning.
Detta ligger också i linje med det tidigare budgetförfarandet.
De ändringsförslag om tidsplanen för anställning vid gränskontrollbyrån, Frontex, som parlamentet hade lagt fram har genomförts.
Parlamentet ökade medlen till denna byrå med 30 miljoner euro under budgetförfarandet och dessa utgör nu de nödvändiga extra medlen.
Det svåraste problemet är satellitnavigeringsprogrammet Galileo.
Parlamentets stora framgång var att det i budgetförhandlingarna lyckades garantera finansiering av programmet genom att öka det belopp som anslås till det med 2,4 miljarder euro under sex år.
Detta möjliggjordes delvis genom en ändring av den fleråriga budgetramen.
Projektet blev alltså helt klart ett EU-projekt.
Nu gäller det att administrera projektet.
Kommissionen föreslår 2 miljoner euro i form av en överföring från driftsanslag till administration.
Administrationen av projektet är dock i en rörig situation.
Projektet har i EU huvudsakligen letts av tillsynsmyndigheten för Galileo (GSA).
Dess uppgift har huvudsakligen varit diskussioner om tillstånd och partnerskap mellan den offentliga och den privata sektorn.
Den privata sektorn var inte delaktig i den inledande fasen, och GSA:s roll är därför oklar, vilket också gäller kommissionens och Europeiska rymdorganisationens (ESA) roll.
Tanken var först att ESA skulle ha ansvaret för genomförandet av projektets tekniska del, som EU skulle övervaka och utrusta.
Arbetsfördelningen mellan de olika aktörerna, såsom kommissionen och särskilda organ, är dock otydlig.
I betänkandet av Etelka Barsi-Pataky föreslår därför utskottet för industrifrågor, forskning och energi att GSA ska avskaffas.
Mot bakgrund av dessa omständigheter kan inte budgetutskottet samtycka till överföring av anslaget till kommissionen, utan föreslår i stället helt enkelt att ett symboliskt anslag införs.
Kommissionen föreslog att den skulle genomföra överföringen inom ramen för sin behörighet innan hela det administrativa systemet för Galileo hade överenskommits.
Att ändra ändringsbudgeten i detta hänseende skulle därför inte försena projektet, utan skulle garantera parlamentets förhandlingsposition.
Jag hoppas att kammaren kan ställa sig bakom utskottets enhälliga ståndpunkt rörande den första ändringsbudgeten.
föredragande. - (DE) Fru talman, herr kommissionsledamot, mina damer och herrar! Föredraganden för 2008 års budget, Kyösti Virrankoski, har verkligen täckt alla viktiga punkter.
Vi talar därför idag om grunden till ett förslag från kommissionen om utnyttjande av EU:s solidaritetsfond i enlighet med punkt 26 i det interinstitutionella avtalet.
Det stämmer att solidaritetsfonden och andra särskilda instrument inte omfattar stora penningsummor jämfört med Europeiska unionens allmänna budget.
De är en utväg för att hjälpa drabbade regioner och befolkningen där i händelse av naturkatastrofer, och som vi alla vet har sådana katastrofer, alltifrån stormar till skogsbränder, blivit ganska vanliga företeelser.
Innan vi fattade beslut tog vi i budgetutskottet initiativ till att hålla en utfrågning till vilken vi bjöd in företrädare för de drabbade regionerna i Storbritannien, lokala organisationer och också företrädare för de statliga myndigheterna.
Vid utfrågningen blev vi mycket tydligt påminda om de utmaningar som de drabbade människorna och regionerna ställs inför och omfattningen av de skador som översvämningarna i juni och juli 2007 orsakade, vilka uppskattades till totalt 4,6 miljarder euro.
Med utgångspunkt från denna utfrågning och våra samtal stödde vi till fullo kommissionens förslag om att 162 387 000 euro skulle ställas till förfogande från solidaritetsfonden i detta särskilda fall.
Låt mig också säga att vi kan förvänta oss ytterligare utnyttjande av solidaritetsfonden under de kommande månaderna.
I sådana fall är det förvisso inte endast Europeiska gemenskapen som uppmanas visa solidaritet. Mot bakgrund av att sådana katastrofer inträffar allt oftare bör medlemsstaterna tänka mer på förebyggande krishantering, dvs. att utvärdera sina civilförsvarssystem, kontrollera hur de lokala brandstationerna är utrustade och undersöka hur de eventuellt kan utveckla olika strategier i framtiden när det t.ex. gäller byggnadsarbeten i områden som riskerar att bli översvämmade.
Sådana åtgärder bör vara en integrerad del av alla långsiktiga strategier om vi vill behålla vår trovärdighet.
Ytterligare ett krav - och vi ligger något bättre till i detta avseende än i andra - är att vi bör göra det till vårt gemensamma mål, en principfråga, att se till att behandling av framtida ärenden till solidaritetsfonden ska avslutas inom maximalt sex månader.
Det är en utmaning för alla. De nationella myndigheterna måste lämna in alla ansökningar och handlingar som krävs inom den föreskrivna tiden, kommissionen måste handlägga det aktuella ärendet på grundval av tillämpliga bestämmelser, och vi i parlamentet måste också behandla ärenden genom snabba överläggningar.
Låt mig slutligen ta upp en punkt som rör ändringsbudgeten.
Med tanke på de svåra förhandlingarna och det pågående slutförandet av lagstiftningsförfarandet om satellitnavigeringssystemet Galileo stöder jag kraftfullt föredragandens villkor att den budgetpost som inrättats för administrativa utgifter bör vara ett symboliskt anslag.
Det är ett steg i rätt riktning om lämpliga administrativa strukturer upprättas inom kommissionen.
Vi är dock inte nöjda med arrangemangen för det framtida samarbetet mellan kommissionen, Europeiska rymdorganisationen och tillsynsmyndigheten för Galileo (GSA).
Under lagstiftningsförfarandet måste det åtminstone fastställas hur man kan undvika dubbelarbete och det bör utvecklas lämpliga administrativa strukturer mot bakgrund av de nya villkoren för satellitnavigeringssystemet Galileo.
Det finns fortfarande ett visst behov av diskussion, vilket jag hoppas att vi kan tillmötesgå så snart som möjligt.
kommissionsledamot. - (EN) Herr talman! Den 18 januari antog kommissionen ett förslag till utnyttjande av solidaritetsfonden för Storbritannien, och vi är nöjda och glada över att budgetutskottet ställer sig positivt till vårt förslag.
Förutom den första ändringsbudgeten för 2008 års budget förslog vi också ett anslag på 162 miljoner euro från solidaritetsfonden till Storbritannien som ersättning för de allvarliga skador som sommarens översvämningar förorsakade.
Som budgetutskottets ordförande redan har sagt har vi nyligen mottagit förfrågningar från två medlemsstater - Grekland och Slovenien - och vi kommer troligen att lägga fram ett nytt förslag mycket snart.
Detta förslag gäller naturligtvis inte endast solidaritetsfonden.
Det är endast solidaritetsfonden som kommer att beröras finansiellt. Andra delar i förslaget är mer tekniska.
Frågan om Galileo är naturligtvis mycket känslig för oss alla och jag förstår till fullo budgetutskottets oro.
Jag måste dock säga att budgetutskottets förslag om att ändra kommissionens förslag kommer att försena medel från solidaritetsfonden med omkring en månad, eftersom frågan måste gå tillbaka till rådet för ytterligare en omröstning, men vi förstår att det är känsligt och vi kan inte motsätta oss budgetutskottets beslut i denna fråga.
Jag hoppas dock verkligen att vårt förslag kommer att stödjas generellt i parlamentet denna vecka.
för PPE-DE-gruppen.- (EN) Herr talman! Jag vill säga att jag stöder ändringsbudgeten, och det är ett par poster som jag vill kommentera.
För det första gäller det solidaritetsfonden. Det var naturligtvis ett anslag med anledning av översvämningarna i Storbritannien i juni och juli förra året.
En stor del av översvämningarna inträffade i min region, och jag kan intyga att många invånare i min region drabbades av förfärliga skador och fick utstå umbäranden.
Det var intressant att notera - men jag är inte förvånad - att detta var det tredje största kravet i historien till solidaritetsfonden.
Kravet uppgick till 4,6 miljarder euro och anslaget motsvarade 162,8 miljoner euro.
Jag är medveten om att min vän och kollega Reimer Böge helt i sin ordning har sagt att detta inte är någon stor summa pengar.
Det kanske det inte är, men som en solidaritetsgest är det mycket uppskattat, tro mig, och jag vill på folkets vägnar i min region rikta ett stort tack främst till ledamöterna i budgetutskottet som enhälligt stödde biståndspaketet - vilket verkligen är en solidaritetsgest.
Men jag vill också visa min uppskattning för kommissionsledamoten och hennes kolleger som handlade detta krav på sju månader.
Jag tyckte att det var en stor insats, fru kommissionsledamot, och jag tackar er för de insatser ni har gjort för att genomföra detta.
Jag kommer naturligtvis att med stort intresse de närmaste veckorna och månaderna följa hur den brittiska regeringen fördelar medlen, men för mig är det helt klart att dessa frågor kommer att väckas alltmer regelbundet i Europeiska unionen med tanke på att det allt oftare framkommer bevis på extrema händelser till följd av klimatförändringar.
Det är också tydligt att det, när det gäller uttryck för solidaritet, faktiskt är hur snabbt svaret kommer som är den viktigaste delen i mekanismen.
Beträffande frågan om Frontex vill jag också säga att jag stöder tilläggsanslaget till Frontex - vi fördubblade anslaget till byrån.
Jag tyckte att det var helt rätt och jag konstaterar att man begär att 25 poster ska inrättas.
Jag anser dock att det är viktigt att vi fortsätter att övervaka fördelningen av medlen för att se till att de ger valuta för pengarna.
På samma sätt stödde jag kraftfullt de Lissabonmål som kommissionen hade upprättat för sig själv, särskilt på området för forskning och utveckling.
Jag erkänner därför behovet av genomförandeorganen för forskning, men jag vill omigen uttrycka min oro för den stora mängden organ som, det måste jag säga, historiskt sett inte har haft rykte om sig att ge valuta för pengarna.
När det slutligen gäller Galileo, kommer den nya budgetposten att göra en hel del för att öka insynen och ansvarsskyldigheten.
Jag är dock överens med mina kolleger i budgetutskottet när vi säger att vi ska gå försiktigt tillväga.
Det är, om jag får säga så, fru kommissionsledamot, ett stort åtagande och - jag lånar lite jargong från rymdåldern -kommissionen är ”djärvt nog på väg dit där ingen kommission tidigare har varit”.
Jag håller därför med min kollega Reimer Böge när han säger att vi stöder detta, men att vi insisterar på att det symboliska anslaget ska införas.
Herr talman! Jag stöder ändringsbudgeten och är glad över att göra det.
för PSE-gruppen. - (EN) Herr talman! Jag ersätter Gary Titley, ledaren för parlamentets socialdemokratiska ledamöter, ikväll, men jag kan tala på alla de socialdemokratiska ledamöternas vägnar och välkomnar ändringsbudgeten och beslutet att bevilja 162 miljoner euro till de regioner i Storbritannien som har drabbats av översvämningar.
Som Richard James Ashworth sa är det ett litet bidrag för att täcka de enorma kostnaderna för de skador som översvämningarna i Storbritannien har orsakat, men vi är tacksamma mot våra kolleger i budgetutskottet, som röstade enhälligt för detta, och också mot kommissionen.
Jag förstår att det var den snabbaste utbetalning som någonsin gjorts; inom sju månader.
Det är därför ett framsteg jämfört med tidigare anslag, även om många människor har fått lida länge.
Vi förstår också att det är en av de största utbetalningar som någonsin gjorts, och vi är tacksamma för det.
Förra veckans översvämningar drabbade 48 000 brittiska hushåll och 700 företag, och de totala skadorna uppskattas till över 4 miljarder euro.
Min egen region Yorkshire var en av de värst drabbade.
Många människor har ännu inte återvänt till sina hem, och därför uppskattas denna hjälp och detta bistånd väldigt mycket.
Jag ersätter Gary Titley, eftersom han har fastnat i London på grund av de mycket allvarliga stormar som har dragit in över Västeuropa ikväll.
Vi kan inte skylla allt dåligt väder på klimatförändringarna, men vi vet faktiskt att antalet extrema väderhändelser ökar.
Vi har sett allvarliga översvämningar, och också bränderna i Grekland och Sydeuropa förra sommaren.
Inga belopp från solidaritetsfonder kan egentligen täcka de skador och de kostnader som vi ser är resultatet av dessa händelser som inträffat på grund av klimatförändringarna.
Vi börjar vårt arbete som parlamentsledamöter om det nya lagstiftningspaketet till följd av klimatförändringarna.
Jag hoppas verkligen att parlamentet kommer att inta en hård hållning och genomföra och enas om en bra lagstiftning som verkligen hanterar klimatförändringarna, så att vi inte behöver komma tillbaks hit och be kommissionen om pengar för att hantera dessa typer av händelser.
för ALDE-gruppen. - (EN) Herr talman! På sätt och vis har jag en lätt uppgift efter de två sista talarna.
Jag vill också tydligt uttala mig för förslaget från våra föredragande Kyösti Virrankoski och Reimer Böge, men i synnerhet vill jag uttala mig för utnyttjandet av solidaritetsfonden till Storbritannien.
En summa på 162 miljoner euro kan tyckas vara okontroversiell men den är oerhört viktig på flera nivåer.
Som parlamentsledamot representerar jag Yorkshire- och Humberområdena som, vilket Linda McAvan sa, drabbats av översvämningar förra sommaren.
Städer och byar i vår region ödelades.
Många människor, till och med i byn i närheten av mig, har fortfarande inte kunnat återvända till sina hem.
Samtidigt som vi vet att utbetalningen kanske inte ändrar dessa regioners situation på en dag kommer den indirekt att lätta trycket på vår regerings egen budget.
För det andra är jag mycket nöjd över att vår regering gjorde denna ansökan som dessutom var framgångsrik.
I början var vi inte alltid säkra på vad som skulle hända, och jag hoppas att vår regering efter denna erfarenhet kommer att bli en stor anhängare till solidaritetsfonden i rådet och att den kommer att övertala andra medlemsstater att göra likadant.
För det sista kommer det brittiska folket, mina väljare, nu att förstå att europeisk solidaritet har en konkret och praktisk betydelse.
Jag tror att det kommer att gälla oss alla i parlamentet.
Eftersom klimatförändringarna går ut över oss kan vi alla komma att representera offren för sådana naturkatastrofer och således kanske tvingas be om europeisk solidaritet.
för UEN-gruppen. - (PL) Herr talman! Solidaritet är EU:s viktigaste och ädlaste princip.
Utan den kan det inte komma på fråga att oberoende stater och nationer handlar gemensamt.
Inrättandet av EU:s solidaritetsfond följde naturligt med denna princip.
I nuläget har vi en summa på en miljard euro tillgänglig varje år.
Det är ingen stor summa, i synnerhet inte förra året och innevarande år, när vi tvingades bevittna en ökning av klimatkatastroferna.
Vi har inte enbart drabbats av översvämningar och stormar utan också av oväntat stora bränder.
Med våra begränsade medel har vi än så länge bara möjlighet att bistå med småskalig hjälp - 3-4 procent av skadorna, eller till och med ännu mindre.
Därför drar jag slutsatsen, samtidigt som jag stöder Reimer Böges betänkande och Kyösti Virrankoskis förslag till ändringsbudget, att solidaritetsfondens resurser gradvis måste ökas.
Två euro per invånare kommer inte att vara tillräcklig hjälp vid enorma förluster.
för IND/DEM-gruppen. - (EN) Herr talman! Det gläder mig att höra att vi i Storbritannien borde få ett ekonomiskt bidrag till kostnaderna efter förra årets översvämningar.
Vi är alla mycket glada över att EU generöst har gett stöd till en medlemsstat som befinner sig i svårigheter. Det är dock inte riktigt så.
För det första täcker bidraget enbart 3.5 procent av skadekostnaderna - en gest som Richard Ashworth säger.
För det andra har det gått nio månader sedan översvämningen inträffade - och det säger man är snabbt!
Det skulle ha varit till större hjälp om vi hade vetat att stödet var förestående.
Då kunde återuppbyggnaden ha planerats därefter.
Om det är något som irriterar oss britter - när vi inser att vi får tillbaka en liten del av de pengar vi har betalat in till EU - så är det att vi är tvungna att be att få pengarna och sedan göra reklam för EU:s generositet.
Snälla, kan vi inte hellre få behålla våra egna pengar och därefter själva bestämma hur vi ska använda dem?
Då skulle de kunna betalas ut snabbare.
(FR) Herr talman! De flesta av våra stater har kreditposter i sin budgetlagstiftning för att kunna ta itu med katastrofer.
I den franska budgetlagstiftningen, till exempel, finns det generella anslag som innebär möjlighet att ge anslag genom dekret i förväg i nödsituationer.
Sedan november 2002 har vi i EU:s budgetlagstiftning införlivat en rätt till finansiering vid katastrofer i solidaritetsfonden.
Vi har också inrättat Europeiska fonden för justering för globaliseringseffekter för att finansiera katastrofer.
När det gäller naturkatastrofer har vi ombetts att ge stöd med mindre än 4 procent för att reparera skadorna efter översvämningen i Storbritannien, skador som kostar mer än 4 miljarder.
Nio månader för att göra anslagsåtaganden är en lång tid, eftersom det per definition handlar om en nödsituation.
Det betyder att sättet anslagsåtaganden antas på i ändringsbudgeten inte är funktionsdugligt.
Ändringsbudgeten borde träda i kraft tidigare så att man kan fastställa att anslagsåtaganden ska göras i förväg genom preliminära och icke-begränsade anslagsåtaganden för katastrofer, översvämningar och bränder.
Mot denna bakgrund är 162 miljoner euro i solidaritet en utmärkt lektion i pragmatik för Storbritanniens medborgare Adam Smith, Ricardo och Margaret Thatcher som bara tror på marknaden, darwinismen och det naturliga urvalet.
När lejonet som ryter i den ekonomiska djungeln drabbas av problem upptäcker han fördelarna med solidaritet.
Det har hänt tre gånger nu - galna kosjukan, mul- och klövsjukan samt översvämningarna - och i morgon kommer de brittiska medlemmarna också att ha chansen att visa solidaritet med de europeiska bönderna som har översvämmats av importer.
- (EL) Herr talman! Ändringsbudgeten visar än en gång det som är självklart: att EU har de mekanismer och den anpassningsförmåga som krävs för att lösa specifika oväntade problem.
Jag skulle vilja ge tre förslag om de två betänkanden vi har diskuterat idag.
Två av dem rör solidaritetsfonden och det tredje gäller Galileoprogrammet.
När det gäller översvämningarna i Storbritannien är tidsintervallet mellan juli och de nuvarande insatserna mycket tillfredsställande.
Det råkar vara den snabbaste insatsen under den tid fonden har tillämpats, åtminstone vad jag kan minnas.
Likväl skapar det ett prejudikat.
I framtiden ska vi förvänta oss sådana omedelbara insatser vid liknande katastrofer, och här syftar jag på miljökatastrofen som vi i Grekland drabbades av förra sommaren bara en månad senare, i augusti.
Jag hoppas därför att kommissionen nästa månad, genom den ansvariga kommissionsledamoten, åtminstone kommer att ge ett förslag om den grekiska begäran att ta solidaritetsfonden i bruk.
Jag behöver inte påminna er om de chockerande bilderna från den stora brandkatastrofen i Grekland.
Vi såg dem alla, överallt i Europa.
Jag hoppas att vi, med vederbörliga ändringar, åtminstone kommer att ha kommissionens förslag i våra händer nästa månad.
Min andra kommentar gäller det åtlöje vi nu gör oss själva till.
Jag har ingen aning om hur parlamentet lyckas med det, men varenda gång vi har goda nyheter är vi de enda som vet det!
Vi är för oss själva och det finns antagligen inte ens en journalist på läktaren!
När ska vi äntligen lära oss att marknadsföra de goda nyheterna på rätt sätt?
Min tredje och sista kommentar gäller Galileoprogrammet.
Jag håller med alla mina kolleger från budgetutskottet, och i egenskap av utskottets föredragande för programmet skulle jag vilja vara tydlig med att vi inte kommer att göra någon utbetalning från det oerhört ansenliga paketet med fonder som vi har inrättat om vi inte kommer överens med rådet om programmets utformning i stort.
Om vi inte vet vem som gör vad - och vi befinner oss fortfarande i oklarhet eftersom vi förhandlar med rådet - ska vi inte göra någon utbetalning.
Vi kommer inte att kasta pengar i sjön.
I morgon bitti har vi en oerhört viktig trepartsdiskussion med det slovenska ordförandeskapet.
Det finns två viktiga centrala frågor.
Jag hoppas att vi kan avsluta förhandlingarna så att vi kan rikta in oss på att göra verkliga framsteg.
- (LT) EU:s solidaritetsfond är ett mycket viktigt stöd till medlemsstater och potentiella kandidatländer vid naturkatastrofer.
Likväl är det, i ljuset av erfarenheterna, uppenbart att solidaritetsfonden måste reformeras och anpassas för att möta nya utmaningar. Man måste även göra den mer effektiv.
För det första är minimitröskeln för skador på 3 miljarder euro eller 0.6 procent av BNP för hög och den utesluter all hjälp till länder som drabbats av katastrofer i mindre skala men som likväl kan få allvarliga konsekvenser för de berörda länderna.
För det andra kan inte medel från fonden betalas ut för att mildra konsekvenserna av terrorism, allmänna hälsokriser och tekniska eller industriella olyckor.
För det tredje uppstår det problem när det gäller medel som kan betalas ut i händelse av uteslutande regionala olyckor.
För dessa är inte användningskriterierna tillräckligt tydligt definierade.
Sammanfattningsvis välkomnar jag reformen av fonden och jag uppmanar rådet att ge en sammanfattning av sin ståndpunkt utan dröjsmål.
(PL) Herr talman! Jag skulle vilja rikta uppmärksamheten mot följande punkter i debatten.
För det första är det beklagligt att kommissionens förslag till Europaparlamentets och rådets förordning om inrättande av Europeiska unionens solidaritetsfond fortfarande inte har antagits av rådet, trots att Europaparlamentet tog ställning i frågan vid första behandlingen för nästan två år sedan, i maj 2006.
För det andra förtjänar utnyttjandet av 162 miljoner euro som en hjälp för att gottgöra de skador (som beräknas till 5 miljarder euro) som översvämningarna under juni och juli 2007 orsakade i Storbritannien och på Irland vårt stöd.
Det är synd att medlen för detta syfte anslås många månader efter att skadorna skett eftersom det kan göra stödet mindre effektivt.
Som det polska ordspråket säger: ”den som ger snabbt ger dubbelt så mycket”.
För det tredje hoppas jag att man, eftersom solidaritetsfondens tak har satts till 1 miljard euro, vid så stora skador som i Storbritannien, snabbt kommer att uppbåda skälig finansiering och att man kommer att tillgodose de nya och de gamla medlemsstaternas behov på lika villkor.
- (EL) Herr talman! Samtidigt som jag vill tacka föredraganden för det mycket goda arbete han har utfört skulle jag vilja göra ett mycket kort påpekande om solidaritetsfonden.
Vi har haft dåligt väder varje år i Europa.
Det är också ironiskt att, just när vi diskuterar dessa viktiga betänkanden, kommer Nordeuropa att drabbas av våldsamma stormar.
Det är verkligen en välsignelse att EU tillhandahåller finansiellt stöd i händelse av sådana katastrofer som i Storbritannien och att man har gjort det tidigare till Cypern.
Trots allt får vi inte glömma att det vid sidan av den finansiella aspekten måste finnas en organisatorisk enhet på gemenskapsnivå som är i stånd att ge omedelbart bistånd till de drabbade områdena.
- (EL) Herr talman, mina damer och herrar! Solidaritet är ett vackert ord och ett ännu vackrare begrepp.
Tyvärr finns det ett mycket stort behov av solidaritet. Verkligheten visar att behovet håller på att bli allt mer trängande på grund av naturkatastroferna, som vi inte längre borde se som någonting naturligt, utan snarare som allt vanligare händelser i våra liv.
Bara under sommarmånaderna 2007 inträffade tre ytterst allvarliga händelser.
Först kom översvämningarna i Storbritannien som vi diskuterar och röstar om idag.
Direkt efteråt följde de hemska bränderna i Grekland, som ni alla känner till, och kort efter detta fler översvämningar i Slovenien.
Allt detta visar oss hur allvarliga fenomenen är och även hur viktigt det är för EU att agera.
Jag blir överraskad när andra medlemmar säger att de inte förstår varför EU skulle tillhandahålla pengar.
Det är inte bara en fråga om pengar, utan också om moraliskt stöd och om en känsla bland invånarna i de drabbade områdena att EU är medvetet om deras tragedi.
I många fall är det en tragedi, och EU gör någonting åt det.
Därför vill jag påpeka, som har nämnts innan, att exemplet med Storbritannien, som vi applåderar, på grund av den relativt snabba insatsen, borde försöka efterliknas i andra drabbade länder.
Det är inte en slump att vårt land, Grekland, är nästa land på listan för bistånd från solidaritetsfonden, och vi hoppas att hjälpen kommer att vara på väg snabbt även i vårt fall.
Jag är dock inte säker på att det kommer att hända och jag undrar om det beror på EU och hur gemenskapen hanterar ansökningar eller på hur Grekland lade fram sin begäran.
Hur som helst: vi hoppas att hjälp kommer att ges snart till Grekland också, för jag försäkrar er att situationen fortfarande är mycket allvarlig hos oss.
Problemet är att de medel till Grekland som sattes in i fonden fortfarande inte har kungjorts.
EU:s solidaritetsfond ses på ett mycket positivt sätt av medlemsstaterna och framför allt av EU:s medborgare, Genom fonden finns det möjlighet att bevilja stöd till de som drabbats av naturkatastrofer som orsakat avsevärda skador.
Fondens syfte är att bidra till att gottgöra de förluster som tillfogats och som väger tungt i många familjers budget.
EU:s finansiella stöd är ett exempel på europeisk solidaritet.
För de europeiska familjer som lider, våra EU-medborgare, utgör stödet det främsta exemplet på de fördelar och förmåner ett medlemskap i Europeiska gemenskapen ger när ett sådant behov uppstår.
Likväl måste vi koncentrera oss på - och hitta de nödvändiga medlen i EU-budgeten - att bekämpa orsakerna till katastroferna och på att inrätta lämpliga arrangemang för krishantering samt lämpliga försäkringssystem.
föredragande. - (FI) Herr talman! Jag skulle vilja tacka alla som har deltagit i debatten för deras utomordentliga, konstruktiva bidrag.
Solidaritetsfonden är oerhört ung och därför har dess gränser satts väldigt högt.
Det har inte varit möjligt att lita på tidigare information om hur mycket pengar som behövs.
Gränserna kanske i viss mån kan ses över i framtiden.
Jag håller med om att snabbhet utan tvekan är en fördel i det här arbetet.
Budgetutskottet har ägnat stor uppmärksamhet åt utnyttjandet av globaliseringsfonden för att övervinna de problem som uppstår på grund av förlorade arbeten.
Det är uppenbarligen ett område som EU kommer att arbeta mycket med i framtiden.
På samma sätt har många tagit upp frågan om krishantering.
I årets budget införlivas ett pilotprojekt för att snabba på förebyggandet av skogsbränder.
Inom det området strävar vi efter nya, goda resultat.
När det gäller Galileoprojektet kommer anslagen inte att öka.
Detta måste givetvis ses som en grundläggande princip.
Den nuvarande finansieringsnivån är tillräcklig, Administrationen måste emellertid vara effektiv.
I synnerhet i nuläget, när finansieringsnivåerna är ansenliga, finns det en risk att projektets administrativa förvaltning också kommer att bli mer byråkratisk.
Den måste vara effektiv och av den anledningen vill vi behålla parlamentets utrymme för förhandling, så att vi tillsammans med kommissionen och rådet kan komma överens om vilken den bästa förvaltningsformen är för att uppnå målet med detta europeiska, mycket ambitiösa och stora projekt.
Jag är övertygad om att vi kommer att uppnå ett tillfredsställande resultat under de kommande veckorna.
Debatten är härmed avslutad.
Omröstningen kommer att äga rum tisdagen den 11 mars 2008.
Skriftliga förklaringar (Artikel 142)
skriftlig. - (RO) Jag anser att Storbritanniens begäran är motiverad och jag stöder utnyttjandet av solidaritetsfonden i det här fallet.
Rumänien har drabbats av stora översvämningar under de senaste åren och de senaste ägde rum nyss.
Liksom i fallet med Storbritannien kunde stora delar av de skador som översvämningarna orsakade ha undvikits genom större förebyggande ansträngningar.
Den befintliga infrastrukturen och de nationella myndigheternas insatser räckte dock inte till inför naturfenomenets kraft. Därför stöder jag de två åtgärder som EU kan vidta för att förstärka nationella och europeiska insatser.
Den första är tilldelning av pengar från strukturfonderna för infrastrukturarbeten som syftar till att lindra naturkatastrofernas effekter och den andra är upprättandet - så snart som möjligt - av en europeisk insatsstyrka, bestående av specialistgrupper från alla medlemsstater som ska ingripa i nödsituationer i alla regioner i EU.
En annan viktig aspekt är omfattningen av de medel som EU anslår i nödsituationer.
Med tanke på att vi planerar en omfattande översyn av EU:s budget anser jag att vi bör överväga att öka de belopp som anslås till EU:s solidaritetsfond.
Högtidligt möte - Högtidlighållande av Europaparlamentets 50-årsjubileum
(Kort framträdande av Europeiska unionens ungdomsorkester, under ledning av Pavel Kotla.)
Det var ett vackert framträdande av Europeiska unionens ungdomsorkester med Pavel Kotla som dirigent.
Tack så mycket.
Mina damer och herrar! Jag hälsar er alla varmt välkomna till kammaren för att fira femtioårsjubileet av Europeiska parlamentariska församlingens konstituerande sammanträde.
Först och främst skulle jag vilja föreslå att vi med acklamation välkomnar alla tidigare talmän som är här i dag: Emilio Colombo, Lord Henry Plumb, Enrique Barón Crespo, Egon Klepsch, Klaus Hänsch, José Maria Gil Robles, Nicole Fontaine och Josep Borrell Fontelles.
Välkomna alla högt aktade tidigare talmän för Europaparlamentet.
(Ihållande applåder)
Dessutom skulle jag varmt vilja välkomna Janez Janša, Europeiska rådets tjänstgörande ordförande, och José Manuel Durão Barroso, Europeiska kommissionens ordförande.
Kommissionsordförande Barroso! Ni är givetvis ett välbekant ansikte här i kammaren, men ni är särskilt välkommen i dag.
(Applåder)
Jag är extra glad att kunna välkomna Lluís Maria de Puig, talman i Europarådets parlamentariska församling, hit till kammaren i dag.
Ni är varmt välkommen.
(Applåder)
Det är ett nöje att kunna välkomna ordförandena och talmännen i de belgiska parlamenten, Herman van Rompuy, det italienska parlamentet, Fausto Bertinotti och den nederländska senaten, Yvonne Timmerman-Buck. De har samlats här i dag i Europaparlamentet tillsammans med andra företrädare för parlamenten i Bulgarien, Tjeckien, Estland, Frankrike, Tyskland, Ungern, Polen, Portugal, Rumänien, Slovakien, Slovenien och Storbritannien.
(Applåder)
Jag välkomnar ordförandena för de övriga EU-institutionerna: ordföranden för EG-domstolens första avdelning, Peter Jann, revisionsrättens ordförande Vítor Caldeira, Europeiska ekonomiska och sociala kommitténs ordförande Dimitris Dimitriadis, Regionkommitténs ordförande Luc Van den Brande och EU:s ombudsman Nikoforos Diamandouros.
Välkomna till Europaparlamentet.
(Applåder)
Det är ett nöje att kunna välkomna följande lokala och regionala företrädare: Strasbourgs borgmästare Fabienne Keller, ordföranden för Alsaces regionala rådsförsamling Adrien Zeller, ordföranden för Conseil Général du Bas-Rhin Philippe Richert och prefekten för regionen Alsace och Bas-Rhin Jean-Marc Rebière.
Välkomna till Europaparlamentet.
(Applåder)
På stol 146 sitter vår kollega Astrid Lulling. Hon är den enda av oss som var ledamot av Europaparlamentet innan det blev en direktvald församling.
(Ihållande applåder)
För nästan exakt 50 år sedan, den 19 mars 1958, sammanträdde den gemensamma församlingen för de tre europeiska institutionerna - Europeiska ekonomiska gemenskapen, Europeiska atomenergigemenskapen och Europeiska kol- och stålgemenskapen - för första gången här i Strasbourg i vad som då hette Maison de l'Europe.
Församlingen bestod enligt Romfördraget, som hade antagits några veckor tidigare, av ”företrädare för folken i de medlemsstater som förenas i Europeiska gemenskapen”.
I dag firar vi detta jubileum eftersom vi, i rakt nedstigande led, är direkta arvtagare till denna parlamentariska församling och dess ursprungliga 142 ledamöter.
Den förste talmannen i denna gemensamma församling var den store Robert Schuman.
I sitt installationstal sa han att församlingen skulle spela en nyckelroll för att utveckla den europeiska andan, som församlingen enligt honom ”hade varit och var en smältdegel för”.
Detta är lika sant nu som då.
Vid det konstituerande sammanträdet varnade samtidigt Robert Schuman sina kolleger för att ett parlamentsarbete med 142 ledamöter - från vid denna tidpunkt sex länder - skulle kräva disciplin från alla.
Detta är som vi alla vet givetvis än mer relevant i dag, med 785 ledamöter från 27 länder!
Inte långt efter det konstituerande sammanträdet började våra företrädare att kalla institutionen ”Europaparlamentet”. Först skedde detta informellt eftersom termen inte fanns i fördragen om upprättandet av Europeiska gemenskaperna.
Det var inte förrän fyra år senare, i mars 1962, som den parlamentariska församlingen fattade ett formellt beslut om att kalla sig för ”Europaparlamentet”.
Trots att det i fördragen om upprättandet av Europeiska gemenskaperna föreskrevs att församlingen ”ska utarbeta förslag till allmänna direkta val enligt en i alla medlemsstater enhetlig ordning” och att ” rådet ska enhälligt fastställa bestämmelserna och rekommendera medlemsstaterna att anta dessa i överensstämmelse med deras konstitutionella bestämmelser” var det inte förrän 1976 som rådet - på grundval av Europaparlamentets rekommendation av den 20 september 1976 - antog en rättsakt om att hålla direkta och allmänna val till Europaparlamentet.
Mina damer och herrar! Den parlamentariska församlingen hade inledningsvis nästan inga som helst egna befogenheter.
Våra företrädare visste att det skulle ta lång tid att utveckla den europeiska parlamentariska dimensionen och att detta skulle kräva en tydlig kompass, engagemang, tålamod och uthållighet från dem och kommande generationer.
Steg för steg har Europaparlamentet tillskansat sig mer och mer egna befogenheter och blivit allt mer medvetet om sina skyldigheter och handlingsutrymme.
Jag tror att jag talar för alla här när jag säger att i dag är parlamentet verkligen värt sitt namn.
(Applåder)
I dag företräder vi nästan 500 miljoner EU-medborgare och vi speglar hela det politiska spektrumet i EU.
Vi är EU:s fritt valda parlament, enat i vår strävan att nå de bästa och mest övertygande lösningarna.
Vi har blivit självsäkra och en central aktör i europeisk politik.
Vi har rätt att vara nöjda.
Denna process inleddes 1958 och det har funnits flera milstolpar längs vägen, på vår gemensamma färd mot europeisk integration.
Europeiska gemenskapen fick sin egen budget 1971och sedan dess har Europaparlamentet spelat en central roll vid antagandet av budgeten.
Det första direkta valet till Europaparlamentet hölls 1979.
Genom enhetsakten 1986 fick namnet Europaparlamentet äntligen rättslig status.
Genom Maastrichtfördragets ikraftträdande för 15 år sedan fick Europaparlamentet äntligen full medbeslutanderätt på vissa områden av gemenskapspolitiken, vilket gjorde det möjligt för parlamentet att verkligen bidra till utarbetandet av lagstiftning, och vid behov dra i nödbromsen, mot rådets vilja.
I Amsterdamfördraget utökades medbeslutandebefogenheterna, medan Lissabonfördraget kommer att göra medbeslutandeförfarandet till normalförfarandet när EU-lagstiftning utarbetas. Det har därför fått det passande namnet ”det ordinarie lagstiftningsförfarandet”.
I dag är vi 785 ledamöter från 27 europeiska länder.
Vi företräder fler än 150 nationella politiska partier, varav de flesta har slagit sig samman i någon av Europaparlamentets sju politiska grupper.
Vi är både en lagstiftande församling och en budgetmyndighet, jämbördig med rådet.
Vi utövar kontroll över kommissionen och utser dess ordförande. Och kommissionen kan inte tillsättas utan vårt godkännande.
Vi förespråkar gemenskapsrättens företräde och vi är EU:s folkvalda församling.
För tre veckor sedan antog vi Lissabonfördraget, som ytterligare kommer att stärka våra befogenheter.
I framtiden kommer beslut i viktiga frågor som rör EU:s medborgare endast att kunna fattas om en majoritet i Europaparlamentet ger sitt samtycke.
Detta gäller även centrala frågor på det rättsliga och inrikespolitiska området.
Vi får emellertid inte slå oss till ro och det är verkligen inte fråga om en oundviklig process.
Vi har varit att tvungna att kämpa hårt hela vägen.
Jag skulle vilja tacka alla som under de senaste fem decennierna, i våra talmäns trygga händer, har arbetat för att stärka den europeiska integrationens parlamentariska dimension och gett ett värdefullt bidrag till denna process.
Ett stort tack till både tidigare och nuvarande ledamöter av Europarlamentet!
(Applåder)
Jean Monnet sa en gång att inget är möjligt utan människor, och inget är permanent utan institutioner.
Jag skulle också vilja ta tillfället i akt för att skänka Paul-Henri Spaak en tanke, den förste talmannen i Europeiska kol och stålgemenskapens (EKSG) gemensamma församling - den institution som föregick Europaparlamentet.
Han gav med sin rapport efter Messinakonferensen i juni 1955 ett viktigt bidrag till utarbetandet av Romfördraget.
Vägen mot parlamentarisk demokrati i EU har följt en logik som vi känner igen från de europeiska ländernas historia.
Vi har skapat en institutionell balans mellan nationell nivå och EU-nivå som har varit en stor framgång och speglar samspelet mellan EU:s olika maktfördelningsnivåer.
Ett viktigt element i denna balans är Europaparlamentets goda samarbete med de nationella parlamenten, som är särskilt viktigt för oss.
Jag är mycket glad att nästan alla medlemsstaters nationella parlament har skickat företrädare på hög nivå för att närvara vid denna sammankomst.
(Applåder)
Jag skulle vilja be er alla - ledamöterna av Europaparlamentet och ledamöterna av de nationella parlamenten - att dra sitt strå till stacken i vår strävan efter att fortsätta detta samarbete i framtiden.
Lissabonfördraget och stadgan om de grundläggande rättigheterna kommer att vara avgörande för att förverkliga demokrati och parlamentarism i EU på alla nivåer.
Vi kan vara stolta över vårt konsekventa och tydliga stöd för reformfördraget och stadgan om de grundläggande rättigheterna.
(Applåder)
Vi behöver en kritisk allmänhet och kritisk granskning av vårt arbete.
Men vi har även rätt till rättvisa.
EU, i all sin mångfald, är mer komplext än någon annan gemenskap i världen.
Jag skulle vilja be medierna - som spelar en viktig roll i kommunikationen med medborgarna - att tänka på det.
EU bör inte göras till syndabock för nationella tillkortakommanden.
(Applåder)
En av de största framgångarna i vår europeiska vision under de senaste 50 åren har varit vårt försvar av demokrati och frihet i hela Europa. I dag är Estland, Lettland.
Litauen, Polen, Tjeckien, Slovakien, Ungern, Slovenien, Bulgarien, Rumänien och det återförenade Tyskland EU-medlemmar - ett resultat som vi bara hade kunnat drömma om och som har förverkligats under vår livstid.
I dag är vi medborgare i Europeiska unionen - enligt Berlinförklaringen av den 25 mars 2007 - ”nu lyckligtvis förenade”. Detta är något vi bör glädjas åt.
När vi ser tillbaka på de senaste 50 åren är det viktigt att även se framåt.
Vi bör självkritiskt påminna oss själva om vilka aspekter i EU:s parlamentariska dimension som fortfarande är otillfredsställande.
Till skillnad från de nationella parlamenten har vi fortfarande inte möjlighet att i budgetprocessen fatta beslut om våra egna finansiella resurser.
Parlamentariskt styre innebär i allmänhet parlamentarisk kontroll över militären. Men EU:s gemensamma säkerhets- och försvarspolitik är fortfarande ofullständig och ger en otillräcklig koppling mellan nationella skyldigheter och skyldigheter på EU-nivå.
Vi saknar fortfarande en enhetlig valordning, vilket innebär att vi fortfarande saknar en viktig förutsättning för effektiva europeiska politiska partier som kan ställa upp i val till Europaparlamentet med gemensamma valsedlar.
Med tålamod, uthållighet och en god kompass har Europaparlamentet ända sedan Europeiska parlamentariska församlingens första session kämpat för att försvara sin position i Europa. Och det måste och kommer det att fortsätta att göra även i framtiden.
Som EU:s direktvalda överstatliga församling visas Europaparlamentet upp som en modell för liknande ansträngningar i andra regioner i världen.
Jag har blivit vittne till detta, och det har ni också, när vi besöker andra delar av världen.
Denna positiva utveckling av Europas parlamentariska dimension hade nästan varit omöjlig att förutse när Rober Schuman installerades som den parlamentariska församlingens första talman den 19 mars 1958.
Men Robert Schuman hade en vision.
Han talade om en Europatanke som måste återuppväckas och beskrev denna som ”la relance de l'idee européenne”.
Vad skulle i dag, efter krisen i samband med misslyckandet med det konstitutionella fördraget, kunna vara ett bättre ledmotiv för den uppgift som vi har framför oss?
Den 19 mars 1958 uttryckte Robert Schuman i sitt korta tal sina farhågor för att en teknokratisk syn kunde få den europeiska integrationen att vittra sönder.
Detta gäller i lika hög grad nu som då.
Robert Schuman var realistisk, blygsam och tydlig i sin beskrivning av möjligheterna för den parlamentariska församling som han ledde till 1960: ”Nous désirons contribuer”, sa han med sin varma och klangfulla röst, ”à créer un noyau de la structure européenne.”
Robert Schuman avslutade sitt första anförande som talman för Europeiska parlamentariska församlingen med ett åtagande om att arbeta för att ena den europeiska kontinenten. Han ansåg att Europa måste betrakta sig själv som en värdegemenskap som förenar kontinentens fria nationer: ”Ainsi seulement l'Europe réussira à mettre en valeur le patrimoine total qui est commun à tous les pays libres.”
Jag skulle vilja bygga vidare på detta.
EU är en värdegemenskap.
Våra institutioner är inte ett mål i sig själva, utan existerar för att tjäna våra värderingar: individens värdighet, mänskliga rättigheter, demokrati, rättsstatsprincipen och ekonomiskt och socialt välstånd.
De tjänar solidaritets- och subsidiaritetsprincipen.
Europa betyder respekt för varandra, respekt för vår mångfald, respekt för våra medlemsstaters värdighet, stora som små.
Denna respekt kan inte påtvingas, men är en viktig grundförutsättning för vår ömsesidiga förståelse och gemensamma verksamhet.
Respekt för EG-rätten, som gör det möjligt för oss att lösa våra tvister i godo och på fredlig väg uppnå en balans mellan olika intressen, måste ständigt förnyas genom de oskrivna regler som styr våra relationer i Europa: omtanke om och respekt för varandra.
(Applåder)
Jag skulle vilja uppmuntra och uppmana alla - oavsett politisk hemvist - att fortsätta visa varandra denna respekt.
Om denna ömsesidiga respekt - som kännetecknas av att visa tolerans för varandras övertygelser, men vara trogen sina egna och samtidigt vara beredd att sluta kompromisser - är framgångsrik, kan EU och Europaparlamentet stå modell för fred i världen.
Vårt europeiska arv bevaras i våra nationers enighet och fredliga samexistens. De har gått samman och bildat Europeiska unionen.
Vi hedrar Robert Schuman och alla ledamöter i den första europeiska parlamentariska församlingen genom att sträva efter att verka i deras anda, och genom att arbeta för ett ansvarsfullt och öppet Europaparlament som finns nära medborgarna, men som om det behövs har kraften att visa politiskt ledarskap.
Om vi fortsätter vårt resoluta arbete har vi inget att frukta vid våra efterträdares bedömning av vårt arbete när de 2058 firar Europaparlamentets hundraårsjubileum.
Kolleger, mina damer och herrar! Låt oss tillsammans glädjas åt den frihet, fred och enighet som präglar den europeiska kontinenten, och som det är ett privilegium för oss att arbeta för.
(Kraftiga och ihållande applåder)
rådets ordförande. - (SL) Mitt anförande kan inte hållas utan känslor, så sa Europeiska parlamentariska församlingens första talman, Robert Schuman, när han för första gången talade i denna respekterade kammare den 19 mars 1958.
Femtio år senare, vid detta festliga jubileum, känner vi precis likadant.
Jag talar här inte bara till 142 nationella ledamöter utan till 785 direktvalda ledamöter av Europaparlamentet.
Om man ser tillbaka på den väg som vi har vandrat och hur den europeiska demokratin har blomstrat de senaste 50 åren blir man stolt och mycket tacksam gentemot dem som skapade Europatanken.
Samtidigt är det vårt ansvar att så bra vi kan fortsätta den europeiska traditionen av fred, samarbete och välstånd.
Låt oss gå tillbaka till 1958. Ett samhälle som led av effekterna av två destruktiva krig, en bipolär värld där väst stod mot öst, det kalla kriget, den kubanska revolutionen, det första chipset, atomexperiment och uppskjutningen av den första rymdsatelliten.
Etthundrasextioåtta miljoner européer i de sex grundarländerna slöt sig samman och bildade Europeiska unionen, vilket läkte krigsår, gav ekonomiskt välstånd och tillsammans med Atlantpakten tryggade fred och demokrati i området.
Tyvärr levde större delen av resten av Europa i en totalitär miljö med civil och ekonomisk stagnation eller till och med tillbakagång.
År 2008 är bilden en helt annan. För att hitta lösningar på dagens utmaningar bryr man sig i vår multipolära värld inte bara om ekonomisk och politisk konkurrens utan även i allt högre grad om samarbete.
Avskaffandet av de gränser som delade Europa längs Berlinmuren, avskaffandet av järnridån och övervakningen av de interna gränserna kommer att fortsätta den här månaden genom att luftrumsgränserna avskaffas inom det utökade Schengenområdet.
Europeiska unionens territorium är mer än tre gånger så stort som för 50 år sedan och unionen har tre gånger så stor befolkning, 23 officiella språk, en starkare inre marknad och en gemensam valuta.
EU-medborgarnas medellivslängd är åtta år längre.
Tjugosju stats- och regeringschefer - en tredjedel av oss levde under totalitära regimer för 20 år sedan - kommer att fatta beslut runt samma bord i morgon.
I dag lever nästan hela Europa i frihet och i demokratier.
Vi bör uppmärksamma denna framgång och fira den.
Europaparlamentets arbete sedan 1958 speglar tydligt de framsteg som har åstadkommits tack vare de senaste 50 årens integration.
Efter er inledande rådgivande roll fick ni under det tidiga sjuttiotalet era första riktiga befogenheter i samband med gemenskapsbudgeten.
Och i slutet av sjuttiotalet höll ni era första direkta val.
Tack vare nya avtal fick ni starkare befogenheter vid antagandet av lagstiftning och vid utnämningen av de högsta europeiska politiska företrädarna.
Den nya Europeiska kommissionen kan inte heller existera utan ert förtroende.
På samma sätt som Romfördraget gav parlamentet nya ansvarsområden 1958, innebär Lissabonfördraget 50 år senare ett stort steg framåt för Europaparlamentet.
Medbeslutandeförfarandet kommer att utvidgas till att omfatta nästan all EU-politik och Europaparlamentets demokratiska kontroll, upprättandet av internationella avtal och utnämningen av de högsta EU-företrädarna kommer att stärkas.
Det gladde mig mycket när ni vid sammanträdesperioden förra månaden antog betänkandet om Lissabonfördraget med stor majoritet.
Jag skulle också vilja gratulera alla medlemsstater som redan har ratificerat detta fördrag. Och jag hoppas att de snart ska följas av de återstående medlemsstaterna.
Medan EU:s första 50 år ägnades åt den europeiska agendan, vår politiska och ekonomiska utveckling och reformer kommer de kommande 50 åren säkerligen även att inriktas på den globala agendan.
Detta framgår tydligt av de ämnen som ska tas upp vid Europeiska rådets möte i morgon.
Det råder ingen tvekan om att vi endast kan hitta godtagbara lösningar på utmaningarna från Lissabon, miljö- och energifrågorna och oron på finansmarknaderna om vi tar hänsyn till globala trender och aktörer och inkluderar dessa i vår verksamhet.
Detta gäller även mänskliga rättigheter och interkulturell dialog, där Europaparlamentet verkligen spelar en ledande roll.
Jag skulle vilja utnyttja detta tillfälle till att på Europeiska rådets vägnar tacka er för er roll när det gäller att uppmärksamma människorättskränkningar och ert valövervakningsarbete och för era delegationers arbete i internationella organ som FN:s råd för mänskliga rättigheter.
Er roll inom de gemensamma parlamentarikerkommittéerna är också viktig och skapar ett mervärde för EU:s politik gentemot tredjeländer och regioner.
Genom er verksamhet och möten med framstående gäster under Europeiska året för interkulturell dialog stärker ni en av de grundläggande europeiska traditionerna, dvs. att ömsesidig respekt och förståelse är grundpelarna för samexistens såväl i Europa som i resten av världen.
Men den styrs av en enda regel. Framgången står i proportion till graden av enighet bland medlemsstater, sektorer, gemensamma intressegrupper och generationer och inom regionala, nationella, europeiska och globala faktorer.
Här måste EU-institutionerna föregå med gott exempel.
”Varje person är en ny värld.
Endast institutioner som bevarar den kollektiva erfarenheten kan mogna.”
Med dessa ord tar Jean Monnet oss ett steg närmare en förklaring till varför EU:s vision fortfarande ofta skiljer sig från verkligheten, och varför många européer, trots de uppenbara framgångarna de senaste 50 åren, fortfarande tvivlar på den europeiska integrationens fördelar.
För att förstå och värdera frihet, fred och mångfald, avsaknaden av gränser och fördelarna med och framtida utsikter till ett enat Europa måste vi alltid vara medvetna om att det finns andra, mycket värre alternativ.
Det är därför som vi måste hålla den europeiska kollektiva tanken vid liv.
Från den kan vi hämta styrka att möta dagens utmaningar.
Gårdagens tankar måste förenas med framtidens tankar.
Hade vi inte slagit oss samman för 50 år sedan skulle vi förmodligen inte ha levt i frihet och välstånd i dag.
Samma sak kan sägas om de kommande 50 åren.
Om vi inte tillsammans försöker hitta lösningar för att minska koldioxidutsläppen och spara energi kommer vi inte att lyckas bromsa klimatförändringen.
Vi kommer att drabbas av fler och fler översvämningar, orkaner, torka, nya sjukdomar, hotade ekosystem och miljöflyktingar.
Det är viktigt att resultaten av EU:s beslut och verksamhet är tillräckligt konkreta och påtagliga för medborgarna för att de ska förstå hur oerhört viktigt EU är för att bevara och förbättra deras livskvalitet.
Herr talman, mina damer och herrar! Jag skulle vilja tacka er för ert bidrag till EU:s utveckling de senaste 50 åren.
Jag vet vad det har inneburit för våra generationer.
Jag föddes faktiskt samma år som Europaparlamentet.
Så länge detta mandat varar, och även efter det, önskar jag er all lycka i ert arbete, massor av nya idéer och ett envist framhärdande i utvecklandet av europeiska värden, demokrati och levnadssätt.
Jag är övertygad om att när vi firar nästa jubileum för denna europeiska demokratiska församling kommer vi ännu en gång att kunna fira synliga framsteg i Europa.
(Applåder)
Ett stort tack till Europeiska rådets ordförande.
Jag ger nu ordet till Europeiska kommissionens ordförande José Manuel Durão Barroso.
kommissionens ordförande. - (FR) Herr talman! Herr rådsordförande, ordförande för de olika EU-institutionerna, tidigare talmän i denna församling, mina damer och herrar, företrädare för de nationella parlamenten, ärade gäster!
Jag är väldigt glad att kunna fira Europaparlamentets första femtio år med er i dag.
Detta jubileum har en stor symbolisk och politisk betydelse för Europa. För femtio år sedan ledde Robert Schuman en ny gemensam församling.
De tre europeiska gemenskaperna hade precis skapat den första versionen av europeisk demokrati.
Sedan dess har detta grundläggande politiska val bekräftats om och om igen i varje stadium av den europeiska integrationen.
Innan någon annan insåg EU:s grundare att det framväxande Europa krävde robusta demokratiska europeiska institutioner för att förkroppsliga de allt starkare banden mellan de sex grundarländerna.
I enlighet med Jean Monnets inspirerade vision var det dessutom nödvändigt att institutioner kunde utvecklas och anpassas till vad EU:s grundare såg som de två viktigaste framtida händelserna: djupare integration och geografisk utvidgning.
Jag måste säga att jag fortfarande är mycket rörd över att se alla er här i denna europeiska demokratiska församling, direktvalda företrädare från länder som fram tills nyligen åtskildes av diktaturer som hindrade Europa från att gjuta liv i friheten.
(Applåder)
Den institutionella triangel som EU:s grundare lämnade i arv till oss är en unik modell i världen och efter 50 år är den fortfarande vital och kraftfull.
Den har anpassat sig till en kraftig utvidgning av de uppgifter som anförtroddes gemenskapen, och nu EU.
Den har även klarat av en stark dynamisk utvidgning av unionen.
Vi har vår sinnrika och balanserade institutionella modell att tacka för denna framgång, en modell som inte följer den klassiska maktfördelningen.
Vi har även vår arbetsmetod att tacka för denna framgång, en metod som respekterar både gemenskapsmetoden och subsidiaritetsprincipen.
Institutionerna är emellertid inte ett mål i sig själva. De tjänar fortfarande ett ideal och mål.
De arbetar i våra medborgares tjänst.
Ju starkare institutionerna är, desto bättre kan de tjäna detta ideal och våra medborgare.
Framför allt ville EU:s grundare bygga Europa för fredens skull.
De ville bygga det nya Europa genom solidaritet.
De valde ekonomi som drivkraften bakom sin politiska vision och sina mål.
Efter femtio år behöver det fredliga Europa, utvidgat till kontinentala dimensioner, starka institutioner för att klara dagens utmaning: globaliseringen.
Ingen medlemsstat kan själv klara denna utmaning.
Tack vare sin erfarenhet av att öppna marknader tillsammans med regler som förkroppsligar värden som frihet, solidaritet och hållbar utveckling är det endast Europa som har de dimensioner, institutioner och instrument som krävs för att hantera och forma globaliseringen.
För att möta denna utmaning måste tjugohundratalets Europa enas för att skörda framgångar i den kunskapsbaserade ekonomin, skapa arbetstillfällen för Europas män och kvinnor och göra sin ekonomi mer dynamisk.
Det måste inta sin rättmätiga plats på världsscenen: en europisk makt, utan arrogans, ett Europa som kan föreslå - inte påtvinga, föreslå - värden som frihet och solidaritet till världen.
Vi kommer att lyckas om vi fortsätter vårt konstruktiva partnerskap mellan våra institutioner.
Inom ramen för detta partnerskap vill jag gratulera Europaparlamentet för dess bidrag till Europaprojektet i alla olika aspekter av våra medborgares dagliga liv.
Under sina femtio år har denna församling fått många befogenheter och en avsevärd makt.
Jag menar makt i betydelsen legitimitet som kommer direkt från europeiska män och kvinnors röster.
Jag menar också makt i dess formella betydelse: medbeslutande, budgetbefogenheter och demokratisk kontroll över EU-institutionerna.
Vad jag egentligen menar är politiskt inflytande.
Europaparlamentet har samtidigt tagit plats som medlagstiftare med delat ansvar inom den institutionella triangeln och i det europeiska politiska livet. Men parlamentet har även knutit allt starkare band med de nationella parlamenten, varav många är representerade här i dag.
Den makt som Europaparlamentet har tillförskansat sig under årens lopp har stärkt EU.
Ett starkt Europaparlament är en viktig partner för de andra institutionerna och - jag måste betona detta - för Europeiska kommissionen.
Jag tror att jag kan säga att förhållandet mellan våra två institutioner blir allt tätare, kraftfullare och mognare. Och det gläder mig mycket.
När Lissabonfördraget har ratificerats kommer detta att stärka gemenskapsinstitutionerna ännu mer.
Det kommer att ge Europaparlamentet mer makt.
Det kommer att främja kommissionens dubbla politiska legitimitet genom starkare band till Europaparlamentet och Europeiska rådet.
Det kommer att ge Europeiska rådet ett fast ordförandeskap, vilket gör att förberedelserna och övervakningen av Europeiska rådets möten kan ske på ett mer konsekvent sätt.
Det kommer att bidra till att utveckla den roll som unionens höga representant för utrikes- och säkerhetspolitiken har, som även kommer att fungera som Europeiska kommissionens vice ordförande.
Genom att stärka våra institutioners legitimitet och göra dem effektivare innebär Lissabonfördraget ett stort steg framåt för EU.
Såväl i dag som i morgon måste vi inse att det inte kan bli tal om något nollsummespel mellan institutionerna.
Ingen av våra institutioner bör stärkas på bekostnad av de övriga.
Tvärtom vill vi alla ha starkare EU-institutioner så att EU kan bli effektivare och mer demokratiskt.
Alla våra institutioner kommer att tjäna på att EU:s institutionella struktur konsolideras.
Mina damer och herrar! I samband med det datum som vi högtidlighåller i dag kom jag att tänka på ett citat från den stora portugisiske författaren Agustina Bessa Luis.
Hon sa att vid 15 års ålder har man en framtid, vid 25 ett problem, vid 40 erfarenhet, men innan femtio har man faktiskt ingen historia alls.
I dag kan Europaparlamentet, denna europeiska demokratiska församling, stolt hävda att det har en lysande historia. Men jag är säker på att ni även har en lysande framtid.
Därför vill jag på Europeiska kommissionens och mina egna vägnar framföra mina hjärtligaste gratulationer och ett stort lycka till med ert arbete för ett enat Europa.
(Applåder)
Stort tack till Europeiska kommissionens ordförande.
Jag skulle nu vilja välkomna Joachim Opitz. Han är här i dag som företrädare för alla tidigare generalsekreterare.
Nu får vi nöjet att än en gång lyssna till Europeiska unionens ungdomsorkester.
(Kort framförande av Europeiska unionens ungdomsorkester.)
(Kraftiga applåder)
(Kammaren reste sig och lyssnade till Europahymnen)
(Sammanträdet avbröts kl. 16.15 och återupptogs kl. 16.20.)
4.
Beskattning av blyfri bensin och diesel (
Röstförklaringar
Muntliga röstförklaringar
(EN) Fru talman! Vad man än tycker om den aktuella debatten om klimatförändringen, och jag tycker mig ana en hel del tomt snack här - tycker jag att vi alla kan enas om behovet av mer energieffektivitet.
Men om vi ska tala om energieffektivitet måste vi se till att vår uppfattning faktiskt till viss del är enhetlig i denna fråga.
Jag ska ge ett exempel: hela vår politik med energisparglödlampor.
Ja, vi vill fasa ut de befintliga glödlamporna, men ändå inför vi avgifter på importen av energisparglödlampor.
Ja, vi talar om att förbjuda kvicksilver i barometrar (även om det faktiskt utgör en mycket liten risk), men ändå uppmuntrar vi samtidigt användningen av energisparglödlampor som innehåller, ja ni gissar rätt, mer kvicksilver.
Inte bara det, utan vi talar om energieffektivitet, men ändå fortsätter vi att resa hit till Strasbourg, vilket släpper ut tonvis med onödigt extra koldioxid.
Om vi verkligen vill gå i täten för energieffektivitet borde vi därför lägga ned parlamentet i Strasbourg.
(PL) Herr talman! Jag röstade för gemenskapens delaktighet i ett forsknings- och utvecklingsprogram i syfte att öka livskvaliteten för äldre människor genom användningen av ny informations- och kommunikationsteknik.
Projektet omfattar utvecklingsmöjligheter inte bara för äldre utan också för funktionshindrade, kvinnor som uppfostrar barn i hemmet och människor på landsbygden.
Enligt min åsikt kommer detta initiativ att hindra en social skiktindelning i Europa på området för tillgången till digitala tjänster, såväl som marginaliseringen av sociala grupper som hotas av en begränsad tillgång till modern teknik.
Det är dock mycket viktigt att komma ihåg att kostnaden för denna teknik måste hållas så låg som möjligt.
(PL) Jag röstade för betänkandet om ”att öka livskvaliteten för äldre människor”, i vilket man hanterar frågor av stor vikt för många EU-medborgare, särskilt den äldre generationen.
Äldre personer är beroende av pensionsförmåner, vilka för det mesta är mycket låga.
Problemet växer med det ökande antalet äldre personer som får dessa förmåner, vilka är begränsade eftersom antalet bidragsgivare minskar.
Vi är alltså på väg mot en situation där en stor grupp äldre personer kommer att ansöka om olika sociala förmåner.
Många av dem kan dock fortfarande utföra olika typer av arbete och kan förbli aktiva på arbetsmarknaden.
Det växande antalet äldre personer, tillsammans med behovet av allt fler tjänster och produkter, ökar efterfrågan på detta område.
(PL) Herr talman! Jag röstade emot betänkandet, eftersom det väcker en rad tvivel.
Jag stöder inte bestämmelserna i direktivet om harmonisering av punktskattesatserna för dieselbrännolja och bensin.
Flera punktskattesatser skapar möjligheter till konkurrens mellan transportföretag från olika EU-länder, vilket tveklöst gagnar konsumenten.
Jag motsätter mig också bestämmelserna om höjda punktskattesatser för bränsle inom hela EU.
Höga oljepriser på de nationella marknaderna och en harmonisering av punktskatterna i alla 27 EU-länder kommer att hindra den ekonomiska tillväxten i länder med låg BNP.
Höjda bränslepriser innebär höjda priser på varor och tjänster.
Jag röstade därför för de ändringsförslag som lagts fram i syfte att låta de nya medlemsstaterna, däribland Polen, bevara olika punktskattesatser.
(PL) Herr talman! Jag röstade emot betänkandet, eftersom den avsevärda höjningen av punktskatter för dieselbrännolja kommer att leda till höjda tullavgifter för varor och tjänster i länder som ska ta ut en lägre punktskattesats än den föreslagna lägsta punktskatten inom gemenskapen, men som ändå är höga med tanke på förhållandena i dessa länder.
Med tanke på att den genomsnittliga inkomsten i de medlemsländer som anslöt sig till EU 2004 och 2007 är relativt låg, är den föreslagna höjningen av punktskatten för stor.
Dess effekt kommer att bli särskilt kännbar i de fattigaste familjerna, eftersom den aktuella höjningen av bränslepriserna redan är en stor börda för deras hushållsbudgetar.
De minst utvecklade länderna, med sina låga inkomstnivåer, borde därför beviljas mycket längre övergångsperioder än de som Europeiska kommissionen föreslår, för att de ska få tid att anpassa sig.
Jag anser därför att den föreslagna ökningen är omotiverad och för stor.
(EN) Herr talman! Det är mycket roligt att se er tillbaka i talmansstolen, varifrån ni lyssnar på dessa röstförklaringar som jag vet att ni verkligen uppskattar.
Jag vill också säga att jag uppskattar vänligheten och förståelsen hos er personal, era tjänsteavdelningar och tolkar denna vecka, när vi har gjort dessa röstförklaringar.
Jag röstade emot detta särskilda betänkande av en massa anledningar.
För det första tror jag på skattekonkurrens.
Jag anser inte att skatteharmonisering eller skatter ska vara en fråga för EU-institutionerna överhuvudtaget.
För det andra har finansministern i mitt land den här veckan infört högre bränsleskatt för brittiska bilar och transportfordon utan att förstå följderna av detta.
Jag vill ta upp ett separat problem.
Jag för en kampanj tillsammans med Northampton Chronicle and Echo för de personer som bor i närheten av min region, där vi får betala mer för vårt bränsle än i alla andra stora städer i närheten.
Jag vill betona att det finns andra problem inom bränslemarknaden, förutom skatteproblemen.
(EN) Herr talman! Jag vill upprepa kommentarerna från min kollega och tacka er, personalen och tolkarna för ert vänliga tålamod när vi försöker lämna dessa röstförklaringar, som ibland kan vara underhållande och ibland tämligen trista för er.
Det förstår jag.
Men det är den underbara kontrasten här i parlamentet.
Låt oss nu tala om skattekonkurrens.
Vi talar om att skapa världens största inre marknad här, och vi talar om att göra EU till världens mest konkurrenskraftiga ekonomi, och vi talar om världskonkurrens, men vad gör vi när det gäller skattekonkurrens?
Jo, liksom det faktiskt anges i motiveringen, är det bästa sättet att lösa konkurrensproblemet att införa en fullständig harmonisering.
Så vi betraktar alltså konkurrensen som ett problem, samtidigt som vi talar om behovet av en mer konkurrenskraftig ekonomi.
Detta borde inte vara en behörighet för EU.
Det är en behörighet för medlemsstaterna, och vi borde låta det vara så, eftersom det bästa sättet att garantera en konkurrenskraftig ekonomi är att se till att vi har skattekonkurrens och inte harmonisering.
(PL) Herr talman! Jag röstade emot betänkandet.
Europeiska unionen har inget intresse av att finansiera Irak.
Det finns andra länder i själva Europa som skulle gagnas mer av detta stöd.
Av rapporten från Caritas Europa framgår att ensamma föräldrar, särskilt kvinnor i 14 europeiska länder - däribland Polen, Österrike, Tyskland och Storbritannien - är särskilt drabbade av fattigdom.
Enligt en EU-rapport har Polen den högsta procentandelen barn som lever i fattigdom av alla EU-länder, med 26 procent.
En polack av fem (19 procent) lever under fattigdomsgränsen.
Och 22 procent av de polska barn som har åtminstone en arbetande förälder hotas av fattigdom.
Det är den högsta siffran i Europa.
Tretton procent av de polacker som har en anställning hotas av fattigdom.
I Österrike lever 47 procent av de arbetslösa ensamstående föräldrarna i kronisk fattigdom.
Låt oss inrikta vårt arbete på Europa.
(EN) Herr talman! I går när ni satt i talmansstolen betonade jag att jag alltid njuter av att läsa betänkandena från utskottet för kvinnors rättigheter och jämställdhet mellan kvinnor och män här i kammaren och undrar varför detta utskott finns.
För att visa min poäng har vi i dag ett betänkande vars slutsatser snarare verkar ha dragits av någon som sett för mycket på tv-serien Kvinnofängelset när de var barn i stället för att titta på den faktiska situationen för kvinnor i fängelse - och huruvida det borde vara en behörighet för parlamentet hur som helst.
I skäl Q anges till exempel: ”Det ökade antalet kvinnor på fängelserna beror delvis på kvinnornas försämrade ekonomiska villkor.”
Jag tror, och jag har kontrollerat detta mot statistiken från ett antal EU-länder, att antalet kvinnor i fängelse helt enkelt ökar för att befolkningen växer.
Andelen kvinnor på fängelserna i Europa sjunker faktiskt.
Det anges här att tillgång till all slags hälsovård ska ges av mycket hög kvalitet i fängelserna.
Det är helt korrekt.
Men det finns många äldre kvinnor i min valkrets som skulle älska att få samma hälsovårdsförmåner som kvinnorna på de brittiska fängelserna.
Därför lade jag ned min röst i omröstningen om betänkandet.
(NL) Jag framhöll i går Turkiets oantastliga position som aspirerande medlemsstat och i detta betänkande bekräftas endast denna särskilda status.
Turkiet har i veckor bombat norra Irak och tiotusentals turkiska trupper har invaderat landet.
Och i stället för att tydligt fördöma dessa angrepp, vad gör parlamentet?
Det ber snällt Turkiet att respektera Iraks territoriella integritet.
Alla regler, alla principer, alla riktlinjer och alla kriterier måste åsidosättas för en turkisk anslutning, från Köpenhamnskriterierna till den internationella rätten och dess förbud mot användningen av angrepp.
Turkiet anser sig stå över lagen och all lagstiftning, och stärks ständigt i denna uppfattning av Europa.
En dag kommer Europeiska unionen att få ångra sin inställning.
(DE) Herr talman! Jag var en sträng och tydlig kritiker av och motståndare till Irak-kriget och det är jag fortfarande.
Jag tror dock att vi också måste kompensera för våra misstag där.
Vi i västvärlden - såväl Europa som USA - har därför en plikt att göra vårt bästa för att säkra fred och stabilitet, vilket kommer att vara svårt nog.
Därför är Gomesbetänkandet utomordentligt bra.
Vi måste verkligen ta tillfället i akt att stödja Irena Záborskás initiativ till frigivandet av den kidnappade ärkebiskopen.
Jag beklagar att resolutionen om detta ämne på grund av ett administrativt misstag här i kammaren inte står med på eftermiddagens dagordning.
Det är vår plikt att göra allt vi kan för att hjälpa denna företrädare för en minoritet vars existens hotas, som har levt tillsammans i fred med sina muslimska grannar i århundraden och som hotas med folkmord precis vid en tidpunkt då vi tar vårt ansvar i Irak.
Det är inte acceptabelt och därför måste vi vidta beslutsamma åtgärder här.
(PL) Herr talman! Jag håller med om mycket i Marie Panayotopoulos-Cassiotous betänkande om situationen för kvinnor i fängelse.
Fängelseledningarna måste kunna garantera rimliga förhållanden för personer som avtjänar fängelsestraff eller som är tillfälligt häktade.
Jag vill uppmärksamma situationen för kvinnor som är anställda på fängelser.
I Polen är 5 000 av de 30 000 kriminalvårdarna kvinnor.
Kriminalvårdarnas ersättning överstiger inte 500 euro per månad.
Med tanke på fängelsepersonalens betydelse när det gäller att se till att straffen avtjänas vederbörligen är det viktigt att merparten av de kriminalvårdare som vaktar kvinnliga fångar är av samma kön.
Det minskar de kvinnliga fångarnas obehag och garanterar ett bättre skydd av deras rättigheter.
Utan en avsevärt höjd ersättning och bättre arbetsvillkor i fängelserna kommer vi inte att nå målen i betänkandet.
(EN) Herr talman! Jag röstade enligt partipiskan om detta särskilda betänkande och emot många av ändringsförslagen.
Jag har dock ett problem med innehållet i skälen.
Det anges att ”det är nödvändigt att skapa en nationell styrka som upprätthåller ordningen, som består av representanter för de olika grupperna och som har alla gruppers förtroende”.
Det handlar om Iraks folk, och den nationella styrkan ska skapas av Iraks folk antar jag.
Man undrar faktiskt hur stor beslutsamhet som de enskilda medlemsstater som bildar Europaparlamentet har lagt ned på detta hittills.
Allt man behöver göra är att se på hur många som har ställt sig bakom insatserna i Irak, oavsett om de tror på dem eller inte.
När vi gör det borde vi försöka att undanröja de problem som vi har orsakat.
Jag anser verkligen att denna resolution visar att det kan orsaka oss många problem att försöka att införa en harmoniserad gemensam utrikes- och säkerhetspolitik i framtiden, såväl här i parlamentet som i våra medlemsstaters huvudstäder.
(DE) Herr talman! Liksom majoriteten av min grupp röstade jag emot detta betänkande, inte bara på grund av ämnet, utan för att denna viktiga fråga fortsätter att utnyttjas för ideologiska strider om begreppen sexuell och reproduktiv hälsa och sexuella och reproduktiva rättigheter.
Jag vill vädja till alla grupper i kammaren att upphöra med denna ideologiska dispyt, som skadar den här frågan.
Vi måste klargöra att reproduktiv hälsa är viktigt, men att det inte har något att göra med abort, eftersom det inte faller inom Europeiska unionens ansvarsområde och varje stat har rätt att stifta sina egna lagar på detta område.
Det är förenligt med subsidiaritetsprincipen, och därför får EU-medborgarnas pengar inte användas i syften som några EU-medlemsstater av etiska, moraliska och rättsliga skäl inte ser som acceptabla.
Vi borde därför helt klart utesluta detta ämne ur våra diskussioner och rikta in oss på neutrala begrepp som faktiskt rör hälsa och inte har något att göra med abortfrågan, om vilken åsikterna går i sär här i kammaren och i vilken jag starkt förespråkar att skydda det ofödda barnet.
Skriftliga röstförklaringar
skriftlig. - (EN) Jag stöder Claude Turmes betänkande om den globala fonden för energieffektivitet och förnybar energi.
Denna fond kommer att använda begränsade offentliga medel för att främja privata investeringar i projekt för energieffektiv och förnybar energi i utvecklingsländer och i övergångsekonomier.
Denna fond, som hjälper alla att nå en viss nivå med energieffektivitet och som stöder förnybar energi, har mitt stöd och jag röstade för den.
skriftlig. - (RO) Resolutionen handlar om inrättandet av ett innovativt finansiellt instrument för att stödja genomförandet av vissa projekt som finansieras genom denna fond till stöd för övergången till en ekonomi med låga koldioxidutsläpp och för anpassning till klimatförändringens effekter.
Att utveckla en sådan ekonomi genom projekt som finansieras genom fonden innebär att nya arbetstillfällen och lika villkor för social utveckling skapas och att skillnader avskaffas.
I denna bemärkelse är det särskilda stöd som avsätts för små- och medelstora företag med tillgång till finansiering för deras projekt inom ramen för den globala fonden positivt.
Jag röstade för denna resolution, eftersom jag anser att dessa två typer av åtgärder, nämligen avskaffandet av utsläppen av växthusgaser och anpassningen till klimatförändringens effekter, måste utarbetas samtidigt, genom en sammanhängande och gemensam politik med positiv inverkan på utvecklingen av en arbetsmarknad och skapandet av nya arbetstillfällen och en ökad BNP.
skriftlig. - (PT) Det kan generellt sägas att syftet med detta betänkande är att främja integrationen av de ”nya” medlemsstaterna i EU:s utrikespolitik, särskilt ”politiken för utvecklingssamarbete” och den ”europeiska grannskapspolitiken”.
I betänkandet konstateras också att de ”nya” medlemsstaterna utgör ett tillfälle för EU att ”stärka Europeiska unionens strategiska närvaro i Östeuropa, Centralasien och Kaukasien”, vilka är regioner som de ”nya” medlemsstaterna har prioriterade förbindelser med och som har fått mindre ”EU-stöd” hittills.
Detta innebär att man måste eftersträva att använda den privilegierade förbindelsen med de östeuropeiska länder som anslöt sig till EU 2004 som ett europeiskt interventionsinstrument (med beaktande av de stora makternas och deras stora ekonomiska och finansiella gruppers intressen, särskilt inom energisektorn) i länderna i Oberoende staters samvälde, på västra Balkan och på Kaukasus.
Det vill säga att man måste eftersträva att använda dessa länders ”erfarenhet” av ”övergången” till kapitalism och till ett medlemskap i Nato och EU som en typmodell i dessa regioner.
Detta är i slutändan vad det handlar om: en politik som döljer kapitalismens intresse för ”utveckling”.
skriftlig. - (EN) Jag stöder DanutBudreikaitės betänkande om utmaningen med EU:s utvecklingspolitik för de nya medlemsstaterna.
Samtidigt som EU:s nya medlemsstater, förutom Malta och Cypern, har en unik expertkunskap när det gäller tillämpningen av och inriktningen för utvecklingspolitiken i våra grannländer i öst, måste vi aktivt uppmuntra deras deltagande i Afrika söder om Sahara och i andra minst utvecklade länder.
Våra nya medlemsstater stärker EU:s roll som en världspartner och de borde få fullständigt stöd i den rollen.
Betänkandet och dess rekommendationer har mitt stöd.
skriftlig. - (PT) Blotta det faktum att vi diskuterar de nya medlemsstaternas roll i Europeiska unionens samarbets- och utvecklingspolitik, särskilt med AVS-länderna, är ett tydligt bevis på framgången för utvidgningsprocessen och för integrationen av de länder som har anslutit sig under de senaste åren.
De ”före detta östeuropeiska länderna” hade förvisso en lång tradition av ”samarbete” med Afrika, och det kan hända att förbindelserna kvarstår, om än under helt andra villkor.
Den mest relevanta frågan är dock att dessa länder, som fortfarande tappert kämpar med kostnaderna för sina reformer, nu kan bidra till samarbetet och utvecklingen med sina befolkningars aktiva samtycke.
Detta exemplariska tillvägagångssätt skulle kunna vara en förebild, vilket vi hoppas, för andra länder i stort sett samma omständigheter i andra delar av världen.
skriftlig. - (PL) Jag röstar för Danuté Budreikaitės betänkande om utmaningen med EU:s politik för utvecklingssamarbete för de nya medlemsstaterna.
Betänkandet håller mycket hög kvalitet, och innehåller en detaljerad analys av den nuvarande situationen för de nya medlemsstaternas utvecklingssamarbete, av de berörda institutionerna och programmen, av mottagarländerna och av de berörda finansiella medlen.
I de frågor som tas upp i betänkandet betonas förbindelserna mellan EU:s medlemsstater och deras nya grannar i öst.
De nya medlemsstaterna är viktiga länkar mellan EU och dess nya grannländer.
Jag vill personligen att effektiva samarbetsformer ska utarbetas mellan de gamla och nya givarna till förmån för de minst utvecklade länderna, inom ramen för vilka de nya medlemsstaternas dominerande inflytande i vissa regioner eller länder ska utnyttjas.
skriftlig. - (PT) Jag röstade för Neena Gills betänkande om förslaget till Europaparlamentets och rådets beslut om gemenskapens deltagande i ett forsknings- och utvecklingsprogram.
Detta program syftar till att öka livskvaliteten för äldre människor genom användning av ny informations- och kommunikationsteknik (IKT).
Europeiska unionens deltagande i detta program kommer att öka unionens möjligheter att ta itu med den demografiska förändringen.
Användningen av IKT kan hjälpa äldre människor att bli mer oberoende och att förbli friska, och det kan öka deras livskvalitet.
skriftlig. - (PT) Vi röstade för detta betänkande, som handlar om Europeiska kommissionens förslag om EU:s deltagande i ett forsknings- och utvecklingsprogram som de olika medlemsstaterna har beslutat att inrätta på området för ny informationsteknik (IKT) för att hjälpa äldre människor och ge dem möjlighet att agera effektivt.
Programmet ”IT-stöd i boende” syftar till att nå samverkanseffekter i fråga om förvaltnings- och finansieringsresurser.
Också Portugal deltar.
I betänkandet, som Europaparlamentet nu har antagit, uppmärksammas och läggs konkreta förslag fram för främjandet av kvinnors roll inom vetenskap och forskning, och betoning läggs på små och medelstora företags deltagande och på lika tillgång för alla medlemsstater till kostnadseffektiva lösningar så att man undviker att öka den digitala klyftan och därmed skapa ett Europa med två hastigheter.
Det föreslås också att kommissionen ska göra en etappgranskning senast 2010 för att bedöma kvaliteten och effektiviteten hos programmets genomförande.
skriftlig. - (FR) Jag vill göra två kommentarer om Gillbetänkandet, som i grunden handlar om att utarbeta forskningsprogram i syfte att göra äldre personer mer oberoende genom användningen av informations- och kommunikationsteknik.
Min första kommentar handlar om förslagens innehåll: det är svårt att se vilket mervärde Europeiska unionen skulle tillföra ett förslag som, helt berättigat, initierats av ett antal medlemsstater - förutom att det skulle göra processen mer byråkratisk och förutom att ett nytt gemenskapsorgan skulle inrättas.
Unionens finansiella bidrag, som uppgår till 150 miljoner euro under ett antal år minus driftskostnaderna för det nämnda nya organet, tycks inte vara ett avgörande argument.
Min andra kommentar rör förslagens utformning.
Det är allt vanligare att lagstiftningsförslag läggs fram i kammaren i form av kompromisser mellan parlamentet och rådet - i syfte att påskynda förfarandet genom att underlätta förslagens antagande vid första behandlingen.
Vad vi ser i praktiken är dock ett lagstiftningsorgan som hålls gisslan av en grupp expertförhandlare.
Jag betraktar spridningen av denna praxis som ett hot mot demokratin.
skriftlig. - (FR) Jag röstade för betänkandet med ett förslag om att Europeiska unionen ska delta i forsknings- och utvecklingsprogrammet om IT-stöd i boende, som har initierats gemensamt av ett antal medlemsstater och tredjeländer.
Den åldrande befolkningen är en utmaning för det europeiska samhället och dess ekonomi.
Den genomsnittliga förväntade livslängden är i dag 80 år och antalet personer på mellan 65 till 80 år kommer att öka med ungefär 40 procent mellan 2010 och 2030.
Nya lösningar tillkommer för att hjälpa människor att hantera minnesförlust, nedsatt syn, hörsel eller rörelseförmåga och minskat oberoende, vilket vi löper allt större risk att drabbas av ju äldre vi blir.
Europeiska unionens deltagande i programmet planeras inom ramen för Europeiska kommissionens sjunde ramprogram för forskning och utveckling.
Europeiska unionen kommer att avsätta 150 miljoner euro för att samfinansiera projekt som kommer att ha en hävstångseffekt värd åtminstone 600 miljoner euro mellan 2008 och 2013.
De länder som deltar i programmet för IT-stöd i boende ska också hjälpa till att finansiera programmet genom att bidra med ett lika stort eller större belopp, vilket innebär att varje land ska investera 20 procent av sin nationella forskningsbudget på detta område.
skriftlig. - (PL) Jag röstade för Gillbetänkandet med titeln ”Att öka livskvaliteten för äldre människor”, som syftar till att främja användningen av modern informations- och kommunikationsteknik som ett stödinstrument för äldre personer.
Som vi vet utmärks våra samhällen av en allt högre förväntad livslängd.
Detta är en mycket positiv utveckling.
Genomsnittet i EU är nu 80 år, och andelen personer på över 65 år kommer snart att nå 40 procent.
Den nämnda tekniken kan avsevärt hjälpa dessa personer i olika situationer, däribland förlänga deras yrkesliv och deras sociala aktiviteter och öka deras livskvalitet.
Funktionshindrades särskilda behov måste naturligtvis också beaktas och tillgången till dessa tjänster och denna teknik måste garanteras främst genom tillhandahållandet av Internetanslutningar via bredband i både stads- och landsbygdsområden så att man undviker geografisk diskriminering.
skriftlig. - (DE) Jag förespråkar att Europeiska unionen ska samfinansiera programmet för IT-stöd i boende, eftersom det inte bara skulle gynna äldre personer utan också andra befolkningsgrupper, såsom personer med funktionshinder.
Det är just på grund av den stora demografiska förändringen av den europeiska befolkningen och den ökade förväntade livslängden under de senaste årtiondena som vi måste stödja ny informations- och kommunikationsteknik som kan göra det avsevärt lättare för människor att hantera de vardagliga hinder som de möter.
Vad gäller den allmänna kostnadsbesparingen inom hälsosektorn till följd av användningen av denna nya teknik vill jag också uppmärksamma er på forskningen om system för ”mobil hälsoövervakning”, vars användning skulle kunna minska de årliga hälsokostnaderna med 1 500 miljoner euro enbart i Tyskland.
Låt mig betona att en av fördelarna med samfinansiering vore att det också skulle ha en positiv inverkan på den privata sektorn, eftersom det indirekt skulle hjälpa små och medelstora företag.
Jag stöder beslutsamt programmet för IT-stöd i boende, eftersom den nya tekniken innebär att äldre personers privatliv fortsatt respekteras och gör det möjligt för dessa människor att åldras med värdighet.
skriftlig. - (EN) Jag stöder Nina Gills betänkande om ”att öka livskvaliteten för äldre människor”.
Genom att slå samman resurserna och samordna forskningen och utvecklingen på EU-nivå kan vi på ett lämpligare sätt bedöma hur vi kan öka våra äldre medborgares livskvalitet.
Genom att fastställa ett minimibidrag garanterar vi alla medlemsstaters deltagande i denna fråga.
Jag vill gratulera föredraganden till hennes betänkande och stöder rekommendationerna i betänkandet.
skriftlig. - Vi har valt att stödja betänkandet i sin helhet, då vår uppfattning är att EU måste komma tillrätta med osund skattekonkurrens på bränsleområdet, främst för att EU ska kunna uppnå sina klimatmål.
Förslaget om skatteharmonisering ska inte heller hindra enskilda medlemsländer att höja sina koldioxidskatter på bensin och diesel.
Detta är ytterligare en viktig orsak till att vi stöder betänkandet.
skriftlig. - (PT) Detta förslag till direktiv syftar till att minska prisskillnaderna för bränsle mellan de olika medlemsstaterna, vilket leder till en snedvridning av konkurrensen och till miljöförstörelse inom vägtransporter.
Prisskillnaderna mellan dieselbrännolja som används som motorbränsle och blyfri bensin är förvisso stora.
Därav betydelsen för Portugal, som är ett av de länder där denna situation är kännbar, med tanke på prisskillnaderna mellan vårt land och Spanien: de portugisiska företagen är utsatta för konkurrens från spanska företag eftersom dessa gynnas genom lägre bränslepriser - bränslekostnaderna uppgår till 30 procent av kostnaderna - på grund av en lägre bränslebeskattning (och moms).
De portugisiska företagen har motiverat frysningen av arbetstagarnas löner med detta kostnadstryck, vilket har allvarliga konsekvenser för arbetskraften.
Europaparlamentets förslag är mer positivt eftersom det avskaffar övergångsperioderna i artikel 18, som är en mycket viktig aspekt i den aktuella situationen, med förhoppningen att det kommer att göra det möjligt att minska skillnaden mellan Portugal och Spanien senast 2010, eftersom Spanien kommer att tvingas höja sin bränsleskatt från 302 euro till 330 euro för dieselbrännolja.
Tillnärmningen kommer att fortsätta 2012 och 2015.
Vad gäller blyfri bensin kommer det tyvärr inte att ske några förändringar på detta sätt.
skriftlig. - (FR) Jag röstade emot Schmidtbetänkandet eftersom Europaparlamentet i detta sammanhang, i stället för att stödja kommissionens initiativ, har utfört ett slags trolleritrick genom att spela ut de gamla medlemsstaterna mot de nya.
Hur som helst kommer beslutet i slutändan att ligga hos enbart ministrarna och måste vara enhälligt.
skriftlig. - (FR) Högre beskattning och fler kontroller: det är Bryssels recept för Europa!
Att harmonisera punktskatter och att harmonisera momsen genom att införa bindande minimisatser som de som vi nu haft i 15 år är bevisligen ineffektivt, helt onödigt och i vissa fall till och med skadligt.
Behöver jag påminna er om att åtgärder som denna hindrar medlemsstaterna från att till exempel sänka momsen inom cateringindustrin, trots att det är en sektor där argumentet om snedvridande gränsöverskridande konkurrens är särskilt svagt och där sänkt moms skulle kunna bidra till att skapa tusentals arbetstillfällen?
Måste jag påminna er om att de nya medlemsstaterna för att följa EU-reglerna tvingas tillämpa skattehöjningar som deras befolkning uppfattar som helt skandalösa - samtidigt som de enligt andra EU-regler måste minska sin inflationstakt?
Det nuvarande förslaget är att öka skatten på dieselbrännolja i enlighet med skatten på blyfri bensin, med förevändningen att man vill skydda miljön och på grund av ett påstått behov att bekämpa ”skatteturism” - med vilket vi menar att vanliga människor drar nytta av konkurrensen!
Det är desto mer skandalöst, eftersom bilförarna i ett land som Frankrike har uppmuntrats att köpa dieseldrivna fordon - förmodligen för att vi nu ska kunna skinna dem mer än någonsin!
skriftlig. - (PT) Genom denna röstförklaring vill jag betona att vi återigen slösar bort ett tillfälle på EU-nivå - eftersom mekanismen finns - att vidta åtgärder för att skydda det småskaliga kustfisket genom att underlåta att tillämpa åtminstone samma skattevillkor för bensin som användare av dieselbrännolja åtnjuter inom jordbruket och fisket.
Vi bör komma ihåg att bensin är det bränsle som används för fartygen inom detta viktiga och största segment i de olika medlemsstaternas flottor, framför allt Portugals.
I sin resolution av den 28 september 2006 om förbättring av fiskerinäringens ekonomiska läge antog Europaparlamentet en rad förslag för att stödja sektorn så att den kan klara de höjda bränslepriserna, med tanke på att de höjda bränslepriserna har en särskilt negativ effekt på fiskerinäringen genom att avsevärt förvärra den befintliga socioekonomiska krisen och drastiskt minska yrkesfiskarnas inkomster, och eftersom det finns en allvarlig risk för att tusentals fiskeriföretag och tusentals arbetstillfällen försvinner.
Ett och ett halvt år senare har praktiskt taget ingenting gjorts på EU-nivå, förutom höjningen av de minimis-stödet.
skriftlig. - (EN) Syftet med Olle Schmidts betänkande om ”beskattningen av blyfri bensin och dieselbrännolja” är att hantera skillnaderna i fråga om bränslepunktskatterna inom unionen.
Den nuvarande obalansen har uppmuntrat till bränsleturism, vilket har ekonomiska och miljömässiga följder.
Avskräckande åtgärder måste vidtas för denna praxis.
Jag erkänner inte desto mindre behoven hos de nya medlemsstaterna, som fortfarande är inne i processen med ekonomisk utveckling och som kommer att behöva tid för att anpassa sig till de föreslagna åtgärderna.
Jag röstade för detta betänkande.
skriftlig. - (FR) Syftet med kommissionens förslag var att införa åtgärder för att minska koldioxidutsläppen i enlighet med de angivna målen i energi- och klimatförändringspaketet.
Varken i kommissionens förslag eller i det betänkande som antagits i dag tas dock upp det brådskande behovet att ta fram ett bränsle som verkligen kan gynna kampen mot koldioxidutsläppen.
Skillnaderna i de planerade anpassningarna och deras spridning, både tidsmässigt och geografiskt inom unionen, kommer att göra de föreslagna åtgärderna ineffektiva.
Om vi verkligen vill gå mot en ”era med ren luft”, borde vi vara mer miljömässigt fantasirika och stödja åtgärder som kommer att göra det möjligt för oss att hantera klimatstörningen effektivt.
Den strategi med ändrad beskattning som föreslås av kommissionen och i Schmidtbetänkandet lyckas varken främja forskningen eller det nya konceptet med ett nytt alternativt bränsle för att bromsa koldioxidutsläppen.
Jag vill i dag beslutsamt ta ställning mot tankesättet bakom detta betänkande och därför röstade jag emot vad som helt enkelt är en kompromiss som undergräver det fastställda syftet.
skriftlig. - (IT) I Gomesbetänkandet redogörs för den dramatiska och svåra situation som Irak befinner sig i.
De icke-statliga organisationerna och de olika organ som ansvarar för återuppbyggnaden av regionen lyckas i praktiken inte lösa de problem som beror på årtionden av krig, diktatur och sanktioner.
Det är i detta sammanhang EU-institutionernas plikt att stödja en mångfasetterad strategi för Irak som ökar EU:s direkta stöd för tekniskt bistånd i syfte att främja rättssäkerheten, rättvisan och en sund ekonomisk förvaltning för att skydda de grundläggande rättigheterna genom att skapa regional stabilitet och säkerhet.
Parlamentet uppmanar därför rådet att främja europeiska företags investeringar i Irak och att föra förhandlingar om handelsavtalet mellan EU och Irak så att den irakiska marknaden i högre grad kan anpassas till EU-reglerna.
I Europaparlamentets förslag, som jag instämmer i fullt ut, föreslås i huvudsak en ny strategi för Irak som innefattar en lämplig användning av Europeiska instrumentet för demokrati och mänskliga rättigheter och stöd för ett pluralistiskt och oberoende informationssystem.
Som utvecklingsutskottets föredragande för Erasmus Mundus-rapporten 2009-2013 kommer jag nu att arbeta för att öka de ekonomiska anslagen för Irak: spridningen av kultur är ett grundläggande steg mot att skapa en verklig rättssäkerhet.
skriftlig. - (PT) I den resolution som antagits lyckas man med den ”förbluffande” bedriften att inte en enda gång hänvisa till USA:s och dess allierades brutala och olagliga angrepp på och ockupation av Irak.
I resolutionen slätas hela dödssiffran på många hundratusentals irakier över, och likaså förstörelsen av ett helt land och den överlagda och omfattande kränkningen av de mänskliga rättigheterna till följd av angreppet och ockupationen.
I resolutionen sägs ingenting om det främsta skälet till de enormt allvarliga problem som Iraks folk och Irak nu står inför, och därmed om hur de ska lösas: nämligen genom det omedelbara tillbakadragandet av alla ockupationstrupper.
I resolutionen stöds i grund och botten status quo, vilket beskrivs som ett fait accompli, och man försöker att främja ett större EU-deltagande i ingripandet i Irak, vilket man betraktar som ytterligare en ”stat som övervakas” av USA/Nato/EU, som t.ex.
Afghanistan och Kosovo. Detta är förbluffande, eftersom man i resolutionen samtidigt anser att grannländerna måste avstå från att ingripa i Irak och måste respektera dess självständighet, suveränitet och territoriella integritet och det irakiska folkets önskan att bygga upp landets konstitutionella och politiska system på egen hand.
Därför röstade vi emot betänkandet.
skriftlig. - (EN) Jag röstade för detta betänkande, trots att det i ett av skälen anges att alla problem i Irak beror på den tidigare regimen.
Det råder inga tvivel om att Saddam Hussein var en brutal diktator som orsakade många av sina landsmäns död, inte minst genom det systematiska försöket att utrota kurderna.
De ockuperande styrkornas totala brist på eventuella strategier för att hantera landets återuppbyggnad har dock också lett till en oändlig misär.
Det gläder mig dock verkligen att parlamentet anser att inget land ska tvingas att återsända människor till Irak.
Landet är inte säkert, inte ens det irakiska Kurdistan, vars gräns turkiska stridsvagnar nyligen korsade, vilket orsakar ytterligare rädsla och instabilitet.
Medlemmarna i många partier i det irakiska parlamentet har talat om för oss att det är farligt att återvända och att det skulle kunna destabilisera själva landet.
I underutskottet för mänskliga rättigheter har vi också informerats om den svåra situationen för de miljontals irakier som lever som flyktingar i grannländerna med lite stöd från det internationella samfundet.
Vi borde stödja de offentliga organen i dessa stater och åtminstone utbilda barnen.
Företrädarna för Mouvement pour la France (MPF) i Europaparlamentet har intagit en konsekvent ståndpunkt sedan början av USA:s ingripande i Irak.
Vårt lands egna erfarenheter och dess band med det irakiska folket gjorde oss uppmärksamma på den mänskliga, militära och moraliska katastrof som ingripandet skulle innebära.
Nu är skadan skedd och det är upp till medlemsstaterna att agera, antingen ensamma eller kollektivt, och rädda och återupprätta vad som nu kan räddas.
Före USA:s ingripande var Irak det enda muslimska landet med ett stort och välmående kristet samfund - ett samfund som hade levt där till och med innan islam kom dit.
En av de mest tragiska konsekvenserna av USA:s ingripande har varit flykten av delar av detta samfund, vilka drivits bort på grund av terror och hotelser.
Det är en katastrof för Irak, nu och i framtiden.
Om man ser till helheten är det snabba urholkandet av en religiös befolkningsmix i Mellanöstern en mänsklig och ekonomisk utarmning som hotar hela regionens stabilitet och välstånd.
Historikern Fernand Braudel ansåg att historien började i Sumarien, men i dag tycks det som om den långa historien med de kristna minoriteterna i Irak har kommit till slutet.
Vi, Europas nationer, kan helt enkelt inte tillåta denna enorma orättvisa genom att underlåta att agera.
De irakiska kristna samfunden var en gång öppna för och välkomnade islam, och tillsammans med sina muslimska grannar byggde de ett land som blomstrade innan det härjades av fanatism och krig.
(Röstförklaringen kortades ned i enlighet med artikel 163 i arbetsordningen.)
skriftlig. - (EN) Det gläder mig att Ana Gomes i sitt betänkande om EU:s roll i Irak ser framåt och formulerar en strategi för att skapa en stabil demokratisk irakisk stat som respekterar de mänskliga rättigheterna och landets rika etniska och religiösa sammansättning.
Irak behöver Europa för att bygga vidare på de aktuella säkerhetsförbättringarna som kommer att räcka långt när det gäller att främja investeringar och öka de icke-statliga organisationernas deltagande i återuppbyggnaden av landet.
Hela Europa har ett intresse av ett stabilt och säkert Irak och jag anser att detta får stöd i betänkandets rekommendationer.
Betänkandet syftar till att garantera att EU får en större andel av det imperialistiska bytet från kriget mot Irak och ingripandena i den vidare Mellanösternregionen.
I detta sammanhang
eftersträvar man i betänkandet sätt och verktyg för att etablera en långsiktig EU-närvaro i Irak för att ”hjälpa europeiska företag att lämna in anbud på kontrakt för att återuppbygga Irak”, dvs. att öka EU-monopolens andel av bytet,
krävs i betänkandet ett villkorslöst stöd för Iraks kollaboratörs-”regering”,
läggs strategier fram för ett aktivt deltagande i den imperialistiska ockupationen.
För att de militära och polisiära styrkorna ska kunna delta i de ockuperande arméerna är allt som behövs att de bär andra huvudbeklädnader och att namnet ändras till ”FN-styrkor”.
Medan man i betänkandet cyniskt medger de katastrofala konsekvenserna av kriget och massakern på det irakiska folket, anges det kort att dessa händelser är avslutade.
Genom betänkandet legitimeras inte bara de ockuperande arméerna, som kallas en ”multinationell styrka”, utan även de privata företagen med mördare som är aktiva i Irak, under förutsättning att regler ställs upp för deras brottsliga verksamhet!
Greklands kommunistparti fördömer betänkandet.
Kommunistpartiet framför sin solidaritet med irakiernas motstånd och med folket i regionens kamp för att bli fria från det imperialistiska oket och för sin okränkbara rättighet att bestämma över sitt eget öde.
skriftlig. - (PT) Det faktum att parlamentet har beslutat att diskutera Europeiska unionens roll i Irak, snarare än att insistera på en meningslös debatt om tidigare frågor, är positivt.
De fem år som nu har betydelse för oss är de kommande fem åren snarare än de gångna.
Utgångspunkten för alla debatter om denna fråga måste nu vara att erkänna att situationen på plats har förbättrats avsevärt, även om den fortfarande är mycket allvarlig.
Vad denna förbättring i synnerhet visar på är att det finns en gångbar väg framåt i form av målet att bygga en demokratisk och säker stat.
Vårt mål kan nås.
Erfarenheterna under de senaste åren visar dock också att målet endast kommer att nås genom ett större engagemang, genom ökad säkerhet, genom att investera i utbildning för de irakiska myndigheterna och genom att aktivt bidra till skapandet av infrastruktur som kommer att göra landets ekonomi livkraftig, vid sidan av oljan, vilket är mycket viktigt.
I Europeiska unionens särskilda fall innebär detta stora investeringar i den ekonomiska återuppbyggnaden av Irak och i skapandet av demokrati i landet.
Ett demokratiskt och säkert Irak som respekterar de mänskliga rättigheterna är av avgörande vikt för regionen och för världen.
skriftlig. - (DE) Jag vet såklart att vi röstade i kammaren om förslaget till betänkande från min kollega Ana Gomes om Europeiska unionens roll och inte om hennes motivering till betänkandet.
Men jag tycker ändå att det är viktigt att föredraganden i sin motivering återigen betonar att invasionen av Irak var en strategisk och humanitär katastrof och att det irakiska samhället återigen traumatiserades av kriget och det åtföljande kaoset och våldet.
Jag välkomnar att föredraganden, utöver alla sina övriga viktiga punkter, uttryckligen konstaterar att kvinnorna måste få en starkare roll och att respekten för kvinnors, minoriteters och barns rättigheter måste främjas om ett gott arbete ska kunna utföras i Irak.
skriftlig. - (NL) Jag beklagar att Europaparlamentet hittills inte har gjort någon som helst analys av kriget i Irak.
Parlamentet har under senare år faktiskt upprätthållit en bedövande tystnad och har inte ens utmanat Bushregeringens lögner.
För ett demokratiskt organ som parlamentet spelar detta stor roll!
Det blir svårt för oss att bevara vår trovärdighet om vi inte ens vidtar åtgärder mot FN-medlemmar som struntar i FN-stadgan.
Ana Gomes gör en bedömning av situationen i Irak.
Hennes betänkande om Europeiska unionens roll i Irak innehåller ett antal goda rekommendationer om hur landet bör återuppbyggas.
I betänkandet behandlas en rad ämnen och jag uppfattar alla föreslagna åtgärder som genomförbara.
Jag välkomnar särskilt förslagen till multilaterala insatser, under FN:s överinseende, för att inleda intensiva diplomatiska samtal mellan USA och Iraks grannländer.
Syftet måste vara att upprätta demokrati i Irak, utifrån principerna med rättssäkerhet, goda styrelseformer och mänskliga rättigheter.
Jag stöder därför betänkandet.
, skriftlig. - (FR) I fjärde Genèvekonventionen angående skydd för civilpersoner under krigstid anges att humanitär, medicinsk och religiös personal ska respekteras och skyddas.
Det är mycket viktigt att vi stöder fallet med Monsignor Paulos Faraj Rahho, den kaldeiska katolska ärkebiskopen som föddes och bor i Mosul, som kidnappades fredagen den 9 februari 2008.
De tre personer som var med honom vid hans bortförande dödades av kidnapparna.
Det var i ett muntligt ändringsförslag till Gomesbetänkandet inte möjligt att nämna Monsignor Rahho vid namn.
Därför vill jag be talmannen att uttryckligen sända två brev med parlamentets stöd och uppmuntran:
Ett till Iraks shiitiska premiärminister Nouri al-Maliki, som har fördömt attackerna på kristna präster och som på den irakiska regeringens vägnar har erbjudit ”skydd och rättvisa” för kristna, med en försäkran om att de som är ansvariga för våldet ska tas fast och straffas.
Det andra till Iraks vice president Tareq al-Hashemi, som är medlem av sunnisamfundet, som också har fördömt terroristattackerna på kristna samfund klart och tydligt och som efter kidnappningen framförde sin solidaritet med vad han kallade sina ”kristna bröder”.
Det är av avgörande vikt att vi uppmuntrar de nationella myndigheterna att göra allt de kan för att garantera att Monsignor Paulos Faraj Rahho friges omedelbart och ovillkorligt.
skriftlig. - (EN) Jag kommer att stödja denna resolution.
Som jag sa i mitt betänkande för över tio år sedan är det grundläggande att vi har en bindande rättslig grund för vår uppförandekod för vapenexport.
Ändå drivs nödvändigheten att exportera av en splittrad europeisk industri som gärna vill ha en lång produktion så att de kan konkurrera med massproducerade vapen från USA med en inhemsk efterfrågan på endast serieproduktion.
Därför behöver vi en inre marknad för försvarsutrustning som kan göra det möjligt för EU att först och främst konkurrera, för det andra att upphöra med att ge näring åt regionala krig världen över och för det tredje att föra in några av sina mest kvalificerade vetenskapsmän och ingenjörer i morgondagens avancerade teknikindustri.
skriftlig. - Vissa medlemsstater har starka egenintressen för att främja en ökad vapenexport.
Vid ett skapande av en gemensam uppförandekod för vapenexport är det därför troligt att vissa medlemsstater med en mer restriktiv policy kan komma att tvingas till att kompromissa.
Vi är av den uppfattningen att övervakningen av vapenexport ska skötas av respektive medlemsland genom landets nationella lagstiftning.
Sverige ska ha fortsatt rätt att kunna bedriva en restriktiv vapenexport om så önskas.
Ett samarbete är önskvärt för att driva på det globala nedrustningsarbetet, men detta sker bäst internationellt, inom Förenta nationernas ram, med tanke på FN:s erfarenhet, kunskap och globala räckvidd.
skriftlig. - (PT) En verkningsfull EU-uppförandekod för vapenexport blir tveklöst allt mer viktigt i sammanhanget med EU:s snabba militarisering, som återspeglas i utkastet till fördrag som nu ratificeras i varje medlemsstat.
Det är inte utan viss ironi som det i själva resolutionen specifikt hänvisas till att ”utvecklingen av den europeiska säkerhets- och försvarspolitiken (ESFP) har gjort att EU genomför allt fler militära och civila uppdrag ... och att EU-anställda i samband därmed kan hotas med vapen som tidigare har levererats av EU:s medlemsstater”.
”Marknaden för militär utrustning” växer inom EU, ”flera initiativ ... för att harmonisera nationella upphandlingsregler avseende vapen samt vapenöverföring och vapenförsäljning inom gemenskapen” uppmuntras och det finns ”en vilja att öka vapenexporten för att främja ekonomiska intressen”.
Lösenordet har fastställts: kapprustning och militarisering av de internationella förbindelserna.
Initiativ och åtgärder för att åtminstone mildra en sådan upptrappning är därför positivt och nödvändigt.
Liksom vi tidigare angav kommer dock regleringen av vapenhandeln att få mycket större betydelse om den åtföljs av en process med multilateral och ömsesidig nedrustning, som i synnerhet borde börja med nedrustningen av de enorma kärnvapenarsenalerna.
skriftlig. - (EN) Den brittiska konservativa delegationen röstade emot resolutionen eftersom den inte accepterar hänvisningarna till Lissabonfördraget eller till utvecklingen av den europeiska säkerhets- och försvarspolitiken, som den motsätter sig.
Vidare är den brittiska konservativa delegationen, trots att den starkt förespråkar en ansvarstagande politik för vapenöverföring, inte övertygad om förtjänsterna med en rättsligt bindande uppförandekod som påförs av EU före antagandet av ett internationellt bindande vapenhandelsfördrag.
skriftlig. - Vi svenska socialdemokrater röstade för betänkandet, då det är viktigt att fängelseförhållandena förbättras på vissa anstalter i Europa och fångars mänskliga och grundläggande rättigheter respekteras.
Dessutom måste ett jämställdhetsperspektiv integreras i kriminalvården och på fängelserna.
Vi har dock vissa invändningar mot delar av innehållet i betänkandet.
Vi önskar inte en harmonisering av fängelseförhållandena i Europa, och vi ifrågasätter starkt skrivningarna i betänkandet om särskilda brottspåföljder eller alternativa straff för kvinnor, gravida kvinnor och kvinnor som lever med små barn.
Vad gäller barnets kontakt med föräldrarna under fängelsevistelsen och tiden därefter måste det, med barnets bästa i fokus, gälla båda föräldrarna och inte bara mamman eller den ena föräldern.
skriftlig. - (EN) Jag och mina konservativa kolleger anser att man alltid bör fundera över hur man kan förbättra situationen för kvinnor i fängelse.
I betänkandet föreslås ett antal möjligheter som kan undersökas vidare, däribland tillhandahållandet av hälsotjänster.
Betänkandet är dock överdrivet preskriptivt när det gäller vad medlemsstaterna bör göra på detta område.
Det är upp till medlemsstaterna att besluta om detaljerna för fängelsepolitiken.
Vi kan i synnerhet inte hålla med om antagandet i skälen C och Q, som vi anser snedvrider andra aspekter av betänkandet som kan vara av värde.
Därför har vi beslutat att lägga ned våra röster.
skriftlig. - (PT) Jag röstade för Marie Panayotopoulos-Cassiotous betänkande om kvinnors speciella situation i fängelser och hur det sociala livet och familjelivet påverkas av att föräldrar sitter fängslade, eftersom det finns bevis för att de europeiska fängelserna i hög grad är anpassade till manliga fångar och bortser från kvinnors särskilda behov.
Jag anser därför att åtgärder bör vidtas för att möjliggöra en förbättring av situationen för kvinnor i fängelse, särskilt i fråga om deras sociala och yrkesmässiga återintegrering, hälsovård och hygien, psykologiska stöd och bevarandet av familjeband.
skriftlig. - (PT) Även om kvinnor utgör ca 4,5 till 5 procent av fångarna i Europeiska unionen fortsätter fängelserna att i grunden vara anpassade till manliga fångar och man tenderar att bortse från det specifika problemet med den begränsade men växande andelen kvinnliga fångar.
De viktigaste områdena är hälsovård, situationen för fängslade kvinnor med barn och yrkesmässig och social återintegrering.
Särskild uppmärksamhet bör riktas på kvinnors hälsovård och hygienbehov.
I synnerhet gravida kvinnor i fängelse kräver specialiserade resurser och särskild uppmärksamhet när det gäller kosthållning, träning, kläder, läkemedel och läkarvård av specialiserad personal.
Barn som vårdas av sina fängslade mödrar behöver lämpligt skydd och lämplig omvårdnad och får inte utsättas för någon typ av diskriminering.
Fängelsestraff för kvinnor har särskilt allvarliga följder när de har varit den enda vårdnadshavaren för barn före fängslandet.
Den sociala integrationen av fångar måste förberedas under och efter fängelsestraffet i samarbete med socialtjänsten och andra relevanta organisationer för att garantera en smidig övergång från fängelse till frihet.
skriftlig. - Vi stöder det arbete som görs i medlemsländerna för att modernisera och anpassa kriminalvårdspolitiken för att bättre tillgodose fångars behov, och som ett led i detta ta hänsyn till kvinnors specifika behov.
Eftersom kriminalvård inte är en EU-kompetens har vi valt att rösta emot betänkandet.
Åtgärder som rör besöksregler, drift av anstalterna, utbildning för anställda i kriminalvården, fångarnas fritidsaktiviteter eller sociala stödåtgärder är och bör förbli medlemsstaternas kompetens för att kunna anpassas och utvecklas efter nationella och lokala behov.
skriftlig. - Vi stödjer det arbete som görs i medlemsländerna för att modernisera och anpassa kriminalvårdspolitiken i syfte att bättre tillgodose fångars behov, och som ett led i detta ta hänsyn till kvinnors specifika behov.
Eftersom kriminalvård inte är en EU-kompetens har vi valt att rösta emot betänkandet.
Åtgärder som rör besöksregler, drift av anstalterna, utbildning för anställda i kriminalvården, fångarnas fritidsaktiviteter eller sociala stödåtgärder är och bör förbli under medlemsstaternas kompetens för att kunna anpassas och utvecklas efter nationella och lokala behov.
skriftlig. - (EN) Jag instämmer i slutsatserna i Marie Panayotopoulos-Cassiotous betänkande om kvinnors speciella situation i fängelser och hur det sociala livet och familjelivet påverkas av att föräldrar sitter fängslade.
Fängelserna är fortfarande anpassade till manliga fångars behov och jag välkomnar betänkandets syfte att lyfta fram de skillnader som kvinnor upplever.
Jag stöder betänkandet.
skriftlig. - (FR) Jag röstade för betänkandet, eftersom det finns ett stort behov av att anpassa förhållandena i fängelserna efter kvinnornas särskilda behov.
Förhållandena i fängelserna i många medlemsstater är fortfarande i dag mycket dåliga och kan verkligen inte ge det speciella stöd som kvinnor behöver.
Kvinnliga fångar har särskilda problem som kräver särskild uppmärksamhet. Framför allt gäller det tillgången på hälsovård.
Därför stöder jag socialistgruppens ändringsförslag med krav på att kvinnliga fångar ska få samma tillgång till screening för bröstcancer och livmoderhalscancer som andra kvinnor.
En tidig diagnos av dessa sjukdomar förbättrar möjligheterna att bota dem. Att vägra kvinnliga fångar tillgång till sådana screeningprogram kan i själva verket innebära ett ytterligare straff.
Kvinnorna är dessutom fortfarande centrala för familjen.
För mödrar bör vi därför om det går försöka underlätta andra påföljder än fängelse under förutsättning att de inte innebär något hot mot den allmänna ordningen.
skriftlig. - Detta är ett område för vilket det inte finns någon kompetens på EU-nivå.
Trots positiva förslag är betänkandet alltför detaljreglerat.
Därför lägger jag ned min röst.
skriftlig. - (EN) När vi röstar om en politik som omfattar ”sexuell och reproduktiv hälsa” så tolkar vi det så, att det innebär att skydda och stärka moderns och det ofödda barnets liv och hälsa.
Vi accepterar inte någon annan definition som antyder att abort skulle inrymmas i det begreppet. Dessutom anser vi att all vård, information, politik eller andra tjänster som ingår i begreppet sexuell och reproduktiv hälsa på samma sätt utesluter abort.
Vi kommer att arbeta på att få denna definition accepterad i alla forum och organ vi kan påverka.
Vi konstaterar att svaret som rådets ordförandeskap gav i parlamentet den 4 december 2003 inte innebar att begreppet reproduktiv hälsa inkluderar ett främjande av abort. Abort får till exempel aldrig framställas som en metod för familjeplanering, i motsats till vad Världshälsoorganisationen säger om fertilitetskontroll.
Det står därför klart att WHO:s definition inte är bindande för eller ens accepterad av statliga och parlamentariska institutioner.
Vi kommer att fortsätta stödja politiska program som främjar ansvarsfulla sexuella beteenden och som skyddar och främjar moderns och det ofödda barnets liv och hälsa, inklusive att tillhandahålla resurser för att uppnå dessa mål.
skriftlig. - Initiativbetänkandet syftar till att integrera jämställdhetsperspektivet i EU:s utvecklingssamarbete.
Junilistan är emot bistånd på EU-nivå och röstar därför nej till betänkandet.
Däremot är flera av de ändringsförslag som har lagts fram av vissa ledamöter av mindre sympatisk karaktär.
Kvinnors rätt till sexuell och reproduktiv hälsa är en viktig komponent för att skapa utveckling.
I detta fall har vi valt att stödja ursprungsförslagen som en motkraft till de olustiga strömningarna i detta parlament.
Arbetet för dessa frågor och utvecklingssamarbete bör dock principiellt ske på den globala nivån genom FN, och inte EU.
skriftlig. - (PT) Vi anser att det här betänkandet har flera förtjänster. En av dem är att det riktar uppmärksamheten på ett stort problem, både i EU och i utvecklingsländerna, nämligen behovet av att garantera tillgången på information om sexuell och reproduktiv hälsa, möjligheten att fritt fatta beslut och att skapa och främja offentliga tjänster som skyddar och tillämpar allas rättigheter, framför allt kvinnornas.
Vi tycker emellertid att man måste understryka att det viktigaste bidraget till ”jämställdhet och ökat medinflytande för kvinnor i utvecklingssamarbete” inte kommer från en politik som bygger på beroende och dominans, avreglering av marknader (se EU:s ekonomiska partnerskapsavtal), utnyttjande av arbetare, ojämlikhet och sociala orättvisor och bristande respekt för mänskliga rättigheter och som framför allt drabbar miljontals och åter miljontals barn och kvinnor.
skriftlig. - (EN) Jag röstade för ändringsförslaget, eftersom jag är fast övertygad om att kampen mot våld, i detta fallet våld mot kvinnor i kris- och konfliktområden, måste få högsta prioritet.
EU kan inte tolerera någon form av våld och därför anser jag att tyngdpunkten bör ligga på att bekämpa sexuellt våld riktat mot kvinnor.
Dessutom anser jag att traditioner inte ska betraktas som något ont.
Sexuell och reproduktiv hälsa och rättigheter är känsliga frågor med både sociala och religiösa dimensioner. Därför får man inte generalisera eller tvinga på samhället några lösningar, framför allt inte ömtåliga samhällen där drastiska förändringar av den traditionella livsstilen kan stjälpa, snarare än hjälpa.
skriftlig. - (DE) Jag röstar för jämlikhet mellan kvinnor och män och för att ge kvinnorna en starkare ställning i utvecklingssamarbetet.
Det sätt på vilket kvinnor i utvecklingsländerna hålls nere av religiösa regler, kulturella rutiner och fattigdom förvärras ofta ytterligare av bristen på utbildning.
I det sammanhanget vill jag särskilt rikta uppmärksamheten på det potentiellt enorma sociala tryck som kan uppkomma om man ökar allmänhetens kunskaper om kvinnornas grundläggande rättigheter. I slutändan skulle detta kunna förbättra kvinnornas situation i de berörda regionerna.
Jag stöder dessutom idén att betrakta ”våld mot kvinnor” inte enbart utifrån de kvinnliga offrens synvinkel. Snarare bör man utveckla praktiskt tillämpbara program som riktar sig till ”den manlige missbrukaren”, så som Feleknas Uca föreslår i sitt betänkande.
Jag är också mycket kritisk mot kommissionens underlåtenhet att inkludera en strategi mot kulturellt eller religiöst våld mot kvinnor i förteckningen över åtgärder.
Dålig tillgång på utbildning skapar handikapp inom andra områden i livet av den enkla anledningen att man har brist på information.
Att vara dåligt informerad i detta avseende kan få dödliga konsekvenser i utvecklingsländer där tillgången på hälsovård och den hygieniska standarden många gånger är under all kritik.
Jag behöver bara nämna den oroväckande höga andelen hiv-infekterade kvinnor - söder om Sahara är den siffran 57 procent.
En mycket positiv punkt är kravet på att utveckla ”könsuppdelade resultatindikatorer”, vilket också skulle göra den kontroversiella frågan om kvotering mindre laddad.
skriftlig. - (EN) När vi röstar om en politik som omfattar ”sexuell och reproduktiv hälsa” så tolkar jag det så, att det innebär att skydda och förbättra moderns och det ofödda barnets liv och hälsa.
Vi accepterar inte någon definition som antyder att abort skulle inrymmas i det begreppet. Och dessutom anser vi att all vård, information, politik eller andra tjänster som ingår i begreppet sexuell och reproduktiv hälsa på samma sätt utesluter abort.
Vi måste arbeta på att få denna definition accepterad i alla forum och organ vi kan påverka
Jag konstaterar att svaret som rådets ordförandeskap gav i parlamentet den 4 december 2003 inte innebär att begreppet reproduktiv hälsa inkluderar ett främjande av abort och att abort till exempel aldrig får framställas som en metod för familjeplanering, i motsats till vad Världshälsoorganisationen säger om fertilitetskontroll.
Det står därför klart att WHO:s definition inte är bindande för eller ens accepterad av statliga och parlamentariska institutioner
Jag kommer att fortsätta stödja politiska program som främjar ansvarsfulla sexuella beteenden och som skyddar och främjar moderns och det ofödda barnets liv och hälsa, inklusive att tillhandahålla resurser för att uppnå dessa mål.
skriftlig. - (EN) I sitt betänkande ”Jämställdhet och ökat medinflytande för kvinnor i utvecklingssamarbetet” välkomnar Feleknas Ucas kommissionens strategi i frågan.
Jag upprepar hennes stöd för en strategi som försöker integrera jämlikhet mellan kvinnor och män i utvecklingssamarbetet.
Jag röstade för betänkandet.
skriftlig. - (FR) Även om jämlikhet mellan kvinnor och män har varit en integrerad del av Europeiska unionens program för utvecklingssamarbete under flera år, så är de faktiska framstegen fortfarande för obetydliga.
Europeiska kommissionen måste därför bestämma mål i termer av siffror och tidsfrister, så att utveckling kan bli en viktig pådrivande faktor för förbättrade levnadsförhållanden för kvinnor.
Därför måste unionen fokusera på tre prioriteringar i sina partnerskap: grundläggande friheter, kvinnors status i det offentliga livet och deras tillgång på hälsovård.
Å ena sidan måste kommissionen vara vaksammare än någonsin tidigare när det gäller våld mot kvinnors fysiska integritet och mänskliga värdighet (i form av tortyr, traditionella former av stympning och tvångsäktenskap).
Å andra sidan måste samarbetet omfatta ett erkännande av kvinnans plats i samhället, vilket påverkar allt från tillgången på kunskap till ekonomiskt oberoende.
Dessutom krävs det insatser så att förebyggande och behandling av aids i utvecklingsländerna blir en realitet till 2010.
Den europeiska utvecklingspolitiken kommer att bli ett totalfiasko om den inte kan radikalt förändra kvinnornas villkor.
Trots betänkandets korrekta slutsatser om kvinnornas tragiska ställning i utvecklingsländerna döljer det själva orsaken till detta: kapitalistiska produktionsmetoder och brutala imperialistiska ingrepp från EU, Förenta staterna och andra imperialiststater och organisationer.
De suger ut dessa länder och plundrar deras källor till välstånd, vilket resulterar i hunger och fattigdom för miljontals människor.
De lösningar som föreslås ligger inom ramen för en kapitalistisk utveckling och EU:s utvecklingsstöd.
En annan typisk aspekt av denna strategi är förslaget att öka antalet kvinnliga egenföretagare för att öka sysselsättningen.
I det sammanhanget är förslagen om rättvisare och mer demokratiska samhällen, flickors och kvinnors tillgång till utbildning och hälsovård, utrotandet av fattigdom och sjukdomar etc. bara tomt prat.
Det är fromma önskningar som avleder uppmärksamheten från sanningen. Att uppfylla människors behov är nämligen oförenligt med kapitalistisk utveckling och strävan efter profit som överordnad princip.
För varje euro som Europeiska unionen ger, så stjäl den tusentals från dessa länder.
En förbättring av kvinnornas ställning och befolkningens levnadsstandard i dessa länder kommer inte att uppnås genom den legaliserade stöld som kallas ”EU:s utvecklingsstöd”, utan genom motstånd mot imperialistisk intervenering, strävan efter jämlika internationella relationer och kamp för en annan utvecklingsstrategi, baserad på befolkningens behov.
skriftlig. - (DE) Betänkandet om jämlikhet och deltagande, om kvinnors roll i utvecklingssamarbetet, täcker ett stort antal olika aspekter och inkluderar också viktiga praktiska frågor.
Som helhet bör det med andra ord absolut få stöd.
En fråga som löper genom hela betänkandet är sexuell och reproduktiv hälsa och våld mot kvinnor, jämte främjandet av kvinnors rätt till självbestämmande.
Det är viktigt att utöka nätverken för mikrofinansiering, eftersom mikrokrediter kan bidra till att förbättra kvinnornas ekonomiska situation.
Jag kan inte förstå varför vissa försöker lägga fram olika ändringsförslag som försvagar betänkandet och helt enkelt bortser från de dokument från FN som finns tillgängliga.
skriftlig. - (PL) Feleknas Ucas betänkande om jämställdhet i utvecklingspolitiken är ett uttryck för europeisk moralisk imperialism gentemot utvecklingsländerna.
Den går ut på att exportera de rika europeiska ländernas sjuka sociala modell till länderna i Afrika och Asien.
De upprepade hänvisningarna till reproduktiva rättigheter betecknar stöd för allmänt tillgänglig abort.
Jag kunde därför inte rösta för betänkandet.
skriftlig. - (FR) Jämlikhet mellan kvinnor och män är en prioriterad fråga i utvecklingsländerna.
Jag uppskattar verkligen Feleknas Ucas grundliga och grannlaga arbete med denna viktiga fråga.
Trots detta röstade jag emot betänkandet, eftersom innehållet i vissa avsnitt i slutversionen, som behandlade sexuell och reproduktiv hälsa på ett oklart sätt, fortfarande är tvetydigt.
Det finns motstridiga tolkningar och några av dem innebär ett hot mot ofödda barns liv.
I nästa betänkande i ämnet bör kvinnors hälsa inte enbart sättas i relation till reproduktion, för alla kvinnor har rätt till en miljö som ger dem möjlighet att njuta fortsatt god hälsa.
Det innebär att man måste ägna särskild uppmärksamhet åt tillgången på säkert dricksvatten, proteiner och basläkemedel, vid sidan om traditionella läkemedel.
Mot bakgrund av Gertrude Mongellas besök den 6 mars 2008 för att uppmärksamma Internationella kvinnodagen vill jag också säga att vi har mycket att lära av afrikansk visdom när det gäller jämlikhet mellan kvinnor och män. Detta är en fråga som upplevs starkt där och något som förs vidare genom muntlig tradition bland kvinnor och män som är välsignade med god andlig och mental hälsa.
Där har vi alla något att lära.
2.
Gripande av demonstranter efter presidentvalet i Ryssland (omröstning)
- Före omröstningen:
författare, för UEN-gruppen. - (PL) Jag föreslår en stilistisk ändring.
Orden ”Europeiska domstolen” bör ändras till ”Europeiska domstolen för mänskliga rättigheter”, annars blir texten obegriplig.
(Det muntliga ändringsförslaget beaktades.)
Begäran om upphävande av parlamentarisk immunitet: se protokollet
Avbrytande av sessionen
Jag förklarar Europaparlamentets session avbruten.
(Sammanträdet avslutades kl. 12.20.)
De internationella finansiella redovisningsstandarderna (IFRS) och styrningen av International Accounting Standards Board (IASB) (debatt)
Nästa punkt är ett betänkande av Alexander Radwan, för utskottet för ekonomi och valutafrågor, om internationella redovisningsstandarder (IFRS) och styrningen av (IASB)
föredragande. - (DE) Fru talman! Ämnet för det betänkande vi har framför oss kan vid första anblicken verka mycket tekniskt.
Det handlar om så kallade redovisningsstandarder inom Europeiska unionen och över hela världen, i synnerhet för små och medelstora företag.
Det kan mycket väl vara en typ av ämne som just nu diskuteras i Europaparlamentet men som inte börjar påverka ekonomin eller vanliga människor förrän efter flera år.
Vid det laget höjs röster om att ingen vet varifrån dessa standarder kommer eller vem som bär ansvaret för dem.
Inte heller kommer någon att veta varför de ska tillämpas.
Ändamålet är att nå en enda uppsättning av globala redovisningsstandarder, i synnerhet för aktiebolag.
Vi stöder det syftet.
Det argument som framläggs för detta är att vi behöver ”standarder av hög kvalitet”, och parlamentet anser sig vara det enda forum som är bemyndigat att fastställa dessa högkvalitativa standarder.
Under dessa tider av turbulens på finansmarknaderna är det förvånande att höra att samma personer som tidigare argumenterat för principen om ”verkligt värde” nu ifrågasätter denna princip och dessutom frågar sig om en ”marknad till marknads-strategi" fortfarande är meningsfull om vi inte längre har någon marknad.
Samma personer som släppte anden ur flaskan är de som nu frågar om vi är på rätt spår.
De enda som ansvarar för dessa standarder är de som arbetar på den här privata organisationens kontor i London, som utan tvivel påverkas av önskan att behålla sitt arbete när de utarbetar sina standarder.
Mitt betänkande, som vi ska rösta om idag, rör därför inte bara hur små och medelstora företag påverkas utan också den grundläggande frågan om vilka som gör upp regler för vem, och vem som övervakar reglernas tillämpning.
Den första frågan vi ska ta itu med är styrningen: hur insynsvänlig är organisationen?
Med andra ord hur insynsvänlig är dess finansiering?
Här finns säkert dolda intressen.
Ledamöterna i detta utskott, som kräver öppenhet och alltid försöker ge en bild av marknaden som insynsvänlig, bör anstränga sig åtminstone en smula för att följa de krav på öppenhet som de fastställer för marknaden!
Mitt intryck så här långt är att denna organisation kämpar med alla tillgängliga medel för att undvika öppenhet i alla former.
Vem fattar besluten om finansiering och väljer ut personal för specifika befattningar?
Varför utnämns dessa personer?
Handlar det om regional balans?
Handlar det om balans mellan sektorerna?
Det aktuella projektet gäller internationella redovisningsstandarder (IFRS) för små och medelstora företag, och det är därför rimligt att fråga vem som representerar de små och medelstora företagen.
Vem vet något om små och medelstora företag?
Och en sak till: varför har internationella redovisningsstandarder för små och medelstora företag kommit upp på dagordningen just nu?
Vem fastställer dagordningen?
Kommissionsledamot Charlie McCreevy and Sir David Tweedie har också många gånger under flera år fått svara på frågan om varför vi egentligen sysslar med detta.
Flera år efteråt vet vi nu varför vi diskuterar internationella redovisningsstandarder för små och medelstora företag i Europa: det är på begäran av Sydafrika och Brasilien.
Vilket underbart svar!
Vi vet mycket väl att fokus här inte ligger på Sydafrika eller Brasilien, utan istället på den europeiska marknaden, där det finns mycket pengar att tjäna om de små och medelstora företagen åläggs att införa något sådant.
Det här är alltså de viktigaste frågorna när det gäller styrning - och några inledande, positiva steg har tagits.
Men alla de organ som ska inrättas i framtiden kommer att bedömas beroende på huruvida de personer som tillhör denna tillsynsorganisation och måste svara på frågor om den på politisk nivå - och det kan vara en kommissionsledamot - också kommer att få makt att utforma nya utvecklingar.
Det är inte tillräckligt för dem att bara bli underrättade om förslag.
Ett av våra syften är konvergens.
Men vi måste se upp så att tolkningen av konvergensbegreppet inte går Europa ur händerna och ersätts av den tolkning som görs av den amerikanska finansinspektionen Securities and Exchange Commission.
I Europa är vi numera ganska väl införstådda med hur den amerikanska fondbörsen kontrolleras.
Vi får inte vara så naiva att vi överlåter kontrollverksamheten till amerikanerna.
Vad vi vill ha är därför det som vi redan har begärt: internationella redovisningsstandarder ur Europas synvinkel och inte så som denna styrelse föreskriver.
Det är de små och medelstora företagen som påverkas här och, utan att skräda orden måste jag säga att de idéer som vi har framför oss idag är alltför komplicerade och svåra.
Jag vill också varna för den frivilliga vägen.
Idag har jag på mig den bayerska nationaldräkten och ett gammalt bayerskt uttryck dyker upp i mitt huvud: det är ”hinterfotzig” och det betyder nåt i stil med ”bakvägen”.
Trots förnekanden och tysta medgivanden vet vi mycket väl att internationella redovisningsstandarder för små och medelstora företag kommer att införas på EU-marknaden bakvägen, via ett litet antal medlemsstater.
Då kommer samma röster att efterlysa en enda uppsättning standarder och de kommer att fortsätta att smussla in sina standarder på marknaden - standarder som är alltför komplicerade, som ingen förstår och som ingen vill ha - bara för att det finns en marknadsmöjlighet.
Det här är ett fall där en minoritet försöker tvinga sin vilja på en majoritet på global nivå, och det är oacceptabelt!
ledamot av kommissionen. - (EN) Fru talman! Jag vill tacka utskottet för ekonomi och valutafrågor, i synnerhet föredraganden Alexander Radwan, för det ansenliga arbete som lagts ner på detta innehållsrika betänkande.
Betänkandet omfattar viktiga frågor som rör den framtida utvecklingen av de europeiska och framför allt de globala kapitalmarknaderna.
I detta korta inlägg kan jag inte beröra alla de frågor som tas upp i betänkandet.
Jag vill därför koncentrera mig på tre punkter.
För det första, frågor om styrning, för det andra EU:s bidrag till International Accounting Standards Board, IASB, och för det tredje projektet att utveckla en redovisningsstandard för små och mellanstora företag.
När det gäller styrningen av IASB belyser betänkandet mycket riktigt det faktum att vårt gemensamma mål är att utveckla högkvalitativa globala redovisningsstandarder.
EU-beslutet att börsnoterade bolag måste använda internationella redovisningsstandarder var ett djärvt och visionärt steg mot det målet.
En uppsättning globalt accepterade redovisningsstandarder skulle vara till stor nytta för våra företag, våra kapitalmarknader och vår ekonomi.
Vi måste arbeta kontinuerligt med att se till att de internationella redovisningsstandarderna förblir relevanta gentemot de föränderliga ekonomiska omständigheterna och att de på ett balanserat sätt representerar alla aktörers intressen.
För att säkerställa att dessa villkor uppfylls fortsättningsvis bör framsteg prioriteras på tre områden.
För det första måste redovisningsskyldigheten hos International Accounting Standards Committee Foundation (IASC Foundation) förbättras, i synnerhet mot offentliga myndigheter.
De senare bör spela en aktiv roll vid val och utnämning av styrelseledamöter.
I detta avseende går det förslag som jag, tillsammans med mina motparter i USA:s Securities and Exchange Commission, den japanska finansinspektionen och den internationella organisationen av institutioner för reglering av värdepappersmarknader, IOSCO, lade fram i november, i samma riktning som förespråkas i betänkandet.
För det andra måste vi se på hur processen för att fastställa IASB:s dagordning kan förbättras.
Processem för att fastställa prioriteringar måste således bli öppnare och tydligare.
För det tredje bör IASB:s samrådsförfarande (due process) förbättras, huvudsakligen genom att se till att standarderna genomgår en fullständig konsekvensanalys innan de antas.
I betänkandet finns konstruktiva förslag beträffande dessa och närbesläktade punkter.
Under den kommande översynen av IASCF:s konstitution finns det tillfälle att genomföra de nödvändiga reformerna.
Utskottet kommer att följa upp dem i samråd med parlamentet, medlemsstaterna och våra internationella partner.
Nu till EU:s bidrag till IASB.
I betänkandet hävdas att EU måste stärka sin förmåga att göra sina synpunkter på redovisningsfrågor hörda på internationell nivå.
Jag instämmer.
Vi bör närmare bestämt finna metoder för att se till att synpunkter från europeiska aktörer, särskilt proaktiva bidrag till IASB:s förfarande för att fastställa dagordningen IASB, kan framföras till IASB på ett mer lämpligt och enhetligt sätt.
Jag ser det här som en utvecklingsprocess och inte som en revolutionär process.
Vi bör utgå från European Financial Reporting Advisory Group (EFRAG) och jag är beredd att ägna mig åt denna brådskande fråga, inklusive möjligheten att använda finansiering från gemenskapens budget för att stödja en sådan struktur.
Jag måste dock komma med en klar och tydlig varning.
Den här strukturen kommer under inga omständigheter att utvecklas till ett förstadium till europeisk normgivare, och det är inte heller fråga om att utveckla europeiska tolkningar av internationella redovisningsstandarder.
Europa måste och kommer att förbli en del av den rörelse som verkar för en enda uppsättning med internationellt accepterade redovisningsstandarder.
Allt annat skulle skada den internationella konkurrenskraften hos våra företag och vår kapitalmarknad.
Jag går vidare till IASB:s förslag om att utarbeta en redovisningsstandard för små och medelstora företag, och vill börja med att konstatera att kommissionen för närvarande inte har någon rättslig grund för denna standard.
Vi har heller aldrig gjort någon utfästelse om att ta över någon som helst standard som IASB utarbetar.
Vi skulle göra det endast om vi var verkligt övertygade om att IASB utarbetar en standard som motsvarar de europeiska användarnas intressen.
IASB har ännu inte slutfört sitt projekt.
Kommissionens synpunkter i detta skede är emellertid tydliga.
Det aktuella utkastet som publicerats av IASB är fortfarande för komplicerat för att bilda en nöjaktig redovisningsram för europeiska små och medelstora företag, särskilt de små företagen.
Vårt fokus förblir att förenkl lagstiftningen för små och medelstora företag, också inom redovisningsområdet.
föredragande för yttrandet från utskottet för rättsliga frågor. - (DE) Fru talman, mina damer och herrar! Systemet med internationella redovisningsstandarder är meningsfullt för stora börsnoterade företag med världsomspännande verksamhet.
Det var därför vi beslöt att anta IAS-förordningen under parlamentets senaste mandatperiod, på förslag av utskottet för rättsliga frågor.
Det slutgiltiga målet - liksom Alexander Radwan redan sagt - var att uppnå konvergens, åtminstone med USA och om möjligt i hela världen.
Systemet är meningslöst om det är fråga om små och medelstora företag, eftersom de för det mesta inte har behov av internationella finansmarknader, Wall Street och så vidare.
Bara av den orsaken kan behovet av att utveckla internationella redovisningsstandarder för små och medelstora företag starkt ifrågasättas.
Utöver det - och här tror jag att kommissionsledamot Charlie McCreevy har alldeles rätt - är det aktuella förslaget ingenting annat än en nerbantad version av, enligt alla sätt att se, extremt komplicerade internationella standarder, som är helt olämpliga för strukturerna i europeiska små och medelstora företag.
Särskilt olämpliga är de för familjeföretag, som drivits av ägarna under flera generationer och som redan har skrivit av sina tillgångar och där tillämpning av reglerna om korrekt värde skulle uppmuntra till girighet och i slutändan kanske mycket väl skulle kunna äventyra företagens möjligheter till överlevnad.
Å andra sidan måste vi vara realistiska.
Frågan om redovisningsstandarder för små och medelstora företag i Europa kommer slutligen inte att kunna undgå vissa påtryckningar om harmonisering.
Vi kräver jämförbarhet, åtminstone inom den inre marknaden.
Därför anser jag att det är viktigt att vi allvarligt tänker igenom hur vi kan utveckla europeiska alternativ till förslagen från London, för att nå större standardisering också inom detta område - men en standardisering som är förnuftig och lämplig för små och medelstora företag och som är inriktad på långsiktig, istället för på kortsiktig värdering.
Jag har ytterligare en anmärkning om organen för internationella redovisningsstandarder (IAS).
Här finns ett verkligt problem, liksom Alexander Radwan antydde.
Det kan finnas en viss geografisk balans, men det finns ingen balans när det gäller ekonomisk betydelse.
Europa är det ojämförligt största blocket och den största region där reglerna om internationella redovisningsstandarder gäller.
Därför måste vi ha ett inflytande som står i proportion till detta, och vi kan helt enkelt inte jämföras med till exempel Australien.
Australien har samma betydelse som ett medelstort EU-land, eller snarare en stor region som Nordrhein-Westfalen.
I detta avseende måste balansen förbättras.
för PPE-DE-gruppen. - (NL) Fru talman! Jag vill först framföra mina gratulationer till Alexander Radwan för att han har slutfört det här grundliga betänkandet.
Det diskuterades ända in i det sista.
I sin slutliga form är det ett betänkande som är klart och tydligt, men ibland också kritiskt.
Föredraganden är övertygad om att IASB:s demokratiska redovisningsskyldighet måste förbättras och jag är glad att se att IASB tar till sig kritiken.
Styrelseordförande Gerrit Zalm antydde nyligen i Europaparlamentet att han var öppen för förslag och redo att lägga fram förslag om att anta strukturen.
IASB arbetar med internationella redovisningsstandarder för små och medelstora företag.
Jag är överens med föredraganden om att de internationella redovisningsstandarderna är för komplicerade och för dyra för små och medelstora företag.
Jag tror också att om små och medelstora företag uppmuntras till frivillig användning av internationella redovisningsstandarder finns det en risk för att de införs bakvägen i Europa.
Som jag ser det måste det finnas en viss differentiering beroende på företagsstorlek.
Det är bra om stora multinationella företag, banker och försäkringsbolag som har världsomspännande verksamhet använder samma standard i sina årsredovisningar.
Små och medelstora företag i Europa bör dock ha sin egen standard.
IASB har åstadkommit mycket i fråga om internationellt börsnoterade företag och deras redovisningsstandarder.
Om små och medelstora företag nu säger att kostnader och insatser kan hanteras lika bra med mer än en standard, kan vi inte använda en enda standard som påförs uppifrån och ner.
Det är också mycket viktigt att beakta investerarnas intressen liksom öppenheten.
Handlingsreglerna har vi för att underlätta, för att se till att vi får pålitlig, tydlig och kostnadseffektiv information om företagens verksamhet.
Jag tror att den bevisade nyttan av internationella redovisningsstandarder också kan gagna den europeiska aktiemarknaden, helt säkert om man i USA byter ut US GAAP-systemet mot internationella redovisningsstandarder.
Jämförbarhet kan här bli till stor nytta för internationella investerare och aktörer.
Idén bakom de internationella redovisningsstandarderna bör således stödjas av Europaparlamentet.
PSE-gruppen. - (FR) Herr kommissionsledamot!
Tack för att ni har tagit er tid att komma till Strasbourg.
Jag vill också tacka föredraganden, i er bayerska folkdräkt.
Jag anser att vi har samarbetat bra och ett bevis på det är det sätt på vilket olika personers ändringsförslag har kunnat införlivas i betänkandet.
Först av allt vill jag göra tre påpekanden om redovisningsstandarder.
Det tycks mig som om vi befinner oss i en ovanlig situation när det gäller styrningen av och funktionssättet hos det organ som ansvarar för att fastställa dessa redovisningsstandarder.
Det finns många former av standardisering.
Inte alla dessa har en så stark påverkan på den finansiella stabiliteten, eller på sådana frågor, när det gäller makt och styrning, som redovisningsstandarderna.
Det som händer idag är en viktig händelse, en mognad.
När redovisningsstandarderna utarbetades, kanske av revisorer som samarbetade inbördes, beredde de marken mycket väl.
Numera är dessa redovisningsstandarder internationella.
De används och tillämpas av var och en och frågan om styrning är därför avgörande.
Hur är det organ som har ansvaret för att fastställa dessa redovisningsstandarder anpassat till internationella styrelseformer, i förhållande till demokratiska organ, organ som lagligen företräder statsmakten, och i synnerhet EU?
Den andra punkt som vi måste titta på när det gäller styrning är givetvis balansen mellan dessa organ.
Vilken är den geografiska balansen, vilken är balansen i fråga om representationen inte bara av dem som utarbetar standarderna, utan också av dem som måste använda dem?
Den tredje punkten är finansieringen.
Hur ska dessa organ finansieras?
Kan idén om en skatt på näringsverksamhet, som skulle kunna samordnas av tillsynsorgan, vara givande?
Skulle organen kunna finansieras av regeringen, av Europeiska gemenskapen?
Vi hoppas att kommissionsledamot Charlie McCreevy ska komma med några väl underbyggda förslag på den punkten.
Den fjärde frågan beträffande dessa organ är programmet.
Är det rätt att de utvecklar begreppet korrekt värde när vi vet vilka effekter det kan ha på den finansiella stabiliteten?
Är det rätt att detta organ utarbetar ett program för små och medelstora företag om Europa inte behöver ett sådant program?
I denna fråga om standarder för små och medelstora företag - bara för att Sydafrika eller Australien kan behöva dem, liksom vår föredragande har sagt - är det riktigt att kommissionsledamot Charlie McCreevy inte kan garantera att Europa får någon talan i dessa organ.
Som ett första steg är det är absolut väsentligt att Europa ser till att finnas med för att representera styrkan hos samtliga medlemsstater och föra fram samtliga EU-medborgares röst, i IASB, IASCF och IFRIC.
Kommissionsledamot Charlie McCreevy, det är ert ansvar.
På den punkten förväntar vi oss att ni ger oss väl underbyggda förslag.
för ALDE-gruppen. - (EN) Fru talman! Internationella redovisningsstandarder används av allt fler länder och växer i betydelse och värde.
Det gör det nödvändigt att stärka IASB:s redovisningsskyldighet och öppenhet, vilket kanske inte framstod tydligt från första början.
Jag välkomnar åtgärder i den riktningen, men jag beklagar att man i några delar av betänkandet framför negativ kritik, i stället för att bekräfta att förändringar är på gång och peka på vägen framåt.
Flera av mina ändringsförslag syftar därför till att se framåt, och understryka fördelar och goda sidor parallellt med behovet av ytterligare anpassning, både av själva standarderna och av IASB som övervakar dem.
Onödig politisering av tekniska frågor måste dock undvikas.
Internationella redovisningsstandarder är ett viktigt verktyg för att främja jämförbarhet över gränserna och minska betungande krav på att företag ska rapportera under olika system, men det vore bra om årsredovisningarna var lättare att använda för andra jämförande syften.
Men det kan mycket väl vara så att verktyg som XBRL-tagging kan utveckla detta.
Jag måste tacka Ieke van den Burg för att hon förra veckan organiserade en intressant presentation i det här ämnet.
De förslag som gäller små och medelstora företag orsakar oro i många läger.
Jag uppfattar dem mest som verktyg för medelstora enheter, som kanske är på väg mot full offentlig rapportering, och mot bakgrund av detta kan det finnas anledning att hantera dem separat eller göra dem frivilliga.
Men som kommissionsledamot Charlie McCreevy framfört är de alldeles för komplicerade för de flesta vanliga mindre och medelstora företag.
(EN) Fru talman! Jag vill tacka min kollega Alexander Radwan för hans utmärkta betänkande.
Jag hoppas att den bayerska folkdräkten han har på sig idag inte betyder att han har ändrat politiska inriktning.
Antagandet av internationella redovisningsstandarder (IFRS) i januari 2005 har gynnat Europeiska unionen genom att förenkla redovisningskraven över gränserna, göra det lättare att jämföra ekonomiska redovisningar för olika länder, konkurrenter och företag samt förbättra arbetet med reglerad tillsyn, bankverksamhet och kapitalmarknader.
Internationella redovisningsstandarder används nu eller antas i mer än hundra länder, inklusive Australien och Sydafrika.
Jag stöder kravet på ökad insyn, effektivitet och redovisningsskyldighet när det gäller IASB.
I betänkandet uppmärksammas att det hann gå 17 månader innan IASB utsåg en ny ordförande.
Detta är oacceptabelt.
IASB är ett privat, självreglerande organ som har fått rollen som regelmakare och det är inte mer än rätt att vi därför kräver ökad redovisningsskyldighet och tillsyn.
Vi bör också vara försiktiga med att kräva extra EU-strukturer som ska hantera tolkningen och tillämpningen av internationella redovisningsstandarder.
Varför då?
Vilken nytta gör de?
Det har gjorts stora framsteg på detta område i fråga om konvergensen mellan Europa och USA samt för den europeisk-amerikanska färdplanen för samordning och harmonisering av redovisningsstandarder.
Förra året undertecknade Förenta staternas president, Europeiska rådets tjänstgörande ordförande och Europeiska kommissionens ordförande ett gemensamt uttalande om att främja och skapa förutsättningar för erkännande av GAAP, de amerikanska allmänt accepterade redovisningsprinciperna, och av internationella redovisningsstandarder i båda dessa jurisdiktioner.
Detta är mycket välkommet.
När det gäller att tillämpa internationella redovisningsstandarder för små och medelstora företag, kan små och medelstora företag vara små eller mindre.
Jag anser att det kanske kan vara bättre att göra tillämpningen valfri för att garantera flexibilitet, snarare än att förhindra den helt och hållet.
(NL) Fru talman! Jag vill upprepa de tidigare komplimangerna till Alexander Radwan, inte minst eftersom hans betänkande gett oss en väldigt intressant debatt om konflikten mellan lagstiftning och självreglering, särskilt på global nivå.
Jag förstår att våra ambitioner lämnar oss i bryderi.
Å ena sidan vill vi att dessa internationella standarder ska tillämpas över hela världen, å andra sidan insisterar vi på vår auktoritet som medlagstiftare för att kunna bestämma innehållet i standarderna och uppfylla vår skyldighet som medlagstiftare på ett ansvarsfullt sätt.
Jag anser att Europaparlamentet på senare tid har visat att det gör det.
Nyckeln anser jag finns i lägliga samråd, ett balanserat beaktande av samtliga parters intressen, inklusive rättigheter för tredje part som t.ex. anställda, lokala myndigheter, leverantörer och så vidare (eftersom adekvat finansiell rapportering gynnar fler än bara finansieringsinstituten), samt en ordentlig konsekvensbedömning.
Kommissionen har här ett tungt ansvar.
Och i den omedelbara framtiden måste dessa funktioner utföras för små och medelstora företags räkning.
Vi kan göra detta till ett verkligt givande projekt för Europeiska unionen.
Till sist har jag två kommentarer som även är relevanta för ett annat betänkande som vi kommer att rösta om under vår nästa sammanträdesperiod, Klaus-Heiner Lehnes betänkande om ett förenklat företagsklimat.
Här anser jag också att reglerna inte bara gäller företag, finansieringsinstitut och de revisorer som lever på dem, utan också anställda samt andra grupper.
Så vi får inte blanda oss i reglernas kvalitet.
Jag har förespråkat att reglerna hursomhelst bör tillämpas för avregistrerade företag och all extern verksamhet.
Jag hoppas att ni håller med om att det även finns arbete för IASB inom det området.
Slutligen vill jag upprepa mitt stöd till standarden eXtensible Business Reporting Language (XBRL).
Som ni vet är Förenta staternas finansinspektion i färd med att besluta om att göra den obligatorisk.
Jag vill uppmana er att tänka på hur EU ska reagera på detta och uppmuntra er att upprätta en färdplan för Europeiska unionen i enlighet därmed.
(EN) Fru talman! Det finns problem med insynen och styrningen av IASB, International Accounting Standards Board, men organisationen har accepterat kritiken och erkänt att det behövs en förändring.
Åtgärder har vidtagits och fler är planerade: publicering av återkopplingsrapporter, beslutsförklaringar, påtryckningar för kostnads- och intäktsanalyser samt en utvidgad och aktivare delaktighet för styrelsen.
Den gjorde sitt yttersta för att kommunicera med Europaparlamentet.
Alexander Radwans betänkande har förbättrats avsevärt jämfört med de tidigare versionerna och jag tror att de positiva ändringsförslagen från PPE-DE-gruppen och ALDE-gruppen idag kommer att förbättra texten ytterligare.
Jag vill tacka föredraganden, eftersom han trots våra meningsskiljaktigheter varit villig att kompromissa när det gäller vissa aspekter inom styrning.
Tyvärr kan jag inte hålla med honom i frågan om internationella redovisningsstandarder för små och medelstora företag.
IASB ombads utarbeta en förenklad version för små och medelstora företag.
Alexander Radwan vill i sitt betänkande inte erkänna att detta även kunde vara användbart i Europeiska unionen.
Trots att förslaget fortfarande inte är klart tillkännages det redan i betänkandet att det definitivt inte kommer att främja europeiska företag.
Ändå har vi fått veta flera gånger att standarderna kommer att bli valfria och är till för växande små och medelstora företag vars målsättning är att bli börsnoterade företag.
Små företag utan ambitioner utanför de lokala marknaderna behöver inte tillämpa dem.
I en opinionsundersökning som utfördes i september i fjol ansåg en tydlig majoritet bland de små och medelstora företagen i Europeiska unionen, inklusive tyska små och medelstora företag, att fördelarna vägde tyngre än nackdelarna och att de skulle komma att förbättra den finansiella rapporteringen.
IASB:s ansträngningar för att utveckla globala redovisningsstandarder av hög kvalitet är ett viktigt och uppskattat bidrag till EU:s och världens ekonomi och vi bör därför välkomna detta.
(ES) Fru talman! Kravet sedan 2005 om att börsnoterade företag ska använda internationella redovisningsstandarder för sina konsoliderade finansiella rapporter har varit ett vittomfattande och mycket inflytelserikt politiskt initiativ.
Cirka 100 länder använder standarderna och deras globalisering har gett förbättrad jämförbarhet och ökad insyn. Därmed har operatörernas förtroende ökat, vilket skapat mer lika villkor och en starkare marknadsdisciplin.
Betänkandet innehåller två stora utmaningar i fråga om styrning.
Å ena sidan har vi ett privat organ, som har upprättat valfria globala standarder sedan 1973 på företagsmässig och professionell grund och som nu befinner sig i en ansvarstyngd position. Det leder i sin tur till en förändring i dess organisation, förfaranden och sammansättning för att det ska kunna bli ett öppnare och mer kontrollerbart organ, med en behörighet som återspeglar den nya rollen.
Det är nödvändigt att erkänna och samordna verksamheten för samtliga berörda offentliga och privata intressen och samtidigt säkra organisationens finansiering och självständighet när det gäller att fastställa standarder.
Organisationen måste dessutom integreras i internationella ledningsstrukturer.
Det är också nödvändigt att stärka den europeiska redovisningsstyrningen genom att anta en mer aktiv och integrerad strategi för upprättande, antagande, genomförande och bedömning av standarder.
Det är avgörande att förbättra den begreppsmässiga ramen för standarder och man bör beakta att de varken är neutrala eller akademiska och kan skapa både vinnare och förlorare.
Likaledes är det viktigt att bedöma deras effekter, garantera att de kan förenas med en europeisk strategi, lära från finansiella omvälvningar och reglera redovisningsstandarderna för administrativa koncessioner på ett balanserat sätt.
De finansiella redovisningsarrangemangen för små och medelstora företag måste vara enkla och kopplas till den interna och globala marknaden.
Dessa frågor tas upp i Alexander Radwans betänkande, som har samlat en bred enighet och som kommer väldigt lägligt med tanke på den kommande översynen i slutet av 2009. Enligt betänkandet ska det tillsättas ett tillsynsorgan och sammansättningen av Standards Advisory Council ska ändras före nästa år.
(DE) Fru talman, herr kommissionsledamot, herr Radwan, mina damer och herrar! Jag välkomnar varmt detta betänkande och denna debatt, eftersom jag anser att vi tack vare den undersöker några mycket känsliga frågor grundligt och över partigränserna.
Flera punkter avtecknar sig tydligt utifrån det som har sagts.
För det första behöver vi en gemensam uppsättning standarder för börsnoterade aktiebolag, men vi vill inte klumpa ihop alla företag.
För det andra, fastän vi inte förkastar särskilda regler som anpassats för små och medelstora företag, måste ramen för dessa regler fastställas av Europeiska unionen. För det tredje är de åtgärder som för närvarande föreslagits alltför komplexa och dyra.
De gör ingen nytta för små och medelstora företag. Av dessa skäl måste vi avvisa dem.
För det fjärde väntar vi fortfarande på tillfredsställande svar på frågorna om vem som gör reglerna och för vem, samt vem som övervakar processen. Det finns ingen demokratisk legitimitet.
Det finns ingen åtskiljande strategi. Små och medelstora företags berättigade önskningar har inte beaktats och systemet för demokratisk övervakning är otillräckligt.
För det femte, genom att ta ställning i denna fråga eller försöka besvara dessa frågor, glömmer vi ofta bort att två tredjedelar av arbetskraften finns inom den privata sektorn i familjeägda företag och att majoriteten av dessa familjeägda företag är små och medelstora företag som inte söker finansiering från kapitalmarknaderna.
Detta är en punkt som vi måste komma ihåg när vi ställs inför denna typ av förslag som behandlar alla företag lika.
Tack för denna givande debatt!
(EN) Fru talman! I punkt 30 i vårt resolutionsförslag påpekas att resultatrapporter inte bara främjar investerarnas, utan också övriga berörda parters behov.
Eftersom vi också uppmärksammar behovet av ändringar i EU-lagstiftningen i punkt 41 vill jag påminna kommissionsledamoten om att parlamentet har röstat för att samtliga ändringar i det fjärde och sjunde direktivet om bolagsrätt ska omfatta ett krav på företagen om rapportering av sociala och miljömässiga resultat.
Jag vill påpeka att sådana krav redan finns i Sydafrika, i Frankrikes lagstiftning om nya ekonomiska förordningar samt i rekommendationerna från projektet ”Prince of Wales's Accounting for Sustainability” från mitt eget hemland, Storbritannien.
Dessutom vill jag fråga kommissionsledamoten, med tanke på kommissionens rekommendation om miljöfrågor år 2001 i vår nya bokföring, om kommissionen skulle kunna utfärda en liknande rekommendation om sociala frågor i bokföringssammanhang.
Kan kommissionsledamoten förmå IASB att inkludera sociala och miljömässiga aspekter i sin planerade publicering av ledningens kommentarer?
Oavsett om kommissionen vill kalla detta för företagens sociala ansvar, kan vi idag kanske enas om att kalla det för redovisning av ansvarstagande företag.
(ES) Fru talman! Den ekonomiska krisen nyligen har visat på betydelsen av högkvalitativa redovisningsstandarder för väl fungerande marknader.
En annan viktig lärdom att dra av krisen är att det råder en viss asymmetri mellan den fastställda vikten av redovisningsstandarder och de privata organens karaktär och ledningsstrukturer, i fråga om deras ansvar för upprättande, fastställande och tolkning av dessa standarder.
Alexander Radwan gör därför rätt i att påpeka att det första som bör hanteras är styrningen.
Jag anser att han har lagt fram intelligenta och realistiska förslag om behoven hos de institutioner som representerar Europeiska unionen, som att vara mer aktiva i processen med att fastställa standarder som ska införlivas i gemenskapens lagstiftning samt engagera sig i hur dessa privata organ fungerar internt.
Ökad insyn, skydd för att förhindra intressekonflikter och bredare geografisk representation är några av förslagen i Alexander Radwans betänkande.
Den andra aspekten som hanteras i betänkandet handlar om små och medelstora företag.
I denna kammare har vi betonat vikten av att förlika två målsättningar: förenkling och sänkta kostnader för små och medelstora företag i fråga om redovisningsförfaranden och tillhandahållandet av lämplig information för marknadsaktörer.
Den sista punkten i Alexander Radwans betänkande - som jag instämmer i - är behovet av globala standarder i en global miljö.
Därför är det mycket viktigt att nå överenskommelser med de andra stora ekonomiska världsmarknaderna, i synnerhet Förenta staterna.
Detta kräver ett större engagemang samt en utökad roll för EU:s institutioner, inklusive denna kammare och alla de som lyssnar idag.
(DE) Fru talman! Jag kan helt och hållet instämma i vad vår kollega precis sagt.
Den bakomliggande premissen här - och Alexander Radwan sätter fingret på detta i sitt betänkande - är att en institution utan ett politiskt mandat likväl bör vidta ett antal åtgärder som påverkar ekonomin, varav några är bindande.
Det räcker inte att uppmana till bättre styrning eller bättre ramvillkor, de politiska organen måste också bli mer engagerade i denna fråga än tidigare.
Vad vi gör här i Europaparlamentet är att ta ett steg i rätt riktning, men ytterligare steg måste tas.
Det finns också en annan aspekt att beakta.
Det som uträttas här på regional organisationsnivå - i detta fall Europeiska unionen - bör också återspeglas i den globala kontexten.
Så det handlar inte bara om att försöka tillämpa dessa regler i vår egen del av världen.
(LT) Fru talman! Som min kollega tidigare nämnde handlar detta betänkande om vem som ansvarar för vad i redovisningsprocessen.
Europaparlamentets roll är mycket viktig och enligt mig berättigad.
Jag vill dock uttrycka en viss tvekan när det gäller beaktandet av varje teknisk detalj och upprättandet av standarder.
Jag anser inte att beskrivningen av bedömnings- och utvärderingsmetoden för säljbara och icke-säljbara tillgångar är helt tillfredsställande.
Därför är jag tveksam till om vi verkligen ska försöka bedöma om det är en bra eller dålig metod.
Vi bör vänta på att experterna har gjort sin bedömning.
Samtidigt har översynen av standarden om icke-säljbara tillgångar och samråd i denna fråga påbörjats.
Endast därefter bör vi fatta vårt beslut.
Jag föreslår därför att vi inte ska stödja förslaget i artikel 30 e eller det i artikel 42.
(EN) Fru talman! Kan kommissionsledamot McCreevy garantera att den gemensamma uppsättningen globala redovisningsstandarder - med en efterföljande satsning på en ökad standardisering av förfarandena - inte på något sätt kommer att rättfärdiga eller för den delen stärka kravet på en gemensam konsoliderad bolagsskattebas i Europeiska unionen?
ledamot av kommissionen. - (EN) Fru talman! Jag vill tacka ledamöterna för deras kommentarer.
Det var verkligen en bred debatt med många åsikter i flera av frågorna och vi har noterat dem.
Jag vill återigen betona att högkvalitativa internationella redovisningsstandarder är avgörande för att både EU:s och världens kapitalmarknader ska fungera väl.
Processen med att utveckla dessa standarder bör därför styras handfast.
Den bör karaktäriseras av en hög insynsnivå och den bör garantera en balanserad bedömning av de berörda parternas intressen.
IASCF, Accounting Standards Committee Foundation, och IASB har under de senaste åren genomfört viktiga reformer av sina interna förfaranden men jag kan inte förneka att ytterligare förbättringar krävs.
Dessutom är jag den förste att erkänna att Europeiska unionen behöver organisera sig bättre för att kunna vägleda och komma med förslag till IASB i dess process med att fastställa standarder.
Kort sagt, även om IASB:s styrning och rutiner vore perfekta, skulle de internationella redovisningsstandarderna endast kunna vara till hjälp för EU:s behöriga parter om de presenterades på ett sammanhängande, övertygande och lämpligt sätt.
Nästan alla talare hänvisade till frågan om internationella redovisningsstandarder för små och medelstora företag och jag upprepar återigen att det för närvarande inte finns någon rättslig grund för att godkänna sådana i Europeiska unionen.
Om den skulle ändras krävs det medbeslutande av Europaparlamentet.
Låt mig bara upprepa, som jag redan sagt tidigare angående internationella redovisningsstandarder för små och medelstora företag: när IASB utförde detta arbete förklarade jag tydligt i ett antal anföranden att de inte skulle förutsätta ett automatiskt stöd för detta särskilda projekt från Europeiska unionen.
Vi skulle endast rekommendera det om det var enkelt och effektivt och uppfyllde behoven hos små och medelstora företag.
De fick reda på detta när de höll på med sitt arbete.
Deras första samrådsdokument har lagts fram.
Jag tog då tillfället i akt och berättade för dem att det inte uppfyllde kriterierna och att som det såg ut nu kunde jag överhuvudtaget inte ens överväga att rekommendera dem för små och medelstora företag, eftersom de varken var enkla eller effektiva.
Det är fortfarande min ståndpunkt men med tanke på vad andra har sagt, i synnerhet John Purvis, skulle det säkert vara bra om det fanns en enkel och effektiv internationell redovisningsstandard för små och medelstora företag - men endast av det skälet.
Idén är bra.
Jag vill inte alls racka ner på idén, men jag kommer varken nu eller i framtiden att stödja något för små och medelstora företag som bara är mer komplext och som ingen förstår.
Det behövs inte.
Jag vill ta denna chans att återigen upprepa vad jag sagt tidigare om detta.
Ieke van den Burg nämnde frågan om XBRL.
Vi arbetar tillsammans med tillsynsmyndigheten för värdepappershandel för att få enighet kring de tekniska standarderna för affärsuppgifter och som ett resultat av denna dialog kan kommissionen vidta ytterligare åtgärder som syftar till kompatibilitet för system för regleringsinformation.
XBRL kan tillåta investerare att utnyttja de internationella redovisningsstandarderna till fullo.
Samtliga åtgärder som syftar till att kräva att XBRL ska användas i Europeiska unionen bör genomgå en grundlig konsekvensbedömning, inklusive en ekonomisk bedömning av kostnader och fördelar.
Jag diskuterade också frågan med Chris Cox, ordföranden för den amerikanska finansinspektionen, under mitt senaste besök i USA och jag stöder att vi i framtiden behåller denna punkt på dagordningen i vår dialog om tillsyn med de amerikanska myndigheterna.
Dessa standarder måste godkännas internationellt samt bli tekniskt oberoende och kompatibla.
Utvecklingen är mycket spännande och jag vet att Ieke van den Burg nyligen har kommit i kontakt med detta.
Jag tog samma chans för några månader sedan och lät experter visa mig hur det i själva verket fungerar.
Jag anser att det verkligen är revolutionerande och samtidigt något att välkomna. Men vi kommer inte att göra någonting åt det riktigt ännu förrän vi har utfört andra saker.
Gay Mitchell tog upp en viktig punkt.
Vi vill inte att IASB ska komma och säga ”ett EU-organ eller något annat organ, vilket som helst”.
Vi vill vara ett internationellt accepterat organ - eftersom detta mål är väl värt att eftersträva - och det måste vara ett oberoende organ.
Jag anser att det ska antas men med ordentlig input från de berörda parterna.
Jag vill påminna alla om att det var Europeiska unionen som gav IASB denna betydelse.
Vi var den största jurisdiktionen som sa att från och med 2005 skulle de internationella redovisningsstandarderna bli regel för börsnoterade företag.
Det var för några år sedan som detta beslut togs, tillsammans med Europaparlamentet, och det i sig gjorde IASB och processen mer betydelsefull.
Jag skulle säga - och jag har sagt detta tidigare även till IASB - att en provkörning - ni kan kalla det en konsekvensbedömning - bör utföras innan standarderna antas, särskilt av IASB, tillsammans med bidrag från Europeiska unionen och andra organ.
Vi bör inte vänta tills standarderna har godkänts av IASB.
Vår roll var att antingen stödja dem eller förkasta dem, inte att ändra dem.
Jag anser att de ska testas ordentligt i förväg för att upptäcka eventuella problem, istället för att allvarliga problem upptäcks sedan man gått igenom hela IASB:s process.
Vi upprepade detta flera gånger för IASB.
Förhoppningsvis uppskattas de nya styrningsstrukturerna av de flesta av oss.
Jag erkänner att det behövs mer arbete på detta särskilda område, men det i sin tur kan ge färre problem i framtiden.
Förhoppningsvis kommer vi en dag att nå en situation där dessa saker mer eller mindre kommer att ske automatiskt och inte vålla för mycket bekymmer för någon, eftersom allt arbete redan kommer att ha gjorts i förväg.
Då kommer vi inte att ha några problem.
föredragande. - (DE) Fru talman, herr kommissionsledamot, mina damer och herrar! Jag vill verkligen tacka för denna debatt, där målet med betänkandet har fått stöd och alternativ har presenterats på flera områden.
Jag skulle vilja nämna två saker.
Det finns en punkt som jag är säker på att vi alla är överens om, och som dessutom har nämnts upprepade gånger idag av flera talare som helt stöder denna allmänna utveckling, nämligen att organisationen bakom de internationella redovisningsstandarderna nu har vidtagit en del åtgärder, till exempel när det gäller frågor om styrning, som ett resultat av påtryckningar från Europaparlamentet och Europeiska unionen.
Ibland måste vi vara tydliga - och jag vet att en del av mina kvinnliga kollegor har kritiserat mig på den punkten - eftersom vissa personer som har talat inför denna kammare under de senaste åren emellanåt har gett ett intryck av att Europaparlamentet inte betyder särskilt mycket för dem.
Hur få framsteg som har gjorts framgår tydligt av betänkandet om styrning, där det föreslås att framtidens tillsynsmyndigheter endast ska följa råd från personer som de har utsett.
Allt jag kan säga om detta är att alla som i framtiden måste redovisa för parlamentet hur han eller hon har röstat i en särskild fråga ska se till att en del av ansvaret och möjligheten att kunna påverka när det gäller politikens utformning är en del av paketet.
Det var det första jag ville säga.
Hur lite engagemang det finns i frågan om konsekvensbedömningar framgår tydligt av diskussionen. Organisationen bakom de internationella redovisningsstandarderna vägrar fortfarande att utföra dem.
När det gäller frågan om standarder för små och medelstora företag vill jag säga något till er som anser att vi ska införa dem på frivillig basis.
Inspirerad av John Purvis - John, detta riktar jag till dig - vill jag citera en oberoende kommentator.
Peter Holgate, partner i PricewaterhouseCoopers, skrev följande i den tyska utgåvan av Financial Times:
”Jag tar inte EU:s ståndpunkt på särskilt stort allvar.
Även om det slutar med att de inte godkänner standarderna kan flera länder anta dem i sina nationella allmänt accepterade redovisningsprinciper.
Om några stora aktörer antar standarderna kommer deatt införas på ett annat sätt, fastän Europeiska kommissionen inte vill vara med och leka.”
I slutändan innebär det att man måste anta att när väl några stater har antagit dessa standarder kommer de att införas obligatoriskt i hela Europeiska unionen.
Sådan är denna organisations strategi.
PricewaterhouseCoopers har redan sagt att de ser detta som en affärsmodell.
Därför behöver vi vår egen uppsättning europeiska standarder för små och medelstora företag: vi kan bygga vidare på internationella redovisningsstandarder om det är lämpligt, men om det inte är det, då utvecklar vi våra egna standarder.
Det är kommissionens skyldighet att se till att man inte prackar på oss standarder bakvägen, standarder som ingen vill ha men som ändå blir allmänt bindande.
Debatten är härmed avslutad.
Omröstningen kommer att äga rum idag kl. 12.00.
Skriftliga förklaringar (artikel 142)
(Sammanträdet avbröts kl. 11.55 och återupptogs kl. 12.00.)
Rättelser till avgivna röster och röstavsikter: se protokollet
Öppnande av sammanträdet
(Sammanträdet öppnades kl. 09.00.)
3.
Återlämnande av kulturföremål som olagligen förts bort från en medlemsstats territorium (kodifierad version) (
Avslutande av sammanträdet
(Sammanträdet avslutades kl. 23.40.)
13.
2007 års framstegsrapport om Turkiet (
- Före omröstningen om ändringsförslag 11:
(DE) Herr talman! Vi håller med våra ledamotskolleger om att vi bör erkänna rollen för det kurdiska språket i Turkiet på lämpligt sätt.
Punkt 11 kräver emellertid ett visst språkligt klargörande på en punkt.
Jag vill därför föreslå ett muntligt ändringsförslag som vi har enats om med de andra skuggföredragandena och föredraganden.
I den ändrade versionen bör meningen därför lyda som följer:
(EN) ”inklusive verkliga möjligheter att studera kurdiska inom det offentliga och privata skolsystemet och använda detta språk i radio- och TV-sändningar, i det offentliga livet och i kontakterna med offentliga myndigheter.”
(Parlamentet gav sitt samtycke till att detta muntliga ändringsförslag skulle beaktas.)
- Före omröstningen om punkt 19:
föredragande. - (NL) Vi vill stryka ordet ”angränsande” eftersom vi vill att ombudsmannen ska samarbeta med alla europeiska ombudsmän och ombudskvinnor.
(Parlamentet gav sitt samtycke till att detta muntliga ändringsförslag skulle beaktas.)
Debatter om fall av kränkningar av de mänskliga rättigheterna samt av demokratiska och rättsstatliga principer (debatt)
20.
Konkurrens - Branschutredning om banktjänster till privatpersoner och mindre företag (
21.
Grönbok om finansiella tjänster till privatpersoner och mindre företag på den inre marknaden(
°
° °
(SL) Jag skulle vilja kommentera vad som sades i början av omröstningen när flera ledamöter försökte använda sig av incidenten vid kärnkraftverket i Krško för att illustrera kärnkraftsverkens bristfälliga säkerhet.
Jag vill påpeka att det verkligen rörde sig om en incident, att det handlade om ett komponentfel, att kraftverket inte stängdes ner utan att verksamheten snarare tillfälligt upphörde av säkerhetsskäl och att reparationer pågår.
Kärnkraftverket erbjuder insyn i sin verksamhet och ledamöterna kan hitta information om det på den slovenska kärnsäkerhetsmyndighetens hemsida.
Jag vill även tillägga att kärnkraftverket i Krško enligt alla säkerhetsindikatorer hör till de säkraste i världen.
Utskottens och delegationernas sammansättning: se protokollet
Översyn av ramdirektivet om avfall (debatt)
Nästa punkt är en andrabehandlingsrekommendation från utskottet för miljö, folkhälsa och livsmedelssäkerhet om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets direktiv om avfall och om upphävande av vissa direktiv (11406/4/2007 - C6 0056/2008 - (Föredragande: Caroline Jackson).
föredragande. - (EN) Fru talman! Jag rättar mig efter ert beslut om att inte ägna tid åt ordningsfrågor och fortsätter med mitt anförande om ramdirektivet om avfall.
Det är lite svårt att göra det mot denna bakgrund, men jag ska fortsätta.
Eftersom det nyligen har förekommit vissa kommentarer om den här punkten i brittisk press, vill jag börja med att ännu en gång uppmärksamma er på den anmälan av ekonomiska intressen som jag har gjort i registret och där jag uppger att jag är medlem i den rådgivande miljökommittén i företaget Shanks plc.
Företaget är verksamt inom en rad avfallsteknologier i Storbritannien och på kontinenten, och det primära ändamålet för den rådgivande miljökommittén är att genomföra oberoende granskning av verksamheten i dess anläggningar.
Bland mina kollegor i kommittén finns ordföranden i EU:s vetenskapliga kommitté för nya och nyligen identifierade hälsorisker och en medlem i den brittiska frivilligorganisationen Green Alliance.
Som många andra ledamöter värdesätter jag det tillfälle som en sådan här erfarenhet ger att på nära håll få inblick i de frågor och problem som den här industrin och de som arbetar inom den möter.
När det gäller direktivet har det varit en lång och svår väg fram till denna andra behandling, och jag gratulerar dem av mina kollegor som har följt med mig hela vägen fram.
Det är en mycket viktig fråga.
Det har krävts klargöranden av olika domar från EG-domstolen om vilken typ av avfall som ska hanteras i anläggningar för energi från avfall.
Det har krävts nya definitioner.
Två befintliga direktiv om farligt avfall respektive spilloljor har upphävts, och bestämmelserna i dessa har överförts till ramdirektivet om avfall.
Men utskottet var inte tillfreds med de ursprungliga förslagen och fortsatte att omvandla direktivet från ett tekniskt till ett propagerande direktiv.
Jag gratulerar mina kollegor till detta.
Jag måste säga att det rådde en dyster stämning i rådet, möjligen på grund av det aktuella ekonomiska läget.
Det fanns ett stort motstånd till vad vi ville göra och rådet var svårt att blidka, men vi fick igenom följande.
För det första har vi lagt till mål för materialåtervinning i texten.
Det var mycket viktigt eftersom det inte fanns några sådana mål i det ursprungliga förslaget, och detta är första gången som materialåtervinningsmål för hushållsavfall förekommer i gemenskapens lagstiftning.
Det är helt och hållet tack vare parlamentet som de finns med.
Enligt den nya artikel 8a måste medlemsstaterna vidta nödvändiga åtgärder för att den totala graden av materialåtervinning av papper, metall, plast och glas från hushåll och liknande avfall ska uppgå till 50 procent till 2020.
För några medlemsstater, som till exempel Tyskland, är det här ett konservativt mål, men för många är det mycket krävande och vi måste ta hänsyn till dem också.
Enligt samma artikel måste graden av materialåtervinning av byggnads- och rivningsavfall vara 70 procent till 2020.
De gröna och deras anhängare sprider rykten om att målen inte kan tvingas fram.
Kanske tror de till och med själva på dem, men märkligt nog avvisar de sitt eget resultat.
Kommissionen har gjort ett uttalande för att hjälpa dem, vilket Stavros Dimas kan bekräfta.
I sitt uttalande säger kommissionen klart och tydligt att om en medlemsstat inte når målen till 2020 kommer kommissionen att betrakta det som ett allvarlig tecken på att medlemsstaten inte har vidtagit nödvändiga åtgärder för att nå målen.
Mot bakgrund av detta, och med stöd i slutsatserna i de nationella lägesrapporter som medlemsstaterna ska lämna vart tredje år, kan kommissionen dra medlemsstaterna inför EG-domstolen om de inte följer bestämmelserna i direktivet.
Det kanske är viktigt för de gröna att inte vara nöjda, eftersom de gröna är eviga miljökämpar, men de borde ta till sig något av vad kommissionen har sagt i sitt uttalande.
För det andra har vi lagt till nya bestämmelser om förebyggande av avfall i artikel 8 a.
Detta innebär att kommissionen måste rapportera om hur EU:s avfallshantering utvecklas och vilka möjligheter det finns för förebyggande av avfall till 2011.
Det visade sig vara omöjligt att få rådet eller kommissionen att gå med på kvantitativa mål för förebyggande av avfall i det här direktivet, delvis eftersom de uppgifter som krävs för dessa riktmärken saknas, men parlamentet har genom sina ändringsförslag skapat en impuls till en politik som i framtiden kan innehålla mål för förebyggande av avfall.
Den nya artikeln utgör därför ett viktigt framsteg.
Den är något som våra efterträdare kan bygga vidare på.
Vi kan inte göra allt i detta direktiv, utan vi måste lämna över en del till våra efterträdare under nästa årtionde.
För det tredje har vi för första gången placerat EU:s berömda avfallshierarki i gemenskapens lagstiftning.
Vi har talat om det här i åratal, men om ni tittar i gemenskapslagstiftningen finns det inte där.
Men det gör den snart, och vi kan fira en liten seger för att vi fått rådet att gå med på att hierarkin ska gälla i form av en prioriteringsordning för lagstiftning som rör förebyggande och hantering av avfall.
För det fjärde har vi enats om att bättre betona hanteringen av farligt avfall, som flera kollegor ville.
För det femte har vi även sett till att man ska fortsätta att prioritera regenerering av spilloljor, men det fanns inte något stöd för en policy, vilket jag vet att några kollegor önskade, som skulle ha gjort det obligatoriskt med regenerering i alla medlemsstater.
Rådet stöder det ändringsförslag som framlagts av Erna Hennicot-Schoepges och hennes kollegor om att underlätta för små och medelstora företag att använda avfallsförteckningen, och vi har även fått stöd för en ny artikel om biologiskt avfall.
Sammanfattningsvis innehåller direktivet uppgifter om vilka effektivitetskriterier som ska gälla för förbränning av avfall, med energiåtervinning klassad som återvinning snarare än bortskaffning.
Det här är bästa tillgängliga överenskommelse.
Att tro att vi kunde ha fått till stånd något bättre genom att gå till förlikning vore att bedra sig.
För att citera en av Jack Nicholsons gestalter: "this is as good as it gets" (ung. bättre än så här blir det inte).
ledamot av kommissionen. - (EL) Fru talman, mina damer och herrar! Jag vill börja med att tacka och gratulera föredraganden, Caroline Jackson, för hennes utmärkta sätt att bidra till granskningen av ramdirektivet om avfall, och skuggföredragandena och utskottet för miljö, folkhälsa och livsmedelssäkerhet för att de bidragit på ett positivt och konstruktivt sätt.
Med det här direktivet tar gemenskapen sitt första riktiga steg mot att skapa ett återvinningssamhälle.
I direktivet introduceras en modern hållning till avfallshantering genom att man betraktar avfall som användbart råmaterial och tillhandahåller tydligare definitioner, ett förenklat regelverk och nya ambitiösa mål.
Tack vare att bestämmelserna i direktiven om farligt avfall respektive spilloljor införlivats, ingår här direktivet i en bredare insats för att förbättra lagstiftningen och förenkla gemenskapens regelverk.
Nästa steg blir förstås att genomföra direktivet framgångsrikt.
Parlamentet har belönats för sina stora insatser och sin uthållighet.
Det var inte lätt att övertala medlemsstaterna att godkänna de nya materialåtervinningsmålen och samtycka till målen för förebyggande av avfall.
Ändå har detta mål uppnåtts i sin helhet.
Det har hörts vissa tvivel om huruvida medlemsstaterna kommer att genomföra dessa mål.
Jag skulle vilja understryka att nuvarande formulering av de kvantitativa målen ger kommissionen har förmågan och den politiska viljan hos att dra medlemsstaterna inför EG-domstolen, om de inte vidtar de åtgärder som krävs för att nå målen för materialåtervinning.
Parlamentet har införlivat många andra betydelsefulla detaljer i direktivet.
Bland dessa är den femskaliga avfallshierarkin, nya bestämmelser om separat insamling av biologiskt avfall och farligt avfall samt många lämpliga klargöranden.
Dessa ändringar gör att kommissionens ursprungliga förslag berikas och att texten förbättras, så att den blir en ambitiös normativ rättsakt för framtida generationer.
Bara det faktum att det varit möjligt att nå en överenskommelse vid andra behandlingen är naturligtvis särskilt tillfredsställande.
Jag vill ännu en gång betona Europaparlamentets konstruktiva roll i den här processen.
Det här direktivet skapar nya ramar för avfallshanteringen och ger en solid grund för andra gemenskapspolitiska initiativ.
Europeiska kommissionen är benägen att stödja kompromisspaketet för att nå en överenskommelse vid andra behandlingen.
för PPE-DE-gruppen. - (EN) Fru talman! Caroline Jackson hänvisade till ett citat av Jack Nicholson, tror jag.
Eftersom jag känner till hennes skicklighet i golf trodde jag att det kunde ha varit från Jack Nicklaus, men utan tvivel skulle de ha sagt ungefär samma sak: "Bättre än så här blir det inte."
Det är en stor hyllning till vår föredragande och jag gratulerar henne å min grupps vägnar.
Vi måste stödja henne och agera.
Det kanske inte är så bra som vi en gång hade räknat med.
Men vi har haft en enorm framgång.
Herr kommissionsledamot! Det är upp till er nu att se till att det genomförs och att utarbeta de efterföljande bestämmelserna om förebyggande till 2014.
Jag vet att ni kommer att sätta igång med den här processen och det är också viktigt.
Det är viktigt eftersom vi har haft en hel bunt med avfallsförslag under min tid i Europaparlamentet. De har handlat om fordon, elektrisk och elektronisk utrustning, batterier, förpackningar och så vidare.
Men avfallet fortsätter att öka i omfattning. Det ökar fortare än våra ekonomier växer.
Fortast växer det i vissa områden som till exempel kommunalt avfall, och det är därför som vi måste agera.
Mitt hemland är ett av de värsta exemplen när det gäller avfall.
Nederländerna hyllar vi som det bästa exemplet.
Men vi behöver alla komma ikapp.
Vi behöver alla återvinna mera så att vi uppfyller villkoren i hierarkin.
Vi måste nå målen för materialåtervinning och förebyggande av avfall etc. Jag tror att vi genom denna åtgärd åtminstone slår in på en bättre väg än tidigare med vår slösaktiga ekonomi, vårt slösaktiga samhälle och vår slösaktiga politik.
för PSE-gruppen. - (IT) Fru talman, mina damer och herrar! Det har varit till nytta för mig att Caroline Jackson och kommissionsledamot Stavros Dimas redogjort utförligt för huvuddelarna i denna kompromiss, som jag också stöder.
Låt mig därför framföra några i högsta grad politiska tankar.
Jag är en förhandlare och jag överväger alltid huruvida den kompromiss som nåtts gäller eller inte.
Därför läser jag texterna igen med nya ögon efter den kväll när förhandlingarna har ägt rum.
Det vete gudarna varför förhandlingar alltid ska sluta på kvällen.
Är en överenskommelse som träffats på förmiddagen mindre värd?
Det är också något att tänka på.
Ärligt talat - och det här säger jag till våra kollegor i de gröna och europeiska enade vänstern samt till Karl-Heinz Florenz som jag ser har lagt fram en ändring igen från miljöutskottet med min signatur som jag därför inte kan annat än stödja - ärligt talat, om man tittar på både kompromissen och texterna från miljöutskottet, har vi verkligen nått - och det är till största delen tack vare er, fru Jackson - ett fantastiskt resultat.
Är vi medvetna om att det inte stod någonting om materialåtervinning i kommissionens förslag och sedan i den gemensamma ståndpunkten?
Det fanns ingenting utom ett skäl där man nämnde återvinningssamhället utan att närmare förklara det. Det fanns ingenting!
Nu har vi precisa mål.
Vi har en granskning 2014 då annat material, som inte täcks för närvarande, ska tas med. Vi vet säkert, som kommissionsledamot Dimas just bekräftade, att rättsliga åtgärder kan vidtas mot medlemsstater som inte genomför de åtgärder som planeras för att nå de här målen.
Detta framstår som mycket viktigt för mig.
Det är också mycket viktigt att det äntligen har inletts ett politiskt och rättsligt förfarande som tvingar medlemsstaterna att utarbeta verkliga planer för förebyggande av avfall och att det äntligen har införts en hierarki för bortskaffande av avfall för miljöns bästa i gemenskapens lagstiftning, som är juridiskt bindande och som gör att avfall inte längre bara är ett problem utan även en resurs.
Uppriktigt sagt tror jag därför inte att det, om vi ser till hela vårt ansvar, skulle ligga i de europeiska medborgarnas intresse att förkasta denna kompromiss och gå in i en riskfylld förlikning. I stället skulle processen för att uppnå och inrätta dessa mål, som här har fastställts på ett tydligt och absolut oomtvistligt sätt, hamna i en sorts rysk roulette.
för ALDE-gruppen. - (EN) Fru talman! Med den här texten hoppas vi kunna vända trenden att producera mer avfall än vi återvinner.
Den är resultatet av flera års debatter och tar hänsyn till verkligheten i två huvudgrupper av medlemsstater när det gäller system för avfallshantering, nämligen stater som återvinner avfall och stater som deponerar avfall.
Kompromissen måste ses i ljuset av detta.
För första gången har förebyggande och materialåtervinning fått en central plats i direktivet.
I den här texten skapas dessutom förutsättningar för högre mål så väl som mål för nya avfallsflöden.
Det är en väl avvägd, uppnåbar och realistisk kompromiss.
Vi anser inte att ändringsförslagen i sin helhet utgör någon risk för den övergripande överenskommelsen.
När det gäller biprodukter, som behandlas i artikeln i och i artikeln om avfall som upphört att vara avfall, har de flesta kritikerna invändningar om skenbar återvinning.
Eftersom det ännu inte finns någon internationell enighet i denna fråga är rädslan befogad.
Därför måste det klargöras att kommissionen ska använda riktlinjerna från februari 2007 för att förhindra detta.
Jag skulle verkligen uppskatta om Stavros Dimas kunde lova oss i dag att ett ämne eller föremål bara får föras ut ur EU som biprodukt om man först uppfyllt villkoren i artikel 4.1 i EU.
Samma sak gäller för avfall som upphört att vara avfall.
När avfall upphör att vara avfall ska det få föras ut ur EU först när villkoren i artikel 5 har uppfyllts i EU.
Detta skulle göra det lättare för parlamentsledamöterna att rösta för kompromissen.
Sammanfattningsvis vill jag framföra mitt tack till föredraganden och skuggföredragandena för deras fruktbara samarbete som gynnar medborgarna i Europa.
för Verts/ALE-gruppen. - (EN) Fru talman! Jag vill också tacka Caroline Jackson.
Visserligen kan vi ha varit oeniga om skatten, men jag tycker inte det råder något tvivel om att samarbetet har fungerat utmärkt diskussionerna igenom.
Jag önskar att vi vore nöjda i dag, men det är vi inte, och jag vill framföra några av skälen till varför vi inte är nöjda med kompromissen.
Vi har gett vårt stöd till 30 av kompromissändringsförslagen, och vi har lagt fram andra för att försöka stärka kompromissen inom områden som farligt avfall, avfall som upphör att vara avfall, biprodukter och separat insamling av biologiskt avfall.
Men de viktigaste frågorna för oss var redan från början att anta bindande mål för avfallsminskning och materialåtervinning och att invända mot omklassificeringen av förbränning som energiåtervinning.
I den slutliga kompromissen finns inga bindande mål för avfallsminskning.
En undersökning om förebyggande av avfall är inget alternativ till stabiliserande åtgärder. Det är ohållbart att avfallet fortsätter att öka i omfattning, och utan denna åtgärd kommer det bara att fortsätta växa.
Även om målen för materialåtervinning och återanvändning har fastställts till 50 procent respektive 70 procent och medlemsstaterna är skyldiga enligt lag att införa åtgärder för att nå dessa mål, är målen i sig inte bindande.
Jag är tacksam för den förklaring som vi har fått av Stavros Dimas, men varför blev det en sådan debatt om formuleringen av detta?
Det var för att man ville undvika att göra de här målen bindande.
Det finns enorma möjligheter att återanvända och återvinna tillverknings- och industriavfall, men detta har utelämnats helt och hållet.
Förbränning får inte ses som ett avfallshanteringsalternativ jämbördigt med materialåtervinning och återanvändning. Det kommer bara att locka fram fler investeringar i förbränningsanläggningar och direkt undergräva avfallshierarkin.
Om den här svaga kompromissen godkänns har vi gått miste om tillfället att säkerställa verkligt agerande och ledarskap inom EU:s avfallspolitik nu när vi i allra högsta grad behöver det.
för GUE/NGL-gruppen. - (GA) Fru talman! Jag vill tacka Caroline Jackson för hennes insatser.
Vi har arbetat mycket bra tillsammans för att förbättra kommissionens ursprungliga förslag, även om vi inte är överens om allt.
Många människor i hela unionen är oroliga för att förbränningsanläggningar ska omklassificeras i förslaget som en form av återvinning om de uppfyller vissa effektivitetskriterier.
Vi är fortfarande emot omklassificeringen av förbränningsanläggningar och har lagt fram ett ändringsförslag för att få detta borttaget.
I den senaste överenskommelsen om materialåtervinning fastställs mål som kan vara mycket svåra att införa på grund av den vaga formuleringen om att medlemsstaterna ska vidta de åtgärder som är nödvändiga för att se till att nå målen för materialåtervinning.
En god lagstiftning kräver att vi preciserar målen bättre och inte överlämnar tolkningen till EG-domstolen.
Därför vill vi försvara och behålla den formulering som röstades fram i utskottet.
Förslagen om förebyggande av avfall har försvagats till den grad att de i inte kommer att kunna vara en tillräcklig hjälp för medlemsstaterna när de ska stabilisera och minska sitt avfall.
Bristen på hänvisning till mål för förebyggande av avfall innebär att lagstiftningen varken innehåller något initiativ till eller några indikatorer för en harmonisering av förebyggande av avfall.
Följaktligen kan vi vara medundertecknare till en del av det arbete vi har utfört tillsammans.
Vi anser emellertid att vi måste lägga fram ändringsförslag till vissa andra delar.
Jag vill än en gång tacka Caroline Jackson för att hon kommunicerat på ett så öppet och inbjudande sätt med skuggföredragandena.
(Applåder)
för IND/DEM-gruppen. - (NL) Fru talman! Utskottet för miljö, folkhälsa och livsmedelssäkerhet har utarbetat en utomordentlig rapport som andrabehandlingsrekommendation.
Då menar jag särskilt sättet att framhålla avfallshierarkin, förkastandet av kategorin biprodukter, den noggranna behandlingen av konceptet för avfall som upphört att vara avfall, skyddsreglerna för farligt avfall samt målen för förebyggande, återanvändning och materialåtervinning.
Den enda negativa aspekten av rapporten från miljöutskottet är det ändringsförslag som stimulerar till förbränning av avfall genom att förbränningen betraktas som effektiv användning om man bara återvinner tillräckligt med energi.
I det resultat av förhandlingarna som vi har nått på två månader finns inte så mycket kvar av rekommendationen från miljöutskottet, och det beror inte på föredraganden utan på rådets kompromisslösa hållning.
Artikeln om biprodukter har inte ändrats och medlemsstaterna kan besluta på egen hand när avfall upphör att vara avfall med allt vad detta innebär i fråga om snedvridning av konkurrensen.
Dessutom har man inte fastställt några mål för förebyggande av avfall, och målen för återanvändning och materialåtervinning är åtskilligt försvagade.
Det är därför som jag inte stödjer kompromisspaketet.
Men jag hoppas att vi ändå kan anta de bättre delarna i rapporten från miljöutskottet när vi röstar i morgon.
Då tänker jag särskilt på ändringsförslagen från GUE/NGL-gruppen och de gröna.
För miljöns bästa är det viktigt att vi går igenom ytterligare ett förlikningsförfarande, då vi faktiskt får rådet att förbättra det som behövs.
Om vi som parlament är övertygande borde det vara möjligt att under ledning av Caroline Jackson åstadkomma mer än i nuläget.
Jag vill tacka Caroline Jackson och skuggföredragandena för deras utmärkta samarbete, och jag hoppas att morgondagens omröstning ger ett framgångsrikt resultat.
(IT) Fru talman, mina damer och herrar! Jag välkomnar och stödjer de ändringsförslag med vilka man avser att införa riktmärken, som är oumbärliga för förebyggande av avfall när det gäller förbättrad materialåtervinning.
Naturligtvis stödjer jag även att man insisterar på en tydligt definierad och tydligt strukturerad avfallshierarki.
Det är också absolut nödvändigt att kunna hänvisa till solida och jämförbara statistiska uppgifter om man ska kunna göra ytterligare framsteg inom förebyggande och materialåtervinning av industriavfall.
Jag anser att vi i parlamentet måste stå fast vid att avfallshierarkin ska tillämpas som en generell regel, och inte som en vägledande princip enligt rådets önskemål.
Det måste framgå klart och tydligt i direktivet vilka kriterier som ska användas för de eventuella avvikelser som man enligt min uppfattning måste ringa in på ett ordnat och tydligt sätt där det behövs, så att det inte råder några tvivel om vad som räknas som återvinning och vad som räknas som bortskaffning av avfall.
Jag håller med föredraganden om att energi från avfallsanläggningar kan spela en viktig roll för hanteringen av hushållsavfall och att vi nu står inför ett viktigt avgörande när det gäller detta med tanke på att EU är beroende av osäker import av energi från så många andra håll i världen.
Jag avslutar med att säga att jag också välkomnar de ändringsförslag som rör regenereringen av spilloljor, som till en början hade uteslutits.
(DE) Fru talman, herr kommissionsledamot, kära fru Jackson!
Jag är missnöjd med kompromissen, men jag är inte missnöjd med min kollega Caroline Jacksons sätt att sköta förhandlingen, utan för en gångs skull, herr kommissionsledamot, är jag missnöjd med kommissionen.
När det gäller flygplan, industri och motorfordon är kommissionen utomordentligt sträng och köpslår för varje grams minskning av koldioxidutsläppen, och det är helt riktigt.
Men när det gäller avfallspolitiken spelar koldioxiden inte alls någon roll.
Det finns uppgifter som tyder på att vi skulle kunna minska koldioxidutsläppen med 100 miljoner ton.
Det är jättechans som försuttits i det här dokumentet.
Det andra skälet till att jag beklagar kompromissen är att vi har blivit en sorts betongföretag.
Vi cementerar skillnaderna i Europa i stället för att rikta in oss på harmonisering.
Visserligen definierar vi mål men de är inte bindande.
Under de kommande 20 åren får vi inga egentliga harmoniserade mål i Europa.
Det är detta som stör mig i den här rapporten.
Tjugo år är nästan en halv generation.
Här borde vi ha varit mycket mer innovativa, och det hade vi också kunnat vara.
Enligt min uppfattning, herr kommissionsledamot, finns det bara ett stort problem, nämligen artikel 14.
Jag skulle uppskatta om ni kunde säga lite mer om den bestämmelsen.
Det må vara en mycket komplicerad fråga i en federal stat.
Det handlar om frågan om blandat eller icke blandat avfall och hur det hanteras i enlighet med principen om att varje land ska ta hand om sitt eget avfall.
Jag ber er vänligen att ännu en gång yttra er i denna fråga i era kommentarer.
Naturligtvis finns det för närvarande en eller annan som säger att vi får en stor majoritet. Men om de här frågorna inte är utredda kommer en del stora länder säkerligen att våndas inför omröstningen.
Jag ber er tänka på att vi ju inte bara har morgondagens behandling. Vi har ju också en tredje behandling, och det är ganska mycket med 64 ändringsförslag i ett förlikningsförfarande.
Så om ni tar tillfället i akt, herr kommissionsledamot, att förklara ett och annat i dessa olösta frågor, skulle jag tro att vi till slut når ett gott resultat.
(EN) Fru talman! I Europa återvinner vi för närvarande bara 27 procent av vårt avfall och nästan hälften av vårt avfall slutar i deponier.
Det här visar att vi måste förändra vår avfallshantering i grunden.
Det viktigaste är att stimulera till förebyggande av avfall, stärka återanvändning och materialåtervinning samt minimera mängden deponerat avfall.
Därför välkomnar jag att avfallshierarkin fick vara kvar i den nya kompromissen efter diskussionerna.
När det gäller förebyggande, som är lagstiftningens huvudsyfte, saknar jag stabiliseringsmålen i den senaste texten, men vi hade redan antagit dem vid första behandlingen.
I de gamla medlemsstaterna genererar en person nästan dubbelt så mycket hushållsavfall, 570 kg per år, som en person i de nya medlemsstaterna, 300-350 kg per år.
De rika länderna borde därför börja minska sin avfallsgenerering först.
Mängden avfall ökar om man ser till hela Europa. Därför räcker det inte med de program för förebyggande av avfall som föreslås i kompromissen.
Vi måste slå fast bindande mål för att stoppa den växande avfallsmängden. Det är därför som jag överväger att stödja ändringsförslag 48 som återinför stabiliseringsmålet för avfall.
Jag välkomnar det obligatoriska målen för återanvändning och materialåtervinning, men jag är rädd att den nya texten, enligt vilken medlemsstaterna "ska vidta de åtgärder som är nödvändiga" för att nå målen, inte räcker till.
Vi behöver konkreta, genomförbara och bindande mål både för hushålls- och industriavfall.
Därför föreslår jag att vi stödjer ändringsförslag 82 för att se till att målen för materialåtervinning drivs igenom.
Nu när jag har framfört de här kommentarerna välkomnar jag rapporten och insatserna från Caroline Jackson, min vän Guido Sacconi med flera.
(EN) Fru talman! Den här överenskommelsen blir inte bättre än så här, säger föredraganden, och det hon har åstadkommit är berömvärt.
Klockan tre på natten under en förlikning går det att göra framsteg som inte hade varit möjliga vid andra tillfällen under förhandlingsprocessen.
Vi är alla överens om att sopberget måste bli mindre.
Från en brittisk butikskedja meddelade man nyligen att man till år 2012 avser att minska förbrukningen av förpackningar med 25 procent och förbrukningen av påsar med 33 procent.
I butikskedjan vill man också se till att livsmedelsavfall omvandlas till energi genom anaerob biologisk nedbrytning.
Dessutom vill man begränsa antalet material som finns i förpackningar till fyra, vilket gör förpackningarna lättare att återvinna eller kompostera, och man vill trycka enkla symboler på alla förpackningar för att underlätta för konsumenterna att återvinna eller kompostera sitt avfall.
Allt detta är nu en fråga om politisk vilja.
Att minska avfallet är en fråga om politisk vilja och den kan stärkas genom EU:s lagstiftning.
Jag misstänker att vi åtminstone kunde ha fått rådet att gå med på att offentliggöra förslag till avfallsminskning några år tidigare än 2014.
Parlamentet har skött sig bra.
Men kanske kunde det har gjort ännu bättre ifrån sig.
(DE) Fru talman, mina damer och herrar! Förslaget är en besvikelse.
Det är näst intill ett misslyckande när det gäller att möta behovet av insatser för att skydda klimatet och spara resurser.
Vi vet att Europeiska miljöbyrån har förutspått att mängden avfall kommer att öka med 50 procent till 2020.
I detta perspektiv är det ett uppenbart misslyckande att man gett efter för medlemsstaternas påtryckningar och inte lyckats faställa bindande mål för stabilisering och materialåtervinning.
Detta har klart och tydligt urholkat det förslag som hade behövts.
Det är också en besvikelse att förbränningen av avfall i allt högre grad blir den sista utvägen, medan förebyggandet av avfall hamnar i bakgrunden.
Det var just för att återställa balansen som vi hade behövt dessa kvoter för materialåtervinning och denna stabilisering av avfallsmängden.
Jag hoppas att vi fortfarande kan förbättra förslaget genom att anta ändringsförslagen och verkligen göra det som behövs, nämligen forma den ambitiösa avfallspolitik som vi behöver i EU.
(IT) Fru talman, mina damer och herrar! Jag beklagar, men jag måste kritisera några av kompromisserna, eftersom de i vissa fall riskerar att undergräva det som parlamentet helt riktigt röstade för vid första behandlingen.
Det är också beklagligt att dessa ändringar till det sämre har införts av rådet och är missriktade och farliga.
Jag säger det här av egen erfarenhet, eftersom jag bor i Italien.
Italien är i det här fallet tyvärr ett exempel på dålig avfallshantering med bristande respekt för gemenskapslagstiftningens anda och bokstav. I gemenskapslagstiftningen finns det ju sedan en tid tillbaka en rättmätig hierarki från minskning till materialåtervinning.
Denna hierarki måste stärkas genom kvantifierade och angivna mål för minskning och materialåtervinning även när det gäller industriavfall. Den får inte försvagas, vilket i viss utsträckning har skett, för att lämna utrymme för en bortskaffningspolitik som undergräver grundtanken med hierarkin.
I Italien har man under de senaste åren till exempel erbjudit miljarder euro som incitament för förbränning av avfall med följder som är uppenbara för alla och som inte på något sätt kan ses som positiva.
(EN) Fru talman! I hela Europa kämpar medlemsstaterna med skenande energipriser.
Därför är det både klokt och nödvändigt att betrakta avfall som ett potentiellt viktigt bränsle.
Det är säkerligen en situation som gynnar alla parter om vi både kan hantera våra stora avfallsmängder och skapa en alternativ källa för energitillförsel, särskilt eftersom vi står inför en energikris och ett ökat beroende av osäker tillförsel av importerad olja.
Därför förstår jag inte att vissa är så förbehållsamma när det gäller att inse det fördelaktiga i att främja energi som utvinns ur avfall.
Jag befarar att vissa kollegor är så starkt bundna vid sina dogmer för materialåtervinning och mot förbränning att de skulle gå miste om tillfället att utvinna värme och el från avfall.
Jag måste säga att jag tror att de har alldeles fel.
I samband med detta kan jag säga att jag tydligt föredrar en maximering av definitionen av "återvinning" i direktivet och att man gör det obestridligt klart att energi från avfall är återvinning och inte bortskaffning av avfall.
Vi borde tillämpa det här särskilt på jordbrukssektorn, där det finns en stor potential.
(FR) Fru talman! Först vill jag framföra ett varmt tack till föredraganden, Caroline Jackson, för hennes utomordentliga arbete som visar prov på hennes gedigna kunskaper inom det känsliga området avfallshantering.
Jag vill också gratulera henne till att hon lyssnat så uppmärksamt under hela förhandlingsskedet. Tack vare detta har vi nått den här svåra kompromissen med rådet och kommissionen.
Vi har ett nytt direktiv med strävan efter att klargöra ett antal punkter.
Vi välkomnar avfallshanteringen och hierarkin och de ambitiöst satta materialåtervinningsmålen för medlemsstaterna, som är 50 procent för hushållsavfall till år 2020.
Avfallshantering måste bygga på förebyggande, återanvändning, materialåtervinning, återvinning och till sist bortskaffning, och denna hierarki måste vara en vägledande princip.
Det är också viktigt att energieffektivitetskriterier införs för förbränningsanläggningar, enligt vad som står i texten, naturligtvis under förutsättning att förbränning endast sker när det inte går att använda någon annan metod.
Mot bakgrund av detta är det mycket positivt att man med den här texten också tillför en mycket noggrann kontroll av farligt avfall och strängare spårningsåtgärder.
Det är förstås en kompromiss och vi önskar att vi hade kommit mycket längre på vissa punkter, exempelvis när det gäller att lägga till miljökriterier i definitionen av återvinning och ställa upp strängare villkor för avvikelser från vad som är avfall och inte. Sedan har vi frågan om biprodukter, som det är problematiskt att definiera.
Hur som helst måste vi absolut stödja den här kompromissen. Vi vet mycket väl att det har varit svårt att komma fram till den, och om vi vill gå vidare till förlikning skulle vi löpa risken att förlora och orsaka enorma förseningar i dessa ärenden.
Vår gemensamma avfallspolitik har hittills varit ett misslyckande, och vi måste inse att det är mycket bättre komma överens om en rimlig lösning, och Europeiska kommissionen måste bevaka mycket noggrant att detta direktiv genomförs ordentligt.
Vi får se om vi kan komma längre om några år.
(FR) Fru talman, herr kommissionsledamot, mina damer och herrar! För egen del är jag varken nöjd med formen eller innehållet i den här kompromisstexten.
När det gäller formen tycker jag inte att vi har gjort vårt jobb ordentligt när vi efter att ha ägnat två år åt att utarbeta en text får veta att de slutliga besluten, som är mer än bara ändringar, har fattats i det tysta och skiljer sig markant från vad som antogs i miljöutskottet och kommer ledamöterna till handa bara några timmar före omröstningen.
När det gäller innehållet är den här kompromisstexten en undanflykt i vilken man inte lyckas ge någon tydlig definition av återvinning, inte längre försöker stabilisera avfallsmängden och inte längre sätter upp några ambitiösa mål för materialåtervinning. Texten är tyvärr ett exempel på kommissionens och rådets oförmåga att överföra de högst ambitiösa tillkännagivanden som görs i europeiska och internationella sammanhang till handling.
Nej, jag är inte nöjd, och jag är faktiskt orolig för vår politiska oförmåga att verkligen agera för miljön och för att förbättra folkhälsan, vilket också är ett skäl till att jag har röstat emot texten.
(FR) Fru talman, herr kommissionsledamot, mina damer och herrar! Till att börja med skulle jag vilja ha gratulera vår föredragande Caroline Jackson, och ALDE-gruppens föredragande Mojka Drčar Murko, till det fina arbete som ni har utfört.
Frågan om farligt avfall omfattar viktiga frågor som spårbarhet, icke-utspädning, harmoniserad lagring av information om avfallsrörelser under lång tid, dvs. fem år för alla delar i kedjan. Trots detta har ingen av dessa frågor behandlas särskilt ingående.
Detta är beklagligt, både för människors hälsa och för miljöns skull.
Jag är mycket besviken när det kommer till biprodukter. Jag är inte emot själva biprodukterna.
Tvärtom inser jag deras betydelse. Men jag anser att det sätt som de definieras på i rådets gemensamma ståndpunkt inte ger tillräckliga garantier och att själva begreppet i slutändan riskerar att missbrukas så mycket att det blir värdelöst.
Andra frågor, exempelvis när avfall upphör att vara avfall och återvinning av avfall, verkar ha offrats för att nå en överenskommelse vid andra behandlingen.
(DE) Fru talman, herr kommissionsledamot, fru Jackson! Vi kommer att lägga fram ett partiöverskridande ändringsförslag som stöddes av en majoritet hör i kammaren vid första behandlingen.
Det tar upp följande problem: I många EU-länder ges obehandlat, osteriliserat matavfall till djur eller dumpas.
Om och om igen riskerar detta beteende att sprida sjukdomar som mul- och klövsjuka.
Därför är det viktigt att se till att matavfall steriliseras och avfallshanteras på ett säkert sätt av godkända bolag och med hjälp av lämpliga metoder.
Medlemsstaterna bör endast kunna tillåta att det används för att utfordra grisar om det har steriliserats i 20 minuter vid en temperatur på 133°C och ett tryck på 3 bar, och om alla övriga villkor i förordning 1774/2002 till fullo har uppfyllts.
Jag är övertygad om att om parlamentet antar detta ändringsförslag kommer rådet att införliva denna regel i kompromissen.
(IT) Fru talman, mina damer och herrar! Den kompromiss som har nåtts är ett steg tillbaka jämfört med den text som antogs i miljöutskottet.
I ursprungstexten angavs det att avfallsproduktionen skulle minska till 2009 års nivåer från och med 2012. Dessutom infördes en ordentlig politik med förebyggande åtgärder som successivt skulle skärpas.
Detta mål har försvunnit i kompromissen, till förmån för vaga skrivningar.
Miljöutskottet hade fastställt minimimål för materialåtervinningen av hushålls- och industriavfall, som skulle nås vid en fastställd tidpunkt - om än långt i fram i tiden.
Även dessa mål har urvattnats. Nu begränsas de till endast vissa typer av material och industriavfall exkluderas.
En annan negativ aspekt är att förbränningsanläggningar över en viss effektivitet gynnas från anläggningar för bortskaffande till återvinningsanläggningar.
Direktivet tycks böja sig för mäktiga lobbyister.
Resultatet i den irländska folkomröstningen har visat att man antingen är på medborgarnas sida, och delar deras oro, eller så riskerar man att EU-tanken förkastas och integrationsprocessen paralyseras.
Parlamentet måste hörsamma de tusentals e-postmeddelanden från EU-medborgare som kräver större engagemang och bindande mål. Annars riskerar vi att gå miste om en utmärkt möjlighet att öka EU-institutionernas trovärdighet.
(HU) Tack så mycket fru talman!
Jag välkomnar kompromisspaketet. Men samtidigt skulle jag vilja understryka hur skör kompromissen är.
Därför är det oerhört viktigt att alla medlemsstater visar ansvar och inte börjar leta efter eventuella kvarvarande kryphål i lagstiftningen.
I Ungern står sorterade sopor för närvarande för 2 procent av den totala avfallsmängden.
Det finns inte mer att säga om det än att hoppas att direktivet kommer att göra att situationen förbättras och att denna låga siffra kommer att öka.
I Östeuropa har investeringarna i avfallshantering ökat de senaste åren, mycket tack vare det strukturpolitiska föranslutningsinstrumentet (ISPA) och Sammanhållningsfonden.
Byggandet av deponier har varit en viktig verksamhet. Men i en rad samhällen har man inlett sopsorteringsprogram, inklusive i vissa fall åtgärder för separat insamling av organiskt avfall.
Å andra sidan har vi inte alls sett några verkliga åtgärder eller investeringar i syfte att minska avfallsmängden och vi väntar fortfarande på en särskild industri för bearbetning av återvunnet material.
Inte minst för Ungern kommer därför EU:s riktlinjer att bli oerhört viktiga.
Enligt statistiken skulle varje samhälle i princip minska sin avfallsmängd med 50 procent så snart det inför pappersåtervinning och separat insamling av organiskt avfall vid dörren.
När vi inför nya skyldigheter måste vi emellertid även ta hänsyn till deras genomförbarhet och de kostnader som är kopplade till dem.
Kan exempelvis ytterligare investeringar göras på samma områden som ISPA-projekt?
Kan de ursprungliga kontrakten ändras?
Om så inte är fallet spelar det mindre roll om det finns en efterfrågan på mer sopsortering eller om det finns lagstiftning på plats för att minska den mängd avfall som deponeras. Enligt de 20-åriga kontrakten måste det insamlade avfallet köras till de deponier som har byggts.
Förutom att anta detta direktiv måste vi därför utan dröjsmål börja arbeta på hur vi kan ändra de befintliga kontrakten.
Jag gratulerar föredraganden till hennes fantastiska arbete.
Tack så mycket.
(DE) Fru talman! Jag tycker vi kan gratulera föredraganden.
Hon har verkligen lyckats nå en godtagbar kompromiss med rådet.
Jag vill framför allt betona inkluderandet av en avvikande avfallshierarki.
Det finns emellertid sämre bitar, som är helt obegripliga och som rådet har infört i dokumentet.
Det handlar bland annat om animaliska biprodukter.
I utskottet hade vi kommit överens om att animaliska biprodukter skulle strykas från detta ramdirektiv om avfall.
Nu har rådet uppfört ett slags byråkratiskt hinder som kommer att leda till protester från jordbrukarna.
Det fastställs att flytgödsel som förädlas till biogas plötsligt blir en avfallsprodukt.
Förstår ni vad detta betyder?
Det betyder att jordbrukare måste ha en avfallshanteringslicens och kommer att bli tvungna att precisera exakt hur mycket avfall och vilken typ av avfall som ska hanteras, och var hanteringen ska ske.
I förordningen om animaliska produkter anges det uttryckligen att flytgödsel ska undantas.
Nu blir det istället enklare för jordbrukaren att sprida flytgödsel på åkrarna än att förädla det till biogas.
Vi skapar med andra ord byråkratiska hinder som försvårar en verksamhet som vi faktiskt uppmuntrar.
Den andra punkten rör spilloljor.
I direktivet om spilloljor - som nu ska upphävas - anges att spilloljor ska behandlas och regenereras.
Stora volymer behandlas i enlighet med detta direktiv.
Det har redan tidigare konstaterats att spilloljor inte behöver regenereras när detta inte är ekonomiskt försvarbart eller tekniskt omöjligt.
Nu fastställs det att det är upp till medlemsstaterna att avgöra detta.
Är vi verkligen en europeisk union eller har vi gått tillbaka till att vara en samling medlemsstater?
Vi styckar helt klart upp marknaden igen.
Det gör mig mycket besviken.
Låt mig gå vidare till frågan om självförsörjning.
De lokala myndigheterna ska nu avgöra vem som får göra sig av med vad och när.
Självklart förekommer det kraftiga påtryckningar från lokala myndigheter med förbränningsanläggningar med överkapacitet.
Detta är emellertid fel väg att gå.
Det är inget alternativ och denna utvidgning får marknadsekonomin att helt sluta fungera på avfallshanteringsområdet.
(NL) Fru talman! Denna kompromiss är helt klart ett betydelsefullt fall framåt för EU:s miljölagstiftning.
Samtidigt är jag inte helt nöjd med kompromissen.
Varför inte?
Min egen region, Flandern, tillsammans med exempelvis Nederländerna, har den bästa avfallspolitiken och är fantastiskt duktig på sopsortering och materialåtervinning. Vi tycker därför att de föreslagna sopsorterings- och materialåtervinningsmålen är totalt inadekvata.
De uppmuntrar oss verkligen inte alls till att bli bättre i framtiden.
Vi är inte heller helt nöjda med att förbränningsanläggningar för hushållsavfall ska kunna betraktas som effektiv användning på grundval av energieffektivitetsformeln. I praktiken tror vi att detta kommer att skapa en hel del förvirring.
När allt kommer omkring är jag säker på att det samlade resultatet måste ses som mycket positivt. Jag vill därför tacka Caroline Jackson så mycket för hennes stora bidrag.
Vi ställer oss bakom kompromissen.
(HU) Fru talman! I sin nuvarande form försvårar tyvärr ramdirektivet om avfall en ökad användning av biogas.
Jag håller helt med vår kollega Horst Schnellhardt från PSE-DE-gruppen om att det nuvarande direktivet är helt inadekvat när det gäller biogasproduktion, och även när det gäller användningen av flytgödsel eller kommunalt avfall.
I sin nuvarande form kommer avfallsdirektivet tyvärr att försvåra en utökad användning av biogas.
Det gör att man måste ifrågasätta Caroline Jacksons betänkande.
Inom ramen för avfallsdirektivet är definitionen av stallgödsel som används för framställning av biogas tvetydig.
Om direktivet syftade till att inkludera detta skulle det bli omöjligt att framställa biogas från stallgödsel, trots att detta skulle ha stora fördelar för energieffektiviteten, miljön och klimatskyddet.
Vi måste skapa ordning och reda på detta område och så snabbt som möjligt se till att vi åter får en konsekvent lagstiftning. När det gäller biogas måste vi därför anta kommissionens ståndpunkt om direktivet.
(PL) Fru talman! Jag gratulerar föredraganden till en realistisk bedömning av det växande avfallsproblemet.
Grundantagandena i de föreslagna bestämmelserna är att förhindra att avfall uppstår och materialåtervinning.
Energiåtervinning är enklare, men bör inte ersätta den svårare materialåtervinningen.
Därför är det nödvändigt att skapa bra villkor som möjliggör materialåtervinning och mer exakta lagstiftningsdistinktioner, exempelvis när metallskrot inte längre ska betraktas som avfall utan som råmaterial.
Vi behöver bättre och billigare materialåtervinningstekniker.
Produkter ska utformas så att de blir lättare att återvinna.
Avfallet måste sorteras och sorteringen måsta anpassas till marknaden på ett sätt som gör att både hushållen och potentiella användare av det återvunna materialet gynnas.
Utan dessa lösningar riskerar vi att upprepa den nuvarande situationen i Neapel, där tyvärr förbränning av avfallet kan visa sig vara den enda lösningen.
ledamot av kommissionen. - (EN) Fru talman! Jag skulle vilja tacka alla talare i debatten för deras positiva bidrag.
På grundval av den text vi har enats om kommer medlemsstaterna nu att göra en rad ändringar för att förbättra sin avfallshantering.
I direktivet fastställs tydliga definitioner och principer för avfallshantering och jag är säker på att detta kommer att lösa de nuvarande tolkningsproblemen, minska antalet mål vid domstolarna och lägga en bra grund för en väl fungerande avfallshanteringssektor.
Några centrala element har inkluderats i det övergripande kompromisspaket som nu föreslås.
De viktigaste är följande:
För det första finns det nu ett klart och ambitiöst miljömål i direktivet.
Graden av miljöskydd har inte bara bibehållits utan i flera fall ökat, exempelvis i samband med farligt avfall.
Medlagstiftarna har enats om flera grundläggande definitioner, inklusive definitioner av avfall, förebyggande åtgärder, materialåtervinning och återvinning.
Definitionerna är tydliga och lätta att förstå.
Dessutom införlivas bestämmelser från två andra direktiv i direktivet för att göra lagstiftningen mer tillgänglig och samtidigt se till att en hög grad av miljöskydd bibehålls.
Man gör en tydlig skillnad mellan återvinning och bortskaffande och kommissionen ges möjlighet att göra distinktionen ännu tydligare om detta skulle behövas.
En tydlig avfallshierarki i fem steg har införts. I denna främjas förebyggande åtgärder och bortskaffande av restavfall ska bara användas som en sista utväg.
Samtidigt ges tillräckligt med flexibilitet för att man ska kunna ta hänsyn till motiverade livscykelöverväganden.
Jag skulle vilja upprepa den vikt som parlamentet under förhandlingarna lade vid att stärka de högre nivåerna i avfallshierarkin genom att införa materialåtervinningsmålen.
Om dessa mål inte har uppfyllts 2020 kan domstolen väcka talan mot medlemsstater för underlåtenhet att uppfylla kraven i direktivet.
Genom den nya skrivningen införs dessutom en mer regelbunden och omfattande process för att övervaka de åtgärder som medlemsstaterna vidtar för att uppfylla målen redan före fristen 2020, i stället för en ren kontroll av att nivåerna verkligen har uppfyllts 2020 när det redan finns befintliga avfallshanteringssystem.
Tack vare ett sådant förfarande med tidiga kontroller kan man undvika obehagliga överraskningar 2020.
Sist men inte minst införs en helt ny dimension på avfallshanteringsområdet i och med detta direktiv. Detta är något som kommissionen gärna går vidare med så snart direktivet har antagits och införlivats.
Det överlåts nu åt medlemsstaterna att fastställa sina nationella planer och nät för avfallshantering. Dessa måste spegla de principer och nya skyldigheter som anges i det reviderade direktivet.
I artikel 14 i ramdirektivet om avfall anges inte om privata eller offentliga myndigheter ska inrätta eller driva sådana nät. Det sägs inte heller något om avfallshanteringen eller avfallsanläggningarna ska vara privat eller offentligt ägda.
Ansvarsfördelningen mellan den privata och den offentliga sektorn kan endast avgöras av medlemsstaterna.
Om det redan finns ett adekvat nät av anläggningar för bortförskaffande och återvinning av avfall - oavsett om detta är privat, offentligt eller en blandning av båda - behöver man inte vidta ytterligare åtgärder.
När det gäller oron för att det saknas materialåtervinningsmål för avfall från tillverkningsindustrin och annat industriavfall kommer kommissionens tjänsteavdelningar att prioritera en undersökning av om det går att fastställa sådana mål inom ramen för översynen 2014, vilket föreskrivs i artikel 8a (punkt 4).
När det gäller frågan om att utfordra djur med animaliska biprodukter som matavfall regleras detta i förordningen om animaliska biprodukter. Även denna är föremål för översyn just nu.
Frågan bör tas upp i den förordningen eftersom ramdirektivet om avfall inte är rätt forum för att reglera hur matavfall används.
På frågan om biproduktskrav och slutavfallskriterier måste uppfyllas i EU innan leverans till tredjeland kan kommissionen bekräfta att så är fallet.
På frågan om stallgödsel ska undantas från räckvidden för ramdirektivet om avfall är svaret att stallgödsel inte betraktas som avfall när det används som gödsel.
Det betraktas emellertid som avfall när det är avsett att bearbetas ytterligare eller bortskaffas, exempelvis genom förbränning, framställning av biogas eller kompostering och deponering.
Om vi skulle undanta stallgödsel från avfallslagstiftningens räckvidd skulle detta leda till en allvarlig lucka i miljöskyddet eftersom vi skulle sakna rättsliga medel för att kontrollera frågor som utsläpp i luft och vatten, deponeringskrav, buller, lukt etc.
Avslutningsvis bör EU främja framställningen av biogas och kompostering av avfall.
Men biogas- och kompostanläggningar är inte miljöneutrala.
Även dessa anläggningar släpper ut föroreningar i luften och i vattnet och kan vara en källa till störningar, exempelvis genom buller eller dålig lukt.
Att undanta stallgödsel avsett för framställning av biogas eller kompostanläggningar från räckvidden för ramdirektivet för avfall skulle innebära att sådana anläggningar undantas från räckvidden för IPPC-direktivet.
För att sammanfatta skulle jag än en gång vilja gratulera Caroline Jackson till hennes utmärkta arbete.
Kommissionen är mycket nöjd med resultatet av förhandlingarna och kan till fullo godta de föreslagna kompromissändringsförslagen.
föredragande. - (EN) Fru talman! Låt mig kort tacka alla kolleger som deltog i debatten.
Det är bara en kollega som jag vill besvara och det är Chris Davies - hädanefter känd som ”Chris Newsnight Davies”, efter det programs om han tycker om att medverka i - som sa att jag gav med mig för lätt gentemot rådet.
Jag hoppas mina kolleger stöder mig när jag säger att jag inte gav med mig för lätt, och att jag aldrig har gett med mig lätt vad det än har gällt.
Anne Laperrouze kan bekräfta att i vattenfrågan blir rådet svårare och svårare att förhandla med.
När den ekonomiska nedgången börjar få konsekvenser inser rådet att denna lagstiftning kommer att kosta pengar och vill därför inte gärna anta parlamentets ändringsförslag.
Vi har ett val i morgon bitti.
Vi kan säga ja till hela paketet med ändringsförslag, och jag hoppas verkligen att vi gör det.
Vi kan rösta ja till vissa centrala ändringsförslag, exempelvis om biprodukter, vilket innebär att paketet faller och vi går vidare till förlikning.
Hur kul skulle inte det vara?
Eller vi kan säga ja till några mindre ändringar, eller ändringar som de som lägger fram ändringsförslaget anser är mindre, exempelvis ändringsförslag 88 som jag väntar på att kommissionen ska yttra sig över. Yttrandet kanske hinner komma till i morgon.
Jag är mycket tveksam till om rådet kommer att godta några ändringar alls, hur små de än må vara. Jag är därför för hela paketet, utan ändringar.
Paketet måste betyda något. Varför kämpade annars rådet så starkt för det?
Det är inte något meningslöst paket som De gröna vill få det till. Det är ett paket med tänder.
Avslutningsvis skulle jag vilja tacka skuggföredragandena - ”Caroline Jackson and the Shadows”, det låter som ett 60-talsband - för deras samarbete, utan att jag för den skull har någon större önskan att se dem om och om igen under förlikningsförfarandet.
Vi borde se till att avsluta denna fråga i morgon.
Debatten är härmed avslutad.
Omröstningen kommer att äga rum i morgon, tisdagen den 17 juni.
Skriftliga förklaringar (artikel 142)
skriftlig. - (DE) Genom det nya ramdirektivet om avfall har parlamentet fått igenom höga och bindande materialåtervinningskvoter.
Det fanns ett akut behov av sådana kvoter och jag ser fram emot när materialåtervinning och sopsortering i allt högre grad kommer att praktiseras i hela EU.
Jag anser att målen om att senast 2020 återvinna 50 procent av hushållsavfallet och 70 % av bygg- och rivningsavfallet är mycket bra mål som har lagt grunden till ett fungerande miljö- och klimatvänligt avfallshanteringssystem i hela EU.
Just på grund av att österrikarna redan är exemplariska när det kommer till sopsortering och materialåtervinning är jag mycket glad att resten av medlemsstaterna nu kommer att delta i denna verksamhet. Härigenom tar vi ännu ett steg mot effektivt miljöskydd.
Vi får inte glömma att avfallsprodukter även är råmaterial och att en effektivare användning av dessa material även kan bidra i kampen mot klimatförändringarna.
Vi måste nu invänta kommissionens specifika förslag om hur vi ska garantera att ekonomisk tillväxt inte leder till större avfallsmängder.
Förberedelser för Europeiska rådets möte efter folkomröstningen på Irland (19-20 juni 2008) (debatt)
Nästa punkt är rådets och kommissionens uttalanden om förberedelserna för Europeiska rådets möte efter folkomröstningen på Irland.
rådets ordförande. - (SL) I morgon inleds Europeiska rådets andra möte under det slovenska ordförandeskapet.
Jag vill gärna redogöra för de huvudsakliga diskussionsämnen som stats- och regeringscheferna kommer att ta upp.
Den första debatten kommer med all säkerhet att ägnas åt att analysera situationen efter folkomröstningen om Lissabonfördraget, som hölls i torsdags på Irland.
Jag vill börja med att återge uttalandet från rådets ordförande Janez Janša: ”Ordförandeskapet beklagar det beslut som fattats av de irländska väljarna och är därför besviket.
Vi kommer självklart att respektera det irländska folket vilja.”
Efter det att det officiella resultatet av folkomröstningen hade offentliggjorts talade Europeiska rådets ordförande med ett antal ledare från de medlemsstater som ännu inte har slutfört ratificeringsförfarandet.
Det är uppmuntrande att veta att dessa medlemsstater är beslutna att fortsätta med ratificeringen.
Som Europeiska rådets ordförande har betonat är Lissabonfördraget absolut nödvändigt för Europeiska unionen och EU-medborgarna, eftersom det leder till ökad effektivitet, mer demokrati och större öppenhet.
Det är ett faktum att de problem och utmaningar som unionen står inför i dag finns kvar.
Det står lika klart att det negativa resultatet av den irländska folkomröstningen inte kommer att bidra till att lösa dessa problem.
Vid morgondagens möte i Europeiska rådet kommer stats- och regeringscheferna att diskutera hur man kan råda bot på denna situation på bästa sätt.
Målsättningen kommer att vara att fastställa en tidsplan för det fortsatta arbetet.
Ordförandeskapet är övertygat om att det är möjligt att finna en lösning i samarbete med Irland, och att situationen från 2005 inte kommer att upprepas.
Vid Europeiska rådets möte kommer vi först och främst att lyssna till Irlands premiärminister (Taoiseach) Brian Cowen, som kommer att förklara omständigheterna kring folkomröstningsresultatet och skälen till resultatet.
Europeiska rådet kommer naturligtvis inte att åsidosätta de andra viktiga utmaningar som vi har framför oss.
EU fortsätter att fungera.
Stats- och regeringschefernas andra stora debatt kommer därför att inriktas på frågan om de stigande livsmedels- och oljepriserna.
Det är ett faktum att de stigande priserna på basvaror har spelat in i den eskalerande inflationen i livsmedelspriserna och den allmänna inflationen inom EU.
Låginkomstfamiljer har drabbats mest direkt av de höga priserna.
Globalt sett är det utvecklingsländerna som är värst drabbade som nettoimportörer av livsmedel.
Det är mycket viktigt att EU spelar sin roll i arbetet med att utforma ett lämpligt gensvar och att EU står enat i sina åtgärder för att hantera konsekvenserna, inte bara med inriktning på de fattigaste segmenten av EU:s befolkning, utan även i utvecklingsländerna.
Därför förväntas Europeiska rådet stödja de nödvändiga åtgärderna inom EU och på internationell nivå.
Jag kommer kortfattat att redogöra för dessa.
EU har redan vidtagit åtgärder för att lätta på trycket på livsmedelspriserna genom att sälja interventionslager, sänka exportbidragen, upphäva kravet på arealuttag för 2008, höja mjölkkvoterna och tillfälligt upphäva importtullarna för spannmål, för att på så vis förbättra försörjningen och bidra till att stabilisera jordbruksmarknaderna.
Med tanke på att det är låginkomstfamiljerna som drabbas hårdast är det helt naturligt att medlemsstaterna planerar kortsiktiga åtgärder för att lindra pressen av de höga priserna särskilt för dem.
Europeiska rådet måste emellertid tänka mer långsiktigt.
Det är egentligen ingen som förväntar sig att livsmedels- eller oljepriserna ska återgå till de tidigare nivåerna inom den närmaste framtiden.
Jag är övertygad om att nästa ordförandeskap i nära samarbete med Europaparlamentet kommer att nå en lämplig överenskommelse om hälsokontrollen av den gemensamma jordbrukspolitiken, som kommer att bestå av åtgärder för att stärka jordbruksproduktionen och garantera en säker livsmedelsförsörjning.
Vi måste även uppmärksamma politiken för biobränslen och hitta ett sätt att garantera deras hållbarhet, både inom EU och i andra länder.
Det kommer att vara viktigt att främja utvecklingen av andra generationens biobränslen.
Mer generellt måste vi fortsätta arbetet med innovation och forskning och utveckling inom jordbrukssektorn för att förbättra effektiviteten och produktiviteten.
Bland de initiativ som vi bör gå vidare med på internationell nivå kommer Europeiska rådet att framhålla unionens bidrag till de globala insatserna för att mildra effekterna av de stigande priserna på dem som lever i fattigdom.
Europeiska rådet kommer bland annat att efterlysa bättre samordning av det internationella gensvaret på den kris som har orsakats av de stigande livsmedelspriserna, särskilt inom ramen för FN och G8-gruppen, stöd till en öppen handelspolitik, snabba reaktioner på omedelbara kortsiktiga humanitära behov och främjande av målinriktat stöd för att stimulera jordbruket i utvecklingsländerna.
Förutom de höga livsmedelspriserna ställs EU inför stigande oljepriser.
Detta kräver en anpassning av EU-ekonomin, och en särskild debatt om den frågan är planerad till i dag.
En ytterligare prioritering för ordförandeskapet är att Europeiska rådet bör se på de åtgärder som har vidtagits för att stärka det europeiska perspektivet för västra Balkan.
Jag vill särskilt betona att en rad stabiliserings- och associeringsavtal har slutförts, dialogen om viseringslättnader för alla länder i regionen har inletts och färdplaner har inlämnats.
Dessutom kommer stats- och regeringscheferna att betona vikten av att involvera alla länder på västra Balkan i regionalt samarbete samt välkomna en rad sektorsavtal.
Västra Balkan är en region som omges av EU-medlemsstater och är därför i stort behov av en bekräftelse på sitt europeiska perspektiv och behöver hjälp med att genomföra reformer.
Ordförandeskapet sätter högt värde på Europaparlamentets stöd i detta avseende.
En annan viktig fråga på dagordningen kommer att vara framstegen mot att nå millennieutvecklingsmålen.
År 2008 är halvtid för tidsgränsen för att nå dessa mål.
Som den största biståndsgivaren är EU medvetet om sitt ansvar och vill spela en aktiv roll för att uppmana världssamfundet att sträva efter att nå millennieutvecklingsmålen.
Europeiska rådet kommer därför att lyfta fram EU:s centrala roll vid internationella konferenser och EU:s åtaganden.
Den tredje uppsättning frågor som ska diskuteras av Europeiska rådet kommer att beröra ekonomiska, sociala och miljömässiga punkter.
Först och främst vill jag ta upp översynen av det arbete som har uträttats med klimatenergipaketet.
Det slovenska ordförandeskapet har nått alla de fastställda målen för detta paket.
Det politiska beslut som antogs vid Europeiska rådets marsmöte var ytterst viktigt.
Europeiska rådet kommer även att ta del av de överenskommelser som nåtts om avregleringen av energimarknaden, som diskuterades i parlamentet i går.
På grundval av slutsatserna från december 2007 kommer Europeiska rådet även att granska de framsteg som har gjorts i viktiga frågor inom områdena migration, rättvisa och terrorism.
Slutligen kommer stats- och regeringscheferna att behandla frågor som rör den europeiska grannskapspolitiken.
Att bygga vidare på och förstärka tidigare framgångar, ”Barcelonaprocessen: en union för Medelhavsområdet” kommer att skapa ytterligare drivkraft i unionens förbindelser med länderna i Medelhavsområdet.
Barcelonaprocessen kommer att komplettera de pågående bilaterala förbindelserna som kommer att fortsätta inom de befintliga politiska ramarna.
Europeiska rådet förväntas välkomna de senaste förslagen om att utveckla ett östligt partnerskap inom ramen för den europeiska grannskapspolitiken.
Under mötet kommer stats- och regeringscheferna även att diskutera kommissionens förslag om Slovakiens anslutning som den sextonde medlemsstaten i Ekonomiska och monetära unionen (EMU) den 1 januari 2009.
Jag vill därför särskilt gratulera Slovakien.
Kort sagt har parlamentets åsikter och debatter bidragit stort till att formulera dagordningen för Europeiska rådets möte.
Den debatt som nu kommer att hållas, och som vi kommer att följa mycket noggrant, kommer också att utgöra ett användbart och viktigt bidrag till diskussionen mellan stats- och regeringscheferna, så jag kommer att lyssna till den med stort intresse.
(Applåder)
kommissionens ordförande. - (EN) Fru talman! Europeiska rådets möte som inleds i morgon har en diger dagordning som omfattar många områden där medborgarna förväntar sig att EU ska agera.
(Några ledamöter till höger, som bar gröna t-tröjor, reste sig för att hålla upp banderoller och affischer med krav på respekt för nejrösten på Irland.
Talmannen uppmanade dem att ta bort banderollerna och affischerna.)
De frågor som ska diskuteras är de plötsliga ökningarna av olje- och livsmedelspriserna, klimatförändringen och energisäkerheten, migration och asyl, för att bara nämna några.
Men det som alla naturligtvis främst tänker på är nejrösten på Irland.
Detta nej till Lissabonfördraget var en besvikelse för alla som vill ha ett starkare, effektivare och mer ansvarsskyldigt EU.
Lissabonfördraget förblir av grundläggande vikt för att vi ska kunna bemöta de utmaningar som Europa ställs inför i dag, att ha en mer demokratisk union, utöka Europaparlamentets befogenheter och erkänna de nationella parlamentens roll i EU-politiken, att stärka EU:s kapacitet att agera på områden som migration, energi, klimatförändringar och inre säkerhet, och slutligen att se till att EU agerar mer samordnat och effektivt på internationell nivå.
Dessa utmaningar har inte försvunnit.
Sanningen är att nejrösten inte löste de problem som det är meningen att fördraget ska bidra till att hantera.
Under de senaste sex åren har vi ägnat mycket energi åt institutionella frågor.
Vi har inte råd att låta den energin gå till spillo med tanke på de många viktiga frågor som kräver snabbt ett agerande i dag, och världen stannar inte och väntar på EU.
Som jag sa förra veckan respekterar kommissionen fullständigt resultatet av den irländska folkomröstningen.
Vi måste nu visa samma respekt för alla nationella ratificeringar ...
(Applåder)
... vare sig de har valt att genomföra folkomröstningar eller parlamentarisk ratificering.
Nitton demokratiska beslut har fattats i processen hittills: 18 för Lissabonfördraget, ett emot.
Åtta andra medlemsstater har ännu inte tagit ställning.
Den irländska regeringen har tydligt förklarat att den respekterar andra länders rätt att fortsätta med sina ratificeringsprocesser.
Det anser jag är en självklar sak.
Alla länder i EU är likvärdiga, alla länder har rätt att uttrycka sin åsikt.
(Applåder)
Det står klart att Lissabonfördraget inte kan träda i kraft innan det råder enhällighet om ratificeringen, men det står lika klart att det irländska valresultatet är ett beslut om Irlands ståndpunkt, och att det inte kan avgöra andra länders ståndpunkter.
Jag förväntar mig att de medlemstater som inte har ratificerat Lissabonfördraget kommer att fortsätta sina egna ratificeringsprocesser.
(Applåder)
Europeiska rådets möte ger oss alla en möjlighet att lyssna mycket noga till vad premiärminister Brian Cowen har att säga.
Sedan måste vi föra ett mycket nära samarbete med den irländska regeringen för att hjälpa till att lösa detta problem.
Jag vill klargöra att Irland har ett ansvar för att bidra till att finna en lösning.
När regeringarna undertecknar fördraget tar de ansvar för att se till att det ratificeras.
Jag vill emellertid att det ska framgå lika klart att det är dags att vi talar allvar om solidaritetsaspekten.
Det var 27 medlemsstater som undertecknade fördraget, och vi måste göra allt vi kan för att se till att alla 27 medlemsstaterna finner en väg framåt.
Alla medlemsstater är lika mycket värda och det måste vi ha klart för oss.
Detta kommer att ta tid och kraft för irländarna, men också för oss alla.
Jag anser att det är viktigt att vi inte fattar några förhastade beslut om nästa steg.
Vi måste ta tid på oss för att finna ett verkligt samförstånd och se vilka möjligheter Irland har.
Men det får inte heller ta alltför lång tid.
Jag vet att det är viktigt för parlamentet att kunna klargöra det framtida agerandet för väljarna i tid till valet till Europaparlamentet.
Europeiska kommissionen är redo att göra sin del - vilket även parlamentet är, det är jag övertygad om - men man kommer inte ifrån det faktum att regeringarna har ett särskilt ansvar i det här avseendet, ansvar för att underteckna fördraget, se till att det blir ratificerat och att främja det europeiska projektet i diskussionerna i den nationella allmänna opinionen.
När det gäller det sistnämnda vill jag generellt påpeka att jag anser att det kan vara bra för den pågående debatten.
Efter att ha utpekat EU-institutionerna som en bekväm syndabock i åratal skapas en stark grogrund för populistiska kampanjer.
(Applåder)
Som jag har sagt flera gånger tidigare kan man inte klaga på Bryssel eller Strasbourg från måndag till lördag och förvänta sig att medborgarna ska rösta för dem på söndag.
(Applåder)
I morgon kommer Europeiska rådet även att betona att nejrösten inte får leda till att EU frestas till institutionellt navelskåderi.
Vi har gjort stora framsteg sedan ett par år tillbaka på grund av våra beslutsamma insatser för att utforma politik i EU-medborgarnas intressen.
Nu när de stigande livsmedels- och oljepriserna leder till stora förväntningar på agerande från EU:s sida har vi inte råd att överge den vägen.
Därför välkomnar jag varmt premiärminister Janez Janšas och det slovenska ordförandeskapets beslut att vika debatten om Lissabon för middagen på torsdag kväll och ägna den övriga tiden av Europeiska rådets möte till att gå vidare med vår politiska dagordning.
I dag känner alla av trycket från prisökningarna på livsmedel och bränsle, men en del har en extra börda.
För de fattigare hushållen utgör dessa kostnader en större andel av hushållsbudgeten, vilket gör att prisökningarna slår ännu hårdare mot dem.
Detsamma gäller vissa ekonomiska verksamheter, eftersom vissa industrier är ytterst beroende av bränsle.
Kommissionen har i två meddelanden om livsmedels- och oljepriserna gjort en noggrann analys av orsakerna till prishöjningarna, om var pressen är starkast och vad vi kan och bör göra.
Vi i EU måste visa att vi vidtar alla åtgärder vi kan på EU-nivå och nationell nivå.
Vi måste analysera de redskap vi har till vårt förfogande på ett dynamiskt och fantasifullt sätt - och fundera över vilka åtgärder som kommer att ha en verklig effekt på kort, medellång och lång sikt.
Vi får inte glömma bort tidigare oljechocker, där EU inte lärde sig de långsiktiga läxorna.
Vi får hoppas att det inte blir likadant den här gången som tidigare, då vi bara fortsatte som vanligt efter alla oljechockerna, och jag hoppas även att vi verkligen lyckas förändra saker och ting den här gången, och förändra mönstret för energiförbrukningen i Europa och i världen.
För att lindra livsmedelsproblemen inom EU kommer vi att lägga fram förslag om att utöka vårt system för livsmedelsdistribution till de mest behövande innan begär en höjning på två tredjedelar av budgeten för detta särskilda område.
Dessutom har EU redskap som kan och kommer att användas. Det handlar om att övervaka priserna, utnyttja våra befogenheter på konkurrensområdet för att kontrollera livsmedelsförsörjningskedjan, öka reserverna och garantera att den gemensamma jordbrukspolitiken är väl anpassad till den nuvarande situationen på jordbruksmarknaden.
När det gäller oljepriserna är omedelbara åtgärder motiverade för att hjälpa de hårdast ansatta hushållen.
Det är emellertid meningslöst att regeringarna använder offentliga medel för att utjämna ökningarna av energipriserna, som med all sannolikhet är här för att stanna.
Vi bör även se på vad som kan göras på EU-nivå inom områden som konkurrens och beskattning.
Kommissionen kommer att lägga fram förslag för att öka insynen i reservlager av olja och kommersiella oljelager.
Vi kommer även att lägga fram förslag om beskattning för att stödja och underlätta övergången till en koldioxidfattig ekonomi, nämligen inom området för energieffektivitet.
Vi kommer vidare att stödja ett högnivåmöte mellan producenter och konsumenter av energi från olja och fossila bränslen.
När det gäller fisket kommer vi att lägga fram ett paket med nödåtgärder för att hantera ekonomiska och sociala problem i syfte att ge medlemsstaterna möjlighet att bevilja kortsiktigt stöd i nödsituationer, och vi kommer att se över reglerna för småskaligt statligt stöd igen.
Jag har tre påpekanden om detta.
För det första måste stödet samordnas för att undvika en våg av nationella initiativ som bara leder till att problemen flyttas runt i unionen.
För det andra måste vi inrikta våra lindringsinsatser på de värst drabbade segmenten av flottan.
För det tredje måste vi finna strukturella lösningar på överkapaciteten inom fiskeindustrin.
De påfrestningar som belastar européerna i dag visar varför EU:s mål för energisäkerhet, energieffektivitet och klimatförändringar är så viktiga för det europeiska samhällets välfärd, och de är därför mer angelägna än någonsin.
Eftersom efterfrågan fortsätter att överstiga tillgången på olja och gas utgör de mål som överenskoms förra året en färdigförpackad lösning för att minska EU:s sårbarhet och den ekonomiska bördan av framtida prishöjningar.
De centrala aspekterna i det paket med förslag som vi har lagt fram och som nu övervägs av parlamentet kommer att utgöra ett avgörande bidrag.
Den grundläggande tanken är att energipriserna sannolikt aldrig kommer att gå tillbaka till de tidigare nivåerna, vilket innebär att vi har ett strukturellt problem.
Vi kan och måste ha kortsiktiga svar för de mest sårbara i våra samhällen. Ett strukturellt problem kräver dock ett strukturellt svar, en strukturell reaktion.
Den strukturella reaktionen är vårt paket för klimatförändring och förnybar energi, att inte vara beroende av fossila bränslen utan i stället främja förnybara energikällor och göra mer när det gäller energieffektiviteten.
Det är den allmänna linje som vi bör följa.
(Applåder)
Därför hoppas jag att de i EU som fortfarande tvivlar på vikten av att förändra våra energimönster och behovet av att bekämpa klimatförändringen till slut, om så inte av dessa anledningar utan på grund av energisäkerheten och behovet av att öka vår ekonomis konkurrenskraft, kommer att inse att vi verkligen måste infria våra åtaganden för klimatförändring och förnybara energikällor.
Den strukturella reaktionen på de strukturella utmaningar vi står inför är i stort sett att spara och diversifiera.
Med spara menar jag att öka energieffektiviteten där vi har en enorm outnyttjad potential.
Diversifiering omfattar både energins källor och geografiska ursprung.
Båda målen handlar om att öka EU:s energisäkerhet.
Det är därför mycket angeläget att vi antar vårt åtgärdspaket för klimatförändring och energisäkerhet.
Europeiska rådets uppgift kommer att vara att ge en signal om detta och förbereda allt för att nå en politisk överenskommelse, senast i december hoppas vi.
Jag anser att det är en viktig uppgift för Europeiska rådet att visa att nejet till Lissabonfördraget inte är en ursäkt för att låta bli att agera.
Det får inte leda till att EU förlamas.
Vi måste visa att vi kommer att finna det rätta sättet för att säkra ett effektivt och demokratiskt fördrag som EU har fått i uppdrag att utforma.
Jag vill gärna avsluta med en mer politisk kommentar.
Jag anser att vi - de som har stött och stöder Lissabonfördraget, parlamentet och kommissionen - inte ska be om ursäkt för detta på något sätt, eftersom konkurrensen utifrån är starkare än någonsin, den kommer att vara hårdare än någonsin.
Vi behöver ett EU som fungerar bättre för våra medborgare, som bemöter de verkliga utmaningar som vi står inför.
Dessa utmaningar kommer att kvarstå: problemen med energisäkerheten, klimatförändringen, problemen med internationell terrorism, ökad konkurrens från utvecklingsekonomier och problemen med migration.
Dessa utmaningar är här, och vi måste hantera dem på ett effektivare sätt.
Därför får vi inte skylla på EU.
Vi måste vara ärliga när det gäller detta.
Det är sant att resultatet av de folkomröstningar som vi håller om EU mycket ofta har blivit ett nej till EU.
Men vi måste vara fullständigt ärliga.
Skulle resultatet alltid bli ja om vi skulle hålla folkomröstningar om de flesta nationella politikområden och de flesta av våra alternativ?
Därför får vi inte skylla på EU eller EU-institutionerna.
Sanningen är att det i dag är mycket tufft att fatta beslut på EU-nivå, nationell nivå eller regional nivå.
Vi måste följaktligen agera klokt, försiktigt och seriöst i detta avseende.
Vi får inte alltid skylla på EU.
Tvärtom måste vi arbeta för att förbättra EU, vara ödmjuka när det gäller bakslagen, förstå vad som inte fungerar bra, göra förbättringar och inte ge upp våra åtaganden.
Jag anser att det bästa sättet att göra detta är att undvika pessimism och inte gå tillbaka till en situation av ”krisfilosofi”, en kris för krisens egen skull.
Pessimism kommer inte att lösa problemet.
Det är sant att vi har ett allvarligt problem, men vi måste lösa det och inte falla tillbaka i depression.
Det bästa sättet att visa att vi är engagerade i vårt projekt - och jag välkomnar även det franska ordförandeskapets avsikter i detta avseende - är att arbeta konkret med de viktigaste områdena där EU kan skapa resultat och hjälpa våra medlemsstater att lösa de problem som verkligen bekymrar våra medborgare mest.
Jag hoppas att vi inte kommer att bli missmodiga av detta och att vi kommer att hålla oss till vår linje.
Vi behöver naturligtvis sjömän och navigatörer vid fint väder, men även för stormiga tider.
Jag anser att vi bör hålla kursen och fortsätta med vårt projekt, så att EU blir nödvändigare än någonsin.
(Applåder)
för PPE-DE-gruppen. - (FR) Fru talman, herr rådsordförande, herr kommissionsordförande, mina damer och herrar! Majoriteten av det irländska folket som gick till val uttryckte sitt motstånd mot Lissabonfördraget.
Min grupp respekterar det beslutet, precis som vi även respekterar de 18 medlemsstater som hittills har uttryckt sitt stöd för fördraget och har ratificerat det.
EU grundas på yttrandefrihet och demokrati.
Vi är demokrater, och därför vill vi att alla medlemsstater ska uttrycka sin åsikt om ratificeringen av fördraget.
Det är först i slutet på den processen som Europeiska rådet kommer att kunna besluta vilken väg vi ska välja, med andra ord - utan att förta vikten av Irlands beslut - får inga medlemsstater hindra de andra från att fritt uttrycka sin åsikt.
Vi hoppas att Europeiska rådet den här veckan kommer att göra en lugn, ansvarsfull och konstruktiv analys av den situation som har uppstått till följd av detta folkomröstningsresultat.
PPE-ledamöterna i min grupp hoppas att Europeiska rådet kommer att uppmana de medlemsstater som inte redan har gjort så att fortsätta med sina ratificeringsförfaranden, vilket inte är mer än rätt.
Mina damer och herrar, det irländska folket har talat.
Det har uttryckt sin oro över syftet med den europeiska integrationen, hur EU styrs, om framtiden för den gemensamma jordbrukspolitiken, om WTO-förhandlingarna, om skattepolitiken.
Det irländska folkomröstningsresultatet avspeglar även det faktum att många inte förstår EU:s komplexitet, och att EU:s relevans inte alltid är så uppenbar för dem.
Det är ett uttryck för den fråga som många medborgare ställer sig om själva syftet med den europeiska integrationen.
Min och min generations motivation - med andra ord att säkra fred på vår kontinent - förstås inte längre av de yngre generationerna.
Det irländska nejet är en vädjan till EU att definiera sina mål bättre och förklara skälen till att fortsätta med integrationen.
Europaparlamentet, som ofta antar svårlästa texter, måste spela sin roll fullt ut i det här arbetet.
Menar irländarna med sin nejröst att våra länder klarar av att lösa klimat- eller energifrågorna, den nya livsmedelsordningen, den personliga säkerheten, invandringen eller utrikespolitiken på egen hand och att de kan agera på likställda villkor med Förenta staterna, Kina, Indien eller Brasilien?
Jag tror inte det.
Menade irländarna med sin nejröst att solidariteten med de fattigaste länderna, den solidaritet som de avsevärt och med all rätt har dragit nytta av under de senaste årtiondena, inte är relevant och att regeln från och med nu är att ”rädda sig den som kan”?
Jag tror inte det.
Ville irländarna slutligen genom att rösta nej lägga den europeiska integrationen åt sidan och uttryckte de en negativ åsikt om anslutningen av ett land som Kroatien?
Jag tror inte det.
PPE-ledamöterna i min grupp är fast övertygade om att Lissabonfördraget, som var föremål för långa förhandlingar och undertecknades av samtliga 27 medlemsstater, är ett stort steg framåt jämfört med Nicefördraget.
Det gör att EU kan fungera bättre och ger oss de redskap vi behöver för att hävda oss i högre grad på världsarenan.
Jag har bara en önskan och det är att EU slutar med sin själviakttagelse så snabbt som det bara är möjligt.
Det är dags att våra länder - om jag får uttrycka det så - slutar med navelskåderiet och börjar arbeta tillsammans för att övervinna de verkliga problemen och utmaningarna.
Dessa utmaningar måste sporra oss till aktion och de ger även upphov till allvarlig oro och ibland vrede, vilket vi kommer att se igen i Bryssel på torsdag, bland dem som är försvagade och belastas av den rådande situationen.
Herr rådsordförande, min uppmaning till er är att ni tar hänsyn till de verkliga problemen i morgon i Europeiska rådet, värnar om alla EU-medborgares välfärd, och utan omsvep tar itu med alla de prisökningar som oroar våra medborgare.
PPE-ledamöterna i min grupp manar till lugn och förnuft i denna upphetsade debatt.
Vi måste lyssna till irländarna, vi måste lära oss av deras röst och vi måste behandla folket i de andra EU-länderna med samma respekt.
(Applåder)
för PSE-gruppen. - (DE) Fru talman! Vi har varit konstant upptagna med att ratificera ett eller annat fördrag i åtta år vid det här laget.
Vi har ratificerat oss själva till döds.
Under dessa åtta år har EU genomgått en period av själviakttagelse och har inriktat sig på sina egna institutionella reformer, om än utan särskilt lyckat resultat.
Detta är samma EU som kräver att anslutningskandidaterna ska genomföra förändringar, och ändå är det uppenbarligen oförmöget att klara av detta själv.
Hur stor trovärdighet ger det oss?
Herr kommissionsordförande, ni påpekade helt korrekt att detta inte är EU-institutionernas fel och att vi inte alltid ska göra dem till syndabockar.
Ni har helt rätt i det, men vem är det exakt som gör dem till syndabockar?
Det finns väldigt många människor i Europas huvudstäder som kommer att samlas för att diskutera fördraget på torsdag, och varje gång de reser hem igen och om rådets möte i Bryssel har varit framgångsrikt, säger de: ”Det var vi, stats- och regeringscheferna, som klarade av alltihop”, och om mötet inte blev lyckat säger de: ”Det var deras fel, allt är Bryssels fel!”
Ni upprepa det ni har sagt här för rådet.
För övrigt genomförs den här debatten med er offentligt, men stats- och regeringscheferna kommer återigen att mötas bakom stängda dörrar på torsdag.
Det måste också upphöra.
Det är medlemsstaterna som bär ansvaret!
(Applåder)
Vi har en nedåtgående spiral, en negativ spiral, och det är mycket farligt.
Det är den europeiska integrationen som står på spel.
Irländarna har hållit sin folkomröstning och vi måste respektera resultatet, men det fanns en faktor som oroade mig djupt.
Med undantag för Sinn Féin - och jag kommer inte att slösa några ord på dem här - manade alla de irländska partierna, PPE-DE, liberalerna och vårt eget parti - till ett ja och det irländska folket röstade nej.
Detta är en varningssignal och alla, även vi här i parlamentet, berörs av det faktum att det finns en förtroendekris, en kris av misstroende gentemot de nationella och naturligtvis även de överstatliga institutionerna.
Jag klarar mig utan era applåder.
Att det är UKIP:s ideologi som företräder den irländska suveräniteten är diskutabelt enligt min mening.
Irländarna klarar sig utan ert skydd.
Jag vill klargöra detta mycket tydligt: vi måste stå enade i vårt gensvar på förtroendekrisen och vi måste ta den på allvar.
Herr kommissionsordförande, jag väntat på att ni äntligen skulle säga ett par ord om kommissionsledamot Charlie McCreevy i dag.
(Applåder)
Det är han som är ansvarig för inremarknadspolitiken i EU: samma inre marknad som alltfler medborgare helt förståeligt ser som ett hot, inte som en möjlighet, till följd av de sociala skillnaderna.
Denna man, som har ansvar för den inre marknaden i er kommission, reser till Irland och förklarar att han inte har läst Lissabonfördraget och att han inte förväntar sig att väljarna ska göra det heller.
Hur kan detta rimligtvis öka allmänhetens förtroende?
(Applåder)
Låt mig säga detta: den bästa socialpolitiska åtgärden för EU som ni kan föreslå den 3 juli är att ta ifrån Charlie McCreevy detta ansvarsområde, för han har bevisat att han inte klarar av uppgiften.
Jag kan inte acceptera en kommissionsledamot med ansvar för den inre marknaden som står för en så skev politisk inställning.
Det Charlie McCreevy vill göra är att avreglera den inre marknaden till bristningsgränsen, oavsett följderna, utan kompletterande sociala åtgärder på EU-nivå eller i medlemsstaterna.
Det är den kris som EU-medborgarna känner av!
Ni måste agera när det gäller denna särskilda kommissionsledamot!
(Applåder)
Jag skulle även gärna ha velat höra er säga något om finansmarknaderna.
Ni har inte sagt ett enda ord om oron på finansmarknaderna ännu.
Jag vill även rikta en kommentar till Joseph Daul: det finns 21 regeringschefer inom EU som tillhör er politiska familj eller liberalerna, och ett lika stort antal ledamöter av kommissionen.
Jag medger gärna att PPE-DE-gruppen i parlamentet är öppen för nya idéer när det gäller vissa socialpolitiska åtgärder.
Jag uppmanar er att äntligen tala med era regeringschefer och med era kolleger i rådet!
EU behöver ett gemensamt agerande på det sociala området.
Ni har majoritet i EU, i rådet, i kommissionen och även här i parlamentet.
Visa för en gångs skull det sociala ansvar som ni just har efterlyst.
Jag uppmanar er att göra detta, till exempel när det gäller min kollega Paul Nyrup Rasmussens betänkande om kontroll av de internationella finansmarknaderna.
Jag uppmanar er att följa upp era storslagna uttalanden om ansvar med konkreta åtgärder.
Ett varmt välkommen till er, herr Daul!
(Applåder)
Vi kommer att finna en väg ut ur denna återvändsgränd, det är jag säker på.
På ett sätt eller annat kommer vi helt klart att få ombord irländarna igen.
Det kommer dock inte att hjälpa oss!
Vi måste erkänna att det fanns en tid då den proeuropeiska rörelsen hade en själ och ett hjärta.
Som Joseph Daul påpekade var detta efter kriget, när Europas fredsskapande kult svetsade samman människorna.
Nu är det den antieuropeiska rörelsen som har hjärta och själ, och ni ser att de är extremt aktiva.
De rusade runt på Irland, sprang i trappor, ringde på dörrar, värvade röster och delade ut sitt kampanjmaterial.
De fanns överallt.
Var höll EU-vännerna hus?
Var finns den rörelse som kampanjade för den europeiska integrationen?
Var finns den passion som vi en gång kände?
Den har flyttat över till den andra sidan, de som talar illa om EU, till högerkanten av det politiska spektrat.
Den finns hos dem som talar illa om EU, och de som helt enkelt gör det för att de är rädda.
I Europa har denna blandning av socialt förfall och rädsla emellertid alltid öppnat dörren för fascism.
Jag vädjar därför till alla konstruktiva demokratiska krafter i EU att ta denna rörelse på allvar!
Låt oss äntligen förena oss igen med en enda målsättning för ögonen: att påminna oss själva om att det aldrig har funnits ett mer framgångsrikt projekt för att trygga freden i Europa och i världen än den transnationella, interkulturella, interreligiösa rörelse som bygger på en balans av sociala intressen och kallas för Europeiska unionen.
Det är ett projekt som är värt att kämpa för, eftersom vi inte får låta dessa människor få övertaget.
(Applåder)
för ALDE-gruppen. - (EN) Fru talman! När den irländske premiärministern ger sig i väg till Bryssel i morgon kan han mycket väl fundera på den irländska popgruppen U2:s hit: ” Where did it all go wrong?”
De andra stats- och regeringscheferna bör även fundera på vad det betyder att vi, på tröskeln till det nya franska ordförandeskapet, har gått hela varvet runt sedan sist: från Nice till Nice.
Det finns tydliga bevis för att en majoritet i alla medlemsstater stöder EU.
Det finns få bevis för att en majoritet i någon av medlemsstaterna är för ett fortsatt uppbyggande av EU.
Vi kan inte säga med säkerhet att något fördrag skulle få majoritet i något av länderna.
Förtroendet för institutionerna ebbar ut.
För att muntra upp stämningen i Berlin kunde man vissla på en annan U2-hit, ”With or without you”, eller tvinga Irland att rösta igen i Paris.
Som Brecht påpekade kan man inte upplösa folket.
Trots att mindre än en miljon personer röstade mot i en opinion som var full av lögner, är folket inte övertygat.
Varför?
För det första för att vi har gjort för lite för att övertyga dem om de förändringar som vi kämpar för.
Kommissionen har en ”plan D” för dialog, men våra medlemsstaters regeringar har ingen motsvarighet till detta.
Här har parlamentet och kommissionen verkligen en roll att spela för att förklara vad EU betyder - men det gäller även alla de nationella regeringarna, varje dag, inte bara när det är dags att ratificera det senaste fördraget.
Och här har vi också en uppgift, inte bara för de politiska partierna på EU-nivå, utan för de politiska partierna i alla medlemsstater.
För det andra har EU visserligen skapat stort välstånd, men nu är det samlat på ett mindre öppet sätt och sprids mindre rättvist.
Våra ledare i politiken och näringslivet har enorma etiska frågor att ge sig i kast med.
Och herr Schulz, jag är ledsen att ni endast har fem stats- och regeringschefer nuförtiden, men dessa frågor väger inte mindre i de länder som styrs av socialisterna än de är i andra!
(Applåder)
För det tredje är fri rörlighet för varor och kapital - och även för tjänster - mycket viktigt, men vår union är inte känd för att ge friheter till folket.
Gränsöverskridande komplikationer i civilrättsliga frågor - vårdnadstvister vid skilsmässor, problem med egendomar utomlands - fyller Europaparlamentarikernas inkorgar.
En brist på garantier i gränsöverskridande brottmål och en nonchalant inställning till dataskydd ökar olustkänslan.
Det som EU lovar i teorin misslyckas man alltför ofta att genomföra i praktiken.
Det är mot denna bakgrund som vi bör avväga vårt svar till Irland.
Här i parlamentet vill vi ha ett nytt fördrag.
Vi vet att det kommer att bidra till att ställa dessa saker till rätta.
Men bortom denna skog av metall och glas är förståelsen alltför liten.
Min grupps rekommendationer till rådet är följande.
Fortsätt med de verkligt viktiga frågorna för EU: öka handeln, bekämpa klimatförändringen och prishöjningarna på livsmedel och bränsle.
Låt dem som vill fortsätta att ratificera fördraget.
Om nödvändigt får vi klara oss med Nicefördraget.
Använd övergångsklausulen för att öka EU:s problemlösningspotential.
Glöm heltidsordföranden till dess att ni har bestämt er för vad sexmånaderspraktiken ska leda till.
Inled en omfattande kampanj för att påminna folket om varför EU finns, informera dem om hur EU fungerar och förklara varför, precis som den legendariska Guiness-reklamen, ”EU är bra för dig”.
EU betyder alltför mycket för alltför många för att denna kris ska kunna ändra den inslagna kursen.
(Applåder)
för Verts/ALE-gruppen. - (IT) Fru talman, mina damer och herrar! Vi har alltid sagt att EU behöver en kortfattad konstitution med en stadga med bindande rättigheter, demokratiska och öppna beslutsförfaranden, begränsade men verkliga befogenheter och de nödvändiga ekonomiska resurserna.
En sådan konstitution borde utarbetas av parlamentet eller en konstituerande församling, upprätthållas strikt och med övertygelse, utan hyckleri, och ratificeras genom den parlamentariska metoden eller i en EU-folkomröstning.
Jag har stor respekt för det irländska folkets vilja, men ingen kan någonsin övertyga mig om att en folkomröstning där halva väljarkåren stannade hemma är mer demokratisk än en parlamentarisk ratificering.
Om majoriteten av stater och folk röstar ja går man vidare och de som röstar nej kan gärna fortsätta att stå utanför och förhandla fram ett system med nya, lösare förbindelser, som det uttrycks i Spinelli-fördraget från 1984.
Vad har hänt de senaste åren?
Medlemsstaterna och kommissionen har valt en väg med komplicerade och motstridiga fördrag som är svåra att sälja och som i slutskedena förhandlades fram i hemlighet i all hast, och gjordes ännu mer oläsliga med sina undantag och protokoll.
Under tiden beslutade de att fördraget måste ratificeras enhälligt, precis som trädgårdsmästarens hund som varken äter kålen själv eller låter någon annan göra det.
Och som om detta inte var tillräckligt fortsätter EU att anta missledd och svag politik, som Jacksonbetänkandet om direktivet i går och Weberbetänkandet i dag, som inte kan erbjuda oss några positiva framtidsutsikter eller förhoppningar.
Detta är en union där mindre och mindre hänsyn tas till allt från arbetstagarnas rättigheter till miljöskyddet och migranters rättigheter, där lobbygrupper från näringslivet är mer värda än medborgarna, där det europeiska intresset har gått förlorat och överröstats av ramaskrin från en regering eller en annan, där valfriheten och de individuella rättigheterna eller nya européers ankomst betraktas som en outhärdlig attack mot folkens identitet, folk som Italiens och Irlands, som har migranter utspridda överallt i världen.
Det är möjligt, och kanske till och med önskvärt, att de länder som inte har ratificerat ännu gör det.
Den irländska regeringen kanske kommer med ett genialiskt förslag.
Men en diplomatisk lösning är inte tillräckligt!
En diplomatisk lösning räcker helt enkelt inte.
Nu mer än någonsin måste vi tydligt och högt förklara att regeringarnas Europa - grumliga och otydliga - är det EU som har misslyckats.
Det EU som förkastade konstitutionen och fortsäter att föra en missriktad, konservativ, trångsynt, nationalistisk och egoistisk politik, som tar andan från Europeiska konventionen från 2003 och i stället får en överenskommelse om en positiv, men minimalistisk och själlös text.
Inget av detta gör emellertid ett mer demokratiskt, aktivt och enat EU mindre viktigt.
Det som behövs i dag är ett initiativ som härrör från vår politiska styrka och från de medlemsstater som är övertygade om att vi måste skapa ett effektivare, mer demokratiskt och mer sammanhållet EU, med tanke på att det nu varken är nödvändigt eller möjligt att fortsätta med Nicefördraget längre.
I ett sådant initiativ kommer det inte att finnas något utrymme för dem som är ovilliga att gå framåt.
för UEN-gruppen. - (EN) Fru talman! Jag vill tacka rådets ordförande, kommissionens ordförande och mina kolleger för deras inlägg hittills i debatten.
Det som har skett var uppenbarligen oväntat.
Nejrösten på Irland är en helomvändning när det gäller åsikten om EU-projektet från en grupp väljare inom EU.
På grund av meningsskiljaktigheterna bland dem som motsatte sig fördraget i folkomröstningen på Irland, på grund av de olika ståndpunkterna - som var både politiskt och ideologiskt motsatta vid många tillfällen - är det svårt att dra några exakta slutsatser om skälen till att folket röstade nej.
Det vi har begärt är att få tid på oss för att begrunda och analysera detta resultat, finna lösningar för att gå vidare och se vad som kan göras.
Detta var nämligen inte - vilket även personer från nejsidan hävdar - en röst mot EU, trots att en del på nejsidan har röstat nej i varenda folkomröstning som har hållits om EU-frågor sedan Irland anslöt sig 1972.
Men de hävdar att detta inte är en röst mot Europa.
De hävdar vidare att det inte är ett sätt att förringa det som EU gör.
Men deras viktigaste slagord under kampanjen var att ”rösta nej till ett starkare Europa”.
Nu kanske de på nejsidan kan tala om för oss vilket slags starkare EU de vill se och vilka lösningar de har att komma med om hur vi ska gå vidare för att hantera de globala utmaningar och svårigheter som vi står inför.
Här i Bryssel har vi i dag jordbrukare och åkare som protesterar mot de höga bränslepriserna.
För ett år sedan kostade ett oljefat 48 US-dollar, i dag kostar det 140 US-dollar.
Den här tiden för ett år sedan hade även de fattiga på Haiti råd att betala livsmedelspriserna, i dag förekommer upplopp på Haitis gator på grund av livsmedelsbristen och de svårigheter den ger upphov till.
Det är dessa utmaningar som vi måste bemöta på EU-nivå, och det är dessa svårigheter som vi måste ta itu med.
Vi får inte glömma att världen inte kommer att gå under.
Vi har varit här förut: både fransmännen och nederländarna röstade nej till det föregående fördraget och man fann en mekanism för att organisera och gå vidare med det europeiska projektet.
Det är inte rätt tillfälle för att skylla på eller peka finger åt varandra.
Tvärtemot vad många som protesterar i parlamentet kan tro är det nu dags att vi visar respekt för varandra, inte bara respekt för de irländska väljarna som uttryckte sin demokratiska åsikt om detta fördrag, utan även respekt för de andra länderna och deras enskilda rättighet att bestämma hur de fungerar och hur de ratificerar fördrag.
Det är inte upp till oss att tala om för någon annan hur man bör gå vidare och hur man inte bör göra det.
Till dem som bär t-tröjor här i kammaren vill jag säga att de inte bara visar en respektlöshet mot parlamentet och parlamentets ledamöter, utan att de inte på något sätt står för eller företräder det irländska folket eller den irländska nationen.
(Applåder)
Jag vill klargöra att det var just dessa flåspatrioter här till vänster om mig, exakt de som hävdar att de försvarar det irländska folkets rättigheter, som kunde ses i irländsk tv när de firade Irlands nej på en pub i Bryssel.
Det dracks naturligtvis, men vilken respekt har de för det irländska folket och den irländska flaggan om de använder den som en bordduk att ställa sina drinkar på?
Det är vad den gruppen står för, det är den slags respektlöshet som de visar gentemot folket.
(Applåder)
Ge oss utrymme att gå vidare.
Det europeiska projektet är värt att bevara.
Det handlar inte bara om fred eller välstånd, det handlar om solidaritet.
För många år sedan skrev den irländske poeten Sean O'Casey följande i Juno and the Paycock: ”Jag såg ofta upp mot himlen och ställde mig frågan - vad är månen, vad är stjärnorna?”
I dag kanske vi själva bör ställa en fråga för vår generation: Vad betyder EU egentligen och hur vill vi att EU ska vidareutvecklas?
(Applåder)
för GUE/NGL-gruppen. - (FR) Fru talman, herr kommissionsordförande, herr rådsordförande, mina damer och herrar! Europeiska rådet skulle göra klokt i att avhålla sig från att visa någon slags arrogans gentemot Irlands folk, som endast utövade en demokratisk rättighet som erkänns i deras konstitution.
I stället för att begära att ratificeringsprocessen ska fortsätta i ett försök att frysa ut detta nya svarta får, skulle det vara bättre att ta itu med en tydlig analys av situationen.
Det var särskilt många ur arbetarklassen på Irland som röstade nej, och jag vill påminna er om att valdeltagandet var mycket högre än tidigare, vilket enligt min grupp visar på att legitimitetskrisen när det gäller den befintliga EU-modellen växer allt djupare.
Denna kris var redan grundorsaken till fransmännens och nederländarnas nejröster, den uttrycks annorlunda på andra håll, men den är alltid en underliggande faktor.
Kom ihåg de omfattande protesterna mot Bolkestein-direktivet, den debatt som uppstod efter Laval- och Vikingaffärerna, särskilt i de skandinaviska länderna, eller i Tyskland efter Rüffert-domen.
I detta avseende vill jag säga min vän Martin Schulz att jag fullständigt håller med om vad han sa om Charlie McCreevy.
Problemet är att dessa beslut - de som jag just har nämnt - inte fattades av Charlie McCreevy utan av EG-domstolen på grundval av särskilda artiklar (artiklarna 43 och 49 i de gällande fördragen som infogas i Lissabonfördraget).
Tänk även på de politiska följderna av den omfattande strejken i Dacia i Rumänien, mot ”lågkostnads-Europa”.
Se på vreden bland jordbrukare och småskaliga fiskare som har stora ekonomiska svårigheter.
Det som ligger till grund för alla dessa situationer är först och främst den nuvarande europeiska ekonomiska och sociala modellen. I stället för att skapa säkerhet leder den till större osäkerhet.
Det är det största problemet.
En annan faktor är EU:s funktionssätt.
Besluten fattas långt ifrån folket och utan deras medverkan.
Vi nöjer oss med att förklara för dem i stället för att rådfråga dem.
Det avsiktliga beslutet att presentera Lissabonfördraget i en form som är fullständigt oläslig för en lekman är i detta avseende en effektfull illustration av vad jag skulle kalla ”elfenbenstornssyndromet”.
Detta har förödande effekter på våra medborgare, särskilt de mindre befolkade nationerna, som tycker att de bollas runt för att tillgodose mäktigare nationers intressen.
Slutligen uppstår alltfler frågetecken i många länder, inklusive Irland, om den roll som EU spelar i världen, där EU förväntas garantera att politikens makt betonas mycket starkare än politiken som maktmedel.
Att undvika dessa diskussioner leder till att krisen i Europa förvärras, att föra diskussionen i ett fullständigt öppet klimat skulle vara det första steget på vägen mot att finna en lösning.
för IND/DEM-gruppen. - (EN) Fru talman! Ingen annan har sagt det, men det kommer jag att göra: Bra gjort Irland!
(Applåder från vissa håll)
Och trots detta, redan innan det officiella resultatet var känt, höll José Manuel Barroso, som såg lömskare och oärligare ut än någon annan jag någonsin har sett, en presskonferens i Bryssel och sa - tvärtemot klubbens regler - att fördraget inte är dött och att vi fortsätter.
Det var uppriktigt sagt en osmaklig uppvisning, det var en förolämpning mot demokratin.
Det står fullständigt klart att ratificeringarna bör upphöra nu och att genomförandet av fördraget bör stoppas.
Efter de franska och nederländska resultaten trodde jag att ni förnekade verkligheten, men nu inser jag att det som ligger bakom detta är ett nytt fenomen, det är ”EU-nationalism”, och att det är det farligaste politiska fenomen som har drabbat Europa sedan 1945.
Ni struntar i väljarna, ni förgör demokratin, och ni har visat att ni inte skyr några medel.
Men ställ er då frågan varför politikerna, varför denna klass, nu är impopulära.
Ja, herr Barroso, senare i dag kommer parlamentet att rösta om en ny kommissionsledamot för rättsliga frågor, och det är sannolikt att en tidigare dömd bedragare kommer att bli kommissionsledamot med ansvar för rättsliga frågor i EU från och med i dag.
I själva verket behöver ni inte UKIP-partiet.
Ni förstör själva EU i väljarnas ögon.
Bra gjort, alla!
(Applåder från vissa håll)
(EN) Fru talman! Jag påminner parlamentet om att rättstaten är viktigare än själva lagarna.
(Högljudda protester)
Lissabon krävde enhällighet.
Att bortse från detta innebär att bortse från rättstatsprincipen i sig.
Irländarna utgör inte bara 10 procent av EU, de utgör 100 procent av dem som har rösträtt och de vet alla, vi vet alla, att andra skulle ha röstat nej om de fått chansen.
(Fortsatta högljudda protester)
Lissabon var obegripligt och irländarna visste varför.
Andra skulle ha röstat nej om de fått chansen.
Att nu föreslå att processen ska fortsätta, tänka ut ännu klyftigare sätt för att återuppliva Lissabon i öppet trots mot allmänhetens vilja, är en arrogant handling av hisnande proportioner och vi har sett allt förut.
Efter det att det tidigare fördraget förkastats stod den österrikiske utrikesministern här och skröt om 36 projekt och institutioner som fortfarande fortsatte. De har fortfarande ingen legitimitet efter misslyckandet med att nå enhällighet om Lissabonfördraget.
Jag har ett budskap till er från Edmund Burke: ”Det är folket som är herrarna och inte ni, och ni ignorerar detta på egen risk.”
(Applåder)
kommissionens ordförande. - (FR) Herr talman! Jag vill lyfta fram det anmärkningsvärda samförstånd som råder i parlamentet om vad vi bör göra härnäst.
Vi anser, med ett fåtal undantag som bara ger färg åt debatten, att alla medlemsstater skulle göra klokt i att slutföra sina ratificeringsprocesser.
Det är också den åsikt som har uttryckts av den irländska regeringen och av ledamöterna, särskilt Brian Crowley, som är irländare och som har förklarat att alla länder har samma rätt att uttrycka sin åsikt.
Om vi kan slutföra denna process kommer vi att kunna diskutera frågan på ett konstruktivt sätt med våra irländska vänner i en anda av solidaritet, för det kan inte råda enighet utan solidaritet.
Jag anser att det är detta samförstånd som håller på att befästas, och jag hoppas att det kommer att befästas av debatten i Europeiska rådet i morgon och senare.
I alla händelser är det den ståndpunkt som kommissionen kommer att lägga fram för Europeiska rådet.
Samtidigt är det, som många av er har påpekat, bland annat Graham Watson och andra, viktigt att vi inte förlamas genom att bara inrikta oss på den institutionella frågan. Det bästa sättet att befästa EU:s demokratiska legitimitet är att skapa resultat och visa att vi verkligen arbetar för våra medborgares bästa.
Världen väntar inte på att EU ska fatta sina institutionella beslut. Det finns brådskande frågor som klimatförändringen, energisäkerheten och migrationen som kräver agerande från EU:s sida, även inom den befintliga institutionella ramen.
Ett annat påpekande, som jag riktar till min gode vän Martin Schulz, är att vi måste undvika att leta efter enkla syndabockar.
Jag tyckte självklart inte att kommentarerna från min kommissionskollega Charlie McCreevy var särskilt välvalda.
Jag skulle emellertid även kunna nämna vissa kommentarer från nationella politiker som inte har varit nyttiga för processen, och även från parlamentets ledamöter, som inte alltid säger det vi vill höra.
Låt oss vara realistiska!
I den valkrets där kommissionsledamot McCreevy kampanjade vann jarösten, och att attackera den irländske kommissionsledamoten nu anser jag inte vara det bästa sättet att garantera en givande dialog med våra irländska vänner.
Vi måste koncentrera oss på de positiva aspekterna utan att försöka hitta enkla syndabockar, det skulle inte vara rättvist.
Om vi agerar i en anda av samarbete med våra institutioner, om vi koncentrerar oss på de resultat som medborgarna förväntar sig av oss, om vi skapar den bästa möjliga atmosfären för denna dialog, anser jag att det kommer att vara möjligt att lösa det här problemet.
Det är ett allvarligt problem, men det kan lösas.
Vi kommer inte att lösa det med ömsesidiga beskyllningar eller med pessimism, ”krisfilosofi” eller tal om en tillbakagång.
Vi kommer att lösa det genom våra ansträngningar, genom våra resultat, för att förstärka vår demokratiska legitimitet och genom att erkänna att vi alla måste agera, i EU-institutionerna och i de nationella regeringarna, och att vi har ett gemensamt ansvar för att hålla våra ideal, vårt europeiska ideal, vid liv.
(Applåder)
(EN) Herr talman! EU som vi känner till det grundas på fyra friheter: fri rörlighet för personer, varor, kapital och tjänster.
Den första av dessa friheter handlar om människor. När Jean Monnet delade med sig av sin vision av Europa för alla dessa år sedan sa han - och jag hoppas mina kolleger har överseende med min dåliga franska - ”Nous ne coalisons pas des États, nous unissons des hommes”.
Det är meningen att EU ska handla om människor, inte om politiker, vilket innebär att EU inte bara måste drivas av människorna, de behöver också se att EU drivs av människor.
I torsdags hörde vi folket tala och deras dom var tydlig, svaret var ett tydligt nej.
Jag vill påminna om bakgrunden till det första konstitutionsfördraget.
Man erkände att EU höll på att bli mer otillgängligt för folket och att man måste göra något åt det.
Den uttalade lösningen var att utarbeta ett fördrag för att göra EU enklare, öppnare, närmare folket.
Men när politikerna var färdiga hade de utarbetat ett fördrag som var mer komplicerat, mer oklart och till och med ännu längre från folket.
Folket anser för övrigt detsamma om detta senaste fördrag.
Vi får inte svara genom att fortsätta som om ingenting hade hänt.
Om folket känner att EU blir mer avlägset och politikerna fortsätter som om ingenting hänt förvärrar det bara problemet.
Vårt problem får inte vara att diskutera hur snabbt EU bör gå fram, utan att diskutera vilken riktning det ska ta.
Lyssna till folket och de kommer att tala om det för er.
Om ratificeringsprocessen fortsätter kommer detta att visa att EU-ledarna inte har lärt sig någonting, att politikerna fortfarande tror att de vet bäst och att det är folket som har fel.
Folket har per definition alltid rätt.
Det kallas för demokrati.
Vi vill ha ett EU som är inriktat på människor och som skapar den demokratin.
Därför får vi inte bortse från det irländska röstresultatet, vi bör bygga vidare på det.
Ratificeringsprocessen bör upphöra och vi måste börja lyssna till folket.
(Applåder)
Avslutningsvis sa Martin Schulz i sitt mycket kraftfulla och eleganta inlägg att det råder en förtroendekris.
Jag håller med honom.
Det är folket som har förlorat förtroendet för politikerna.
Nu har vi ett tillfälle att erkänna detta, att visa att vi har lyssnat, och att återvinna och återuppbygga deras förtroende.
Det räcker inte att vi alla blir storslagna talare, vi måste visa att vi är goda lyssnare också.
(Applåder)
(EN) Herr talman, nej, nej, nej!
Det som den ärade ledamoten just har talat om är inte demokrati.
Demokrati är att säga ”vi respekterar irländarna, precis som vi respekterar alla andra medlemsstaters beslut”.
Därför stöder jag kommissionsordförandens uttalanden.
Det råder samförstånd om processen här i parlamentet, om att vi ska respektera irländarna, men även respektera alla de andra medlemsstaterna.
Låt oss fortsätta processen, det är vad vi måste fortsätta med i dag.
För det andra: inga fler pauser tack!
Inga fler perioder av ”eftertanke”.
Inget mer svammel.
Vi måste inrikta oss på de verkliga problemen.
Det är vad vi måste göra.
Ordförande José Manuel Barroso måste naturligtvis försvara sina kommissionsledamöter, även Charlie McCreevy.
När vi kritiserar Charlie McCreevy är det inte en personlig fråga.
När ordföranden för min grupp nämner Charlie McCreevy rör det hans politik - och hans politik är även José Manuel Barrosos politik.
José Manuel Barroso har sagt många kloka saker i dag, men när han talade om befogenheter på konkurrensområdet hörde jag ingenting om spekulationerna på finansmarknaderna mot livsmedelspriserna.
Jag skulle ha velat höra något om det, och jag skulle ha velat höra det från Charlie McCreevy.
När ordförande Barroso talade om ekonomin hörde jag honom inte säga att vi saknar arbetsillfällen i Europa.
Jag skulle ha velat höra honom säga det, att vi förlorar arbetstillfällen till följd av finanskrisen.
Jag skulle vilja se att kommissionen kom med en ny plan för att blåsa nytt liv i ekonomin - inte en teoretisk plan utan en samordnad investeringsåtgärd.
För det tredje försöker Charlie McCreevy just nu säga att skälet till att vi har en finanskris är finansorganen och finansinstituten - Standard & Poors, FTSE och andra - och att vi ska reglera dem.
Men det är på sätt och vis som att skjuta budbäraren.
Jag anser verkligen att kommissionsledamoten bör säga i dag att, ja, jag håller med om att vi har en finanskris, och ja, jag instämmer i att vi måste genomföra en allmän reglering som är bättre än den vi har, så att vårt svar blir nya arbetstillfällen och ett bättre klimat, inte mer pengar och en ökad inriktning på hur man ska skapa vinster från ingenting, i stället för på produktion och arbetstillfällen.
Ge oss det intrycket i dag, och ni har ett verkligt budskap att förmedla till vanligt folk.
(EN) Herr talman! Som irländsk ledamot företräder jag de 54 procent som röstade nej och de 46 procent som röstade ja.
Verkliga demokrater ser inte bara till resultaten, utan strävar efter att företräda hela folket.
Jag företräder en suverän stat, men man kan inte upprätthålla suveränitet i sin egen medlemsstat - i mitt fall Irland - om man inte upprätthåller alla medlemsstaters suveränitet.
Om en annan medlemsstat bestämmer sig för att utöva sin suveränitet och ratificera Lissabonfördraget eller något annat, kan ingen verklig demokrat, inga av de demokrater som stolt viftar med flaggor i dag och påstår sig vara irländare, rimligen protestera mot detta.
Irland talar för Irland, Slovenien för Slovenien.
Det är verklig demokrati och suveränitet.
En kärnfråga i debatten om Lissabonfördraget på Irland var enhällighetsprincipen.
Vi behöver enhällighet för att kunna ratificera Lissabonfördraget.
Samtliga 27 medlemsstater måste vara överens - det är kärnan.
Detta är det första riktiga testet av enhällighetsprincipen enligt Lissabonfördraget.
Vi får inte underkännas i detta test och däri ligger utmaningen.
Som politiker är det vår uppgift att visa att vi är situationen vuxen och klarar av denna utmaning, att lyssna till våra medborgare, finna lösningar och fortsätta med arbetet att bygga upp ett bättre Europa.
En del på nejsidan på Irland talade om en bättre uppgörelse.
Låt oss vara optimistiska och söka en bättre uppgörelse för alla medborgare.
Vi behöver lite tid och utrymme på Irland för att fundera och agera för att finna lösningar.
Den goda viljan för Europa finns där på Irland.
Vem skulle kunna ha förutsagt 1945, när Europa låg i ruiner, att vi skulle fira 50 år av fred år 2008?
Låt det vara vår inspiration.
EU är ett pågående arbete, en process - visserligen svår, men alltid, alltid värd mödan.
Det är därför vi är här.
Europas medborgare vill ha en union som fungerar.
Det vill irländarna också.
Det är jag hundra procent säker på.
Vi får inte göra dem besvikna.
(DE) Herr talman, herr rådsordförande! Det budskap jag får från regeringarna är att detta är ett irländskt problem.
När jag talar med medborgarna får jag budskapet att detta är ett europeiskt problem, en konflikt med EU.
Regeringarna talar om för oss att det är en diplomatisk konflikt.
Medborgarna säger oss att det är en förolämpning mot deras suveränitet, de anser att de utestängs och är djupt sårade.
Regeringarna talar om för oss att denna nejröst är obegriplig.
När jag lyssnar till medborgarna förklarar de att det är fördraget och processen som är obegripliga.
Regeringarna säger oss att de måste ta itu med de verkliga frågorna på dagordningen.
Medborgarna förklarar att de har försökt uppmärksamma de verkligt viktiga frågorna i åratal, och jag vill påpeka för kommissionsordföranden att de inte menar den militära, polisiära och inre säkerheten.
De talar om socialt ansvar och ett europeiskt svar på globaliseringen.
De talar om mer demokrati och insyn.
Regeringarna planerar att fråga den irländska regeringen vad som orsakade nejsidans seger.
I stället bör regeringarna själva fråga sig följande: Vems fel är det egentligen?
Regeringarna struntade i skriften på väggen efter nejresultaten i Frankrike och Nederländerna.
Har regeringarna tagit itu med de verkliga frågorna?
Bemötte de verkligen de svikna förväntningarna vid översynen av fördraget?
Var inte fransmännen tydliga nog i sina krav på en ny social ordning, ökat socialt ansvar och rättvisa?
Var kraven på mer demokrati helt enkelt inte tillräckligt tydliga?
Så vad gjorde ni?
Ni stuvade om i fördraget och skapade ett oläsligt hopkok av fotnoter, korshänvisningar och undertexter, och ni undrar varför medborgarna förkastar det.
Det finns en stor risk i denna skymf mot suveräniteten.
Den är inte bara en förolämpning mot det irländska folket, det finns en verklig risk för att denna missnöjeskänsla kommer att sprida sig och att européerna i allmänhet kommer att säga: det irländska folket har röstat för oss!
Ansvaret för detta ligger hos er, regeringarna!
Det är verkligen dags ...
(Talmannen avbröt talaren.)
(PL) Herr talman! Det är en väldigt spänd debatt.
Jag vill emellertid mana till försiktighet, stor försiktighet i uttalandena efter den irländska folkomröstningen.
En antydan om att Irland borde skämmas eller till och med uteslutas ur unionen är långt skadligare för EU än själva resultatet av folkomröstningen.
Martin Schulz, som sin vana trogen var något upphetsad, kom tyvärr med en sådan antydan.
Vi måste komma ihåg att Bryssels förmyndaraktiga hållning orsakade irritation på Irland och var ett av skälen till att Irlands folk röstade mot fördraget.
Det är inte sant att EU kommer att bli lidande utan det nya fördraget.
EU kommer att bli lidande till följd av intressekonflikter och medlemsstaternas egoism.
Det har ingenting med Irland att göra.
EU:s utrikespolitik kommer till exempel att bli lidande på grund av Tyskland.
Tyskland vill upprätta goda förbindelser på egen hand med Ryssland på bekostnad av länderna i Centraleuropa.
Frankrike bör ges skulden för att det blundar för Rysslands nyimperialistiska politik i regionen samtidigt som man kommer med plattityder om hur EU, Polen inberäknat, ska kämpa sig fram.
Fördraget får inte utnyttjas som en rökridå för våra egna misslyckanden.
Det beslut som fattats av Irlands folk får inte utnyttjas för att dölja våra egna fel och brister.
(Applåder)
(GA) Herr talman! Det irländska folket har talat.
Det irländska folkets nej till Lissabonfördraget i torsdags var inte en röst mot EU.
Irlands plats är i EU.
Irland har vunnit sociala och ekonomiska fördelar - både nord och syd - till följd av sitt medlemskap, även om några svårigheter fortfarande kvarstår.
Frågan var följande: är Lissabonfördraget bra för Irlands folk, för resten av EU och för utvecklingsvärlden?
Lissabonfördraget lades fram för Irlands folk och har förkastats.
Lissabonfördraget är slut.
Det irländska folket vill, precis som folken i Frankrike och Nederländerna tidigare, ha en bättre uppgörelse.
Nu har vi en möjlighet att blåsa nytt liv i debatten om EU:s framtid.
Vi måste utnyttja denna möjlighet.
Det skulle inte vara godtagbart att EU-ledarna försökte hitta sätt för att undvika eller kringgå folkets demokratiskt uttryckta vilja.
Ratificeringsprocessen måste upphöra, precis som den gjorde efter förkastandet av EU-konstitutionen.
Men den här gången måste vi lyssna till det irländska folket, vi måste lyssna till folket.
Många av de farhågor som tidigare uttrycktes i Frankrike och Nederländerna kom upp även i den irländska folkomröstningen.
Vi måste lyssna till folkets farhågor och bemöta dem.
(EN) Under folkomröstningskampanjen på Irland kom en rad centrala frågor upp gång på gång: det demokratiska underskottet, Irlands förlorade makt i EU, neutralitet och icke-militarisering, arbetstagarnas rättigheter, samhällsservice och fördragets inverkan på utvecklingsvärlden.
Dessa frågor måste bemötas.
Det europeiska projektet genomgår nu ett demokratiskt test i och med gensvaret på omröstningsresultatet på Irland.
Lyssnar EU till folket, respekterar EU deras demokratiska vilja, eller stöter det bort sina medborgare genom att åsidosätta allt detta?
Enligt min åsikt måste demokratin vara förhärskande.
Vi måste lyssna till vad det irländska folket har sagt.
Vi måste glömma talet om att åsidosätta dem eller fortsätta utan dem, isolera dem eller skylla på dem.
Vi måste lyssna mycket noga och lugnt på vad det irländska folket har sagt och till de problem som de har uppmärksammat när det gäller neutraliteten och hela frågan om militariseringen av EU, när det gäller demokrati och Irlands och andra små EU-nationers röst, arbetstagarnas rättigheter, samhällsservice och det sociala Europa.
Vi måste lyssna till detta.
Vi måste nu ta tillfället i akt för att tala med den irländska regeringen, lyssna till det irländska folket och staka ut rätt kurs framåt och en text som alla kan vara nöjda med i framtiden.
(EN) Herr talman! Jag kände att det fanns två förhärskande stämningslägen under kampanjen.
Det första var en allmän känsla av att beslutsprocessen flyttades ännu längre från medborgarna till förmån för en avlägsen byråkrati.
Den andra känslan, som kanske var djupare, var att värderingarna har gått förlorade, eller rättare har förändrats.
Irland satte en ära i sina kristna värderingar, men började bli en materialistisk nation.
Det har talats i mycket nedvärderande ordalag om mitt land sedan i fredags.
Det är som om ni känner er förolämpade.
Det som faktiskt hände var att Irland bestämt sa ”nej tack” till Lissabonfördraget.
Om den reaktion på folkets demokratiska vilja som jag har sett under de senaste fem dagarna är indignation, är det något fel någonstans.
Missta er inte: Irland är EU-vänligt.
Vi anser, vilket ni uppenbarligen inte gör, att projektet har förlorat sin riktning.
EU har förlorat det man behöver mest - demokratin - ur sikte och man glömmer bort det som är viktigast - medborgarna.
Innan ni försöker kringgå vårt demokratiska beslut, ställ två frågor.
För det första: tror ni uppriktigt att Lissabonfördraget skulle överleva folkomröstningar i de andra 26 länderna?
Och för det andra: är det en demokratisk handling att hota ett land för att det är demokratiskt?
(Applåder)
- (NL) Herr talman! Ju längre detta fortsätter desto mer uppför sig de europeiska byråkraterna som ett släkte av politiska autister, fullständigt avstängda från verkligheten, från medborgarna, som de likväl fortfarande hävdar att de tjänar.
Nu säger de att lilla Irland inte har rätt att opponera sig mot ett EU-fördrag, som snart kan ratificeras av 26 av de 27 medlemsstaterna.
Vilken arrogans!
När allt kommer omkring är det bara Irland som har sagt nej eftersom det är det enda landet som har getts chansen att göra det.
Alla vet att Lissabonmonstret, som uppstod från den dödfödda EU-konstitutionen som ett Frankensteinmonster, skulle förkastas genom ett rungande nej av nästan alla de andra medlemstaterna om dessa väljare gavs chansen att rösta.
I demokratins namn buas ett demokratiskt valresultat ut och avfärdas.
Vi är på god väg mot en totalitär euronazistat.
(SL) Det irländska folkets beslut var demokratiskt och vi respekterar det, så det finns inget skäl att vädja till oss demokrater att visa respekt.
Det råder inget tvivel om detta, och ändå är det inte nog att bara respektera resultatet, vi måste även vara medvetna om följderna och måste analysera, ur irländsk och europeisk synvinkel, varför majoriteten i en av EU:s framgångsrikaste medlemsstater vände sig mot ett fördrag som stats- och regeringscheferna - även Irlands - undertecknade förra året i syfte att ta fram en effektiv gemensam strategi för att bemöta de nya och komplicerade utmaningarna, vare sig det handlar om miljö, energi, migration eller hälsa.
Jag håller med om att vi bör ta tid på oss för att begrunda detta, men den fortsatta ratificeringen får inte påverkas.
En fortsatt ratificering kräver ingen vidare eftertanke och processen måste fortsätta.
Frågan gäller inte bara Irland och hela det nuvarande EU, utan även Europas framtid, som ännu inte är helt enat.
I detta sammanhang gratulerar jag det slovenska ordförandeskapet till alla deras framgångar med att knyta länderna på västra Balkan närmare EU, särskilt stabilitets- och associeringsavtalen med Serbien och Bosnien och Hercegovina.
I detta sammanhang måste vi glädjas över alla framsteg som görs i en europeisk framtidsanda, och vi måste bekämpa alla möjliga konfliktkällor, vilket möjliggörs genom det europeiska perspektivet.
Jag uppmanar till outtröttliga insatser på detta område.
Jag hoppas att segern för de EU-vänliga krafterna i Makedonien kommer att bidra positivt till att rådet beslutar om att inleda förhandlingar med detta land, som redan är ett kandidatland och har suttit länge ute i väntrummet.
Jag hoppas även att den nya makedonska regeringen, som har getts ett starkt mandat, kommer att dra nytta av detta nya förtroende genom att föra en politik som stärker utvecklingen mot att inleda förhandlingar.
(DE) Herr talman!
Det jag vill se i Europeiska rådet i morgon är ärlig självkritik, eftersom man uppenbarligen har misslyckats med att kommunicera och informera allmänheten om detta nya EU-fördrag.
Det är häpnadsväckande att regeringarna förhandlar om ett fördrag och undertecknar det vid högtidliga ceremonier, och sedan reser tillbaka till sina huvudstäder och inte tänker mer på den saken.
Det är en stor orsak till den uppståndelse vi har upplevt i det förgångna och som vi nu möter med Irland.
(Applåder)
Nu är det dags att ta lärdom. Rådet måste äntligen gå ifrån sin blockeringstaktik och ta initiativ till en gemensam kommunikations- eller upplysningsstrategi tillsammans med kommissionen och parlamentet så att vi verkligen får med oss medborgarna på vår resa mot EU i stället för att lämna kvar dem vid vägkanten.
För närvarande uppför sig institutionerna som föräldrar som föder ett barn till världen och sedan slänger ut barnet i rännstenen och glömmer bort det.
Det är helt enkelt oacceptabelt.
Nu måste vi ta konsekvenserna och det innebär att vi måste utforma en gemensam kommunikations- och informationspolitik som även den ingår i den demokratiska processen.
Det är grunden för demokratin, så att folk förstår vad EU handlar om och känner att de är delaktiga i processen.
Jag lyssnar gärna till de budskap som sänts av Irlands folk, men när Kathy Sinnott talar om för oss, vilket hon gjorde i går, att majoriteten av väljarna i en stad röstade mot Lissabonfördraget på grund av att en avfallsförbränningsanläggning byggs där och vi har EU-lagstiftning som främjar avfallsförbränning, undrar jag verkligen vad det har med Lissabonfördraget att göra.
Vi har hört många sådana argument, och vi måste vara ärliga: alla argument är faktiskt inte helt relevanta eller värda att övervägas.
Vi måste fundera på ett nytt recept för ratificeringen av EU-fördrag.
Varje land måste få uttrycka sin åsikt och jag hoppas att det brittiska överhuset kommer att ratificera fördraget i eftermiddag och sända en tydlig signal om att processen fortsätter.
(EN) Herr talman! I eftermiddag kommer det brittiska parlamentet vid Westminster att slutföra ratificeringsprocessen av Lissabonfördraget.
Det kommer att vara uppiggande att läsa i pressen i morgon att britterna äntligen säger ja till EU.
Det kommer att göra mycket för att återställa Storbritanniens moraliska anseende och politiska trovärdighet och bör även hjälpa irländarna att nå ett nytt samförstånd som grundas på mindre libertas och mer veritas.
Det är bisarrt att Nigel Farage och hans högertrupper föredrar att låta en folkomröstning i ett främmande land styra och fatta ett beslut i stället för det brittiska suveräna parlamentet.
Det bekräftat min åsikt att en plebiscit - en allmän folkomröstning - är en form av demokrati som möjligen är lämpad för revolutionära omständigheter, men är fullständigt olämplig för informerade och överlagda beslut om en komplex fördragsöversyn.
Därför måste parlamentet hjälpa rådet att kommunicera innehållet i Lissabonstrategin.
(EN) Herr talman! Lissabonfördraget är dött.
Utan enhällighet är detta helt enkelt ett juridiskt faktum.
Väljarna, inte bara på Irland utan även i Frankrike och Nederländerna, har sagt nej till fördragstexten eller dess tvillingbror.
Om vi vill återvinna folkets förtroende måste vi göra mer än att bara ompaketera och döpa om Lissabontexten och försöka få igenom den.
Det nya fördraget var alltför lätt att förlöjliga och alldeles för komplext och svårfattligt för att förklara, vilket gör det svårt för jasägarna i en folkomröstning i vilket land som helst.
Många av ändringarna i Lissabonfördraget är bra, till och med nödvändiga, men de uttrycks på ett så oklart och obegripligt språk att knappast någon kan förstå det.
Det är upp till de övriga åtta medlemsstaterna att besluta om och hur de ska fortsätta med ratificeringen, men jag anser att det skulle hjälpa mycket om till exempel Storbritannien beslutade att göra detta genom en folkomröstning, så vi får se om vi har folkets förtroende för att fortsätta med den här processen.
(IT) Herr talman, mina damer och herrar! Om den irländska folkomröstningen är oviktig och obetydlig, varför hölls den då?
Varför beslutade man att det skulle finnas en möjlighet att hålla en ”plebiscit”, som vi har hört?
Det är allvarligt när ett parlament förnekar vikten av och vägrar ge folket fullständig yttrandefrihet, som det irländska folket har fått.
Detta valresultat är helt enkelt en vacker gravsten, med ett keltiskt kors på toppen, för utsikterna till en europeisk superstat, vilket våra befolkningar ogillar så starkt.
De vill inte att den politiska och även den monetära suveräniteten ska säljas ut.
Detta läge är hoppingivande för oss som, precis som det irländska folket, tror starkt på ett Europa av folk och regioner.
Av detta skäl begär även vi i Padanien en folkomröstning, även om fördraget rättsligt sett nu naturligtvis har förkastats och gått i graven.
Allt detta beror på det otroliga förfarandet att ett fördrag som påverkar våra folks framtid ska godkännas genom en parlamentarisk omröstning, som utestänger folket och medborgarna.
Som tur är finns det en fri nation som har en verklig frihetskänsla i venerna.
Kanske den styrkan kommer från att de har varit tvungna att kämpa för sin frihet.
Det är dags att inse den verkliga innebörden i detta röstresultat: man säger ”nu får det vara nog” till Brysseleurokraterna som vill bygga upp en superstat långt ifrån våra medborgares intressen och själ.
I Padanien känner vi oss alla som irländare i dag.
(CS) Herr talman! Efter den irländska folkomröstningen skäller den socialdemokratiska gruppens ordförande Martin Schulz på oss medborgare i de små medlemsstaterna, särskilt Irland och Tjeckien, med en typisk tysk dryg arrogans.
När så små länder blockerar den gemensamma reformprocessen måste vi enligt honom fråga dem om de vill vara kvar i EU eller inte.
Herr talman, jag kan försäkra er om (och ni kan vidarebefordra det, Martin Schulz) att nu när irländarna har tagit kål på denna sjukliga skapelse från det tyska ordförandeskapet som kallas för Lissabonfördraget, kommer tjeckerna gladeligen att begrava det och ändå fortsätta att vara EU-medlemmar.
De kommer att begrava Lissabonfördraget eftersom stadgan finns med där, och det kommer att leda till att möjligheten till ett återlämnande av Sudetenland-området öppnas för vårt land första gången på 60 år, och till en möjlighet att revidera ett rättvist resultat av andra världskriget i stället för de så kallade Beneš-dekreten. De kommer även att begrava fördraget eftersom de små medlemsstaterna berövas sin vetorätt och Tysklands röstetal i stället ökas från 9 till 18 röster.
Martin Schulz borde snarare fråga sig vilket resultatet hade blivit i Tyskland om tyskarna hade fått folkomrösta om Lissabonfördraget.
Jag gratulerar Irland och oss alla.
(CS) Mina damer och herrar! Att erkänna att Lissabonfördraget är dött och var en återvändsgränd är den enda demokratiska och ärliga lösningen.
I morgon är det hög tid att stats- och regeringscheferna äntligen inser att politiken i demokratier inte förs över gåsleverkanapéer i luftkonditionerade möteslokaler, och att de slutar att försöka styra över andra människors liv från Bryssel.
Den irländska folkomröstningen visar tydligt att folket inte tänker finna sig i beslut från ovan och arrogansen från unionens maktelit.
Rådet måste göra beslutsprocessen tillgänglig för allmänheten och sluta lura medborgarna.
Lär vi oss inte av vår historia?
Efter alla de blodiga händelserna på 1900-talet, vill den politiska eliten verkligen att de stora länderna ska fatta beslut för de mindre igen?
Var det inte tillräckligt för vissa premiärministrar och presidenter att ha levt en stor del av sina liv i en totalitär regim?
I morgon bör rådet friska upp grundkunskaperna: varför unionen skapades och vilka värden den bygger på.
Rådet bör respektera lagstiftningen och bestämmelserna och omedelbart förklara att en fortsatt ratificering av det nu begravda Lissabonfördraget är fullständigt meningslös.
(EN) Herr talman! Om ni tror att jag begriper mig på det irländska folkomröstningsresultatet så har ni fel, det gör jag inte.
Även om jag är djupt besviken på resultatet är jag säker på en sak: vi måste acceptera det som folkets demokratiska vilja och respektera det.
Vilken skräll för historieböckerna, när jag bakom mig här i dag ser en brokig skara av kolleger från extremhögern, inklusive Jim Allister och en gammal brittisk fängelsekund på köpet, alla iklädda grön tröja, som kräver respekt för det irländska röstresultatet.
(Protester från vissa ledamöter av IND/DEM-gruppen)
Hur annorlunda kunde inte historieböckerna ha skrivits om de brittiska kollegerna alltid hade respekterat det irländska folkets vilja!
Hur annorlunda kunde inte allt ha varit!
Hur många liv kunde inte ha sparats!
Jag välkomnar det - trots att det kommer mycket sent.
Vi måste alla respektera det irländska röstresultatet.
(Protester i bakgrunden)
Han hade mycket tid på sig för att öva bakom galler, så han kanske kan hålla tyst ett ögonblick ...
(Applåder)
En av de irländska ledamöterna här i parlamentet, som redan har talat under morgonen, delade ut valreklam med en injektionsspruta på under kampanjen.
Hon kanske kan berätta för parlamentet var dödshjälp förespråkas i Lissabonfördraget, och var i Lissabonfördraget det talas om abort, prostitution, beslut om företagsskatter och risker mot den irländska neutraliteten.
Jag väntar på sanningen.
Den irländska regeringen måste lugnt analysera resultatet för att utröna exakt vad i fördragstexten som våra väljare röstade mot och de måste komma med svar som inte bara är godtagbara för nejsägarna på Irland, utan även för alla de andra medlemsstaternas regeringar och medborgare som, enligt min mening, också har rätt att säga sin mening och uttrycka sin ståndpunkt, vilket vi också måste respektera.
Det krävs en välavvägd reaktion på de irländska väljarnas uppriktigt kända oro, men vi får inte vara undfallande mot extremisterna.
När dammet lägger sig hoppas jag att kollegerna kommer att hålla med mig om att ett Europa i två hastigheter inte är svaret, utan början till slutet för vår union, vår tids framgångsrikaste demokratiska fredsprojekt.
Det har alltid varit lättare att sprida fruktan än hopp.
En berömd irländsk politiker, en av våra egna - James Dillon - sa en gång: ”När en lögn berättas väl och tillräckligt ofta är det förbaske mig omöjligt för sanningen att någonsin hinna i fatt den.”
Jag lyckades inte med det.
Vi misslyckades med att få tillräckligt många av våra väljare att skilja fakta från fiktion, trots de tappra insatserna från vår valgeneral Gay Mitchell och mina kolleger.
Det är nu upp till vår nya Taoiseach, som har fått en olycklig början, att komma med en lösning.
(Applåder)
(EN) Herr talman! Vi får inte bara lyssna till vad som sägs om det irländska resultatet, utan måste fundera över och smälta det.
Men som det redan har påpekats måste vi också lyssna till de andra 26 länderna och ta hänsyn till deras resultat och även den oro som kan uttryckas under ratificeringarna.
Och sedan måste vi växa med uppgiften och ta itu med den enorma utmaningen att överbrygga klyftorna.
Om vi får 26 ratificeringar och ett förkastande är det varken orimligt eller odemokratiskt att fråga den stat som har sagt nej om den kan överväga möjligheten att anpassa reformpaketet, se över det, förklara det bättre och kanske söka en ny kompromiss i stället för att blockera alla reformer.
Det finns inget orimligt eller odemokratiskt med det.
Även en del av nejsägarna på Irland har trots allt erkänt att deras avsikt var att omförhandla för att nå en bättre överenskommelse.
En del - och vi har hört det från vissa håll i kammaren - vill bara lyssna till den ena sidan, till det svar som de vill höra, nämligen ett nej.
Jag vill lyssna till båda sidor och sedan finna en lösning som är godtagbar för samtliga 27 medlemsstater.
Det är den utmaningen vi alla måste visa att vi klarar av.
(FR) Herr talman! Det är självklart aldrig oväsentligt när folket röstar nej när de tillfrågas om EU:s framtid, och vi varken kan eller får nonchalera detta nej.
Vi måste tvärtom se det i vitögat och försöka bemöta det.
Som jag ser det finns det två frågor som vi måste ta itu med.
Den första handlar om demokrati.
Medborgarna förväntar sig att EU ska vara begripligt, synligt och förstående och tillhandahålla information och stöd.
Denna fråga berör alla, inte bara de nationella regeringarna.
Den berör även EU-institutionerna, särskilt kommissionen och rådet.
Det är den första frågan.
Den andra frågan handlar om EU:s känsla och själ, och som Martin Schulz just nämnde, unionens existensberättigande.
Varför byggde vi upp EU?
Unionen får inte bara inskränka sig till marknadsfrågor.
Vi skapade inte bara EU för konkurrensens skull, vi har slutit upp bakom gemensamma värderingar, vi har ett samhällsprojekt, vi har en samhällsmodell - en ekonomisk, social, hållbar och mänsklig samhällsmodell - och den modellen förtjänar att hjälpas fram, föras framåt och försvaras.
Det är vad våra medborgare förväntar sig.
Världen har förändrats en hel del sedan Romfördraget.
Vi måste gå tillbaka till där vi började och lägga en ny grund för det europeiska projektet för att kunna bemöta de kriser som vi för närvarande ställs inför - finanskrisen, livsmedelskrisen, energikrisen - men även hantera de avsevärda problem som vi måste ta itu med.
Hur kan vi skapa och utforma en mer hållbar och rättvis tillväxt av högre kvalitet?
Hur kan vi minska skillnaderna?
Hur kan vi åstadkomma en ny global balans?
Hur kan vi ompröva frågan om utvecklingsländerna och särskilt deras självförsörjning?
Det är dessa frågor som vi måste besvara och jag anser att det nu mer än någonsin är sista chansen för EU att återgå till politiken.
(DA) Herr talman! En ledande populär dansk affärsman skrev följande i gårdagens upplaga av tidningen Berlingske Tidende: ”Européerna stöder fullständigt internationellt politiskt samarbete och ansvar.
När EU-medborgarna förklarar sitt stöd för demokrati på nationell nivå stöder de naturligtvis demokrati på EU-nivå, och det är exakt vad som saknas.”
Vi har fått upprepade försäkringar om att Lissabonfördraget inte kan träda i kraft fast det bara är ett enda land som förkastar det, men vad skrev Hans-Gert Pöttering i sitt uttalande av den 13 juni?
(DE) ”Att ett EU-land har förkastat fördragstexten får inte leda till att de ratificeringar som redan har genomförts av 18 EU-länder inte är värda något.”
(DA) I enväldets tidsålder möttes kungar och kejsare för att dela upp makten mellan sig.
Dessa dagar är nu tillbaka.
Prins Pöttering, kejsare Barroso och härskarna över deras vasallstater har beslutat att EU-medborgarna inte betyder något.
Tjugosex länder fick inte rösta och Irland, det enda land som röstade, har upptäckt att det inte betydde något.
Unionen har inget folkligt stöd.
(DA) Herr talman! I fredags röstade det irländska folket nej till Lissabonfördraget, som är en dålig kopia av den konstitution som även Frankrike och Nederländerna röstade nej till.
Trots detta förklarar kommissionens ordförande att ratificeringen ska fortsätta.
Vi får höra att ett lands skepticism inte får bromsa utvecklingen.
Man får det att se ut som att det finns ett problem med det irländska folket.
Men så är det inte.
Klyftan finns inte mellan det irländska folket och EU, den finns mellan folket och EU:s stats- eller regeringschefer.
Klyftan finns inte mellan vissa EU-länder och de övriga EU-länderna.
Frankrike, Nederländerna och Irland vill inte hejda utvecklingen, de vill ha en annan slags utveckling.
Varför är det så svårt att förstå?
Vad Martin Schulz anbelangar skulle jag vilja säga till honom att han borde skämmas.
Ni jämför de som ni kallar ”antieuropéer” med fascister, men det är er retorik som är fascistisk.
Ni säger att antieuropéerna sprang upp och ned i trappor och gick ut och värvade röster.
Man behöver inte vara så historiskt medveten för att minnas vad som sades om de svarta förra århundradet.
Detta är skandal!
Ni borde skämmas!
(DE) Herr talman! Det irländska folket har sagt nej till fördraget och EU-magnaternas svar gjorde irländarna rasande, eftersom man nu kallar Taoiseach till Europeiska rådet för att ställas till svars för deras ”dåliga uppförande”.
Detta är barnsligt och ovärdigt grundarnas europeiska vision.
Det är emellertid ännu kortsiktigare att kräva att Irland ska uteslutas eller försöka driva igenom fördraget.
Om vi upprepar omröstningarna till det önskade resultatet uppnås kommer detta ohjälpligt att skada bilden av EU.
Vi har hållit 290 folkomröstningar i EU sedan 1990, men ändå har det hittills inte hållits några folkröstningar om mycket viktiga beslut som Turkiets anslutning eller införandet av euron, och vi får inte säga vår mening om något så viktigt som Lissabonfördraget.
Bryssels tolkning av vad demokrati är - att medborgarna endast förväntas ge sin välsignelse till EU:s beslut eller rösta för de parter som EU gillar - leder faktiskt tankarna till Sovjetunionen.
I stället för att ta anstöt måste EU acceptera irländarnas nejröst för vad den är: en chans till en ny inriktning, mot politik som inriktas på folket och EU-medborgarna.
(DE) Herr talman! Som Martin Schulz så vänligt påpekade finns det faktiskt många regeringschefer från PPE-DE, vilket visar att PPE-DE står närmare medborgarna och därför vinner fler val.
Trots detta är det ett faktum att allt fler tecken tyder på att vi måste finna en balans mellan rationell ekonomisk politik och socialpolitik.
Jag respekterar fullständigt resultatet av den irländska folkomröstningen.
Det jag däremot inte respekterar är de lögnkampanjer som vissa personer från vänstern och högern har drivit i ett försök att vilseleda folket och göra dem fientligt inställda till det enade Europa, detta enade EU som är det mest framgångsrika konceptet i vår kontinents historia, som har åstadkommit fred, frihet och välstånd.
(Applåder)
Vi måste erkänna att EU är särskilt gynnsamt för de mindre nationerna.
De sitter med oss runt bordet, de har platser här i parlamentet, och ingenting kan beslutas i EU utan deras medgivande, medan de stora nationerna tidigare kunde trampa ned de mindre.
Det är skillnaden i vårt EU, alla nationer är lika mycket värda, och det är vad ni försöker förstöra med era brittiska imperialiståsikter, herr Farage!
Vi behöver detta fördrag för att utvidgningen ska kunna fungera effektivt och för att skapa mer demokrati genom att överbrygga den demokratiska klyftan och stärka de nationella parlamenten.
Vi behöver det här fördraget för att skydda subsidiaritetsbestämmelsen och kunna övervinna framtidens utmaningar, från energikrisen till den organiserade brottsligheten, och för att ha resurser för att bemöta livsmedels- och oljepriserna och andra liknande utmaningar.
Allt detta kommer att raseras om vi inte förser oss med de instrument som fastställs i Lissabonfördraget, särskilt instrumenten för sociala rättigheter, nämligen stadgan om de grundläggande rättigheterna, och den ”sociala klausulen”, enligt vilken de sociala frågorna måste beaktas i utformningen och genomförandet av all politik.
Tjugosex medlemsstater kan nu ratificera fördraget och samtliga har åtagit sig att göra detta.
Det var Storbritannien som lärde mig att parlamentet talar för folket i en representativ demokrati och jag kommer inte låta UKIP-partiet rasera det jag har lärt mig från Storbritannien.
Dessa 26 medlemsstater kan ratificera fördraget genom en parlamentarisk process, och om den processen slutförs framgångsrikt kan det irländska folket överväga saken på nytt.
Vi förväntar oss förslag från Irland för att bevara sammanhållningen i vår gemenskap av 27, för jag vill inte se ett splittrat EU och jag vill inte se ett inåtvänt Europa.
Jag vill se ett EU som förblir en enhet av likar, med 27 länder, och det är därför jag stöder Lissabonfördraget.
(EN) Herr talman! Jag är mindre diplomatisk än de flesta av mina kolleger här i parlamentet.
Faktum är att lögner, usla lögner och statistik besegrade sanningen i den irländska folkomröstningen.
Lissabonfördraget har inte gått i graven.
Men Irlands vägval är ett suveränt beslut av det irländska solket.
De enda som kan ändra beslutet om fördraget är det irländska folket.
Om det sker eller inte beror på de diskussioner som kommer att inledas i morgon mellan den irländska regeringen och de andra 26 stats- och regeringscheferna.
Det finns inget trollspö.
Det kommer att ta tid att dra slutsatser.
Jag föreslår en ny tidsgräns för ratificeringen av Lissabonfördraget.
Att fastställa ett datum före valet till Europaparlamentet anser jag vara ett rimligt mål.
Om det irländska folket fortsätter att vara missnöjt med Lissabonfördraget i den form som slutligen överenskoms mellan oss och resten av EU, kommer Irland inte ha något annat alternativ än att omförhandla sin förbindelse med unionen.
Det skulle vara ett ödesdigert vägval för ert land.
EU har väldigt lite att förlora om Irland går ur, men Irland har allt att förlora om det går ur EU.
De globala utmaningar som vi alla står inför i denna ständigt föränderliga och sammanlänkade värld är tydliga: klimatförändringen, de demografiska förändringarna, migrationen och energikrisen, svälten och fattigdomen som dödar miljoner människor, osäkerhet för människorna, internationell brottslighet, och en identitetskris i praktiskt taget alla våra medlemstater som grädden på moset.
Problemen kommer inte att lösas genom att någon av medlemsstaterna gömmer huvudet i sanden och hoppas att problemen försvinner av sig själva.
Avslutningsvis vill jag uppmana EU att visa en verklig förmåga att skapa anständiga levnads- och arbetsvillkor.
Detta kommer att förstärka vår enighet och solidaritet och ge en positiv lösning på denna kris.
(Applåder)
(EN) Herr talman!
Om irländarna hade röstat ja, tror någon här att de gröna t-tröjor som syns i kammaren skulle ha haft texten ”Respektera det irländska omröstningsresultatet”?
Sanningen är att de varken respekterar irländarna eller demokratin.
De respekterar endast ett nej, och det är faktiskt ganska unikt.
När Sverige gick med i EU fanns det 12 medlemsstater.
Det var 1995.
I dag finns det 27 medlemsstater.
Det är en stor förändring och jag tror att det är mycket få som kan ifrågasätta att EU har blivit mycket, mycket bättre till följd av utvidgningarna och den starka utvecklingen.
I dag när vi diskuterar den irländska folkomröstningen kan vi säga att de som sa nej hela tiden hade fel hela tiden, och att det har visat sig att vi som förespråkade en framtida utveckling av EU hade rätt.
Låt oss alltså fortsätta på samma sätt som vi har nått dessa resultat på, med uthållighet, visioner, demokrati och respekt för alla medlemsstater.
Låt oss fortsätta med demokrati i varje medlemsstat med en ratificeringsprocess och respektera resultatet i de olika medlemsstaterna, samtidigt som vi fortsätter att vara uthålliga i våra insatser.
Vi måste gå längre när det gäller energimarknaden, den inre marknaden och hur vi ska kunna förbättra resultaten inom alla områden, men vi måste också ha klart för oss att Nicefördraget inte är tillräckligt om den utveckling och de visioner som vi har åstadkommit så mycket med ska kunna fortsätta.
Så låt oss fortsätta och låt oss vara det EU som säger ja.
Vi måste komma ihåg att nejsägarna inte har åstadkommit någonting i EU.
(Applåder)
(SL) Den här diskussionen är inte ny.
Vi hade redan en liknande diskussion när väljarna i Frankrike och Nederländerna förkastade konstitutionsfördraget, och vid den tidpunkten försäkrade kommissionen och rådet oss att ratificeringsprocessen skulle fortsätta.
Men sedan föll båda, tillsammans med parlamentet, för frestelsen att göra ett uppehåll i ratificeringsprocessen.
I dag är jag, trots att vi respekterar de irländska väljarnas beslut, för förslaget att vi inte ska stoppa ratificeringsprocessen, utan slutföra den.
Jag anser att det kommer att bli lättare att finna lösningar för att godta Lissabonfördraget om vi fortsätter än om vi återigen faller för frestelsen att stoppa processen på grund av en folkomröstning.
För det andra måste vi ha en sak kristallklar för oss: det finns en stor klyfta i uppfattningen av vikten av EU mellan den politiska eliten på hemmaplan, i de nationella cirklarna, i EU och bland majoriteten av våra medborgare.
Här måste vi fråga oss själva om parlamentet, rådet och kommissionen kan göra mer för att överbrygga denna kommunikationsklyfta och återigen inspirera våra folk med den europeiska tanken.
Jag välkomnar det slovenska ordförandeskapets planer för morgondagens rådsmöte, men föreslår att även den frågan diskuteras - en ny kommunikationsstrategi för dialog mellan medborgarna och EU - inte bara för att slutföra ratificeringen av Lissabonfördraget, utan även i andra aspekter.
(Applåder)
Herr talman! Det har talats om respekt här i dag och det råder inget tvivel om att vi måste respektera resultatet av den folkomröstning som hållits på Irland, där en del röstade ja och andra röstade nej.
Jag tror att vi alla är eniga om att vi även måste respektera de återstående länderna och därför fortsätta med ratificeringen.
Jag vill emellertid tala om respekt för demokratin och jag vill tydligt klargöra att folkets godkännande har samma värde som ett parlamentariskt godkännande, exakt samma värde.
Vi måste minnas vad ”r” står för, ”r” som i respekt.
För det andra har vi ”e” som i eftertanke.
Vi måste se på skälen till att det blev nej på Irland, vi måste anstränga oss för att förklara varför Lissabonfördraget är bättre än de befintliga fördragen, och det måste vi göra med fakta och siffror.
Vi måste förklara för folket att Lissabonfördraget - precis som den irländska hästen som vann Epsom Derby för några dagar sedan, som heter New Approach - också är en ”ny strategi”, vilket EU behöver för att ge mervärde till folket.
Efter ”e” som i eftertanke kommer ”l” som i lösning.
Vi måste finna en lösning, och i det avseendet vill jag vara fullständigt uppriktig: en del av nejanhängarna använde ett farligt och skamligt argument.
De sa: rösta nej och sedan kommer vi att omförhandla Lissabonfördraget till fördel för Irland”.
I detta sammanhang vill jag klarlägga att EU är en gemenskap av rättigheter, där samhällsmodellen råder och besluten måste respekteras.
Vi i Europaparlamentet förklarar tydligt att det inte kommer att bli någon omförhandling av Lissabonfördraget.
EU-medborgarna och parlamentet anser att den punkten är avgörande för EU:s vidare utveckling.
Vi som är för fördraget vill bygga vidare på det vi har.
Min fråga är: vilka alternativ läggs fram av dem som vill ha en nejröst?
Jag skulle vilja att de förklarade det för mig.
(FR) Herr talman! I dag är det den 18 juni och som fransman är jag uppfylld av uppmaningen från London: gör motstånd, fortsätt, härda ut och ge aldrig upp.
Ordet ”veto” skrivs med samma fyra bokstäver som ordet rösta - ”vote” - men det finns inget veto för de andra och därför måste vi fortsätta.
För övrigt är det sjätte gången det blir nej på nio folkomröstningar sedan Berlinmurens fall.
Det ger upphov till frågetecken.
Det sägs att EU inte är tillräckligt socialt; det kommer aldrig att vara tillräckligt socialt.
Det är inte tillräckligt demokratiskt; det kommer att förbli ofullkomligt.
Det är för byråkratiskt; det kommer alltid att finnas tekniker som kallas teknokrater.
Jag anser att EU genomgår en mycket allvarlig identitetskris.
Det var lättare förr.
I dag finns EU lite överallt, det är inte säkert på vad det betyder, på sin historia, sitt öde, och det är det vi måste tackla.
För att göra det behöver vi ett starkt ledarskap, och det är ur den synvinkeln som vi står lite ensamma.
(Applåder)
(IT) Herr talman, mina damer och herrar! Jag anser - som rådsordföranden och ordförande José Manuel Barroso båda har sagt - att det faktiskt finns ett antal andra punkter på dagordningen för morgondagens möte i Europeiska rådet, och inte bara resultatet av folkomröstningen på Irland.
Den här frågan har dock tagit upp praktiskt taget all tid av morgonens debatt.
Det är en viktig fråga.
Flera skäl har angetts och vi analyserar varför det irländska folkets svar blev som det blev, men i själva verket vann nejsidan endast med en snäv marginal över jasidan.
Mycket har redan sagts, men jag anser att vi måste hantera frågan om varför irländarna röstade som de gjorde på ett praktiskt sätt och diskutera hur vi ska fortsätta.
Mycket har redan tagits upp som sagt, men enligt min mening ligger svaret i det faktum att EU-medborgarna saknar information.
Det är allas fel, vi delar skulden, regeringarna bär skulden.
Generellt sett har det påpekats - och det håller jag med om - att regeringarna tar åt sig äran när saker går bra men när det går dåligt eller finns anledning till kritik, då är det alltid EU:s fel.
Jag håller fullständigt med om det.
Trots detta är ingen tvungen att stanna kvar i EU.
Jag anser att vi måste respektera resultatet av den irländska folkomröstningen.
Men vi måste respektera de andra 26 medlemsstaternas önskningar lika mycket, de är 18 för närvarande men kommer snart att vara 26.
Ingen ska tvingas att stanna kvar om de känner sig instängda.
EU måste gå framåt, det kan inte stå stilla.
Avslutningsvis anser jag att Europeiska rådet i morgon måste fatta ett tydligt beslut om en ny strategi - stats- och regeringscheferna kan göra detta - en ny strategi där de som vill vara kvar kan stanna kvar ombord, men EU måste gå vidare i det allmänna intresset.
(EN) Herr talman! Jag förmodar att UKIP-partiets ledares fixering vid bedragare beror på hans eget partis nära kopplingar till bedrägerier och bedragare.
För att återgå till debattens huvudtema står det klart att Lissabonfördraget inte kan träda i kraft den 1 januari som vi hoppades.
Vi måste vänta på att den irländska regeringen talar om för oss hur den anser att vi bör gå vidare.
Men under tiden bör de andra staterna utöva sin suveräna rättighet att ratificera fördraget.
Min egen medlemsstat kommer att slutföra sin ratificering i dag enligt sin mångåriga och allmänt respekterade parlamentariska tradition.
Under tiden fortsätter globaliseringen och den osäkerhet som den orsakar snabbt, vilket vi såg starka bevis för i den irländska folkomröstningen.
EU är en politisk process som är utformad för att hantera dessa frågor, så det är vad vi bör göra: se på millennieutvecklingsmålen, klimatförändringen och migrationen.
Hur bör vi agera?
Det är skälet till att jag kommer att försöka undvika alltför mycket inåtvänt institutionellt navelskåderi och i stället fundera över åtgärder som förbättrar alla våra medborgares liv.
Jag har emellertid en fråga till det slovenska ordförandeskapet: kan ni tala om för mig vilka följder det irländska folkomröstningsresultatet får för Kroatiens anslutning till EU?
(PL) Herr talman! Vi diskuterar förberedelserna för Europeiska rådet.
Jag anser naturligtvis att alla ledamöter som har talat har rätt om man ser till vissa större eller mindre grupper av medborgare.
Vi måste emellertid tänka på att den här debatten skulle ha sett helt annorlunda ut om den hade hållits i onsdags i förra veckan.
Vi skulle säkerligen inte ha diskuterat problemet med Lissabonfördraget.
I stället skulle vi ha diskuterat det europeiska folkets vardagsproblem.
Som läget är nu är EU-medborgarna inte särskilt oroade över att det irländska folket har sagt nej till Lissabonfördraget.
De är mycket mer oroade över bensinpriset på bensinstationerna och de andra problem som de möter i sin vardag.
Det skulle vara fel av oss att enbart inrikta dagens diskussioner och resultatet av toppmötet på Lissabonfördraget.
Vi måste inse att vi som politiker nu måste hantera två viktiga frågor.
En är hur vi ska tillgodose våra medborgares förväntningar på vardagen, och den andra är Lissabonfördraget och dess genomförande.
Genomförandet av Lissabonfördraget kommer att avgöra vår förmåga att hantera de frågor som engagerar det europeiska folket i framtiden.
Därför måste vi försöka skilja på dessa frågor och inte bara diskutera Lissabonfördraget, utan även de aktuella frågor som är av intresse för våra medborgare.
Vi måste förklara för medborgarna varför det kommer att bli lättare att lösa deras vardagsproblem om vi antar och genomför fördraget.
Vi måste förklara varför de institutionella lösningar som vi föreslår är bra för EU.
De föreslagna arrangemangen kommer att leda till ökad solidaritet och omsorg om varandra, och större respekt för vad vi står för i våra respektive länder.
Jag delar fullt ut synpunkterna att varje medlemsland har rätt att säga sitt.
Det är en demokratisk rättighet.
Jag har också den uppfattningen att Lissabonfördraget i flera avseenden är bättre än nuvarande fördrag.
Det gäller möjligheterna till fortsatt utvidgning och ökad öppenhet, men också arbetstagares rättigheter.
När jag besökte Irland och träffade fackliga företrädare under kampanjen fanns det en berättigad oro över att balansen mellan marknad och sociala rättigheter inte är den rätta i dag.
Också i Irland pekade man på domarna i EG-domstolen rörande Lavalmålet och Rüffertmålet.
De två allvarligaste konsekvenserna är följande: För det första är det inte lika behandling efter domarna.
De som kommer från medlemsländer med sämre löneförhållanden får nöja sig med minimilön och inte med lika lön.
För det andra blev strejkrätten inskränkt på ett sätt som är alldeles oacceptabelt.
De frågorna måste rådet och kommissionen ta sig an.
Det handlar om balansen mellan det sociala Europa och marknadens Europa.
Klarar vi inte av denna balans kommer medborgarna att vända EU ryggen.
Där har vi alla ett ansvar, alla tre institutionerna, och vi måste göra det snart.
(EN) Herr talman! Det finns inget problem med att respektera de irländska väljarna men vi måste respektera de beslut som har fattats av 18 demokratiskt valda nationella parlament i lika hög grad och dessutom visa lika stor respekt för de återstående åtta medlemsstaterna, och även låta dem fritt besluta om reformfördraget.
Med all vederbörlig respekt för det irländska folkomröstningsresultatet kan EU-27 inte tas som politisk gisslan av ett begränsat antal motståndare till Lissabonfördraget.
Det finns inget alternativ till reformen av EU.
Ja, EU kan stanna upp, men omvärlden kommer inte att stanna och vänta på oss, och den mest dramatiska skadan av detta röstresultat kommer att drabba Europas solidaritet: vår gemensamma utrikes- och säkerhetspolitik och energisolidariteten.
Det finns även en etisk dimension som vi bör betänka.
Denna folkomröstning är en varningssignal om att det krävs ett trovärdigt åtagande till våra grundläggande värderingar.
Våra medborgare kanske aldrig blir fullt informerade om detaljerna i fördragen, men de kommer alltid att kunna skilja mellan integritet och verkligt engagemang å ena sidan och halvsanningar och realpolitik å den andra.
I stället för att leva från ett nationellt val till ett annat, i stället för att hänge sig åt konsumentdemokrati som inriktas på att få mer och mer pengar från EU, behöver vi ledare som kan förmedla det budskapet till våra medborgare. ”Först av allt, vad kan ni göra för Europa?”
Och tro mig, om vi har sådana ledare kommer vi att finna medborgare som vill stödja oss.
(CS) Mina damer och herrar! För sex månader sedan åtog sig EU:s 27 stats- och regeringschefer att ratificera reformfördraget genom att skriva under dokumentet.
Jag vill att Europeiska rådet ska minnas det vid sitt möte på torsdag.
Jag vill särskilt att den tjeckiske premiärministern Mirek Topolánek ska påminnas om sin skyldighet att genomföra ratificeringen. Han hävdar, precis som den tjeckiske presidenten, att Lissabonfördraget har gått i graven och att det inte är någon mening att fortsätta med ratificeringen.
Jag vill särskilt uppmana de premiärministrar som hör till gruppen för Europeiska folkpartiet att påminna den tjeckiske ministern om hans skyldighet och det ansvar som tillkommer ett land som snart kommer att överta ordförandeskapet.
Eftersom Tjeckien kommer att ta över EU-ordförandeskapet den 1 januari 2009, det sista kapitlet i ratificeringsprocessen, kommer lösningen på hela problemet med Lissabonfördraget att vila på Tjeckiens axlar.
Jag upprepar att jag skulle vilja att gruppen för Europeiska folkpartiet påminner den tjeckiske premiärministern om hans skyldighet.
(RO) Det möte i Europeiska rådet som vi förbereder i dag är avgörande för EU:s framtid.
Ett av de mest välmående EU-länderna, som är ett representativt exempel på hur ekonomisk framgång kan nås genom EU:s integrationsåtgärder, har sagt nej till Lissabonfördraget.
Samtidigt har 18 EU-länder antagit dokumentet, de flesta av dem hör till samma grupp av 18 länder som också sa ja till det europeiska konstitutionsfördraget.
Jag är lika besviken över resultatet av Irlands folkomröstning som många av de föregående talarna.
Trots detta måste vi fortsätta med de reformer som EU så väl behöver.
Ett EU med flera olika hastigheter, för vilket det har funnits förfaranden ända sedan Amsterdamfördraget, och med väldefinierade undantagsalternativ är den enda vägen framåt för närvarande.
De länder som nyligen har anslutit sig till EU, t.ex. Rumänien, måste få samma chanser till utveckling som Irland har haft.
I tider som dessa måste vi minnas och återigen sluta upp kring de saker som enar oss och finna en anledning att fortsätta framåt.
I sitt berömda tal om ett ”Europas förenta stater” sa Sir Winston Churchill att det inte skulle finnas några gränser för européernas lycka, välstånd och ära om Europa enas kring sitt gemensamma arv.
Jag tror på den visionen, samtidigt som jag är medveten om vilka stora insatser som krävs för att åstadkomma detta.
Men det får inte hindra oss från att fortsätta.
(DE) Herr talman! Vi behöver förbättringar, inte bortförklaringar!
Trots detta måste det klargöras mycket tydligt att det är de nationella regeringarna som bär det största ansvaret för allmänhetens inställning till EU i våra medlemsstater.
EU-toppmötet i morgon och dagen efter måste leda till en sak: stats- och regeringscheferna måste be sina medborgare om ursäkt för den bristande ärligheten när det gäller gemenskapens beslut, för att de har misslyckats med att ge allmänheten lämplig information, för att ha misslyckats med att kommunicera med dem och deras bristande mod och integritet när det gäller deras del av ansvaret för de beslut som fattas i EU.
EU-politik är inrikespolitik.
Den måste därför vara integrerad i regeringarnas informations- och kommunikationspolicy.
Att göra EU till syndabock för alla problem i stället för att ta sitt ansvar och sedan be medborgarna om stöd två veckor före en folkomröstning är oärligt, oansvarigt och lömskt.
Här krävs det förbättringar.
(EN) Herr talman! Irländarnas nejröst visar att EU, ett oöverträffat och framgångsrikt exempel i världspolitiken, har svårigheter.
Men för att en folkomröstning verkligen ska utvisa folkets vilja måste den föregås av en informationskampanj.
I det irländska fallet kan vi mäta en grad av överensstämmelse, eller en total avsaknad av överensstämmelse, mellan Lissabonfördraget och argumenten mot det.
Demokratin kräver naturligtvis att vi tar hänsyn till det irländska resultatet, och det gör vi.
Men demokratin får inte heller utövas på bekostnad av andras rättigheter, nämligen de som redan har ratificerat Lissabonfördraget och, viktigast av allt, den får inte missbrukas av minoriteten för att utpressa majoriteten.
Jag är rädd för att den irländska nejrösten kommer att uppmuntra snarare än motverka de befintliga tendenserna att åternationalisera en del av den gemensamma politiken genom att förlänga det juridiska tomrum som EU har befunnit sig i sedan konstitutionsfördraget förkastades.
Avslutningsvis vill jag, som ledamot från ett före detta kommunistland som gjorde stora insatser för att komma med i EU, säga att jag skulle avsky att se att kommunismen lever längre än EU.
(PL) Herr talman! Det kan verka som att alla avtal som ingås i Lissabon är dömda att misslyckas.
Lissabonstrategin och Lissabonfördraget har båda slutat i fiasko.
Förra veckan förkastade Irland Lissabonfördraget i en folkomröstning.
Detta innebär att dokumentet nu är dött.
Vid det förestående toppmötet kommer man att bli tvungen att bedöma om det finns något hopp om att återuppliva fördraget.
Europaparlamentet bör sända en tydlig signal om att det godtar demokratins regler, även om vissa ledamöter kan vara missnöjda med resultatet.
Att förolämpa och tvinga Irlands folk är oacceptabelt.
Ett sätt att utöva acceptabla påtryckningar skulle vara att fortsätta ratificeringen av fördraget i andra medlemstater.
De extrema och oansvariga kommentarerna om möjligheten att utesluta ett så förmodat arrogant land från unionen är oroande.
Vi hoppas att Europeiska rådet kommer att överväga ett nytt och mer demokratiskt recept för EU.
(FR) Herr talman! Vi vet alla att demokratin inte är en stillaflytande flod, men vi vet också att det är den demokratiska metoden som vi har valt för att organisera vårt samhälle.
Jag anser därför att det irländska nejet inte är annorlunda än fransmännens eller nederländarnas nej, men att vi, precis som 2005, inte lyckades förklara varför EU är bra för våra medborgare.
Vi lyckades inte lugna dem i fråga om den miljökris som har drabbat dem.
Jag ogillar emellertid spekulationer och anser att vi bör vänta till dess att ratificeringarna har avslutas.
Men jag vill ändå uppmana rådet att sända en stark signal till medborgarna för att visa att det finns en verklig önskan om öppenhet och att förstärka demokratin till våra medborgares fördel.
Jag uppmanar rådet att öppna sina dörrar och att kommissionen och rådets ordförandeskap ska utses samtidigt som valet till Europaparlamentet.
Det skulle verkligen vara en stark signal och vi behöver ingen ratificering av fördraget för att göra den typen av ändringar.
(EN) Herr talman! Jag har lyssnat noggrant till den livliga debatten.
Ja, irländarna har talat och de har sagt nej.
Men en av de saker som oroar mig djupt är att de som röstade nej kände att det inte fanns några risker med att göra det, de trodde kanske att läget inte skulle förändras.
Nu framgår det mycket klart av debatten att andra länder anser att deras ratificeringsprocesser genom respektive parlament är lika mycket värda och att de kommer att fortsätta.
Irland kommer alltså att ställas inför ett dilemma och irländarna måste tänka över situationen om de övriga 26 medlemsstaterna ratificerar. Det är viktigt att vår Taoiseach Brian Cowen uttalar sig inom de närmaste dagarna och kommer med en analys av resultatet och eventuellt förslag om hur vi bör gå vidare.
Jag vill särskilt vända mig till Kathy Sinnott, som använde en del ganska förfärliga argument för en nejröst i sin kampanj.
När det gäller oron för att Irland förlorar sina värderingar vill jag påpeka för henne att vi inte kan skylla på EU för att värderingar går förlorade på Irland.
Det har vi åstadkommit själva, så vi måste sluta att vältra över ansvaret för det på EU och i stället se på våra egna materialistiska värderingar på Irland och på andra håll.
(PL) Herr talman! Jag är fast övertygad om att ratificeringsprocessen av Lissabonfördraget bör fortsätta.
För de länder som har undertecknat dokumentet är detta en internationell rättslig skyldighet enligt Wienkonventionen om fördragsrätt.
Fördraget medför en möjlighet till att göra de nödvändiga reformerna av EU.
Det kommer till exempel att bli möjligt att inrätta en gemensam energipolitik för EU.
Denna politik är mycket viktig för unionen och även för mitt land, Polen.
Den skulle garantera energisäkerhet för alla polska medborgare.
Jag företräder Silesien, som har en befolkning på fem miljoner personer.
För min region skulle en energipolitik vara en möjlighet till framsteg och utveckling, eftersom Silesien är rikt på energiresurser.
Jag ställer därför frågan: ska allt detta omintetgöras av det irländska nejet i folkomröstningen?
Jag respekterar resultatet av folkomröstningen på Irland, men samtidigt har jag svårt att godta att 109 964 irländares röster, som utgör skillnaden mellan nej- och jarösterna, ska få avgöra framtiden för mitt land, min region och i själva verket hela EU:s framtid.
Det får inte ske.
(DE) Herr talman! Jag vill tacka Irlands folk och även CAEUC, som kampanjade mot Lissabonfördraget på Irland.
Fördraget har nu förkastats tre gånger: en gång i Frankrike, en gång i Nederländerna och nu förkastandet av en något ändrad version av fördraget av Irland.
Vi måste faktiskt acceptera detta till slut.
Det får mig att tänka på Bertolt Brecht, som en gång sa: ”skulle det inte vara lättare i det fallet om regeringen upplöste folket och valde ett annat”?
Så tolkar jag ett antal av de uttalanden som har gjorts här.
Fördragets innehåll diskuterades faktiskt på Irland, särskilt den nyliberala inriktningen, inriktningen på militarisering och framför allt den odemokratiska karaktären.
Vi måste helt enkelt bara acceptera det här folkomröstningsresultatet.
Fördraget har gått i graven och vi behöver ett nytt.
För vår del kommer vi att mycket noggrant notera och dokumentera det flertal odemokratiska uttalanden som har gjorts här.
rådets ordförande. - (SL) Det ord som har hörts - och lästs - oftast i kammaren i dag har varit ”respekt”.
Här vill jag tillägga att vi även måste respektera vissa fakta, och jag vill lyfta fram följande punkter.
För det första: ratificeringen av ett nytt EU-fördrag faller inom medlemsstaternas exklusiva befogenheter.
Deras exklusiva befogenheter.
Rådet har absolut ingen roll i dessa processer, och ordförandeskapet ännu mindre.
För det andra: varje medlemsstat genomför den här processen enligt sina egna regler, som staten formulerar på sitt eget oberoende och suveräna sätt.
Det leder oss in på en kanske grundläggande punkt.
Vissa medlemsstater har genomfört en parlamentarisk ratificering eller kommer att göra det, och en är bunden av folkomröstning.
Men det betyder inte att det är något fel med parlamentarisk ratificering.
Jag avvisar bestämt påståendena från dem som anser att parlamentarisk ratificering är bristfällig eller mindre demokratisk än en folkomröstning.
Det är inte sant.
Det är inte sant.
Det finns absolut inget fel med parlamentarisk ratificering.
Från EU:s synpunkt är den fullständigt likvärdig andra demokratiska processer.
För det tredje: varje medlemsstat talar för sig själv.
De irländska väljarna talade för Irland.
De talade inte för någon annan medlemsstat.
Detta innebär att alla andra medlemsstater har exakt samma rättighet.
Arton medlemsstater har redan ratificerat Lissabonfördraget, de andra har inte uttalat sig än, och ordförandeskapet anser att ratificeringen måste fortsätta.
De som hävdar att Lissabonfördraget har gått i graven, de som kräver ett omedelbart stopp av ratificeringsprocessen, förnekar medlemsstaternas rätt att tala för sig själva, samma rätt som de så ivrigt försvarar i Irlands fall.
(Applåder)
För det fjärde: vi har redan varit i den här situationen och då fann vi en lösning.
Vi kommer att finna en lösning den här gången också, som bygger på anledningarna till att denna situation uppstod, men ordförandeskapet vill inte spekulera om detta.
Ordförandeskapet vill inte dras in i diskussioner om fördraget kanske är för komplicerat, om det var något fel med kommunikationen, eller kanske, som Proinsias De Rossa betonade, att det ljögs en massa.
Nej, vi kommer att låta våra irländska kolleger analysera skälen till detta resultat och även föreslå sin vision av en möjlig väg ut.
Och vi kommer att finna den vägen ut, det är jag säker på.
Vi kommer att finna den.
Europeiska rådets möte i morgon markerar början på vårt sökande efter en väg ut.
Den sista punkten: punkten på föredragningslistan för morgonens sammanträdessession var inte resultatet av den irländska folkomröstningen, utan förberedelserna inför Europeiska rådet.
Ordförandeskapet kommer att föra diskussionerna i Europeiska rådet enligt denna linje för att klargöra att EU inte har någon anledning att stanna upp, att EU fortsätter att fungera, och därför kommer vi att behandla ett antal frågor i linje med den planerade dagordningen.
Vi kommer att behandla problemen med livsmedels- och oljepriserna, vi kommer att diskutera ekonomiska, sociala och miljömässiga frågor, vi kommer att behandla utmaningarna i samband med den internationella utvecklingen och vi kommer att diskutera frågan om västra Balkan.
I detta sammanhang vill jag också svara Gary Titley - det blir inga direkta följder för EU:s utvidgningspolitik, som kommer att fortsätta, vilket även gäller den europeiska grannskapspolitiken och annan politik.
Tack till alla, och särskilt dem som gav sina åsikter om dessa andra frågor, och jag är säker på att Europeiska rådets möte kommer att bli framgångsrikt.
(Applåder)
kommissionens vice ordförande. - (EN) Herr talman! Jag vill tacka de ärade ledamöterna för deras mycket intressanta inlägg.
Det här är naturligtvis den rätta arenan för en debatt om demokrati och respekt för omröstningsresultat.
Irländarna röstade nej, så varför är detta inte över?
Varför säger inte EU bara: ”Fördraget har gått i graven, låt oss gå vidare?”
Varför insisterar vissa personer och medlemsstater på att genomföra sina egna ratificeringsprocesser?
Varför insisterar vi på att gå tillbaka till skälen till att vi inledde hela den här debatten om ett nytt fördrag för EU?
Jag vill gärna säga ett par ord om detta eftersom vi inte får glömma att EU-ledarna har investerat ett stort politiskt kapital i hela det här förfarandet.
Det har gått mycket tid och energi åt att diskutera de bakomliggande frågor och problem som gör det nödvändigt att utforma ett nytt maskineri för EU, som har förändrats så dramatiskt på så kort tid.
Jag vill bara nämna tre skäl till att vi anser att det krävs ett nytt fördrag.
För det första skulle ett nytt fördrag ge stadgan om de grundläggande rättigheter bindande kraft.
EU handlar inte bara om den inre marknaden - som någon påpekade - utan också människors och arbetstagares rättigheter.
Ett annat skäl är naturligtvis att vi vill kunna visa upp en enad front i världen, vara starkare på den internationella arenan och göra detta på grundval av våra värden.
Vi vill försvara oss på den internationella arenan, kämpa för en hållbar utveckling, diskutera oljepriserna, konfliktförebyggande och andra viktiga frågor.
Det är ett av skälen till diskussionerna om ett nytt fördrag.
Det tredje skälet är naturligtvis att göra EU mer demokratiskt.
Hur ironiskt är det inte med tanke på de som talar om att respektera nejrösten och resultatet, att fördraget i själva verket skulle ge mer makt till det direktvalda Europaparlamentet.
Detta skulle innebära ökat deltagande för de nationella parlamenten och att rådet måste hålla sina överläggningar offentligt, där medborgarinitiativet är en av de viktiga faktorerna i kapitlet om deltagande demokrati, som är en ny förbättring i fördraget.
T-shirt-partyt där borta har texten ”Respektera nejrösten”.
Min tanke om hur vi bör göra detta är bland annat att känna till vad som oroar det irländska folket.
Det är att förstå varför de röstade nej.
De har gjort sina egna tolkningar men jag anser att det är mycket viktigt att den irländska regeringen, med hjälp av opinionsundersökningarna från vår Eurobarometer, bättre förstår problemen och om det finns något vi kan göra åt dem.
Är det inte det som är tanken med demokrati?
Det är vägen framåt - att förstå deras argument, att arbeta tillsammans med de andra medlemsstaterna och även få deras respekt för de problem som vi förhoppningsvis kommer att lyckas lösa tillsammans.
Precis som vi gjorde efter nejrösten i de franska och nederländska folkomröstningarna har vi redan genomfört en Eurobarometerundersökning, som jag tror kommer att bidra till att förbättra förståelsen av utmaningarna i samband med folkomröstningar.
Att hålla en folkomröstning har sina fördelar, men även sina avigsidor - eller snarare utmaningar ur en demokratisk synvinkel.
Efter det att väljarna har förelagts en så komplex och omfattande text som ett nytt internationellt fördrag, finns det självklart rum för olika tolkningar av resultaten.
Vi måste förstå bättre vad irländarna sa, vad de är rädda för och vad de hoppas på.
Jag tolkar redan de preliminära resultaten som att detta inte är ett generellt nej till EU.
Det är också att förstå och respektera deras roll i EU.
Fördelen med att hålla en folkomröstning är att man måste informera och kommunicera med medborgarna, med alla utmaningar som det medför.
Alla inser säkert att vi även måste analysera hur vi kan förbättra kommunikationen och informationen till medborgarna.
Jag har alltid sagt att kommunikation är ett redskap för demokrati.
Detta måste bygga på medborgarnas rätt att veta vad som pågår på EU-nivå, vad som beslutas och hur medborgarna kan säga sin mening.
Detta arbete måste intensifieras ytterligare och det är skälet till att kommissionen kommer att fortsätta med det vi inledde för ett par år sedan, som vi kallar Plan D, som i debatt, dialog och demokrati.
Detta kommer att bygga på tanken att medborgarna ska ha ett egenansvar för EU-politiken ...
Fru kommissionsledamot, mina damer och herrar! Jag förstår att det blir lite stimmigt eftersom många kolleger kommer in i kammaren nu, men jag vill be dem som är på väg in att inte stå och småprata eftersom många eftersom många kolleger gärna vill höra kommissionsledamotens slutsatser.
kommissionens vice ordförande. - (EN) Herr talman! Jag försökte sammanfatta att vi behöver skapa ett medborgerligt egenansvar för EU:s politik, för att göra den begriplig och relevant och se till att EU-institutionerna är ansvarsskyldiga och tillförlitliga för dem som de tjänar.
Vi måste föra en bred och kontinuerlig debatt om EU:s framtid mellan de demokratiska institutionerna i EU och medborgarna, både på nationell nivå och på EU-nivå, och vi måste öka medborgarnas delaktighet genom att ge dem tillgång till information, så att de kan föra en informerad debatt om EU.
Vi har redan föreslagit att en ram ska inrättas för detta, som Jo Leinen redan har påpekat - och tack för att ni gör det.
Jag tackar Janez Lenarčič för att han försöker finna en lösning på detta.
Jag tackar även parlamentet för att det stöder insatserna för att förbättra effektiviteten i kommunikationen med medborgarna, eftersom vi måste ta detta på allvar och anslå de resurser och skapa den ram som vi behöver för att arbeta i partnerskap även med medlemsstaterna, och naturligtvis göra våra texter och beslut så lättlästa som möjligt.
Vi höll en debatt om det konsoliderade fördraget.
Det tog lång tid för rådet att godta det och offentliggöra en konsoliderad version av fördraget, men till slut gjorde rådet det, och detta är naturligtvis ett av de verktyg som vi har för att nå ut på ett bättre sätt till våra medborgare.
Vi måste fortsätta att dra slutsatser och dra lärdom av det irländska exemplet, men vi måste respektera deras nej.
Det gör vi bäst genom att verkligen ta reda på vad som oroade dem, genom att finna lösningar tillsammans och även låta de andra medlemsstaterna säga sin mening.
Jag hoppas att även denna debatt kommer att bli ett positivt bidrag till ledarnas möte i morgon och på fredag.
Ett varmt tack till alla för en bra och konstruktiv debatt.
(Applåder)
Tack, fru kommissionsledamot.
Debatten är härmed avslutad.
Jag vill informera parlamentet om att Hans-Peter Martin har begärt att få göra ett personligt uttalande enligt artikel 145 i arbetsordningen.
Enligt artikel 145 kommer jag att ge Hans-Peter Martin ordet när protokollet för detta sammanträde justeras.
Skriftliga förklaringar (artikel 142)
skriftlig. - (EN) Jag gratulerar hjärtligt väljarna i Republiken Irland för att de på ett övertygande sätt har förkastat den ompaketerade konstitutionen.
Genom att göra detta slog de ett slag för miljoner demokrater i EU, som förvägras rätten att säga sin mening genom ett totalitärt försök från EU-eliten att pracka på oss alla Lissabonfördraget.
Utmaningen för eliten är nu om de har ärligheten och integriteten att erkänna att fördraget är dött.
Lissabon satte upp sitt eget överlevnadstest. Enhällig ratificering.
Fördraget har underkänts i detta test på ett spektakulärt sätt.
Precis som sin föregångare konstitutionsfördraget stupar det över demokratins klippa.
I stället för att se verkligheten i vitögat fruktar jag att vi återigen kommer att utsättas för en konspiration från Bryssel för att kringgå folkets vilja.
Om ni gör detta kommer ni till slut att möta samma öde.
Så bespara er det besväret och erkänn att fördraget har gått i graven, utan några utsikter till att återuppstå.
skriftlig. - (EN) Jag vill hylla Lissabonfördraget i dessa tider av kris och institutionell osäkerhet.
Jag vet inte om det någonsin kommer att träda i kraft, men de som vill undvika populism anser att det är ett bra fördrag.
Det konstruerades och diskuterades naturligtvis inte lika demokratiskt som konstitutionsfördraget.
Det är naturligtvis inte en perfekt text - det finns inga perfekta texter.
Det är naturligtvis för komplext - men vilket EU-fördrag är inte det?
De som säger att de inte förstår Lissabonfördraget visar i själva verket att de inte har något förtroende för sina ledare.
Men det är en text som bidrar till att utveckla demokratin i EU.
Fördraget skulle göra EU öppnare, effektivare och mer socialt lyhört.
Ett enkelt exempel: om stadgan om de grundläggande rättigheterna hade varit i kraft skulle inte EG-domstolen ha kunnat fatta Viking- och Lavalbesluten, som är så skadliga för arbetstagarna.
Så vi behöver mer Europa, inte mindre.
Mer demokrati.
Mer politik.
Som socialister har vi nu en skyldighet att förklara för folket vilket slags nytt och annorlunda EU vi vill ha.
skriftlig. - (HU) Jag hör till dem som anser att saker och ting inte längre kommer att vara desamma i EU som innan irländarna röstade nej.
En sak som vi absolut inte får göra är dock att bortse från resultatet av den irländska folkomröstningen.
Jag hör emellertid även till dem som anser att vi måste fortsätta med ratificeringsprocessen, eftersom alla medlemsstater har samma rätt att uttrycka sin åsikt om EU:s gemensamma framtid.
Vi måste lösa detta komplicerade pussel genom att å ena sidan lyssna till de irländska medborgarna och å andra sidan vederbörligen beakta alla de andra medlemsstaternas inställning, som vill vandra vidare längs den gemensamma europeiska vägen.
Det är en svår ekvation, och vi måste ta varje tillfälle i akt för att bedöma läget.
För att göra detta behöver vi samtliga 27 medlemsstater.
Jag anser att alla de 27 medlemsstaterna måste finna en gemensam lösning och fatta ett gemensamt beslut om nästa steg.
Som kommissionens ordförande José Manuel Barroso sa: ”27 medlemsstater undertecknade fördraget, och vi måste göra allt som står i vår makt för att se till att samtliga 27 medlemsstater finner en väg framåt”.
Vi måste finna en lösning, ett sätt att bryta dödläget.
skriftlig. - (RO) Den europeiska processen måste fortsätta.
De irländska medborgarnas nej till Lissabonfördraget måste respekteras.
Samtidigt måste vi ta hänsyn till EU-medborgarnas intressen i ett bredare perspektiv genom att effektivisera EU:s struktur och fortsätta med utvidgningsprocessen.
De irländska medborgarna har inte bara rättigheter, utan även skyldigheter inom EU.
De måste vara medvetna om följderna av att de förkastade Lissabonfördraget.
De irländska medborgarna kommer att bli tvungna att i en ny folkomröstning besluta om de vill gå ur eller stanna kvar i EU på grundval av Lissabonfördraget.
Att avbryta den europeiska processen genom att åberopa irländarnas ”intakta suveränitet” innebär i själva verket att man sätter stopp för den naturliga önskan som medborgarna från Kroatien, Republiken Moldavien etc. hyser om att närma sig EU.
Precis som Irland och irländarnas politiska företrädare har rätt att kämpa för sina medborgares önskningar har Rumänien rätt att kämpa för Moldaviens anslutning till EU.
skriftlig. - (PT) Efter den segerrika nejrösten i den irländska folkomröstningen om Lissabonfördraget bör EU-ledarna nu erkänna det som är uppenbart: att Lissabonfördraget har misslyckats.
De vet att det bara krävs att en medlemsstat inte ratificerar ett fördrag för att det inte ska kunna träda i kraft.
Så är reglerna.
Det bör även noteras att förkastandet följer på två identiska resultat i Frankrike och Nederländerna om den så kallade europeiska konstitutionen, som var Lissabonfördragets föregångare.
Det enda som kommissionens ordförande har erkänt är emellertid att det kommer att ta tid och vara svårt att lösa det problem som har uppstått i och med den irländska folkomröstningen.
Han försöker lägga skulden på Irland och vägrar erkänna att problemet härrör från den djupa legitimitetskris som har uppstått till följd av den nyliberala, militaristiska och federalistiska politik som förs.
Europeiska rådet måste därför besvara en grundläggande fråga den här veckan: om ratificeringsprocessen av Lissabonfördraget ska avbrytas på grund av att det har gått under, eller om man ska inleda en debatt om de verkliga skälen till folkets missnöje och genomföra de nödvändiga politiska förändringarna för att tackla de nuvarande kriserna, med andra ord främja ökad social rättvisa och ökad anställningstrygghet med rättigheter, bekämpa spekulativa vinster och priser och prioritera kampen för social integration.
skriftlig. - (RO) Irländarnas folkomröstning nyligen har tolkats på olika sätt i EU och inläggen här i kammaren bekräftar de svårigheter som detta omröstningsresultat kan ge upphov till.
Jag vill kort nämna de problem som de irländska medborgarnas nejröst kan orsaka för den allmänna opinionen i de länder som nyligen integrerats i EU, särskilt de östeuropeiska länderna.
Medborgarna i dessa länder kommer att ha mycket svårt att förstå att de tvingas integrera dessa EU-normer, som medför ekonomiska uppoffringar, i den nationella ramen samt en rad offentligpolitiska frågor som medborgarna anser vara alltför restriktiva i det ekonomiska skede som dessa länder befinner sig i nu.
Här vill jag betona att alla försök att införa någon slags specialbehandling inom gemenskapsramen med all säkerhet kommer att ge utslag i det politiska valet 2009, vilket kan ge upphov till att den väljarkår som mycket entusiastiskt röstade för dessa länders anslutning till EU radikaliseras.
skriftlig. - (HU) Den irländska folkomröstningen kan tolkas på många olika sätt.
Den är en seger för folkets suveränitet, vi kan inte förneka detta enkla faktum.
Men samtidigt visste de flesta väljarna inte vad de röstade för, vilket framgår av att nejanhängarna byggde sin kampanj på historiska missnöjesanledningar som faktiskt hade lösts genom EU-medlemskapet.
Vi kan tycka att det är orättvist att 53 procent av väljarna i ett relativt litet land har makten att hindra 26 andra nationer från att fördjupa sitt samarbete och infria den europeiska drömmen.
En sak är dock säker, och det är att i framtiden måste vi diskutera integration med EU-medborgarna på ett mer intelligent, övertygande och lättförståeligare sätt.
Av detta skäl har Europaparlamentets utskott för kultur och utbildning tagit initiativet till ett betänkande med arbetstiteln ”Aktiv dialog med medborgarna om Europa”.
Jag har fått i uppdrag att utarbeta detta betänkande.
Jag ber mina ledamotskolleger att stödja vårt arbete genom att dela med sig av sina tankar, låt oss samla våra tankar, så att vi inte bara lär oss att förstå och stödja frågan om integration och samarbete, utan även ser till att EU-medborgarna gör detsamma.
skriftlig. - (PL) I dag diskuterar vi EU:s framtid.
Vi gör detta i kölvattnet av de känslor som väckts av resultatet av folkomröstningen på Irland.
Jag vädjar till alla berörda, parlamentets ledamöter och kommissionens och rådets företrädare, att avstå från att läxa upp Irlands folk och hota dem med en rad repressalier, inklusive uteslutning från EU.
Faktum är att unionen finns och den irländska nationens röst är inte en röst mot EU.
Enligt min åsikt är den ett uttryck för motstånd mot det dokument som kallas reformfördraget från Lissabon.
Det irländska folket förkastade just denna version av reformen som förelades dem.
Det är högst sannolikt att medborgarna i andra länder skulle ha svarat på exakt samma sätt om frågan hade avgjorts genom en folkomröstning hos dem.
Fördraget är när allt kommer omkring oförståeligt även för utbildade EU-medborgare.
Vi skulle göra klokt i att överväga om detta inte är en ny signal som visar att den så kallade eliten måste försöka överbrygga den avsevärda klyfta som finns mellan medlemsstaternas medborgare och ledarna för de politiska grupperingarna för närvarande, både på nationell nivå och EU-nivå.
I de berörda bestämmelserna i den internationella rätten anges det faktiskt att om en av parterna till ett internationellt avtal inte godtar avtalet är det inte bindande i den formen.
Detta står klart, oberoende av våra åsikter om dokumentet i allmänhet.
Irlands folk valde fritt.
Vi måste respektera deras beslut och söka positiva lösningar för EU:s framtid.
Som ordspråket lyder, vox populi, vox dei.
skriftlig. - (FI) Kris!
Kris!
På nytt ropar man att EU befinner sig i kris eftersom irländarna förkastade Lissabonfördraget i sin folkomröstning torsdagen den 12 juni.
Fördraget kan bara träda i kraft om det ratificeras av alla medlemsstater.
EU-ledarna efterlyser nya lösningar men få har något att erbjuda.
Det finns åtminstone två problem.
Lissabonfördraget är så dunkelt att det nästan är omöjligt att förstå.
Skulle ni vara beredda att underteckna det?
Dessutom verkar EU-eliten uppenbarligen vilja gå fram för fort.
Nu är det dags för de små medlemsstaterna att agera.
De bör insistera på att varje medlemsstat ska ha sin egen kommissionsledamot.
Det var ursprungligen Finlands och många andra länders önskan.
Om Lissabonfördraget fick effekt skulle det leda till en situation där varje medlemsstat skulle vara utan kommissionsledamot under en tredjedel av den tid man har till förfogande från 2014.
Ordalydelsen i fördraget är så vag att de små medlemsstaterna uppenbarligen i praktiken skulle vara utan kommissionsledamot längre tid än de stora medlemsstaterna.
Många tror att Irland förkastade fördraget delvis på grund av kommissionsfrågan.
Finlands kommissionsledamot är särskilt viktig för små medlemsstater, även om det är kommissionsledamöternas plikt att främja hela EU:s intresse.
I Finland är varje region glad om den har ”en egen” minister i regeringen.
Det är nu dags för EU-ledarna att noga tänka över vad som är orsaken till allmänhetens växande misstro mot EU.
Har unionen handlat i alla medborgares intresse på bästa möjliga sätt?
Har den ökat samarbetet på olika områden och expanderat för snabbt?
skriftlig. - (PL) Det beslut som fattats av Irlands folk har försatt EU i en svår situation.
Det visar också att EU bygger på aktiv demokrati.
Lissabonfördragets öde var inte uppgjort på förhand.
Liknande situationer har uppstått i det förflutna.
År 1993, efter ett negativt resultat om ratificeringen av EU-fördraget, beslutade Danmark att hålla ytterligare en folkomröstning.
Likaså beslutade man att hålla en andra folkomröstning på Irland efter katastrofen med ratificeringen av Nicefördraget 2001.
Jag är fast övertygad om att vi även denna gång måste respektera resultatet av den irländska folkomröstningen som ett suveränt beslut.
Unionen grundas på respekt för alla medlemsstaters rätt att uttrycka sin egen vilja.
Det måste tydligt framgå att förkastandet av fördraget inte innebär att det irländska folket motsätter sig unionen.
Det förestående mötet i Europeiska rådet utgör ett tillfälle att fundera över orsakerna till och följderna av den situation som har uppstått.
Detta får inte enbart begränsas till att läxa upp och kritisera Irland.
Rådet, kommissionen och parlamentet måste fundera över vad som kan göras för att européerna ska förstå fördraget och ledarnas avsikter bättre.
Jag är mot ett återinledande av förhandlingarna om fördragsreformen.
EU får inte bli ett Europa med två hastigheter eller mer.
EU måste visa för sina egna medborgare att det är ett gemensamt projekt genomsyrat av solidaritet.
Jag är övertygad om att rådet kommer att finna en lösning som är godtagbar för de länder som redan har ratificerat fördraget, för Irland och även för de medlemsstater som ännu inte har bestämt sig för hur de ska gå vidare.
skriftlig. - (PL) Resultatet av den irländska folkomröstningen skapade oordning i ratificeringsprocessen av reformfördraget.
Folkomröstningen visar oss även hur mycket energi vi faktiskt måste ägna åt vårt storslagna europeiska projekt för att skapa ett EU som kännetecknas av fred och solidaritet, vars främsta intresse måste vara medborgarnas välfärd och som spelar en stark roll på den globala ekonomiska och politiska arenan.
Vi har bevis för det höga pris vi får betala om vi inte engagerar oss i en dialog med våra samhällen för att förklara vad integration egentligen handlar om.
Ratificeringsprocessen måste fortsätta och jag är säker på att Irland kommer att göra allt det kan för att lösa den här situationen.
Jag håller med om de åsikter som uttrycktes av Martin Schulz, ledaren för den socialdemokratiska gruppen i Europaparlamentet, om att det sätt som kommissionen och Europeiska rådet fungerar på är ett av de underliggande skälen till det nuvarande läget.
Att utöka Europaparlamentets befogenheter som en demokratisk institution skulle bidra mer till att rationalisera unionen än storslagna förklaringar och program, eftersom de inte når medborgarnas hjärtan och sinnen.
skriftlig. - (ET) Mina damer och herrar! Dublins nej till Lissabonfördraget kom som en överraskning, eftersom det är med hjälp av EU-stöd som Irland har byggt upp en konkurrenskraftig ekonomi, stabiliserat arbetsmarknaden och skapat ett välfärdssamhälle.
Irländarna skulle kunna ha röstat för ett starkare och mer konkurrenskraftigt EU, som tjänar medborgarnas intressen bättre än tidigare.
Personligen anser jag att det visserligen är demokratiskt att folkomrösta om Lissabonfördraget, men på ett bedrägligt sätt.
Interna problem, som EU inte ingriper i, skapade oundvikligen spänningar som behövde luftas.
Därför är det lätt att skenbart skapa ett tillfälle för att uttrycka sitt missnöje, utan att bry sig om vad frågan egentligen handlar om.
De opinionsundersökningar som genomfördes före folkomröstningen visar även de på den fingerade demokratin och de spänningar som kom till uttryck, eftersom det framgick av undersökningarna att de personer som röstade nej inte kände till det verkliga innehållet eller visste särskilt mycket om vikten av Lissabonfördraget.
Det är upp till de irländska politikerna att besvara frågan ”varför”.
Irland har konsekvent varit en av de medlemsstater som mest har utnyttjat EU-stöden.
Irländarna är kända för sin positiva inställning till EU.
Därför är det ännu mer ironiskt att vi på grund av Irland blir tvungna att sätta stopp för skapandet av en starkare gemensam framtid.
Estland ratificerade Lissabonfördraget en dag före den irländska folkomröstningen.
Detta innebär att Tallinn, till skillnad från Dublin, har bidragit till att bygga upp denna gemensamma framtid.
Jag är en stark anhängare till ratificeringsprocessen, och jag tror på att Irland kommer att göra ett nytt försök att övertyga EU:s 500 miljoner medborgare om att även irländarna är stolta över att vara européer.
Dublins tacksamhetsskuld till EU är uppenbar.
skriftlig. - (EN) Herr talman! Även om resultatet av den irländska folkomröstningen blev en stor besvikelse för EU är det inte rätt tid att få panik och leta efter en syndabock.
Europeiska rådet ska hålla sitt möte den 19-20 juni i Bryssel.
Vi måste först ta oss tid att lyssna till förklaringarna från Taoiseach Brian Cowen och till hans förslag om hur vi bör gå vidare med Irland.
Enligt min åsikt måste de åtta återstående medlemsstaterna fortsätta med ratificeringen enligt planerna, trots Irlands nej.
Lissabonfördraget är absolut nödvändigt för en framgångsrik fortsättning på det europeiska projektet.
Det skulle vara otänkbart att inleda nya förhandlingar, eftersom EU har förhandlat om sin framtid under de senaste nio åren.
Med Lissabonfördraget skapas en mer förståelig, demokratisk och effektiv europeisk union och vi kan inte ge upp om detta ännu.
skriftlig. - (FI) Demokrati betyder bokstavligen folkmakt.
Det kan inte finnas demokrati utan folket och det är inte bra för folket att vara utan demokrati.
Irländarna fick chansen att rösta om den nya konstitutionen, Lissabonfördraget.
Det var demokrati och irländarna röstade nej på alla andra nationers vägnar.
Nejrösten stod för 53,4 procent av rösterna, och 46,6 procent röstade ja.
På Irland ville de inte att EU skulle gå mot en federation eller militariseras eller att det skulle bli ett ytterligare maktskifte till de stora ländernas fördel.
Federationstanken främjas av personer som är dåliga demokrater och dåliga förlorare.
De har börjat återuppliva den döda kroppen med tvång.
De förklarar att de små länderna inte behövs om de inte böjer sig för de större ländernas mycket verkliga makt.
På detta sätt blir de skyldiga till att EU-demokratin missuppfattas.
Irländarna kritiseras för hur de har utövat sina befogenheter, men ingen skrattar åt ungrarna, trots att det ungerska parlamentet röstade ja redan innan det ens hade hunnit granska det oläsliga fördraget.
Det irländska folkets beslut är demokratiskt, medan det ungerska parlamentets beslut inte är det.
Önskan att ha en konstitution för EU härrör inte från folkets behov, utan från elitens vilja att dela upp makten mellan sig.
Utan folkomröstningar kommer det att bli en kupp - både i de små och i de stora länderna.
skriftlig. - (EN) Medan vi håller dörrarna stängda för stater som Kroatien, Turkiet, Ukraina och Moldavien, som kämpar för att bli medlemmar, försöker vi hålla kvar stater som är osäkra på om det är värt besväret att vara medlemmar i en stark union.
Det är orättvist, föga lönande och ohållbart att behandla EU-skeptikerna bättre än EU-entusiasterna.
Lika respekt för alla nationer innebär att varje stat måste ta sitt eget ansvar.
Att försöka att lirka och fresta någon med illusoriska protokoll för att ändra beslut utan att ändra övertygelsen bakom dem, skulle vara en förolämpning och visa på bristande demokratisk respekt.
Det irländska folket bör ta så mycket tid som det behöver på sig för att fundera över sin europeiska framtid.
Den bästa ramen för en sådan demokratisk eftertanke kanske skulle vara ett tidigt val.
Hur som helst, irländarna måste använda sin egen tid och inte ta upp andras.
Därför måste man överväga en tillfällig status för Irland inom EU och låta den europeiska integrationsprocessen fortsätta med ett mindre antal medlemsstater.
Till slut bör det irländska folket genom en ny folkomröstning besvara frågan om de vill stanna kvar i EU på grundval av Lissabonfördraget eller om de vill spela en ”riddarroll” i den stormiga globala ordningen.
skriftlig. - (PL) Med hänsyn till det irländska folkets beslut i den senaste folkomröstningen är det ännu viktigare att Polen avslutar ratificeringen av Lissabonfördraget.
Om Polens president stoppar processen på grundval av argumentet om slutsignaturer, kommer han därmed att alliera vårt land med dem som är mot fördraget, i opposition mot den överväldigande majoritet som har godtagit det.
Detta skulle inte vara till vår fördel.
Tidigare har vi tagit till hot, en del skulle till och med kalla det utpressning, men vi gick med på en kompromiss.
Vi måste stå för följderna av denna kompromiss, särskilt efter resultatet av folkomröstningen på Irland.
Polen har faktiskt ett tillfälle att spela en roll i en viktig insats för att skapa ett starkt EU.
En snabb ratificering av fördraget kommer inte att vara en rutinåtgärd, utan en viktig politisk gest.
Jag anser att man kan ta för givet att innehållet i fördraget kommer att genomföras förr eller senare, med eller utan Irland.
Därför är det viktigt att vi befinner oss på rätt sida vid rätt tillfälle.
skriftlig. - (RO) Europaparlamentet och de andra EU-institutionerna måste respektera det irländska folkets röst i folkomröstningen.
Jag vill att det ska framgå mycket tydligt: de irländska medborgarna röstade inte mot EU, utan mot Lissabonfördraget.
Vi har fått tydliga signaler om att innehållet och grunderna för detta fördrag inte har förståtts, och det irländska folkets oro för beskattningssystemet och bevarandet av neutraliteten har spätts på av vissa politiska partier.
Europaparlamentet måste sända en tydlig signal till stöd för ratificeringsprocessen i de andra medlemsstaterna.
Samtidigt måste vi komma med genomförbara lösningar för de irländska medborgarna och den irländska regeringen så att de kan komma ur denna återvändsgränd.
Till syvende och sist är Lissabonfördraget ett nödvändigt steg framåt för att EU-institutionernas system ska fungera effektivare under de ännu svårare globala förhållanden som varje medlemsstat måste bemöta: den ekonomiska konkurrenskraften, klimatförändringen, prisökningarna på naturresurser och många andra aspekter som påverkar oss alla.
skriftlig. - (CS) Lissabonfördraget har blivit ett dött dokument, precis som när fransmännen och nederländarna förkastade utkastet till konstitution för EU.
Även om Europaparlamentets talman Hans-Gert Pöttering förklarade att syftet med fördraget var att skapa ökad demokrati, ökad politisk effektivitet och ökad klarhet och öppenhet och att ratificeringsprocesserna måste fortsätta i de medlemsstater som inte har ratificerat Lissabonfördraget ännu, är detta bara meningslösa fraser.
Om folkomröstningar hade hållits i andra länder än Irland skulle det irländska nejet säkerligen inte ha varit det enda.
Tänk på de knep som ”EU-eliten” tog till, som presenterade en text som inte var något annat än en avdammad och ändrad version av utkastet till EU-konstitution för ratificering!
Förutom irländarna skulle fransmännen och nederländarna säga nej igen, eftersom de opinionsundersökningar som har genomförts i dessa länder åtminstone visar så mycket.
De som ”styr” EU-politiken skulle äntligen inse att majoriteten av medborgarna förkastar unionen som ett militaristiskt och nyliberalt projekt som är fullständigt antisocialt!
Resultatet av den irländska folkomröstningen är inte en katastrof för EU som vissa vill få oss att tro.
Det är en chans att inleda en ny diskussionsprocess där de vanliga medborgarna äntligen får delta.
Irländarna röstade ju inte mot EU. De röstade mot innehållet i Lissabonfördraget, som skulle rasera den sociala standard som har nåtts hittills, och förvandla unionen till ett militaristiskt konglomerat.
Den så kallade europeiska tanken äventyras inte av dem som förkastar Lissabonfördraget. Den äventyras av dem som nu skriker att vi ska gå vidare eller vill införa ett EU ”med två hastigheter”.
skriftlig. - (FR) I morgon måste Europeiska rådet dra slutsatser från resultatet av den irländska folkomröstningen om Lissabonfördraget.
Det är upp till Irland att genom sin Taoiseach analysera detta folkomröstningsresultat och på nytt upprepa att landet vill att den europeiska integrationen fortsätter.
Jag hoppas att EU-27 enas om att fortsätta ratificeringsprocessen i de medlemsstater som inte har fattat ett beslut ännu, så att vi får veta varje lands exakta inställning till denna text.
Det slovenska och därefter det franska ordförandeskapet måste arbeta tillsammans med Irland för att försöka finna en rättsligt godtagbar situation för att en gång för alla sätta punkt för över 15 års insatser för att reformera det utvidgade EU:s funktionssätt.
Det franska ordförandeskapets ansvar kommer sannerligen att öka med tanke på att den europeiska ramen har rubbats och de globala marknaderna för råmaterial för livsmedel och bränsle rusar i höjden.
Europas folk känner tveksamhet.
Europeiska rådet måste visa dem att EU bidrar till att infria deras förväntningar genom att fatta beslut om de grundläggande frågorna.
Även om detta kanske inte löser den institutionella frågan omedelbart är det ändå det bästa sättet att visa irländarna att de har blivit hörda.
skriftlig. - (HU) Lissabonfördraget har förkastats av just det land som hittills har varit ett gott föredöme för hur man utnyttjar fördelarna med den europeiska integrationen så mycket som möjligt.
Den djupa förtroendekrisen i politiken åskådliggör även detta.
Dålig kommunikation när det gäller att visa på fördelarna med Lissabonfördraget spelade även in mycket i detta misslyckande.
Irland beslutade inte om fördraget, resultatet av folkomröstningen avgjordes av inrikespolitiska frågor.
Folkomröstning som institution har visat sig vara ett olämpligt instrument för att besluta om så komplexa frågor som denna.
Lissabonfördraget handlar inte bara om den institutionella reformen av EU, utan fördraget och stadgan om de grundläggande rättigheterna gör EU till en verklig politisk gemenskap och en värdegemenskap.
Det är en ny nivå i den europeiska integrationens utveckling i kvalitativa termer.
Det irländska folkomröstningsresultatet är ett stort problem, men det beror på oss om EU ska falla tillbaka i kris den här gången eller om det agerar snabbt och beslutsamt.
Det största misstaget i det nuvarande läget skulle vara att omförhandla den uppgörelse som det krävdes så stora ansträngningar för att nå, och därför bör vi behålla Lissabonfördraget som det är.
Nästan två tredjedelar av medlemsstaterna har antagit fördraget, inklusive Ungern, som var det första landet att göra det.
Ratificeringsprocessen måste fortsätta.
Irland måste bestämma sig så snart som möjligt om man vill fortsätta att vara en del av den fördjupade integrationen eftersom ett land inte får stå i vägen för de andra 26 länder som vill gå vidare.
Jag har fullständigt förtroende för att Europeiska rådet kommer att finna en väg ut ur denna situation vid det möte som inleds i morgon.
Arbetet med att bygga upp Europa måste fortsätta, och för att göra det behöver vi Lissabonfördraget.
skriftlig. - (RO) EU behöver en ny institutionell ram efter Nicefördraget, och Lissabonfördraget är en bra text även om det är mindre ambitiöst än den europeiska konstitutionen.
Arton medlemsstater har ratificerat Lissabonfördraget i sina nationella parlament.
Irland beslutade om ratificeringen genom folkomröstning, och irländarna förkastade fördraget.
År 2001 röstade Irland mot Nicefördraget också, för att ett år senare ratificera det.
Det irländska folkets röst visar att detta lands befolkning anser att gemenskapens institutionella uppbyggnad är komplicerad.
Det är vår skyldighet att förklara behovet av och bestämmelserna i detta fördrag för EU-medborgarna.
I fördraget hanteras frågan om klimatförändringen, EU-ekonomin definieras som en social marknadsekonomi, behovet av en gemensam energipolitik betonas, och i synnerhet ges den europeiska stadgan för de grundläggande rättigheterna rättsligt värde.
Detta reformfördrag bidrar till att öka demokratin genom att utöka Europaparlamentets befogenheter och ger hälften av de nationella parlamenten möjlighet att förkasta ett lagstiftningsförlag om de anser att det strider mot subsidiaritetsprincipen.
Det irländska folkets röst är en indikation på att vi måste visa ansvarskänsla och att det krävs mer dialog, att vi måste förklara bestämmelserna i detta nya fördrag för EU-medborgarna på ett mer detaljerat och bättre sätt, och även förklara varför det är nödvändigt.
skriftlig. - (PL) De EU-nationer som längtar efter frihet och suveränitet har nu anledning att tacka den irländska nationen.
Ett budskap av frihet och hopp har sänts ut, högt och tydligt, från lilla Irland.
Det budskapet måste fungera som en väckarklocka för demokratins fiender, som sätter sig över folkets vilja och bryter mot de tidigare överenskomna spelreglerna.
Frågan om vad man ska göra härnäst har uppstått.
Jag hävdar att vi i stället för att drömma om en ouppnåelig europeisk superstat bör inleda en debatt om nationernas rättigheter.
Vi bör först enas om en stadga om nationernas rättigheter och använda den som en grund för att fastställa principerna för den europeiska integrationen.
Mina damer och herrar, ni är EU:s arkitekter.
Jag uppmanar er att sätta stopp för manipuleringen och att låta folket avgöra sin egen framtid genom att ge dem sanningen.
Jag uppmanar er att låta nationerna leva i sina suveräna stater, som kommer att bestämma själva hur och med vem de ska samarbeta och hur och med vem de ska integrera sig.
Det irländska folkets rungande nej har gjort Lissabonfördraget omöjligt att genomföra.
Detta utgör ett avsevärt nederlag för rådet, kommissionen och Europaparlamentet, och även för centerhöger- och centervänsterregeringarna i EU:s medlemsstater (Ny demokrati (ND) och Pasok i Grekland).
Det är ett bakslag för kapitalismens företrädare i allmänhet, som spelade en ledande roll i att tysta ned nejrösten från Nederländernas och Frankrikes folk mot EU-konstitutionen, och genom att undertrycka den ökande rörelsen inom EU som protesterar mot och förkastar Lissabonfördraget.
Det är exakt dessa politiska krafter som bildar den stora alliansen i rådet, kommissionen och Europaparlamentet: gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater, socialdemokratiska gruppen i Europaparlamentet, gruppen Alliansen liberaler och demokrater för Europa, gruppen De gröna/Europeiska fria alliansen och andra anhängare till den europeiska ”monoliten”, med deltagande från Europaparlamentets ledamöter från Ny Demokrati och Pasok.
Vid parlamentets plenarsession den 20 februari 2008 röstade de alla mot förslaget att respektera det irländska folkets utslag och mot att hålla folkomröstningar om Lissabonfördraget i medlemsstaterna.
Rådets och kommissionens hårdhänta politik för att fortsätta ratificeringen av Lissabonfördraget är en autokratisk handling av förakt mot det irländska folkets vilja och folkens vilja i allmänhet.
De politiska gruppernas sammansättning: se protokollet
Anföranden på en minut om frågor av politisk vikt
Nästa punkt är anföranden på en minut om frågor av politisk vikt.
(EL) Herr talman! Konkurrenspolitiken är Europeiska kommissionens exklusiva befogenhet.
Man kan då fråga sig varför kommissionen inte utövar denna exklusiva befogenhet när oljepriset har gått upp med 50 procent sedan början av året.
Anledningen till oro är desto större eftersom kommissionen underlåtit att ta sitt ansvar på två fronter. Det gäller dels externt när det är uppenbart att en oljekartell har medverkat till att fastställa priser som är mycket betungande för de mer sårbara befolkningsskikten i EU, dels internt när en annan kartell på samma sätt upprätthåller extremt höga priser eftersom oljebolagens vinster fortsätter att vara överdrivet höga.
Jag uppmanar därför kommissionsledamoten med ansvar för konkurrensfrågor att ta sitt ansvar inom de särskilda områden där medborgarna förväntar sig detta - dvs. i frågor som rör deras dagliga liv.
(Applåder)
(HU) Tack herr talman! Allergier är vår tids farsot.
Allergierna har spritt sig i Europa efter andra världskriget och i dag är en tredjedel av alla barn allergiska.
Om vi inte gör något kommer i framtiden halva Europas befolkning att drabbas av denna sjukdom.
Kemikalier i livsmedel och förorenad miljö orsakar allergier, men allergiska symptom kan också utlösas av naturliga och syntetiska livsmedelstillsatser, kryddor, pollen och andra naturliga ämnen.
I Ungern är ambrosia det största problemet.
Tyvärr saknar EU för närvarande en allergistrategi, vilket kommissionen på min förfrågan bekräftat.
Civila samhällsorganisationer för allergiska sjukdomar och många miljoner europeiska medborgare som lider av allergier förväntar sig att vi ska agera mot allergier även på EU-nivå och att vi ska göra något för att förebygga och stoppa spridningen av allergiutlösande ämnen samt se till att sådana sjukdomar blir symptomfria.
En insats mot allergier skulle också visa att EU bryr sig om medborgarnas hälsa och problem i det dagliga livet.
Tack så mycket!
(EN) Herr talman! Vid toppmötet mellan EU och Ryssland, som hölls förra veckan i Khanty-Mansiysk, gavs klartecken för förhandlingar om ett nytt partnerskaps- och samarbetsavtal.
Förutom denna viktiga händelse höll president Toomas Hendrik Ilves och president Dmitri Medvedev det första officiella mötet på stats- och regeringschefsnivå mellan de två länderna på över 14 år.
Gränsfördraget mellan Estland och Ryska federationen var en av många frågor som diskuterades.
President Ilves förklarade att den ingress som det estniska parlamentet beslutat lägga till, och som den ryska duman sedan inte ratificerat, var onödig.
Kommissionsledamot Siim Kallas erinrade om att tillägget om fredsfördraget i Dorpat (Tartu) i ingressen endast var en inrikespolitisk provokation betingad av omständigheterna.
Jag kan inte se något skäl till att denna ingress inte skulle tas bort från gränsfördraget, eftersom fredsfördraget i Dorpat fortfarande är ett giltigt internationellt fördrag och man i det nya gränsfördraget bara fastställer kontrollinjen mellan Estland och Ryssland, de två ländernas gränser och EU:s externa gräns.
(PL) Herr talman! I förra veckan föreslog parlamentsledamot Silvana Koch-Mehrin, företrädare för det tyska Freie Demokratische Partei, att om Polen beslutade att inte ratificera Lissabonfördraget skulle landet uteslutas ur unionen.
Detta skandalösa yttrande var en kommentar till den polska presidentens uttalande i samband med frågan om det var någon mening med att skriva under fördraget efter fiaskot med den irländska folkomröstningen.
Enligt EU-lagstiftningen krävs det nämligen enhällighet i detta sammanhang.
Detta absurda yttrande från en kollega kan ses som ett uttryck för Europaparlamentets skamliga vana att inte ta hänsyn till de europeiska folkens vilja, något som innebär ett verkligt hot mot demokratins grunder.
Brist på respekt för resultatet av den irländska folkomröstningen och uppmaningen att utesluta Polen från EU är bevis för detta.
Länder som baserar sina ställningstaganden på gemenskapsrätten ska straffas bara för att de följer lagen.
Det är den sanna bilden av EU i dag.
EU befinner sig bara en hårsmån från totalitarism.
Jag vill uppmana alla mina kolleger här i parlamentet att visa större respekt för dem som valt oss.
Det är vi som förutsätts omsätta deras vilja i handling, inte tvärtom.
Vi får inte glömma det!
Herr Rogalski! Vi är mycket glada över att höra att er president har förklarat att Polen kommer att ratificera Lissabonfördraget.
Det är nämligen vad parlamenten enades om att göra.
(HU) Herr talman! I maj sände ledarna för den rumänska folkgruppen i Ukraina ett öppet brev till Rumäniens president där den lät höra sin röst genom ett enskilt uttalande mot Ukrainas diskriminerande utbildningspolitik som syftar till att helt avskaffa undervisningen i rumänska och med våld assimilera den rumänska folkgruppen.
Ungrare som bor i de ukrainska Subkarpaterna drabbas av samma minoritetsfientliga politik.
Enligt utbildningsministeriets dekret nr 461/2008 ska skolutbildningen för nationella minoriteter hädanefter bedrivas på Ukrainas officiella språk och undervisningen fullständigt anpassas till det ukrainska systemet.
Europaparlamentet och EU-medlemsstaterna, inklusive Rumänien och Ungern, fördömer Ukrainas systematiska försök att assimilera nationella minoriteter och uppmanar Ukraina att fullt ut uppfylla de internationella åtaganden landet har gjort när det gäller mänskliga rättigheter och minoriteters rättigheter samt bestämmelserna i den europeiska stadgan om regionala språk och minoritetsspråk som Ukraina också har undertecknat.
(PT) Herr talman! Jag skulle vilja använda detta tillfälle till att uttrycka vår solidaritet med de anställda i företaget Fapobol mot vilka ett disciplinärt förfarande har inletts med avsikten att avskeda dem för att de krävt att deras innestående löner ska betalas ut.
Efter det disciplinära förfarandet har Fapobols ledning vidtagit den oacceptabla åtgärden att sända ut meddelanden om uppsägning till de anställda, bland vilka många har arbetat i företaget mer än 35 år.
Hela företagsstrukturen berörs, inklusive arbetsgivar- och fackföreningsrepresentanter som deltagit i en demonstration där man krävde utbetalning av innestående löner.
Vi uttrycker vår solidaritet med alla arbetstagare och fackföreningsmedlemmar som drabbats av denna repressiva aktion och även med fackföreningen för de anställda i kemi-, läkemedels-, olje-, och gasindustrin i norra Portugal. Vi anser att företagets åtgärd bör fördömas i starkast möjliga ordalag här i parlamentet, eftersom man försöker skrämma arbetstagare och fackföreningsmedlemmar genom ett agerande som liknar häxjakt och som går stick i stäv med principerna om demokrati och frihet.
(BG) Ärade kolleger! Jag skulle vilja informera er om hur två bulgariska barns och deras föräldrars rättigheter åsidosatts i Nederländerna.
I juni 2006 omhändertog socialkontoret den bulgariska medborgaren Roumyana Ivanovas barn.
Roumyana Ivanova är bosatt i Nederländerna och barnen är fyra och fjorton år gamla.
Det enda tillåtna mötet med barnen avbröts eftersom modern talade bulgariska.
Föräldrarna har sedan dess inte träffat sina barn på ett år trots upprepade framställningar.
Barnen hålls åtskilda från varandra i strid mot lagen.
Flickan befinner sig i ett ungdomsfängelse för problembarn och myndigheterna lämnar inte ut några uppgifter om var pojken befinner sig.
Till och med ambassadören nekas ett sammanträffande och får ingen information.
Det bulgariska statliga organet för skydd av barn och även andra organisationer fortsätter att sända in ansökningar om att barnen ska kunna få växa upp i Bulgarien i enlighet med artiklarna 5, 9 och 20 i FN:s konvention om barnets rättigheter som föreskriver rätt till kontakt med föräldrar och rätt till uppfostran och omvårdnad i hemlandet.
De nederländska myndigheterna har hittills inte uttalat sig.
Jag är övertygad om att den bulgariska och europeiska allmänheten inte passivt kommer att åse hur internationella konventioner överträds och inte heller att den kommer att acceptera ett andra Libyenfall, fast denna gång i hjärtat av Europa.
Jag uppmanar er att klart och tydligt ta ställning i denna fråga och framföra detta ställningstagande till de nederländska myndigheterna.
(BG) Herr talman! Bron är en symbol för förening och den finns på alla sedlar från 5 till 50 euro.
Men det finns en bro i Europa som, även om den kallas vänskapens bro, fortfarande splittrar folk.
Det är den enda bron mellan Bulgariens och Rumäniens 350 kilometer långa flodgräns som utgörs av Donau.
Att korsa bron fram och tillbaka kostar nästan 17 euro.
Avgiften är obefogad och utgör ett hinder för både handel och människors fria rörlighet.
Den avspeglar inte den verkliga kostnaden för underhållet av bron.
Under 2007 uppgick de insamlade avgifterna till tolv miljoner på den bulgariska sidan, medan bara 17 000 euro investerades i brons underhåll.
Jag är övertygad om att om det görs en anmälan till EG-domstolen kommer domstolen att förklara avgiften olaglig.
Men varför skulle invånarna i Rousse och Giurgiu vänta på det?
Jag uppmanar de bulgariska och rumänska myndigheterna att gå medborgarnas förväntningar till mötes genom att avskaffa avgiften för att passera bron mellan Rousse och Giurgiu.
Jag uppmanar också kommissionen att försöka finna en lösning på detta för allmänheten så angelägna problem.
(ET) Min kollega Toomas Savi har redan nämnt Khanty-Mansiysk, en liten stad i Sibirien där toppmötet mellan EU och Ryssland ägde rum i slutet av förra månaden. Det var också platsen för en annan mycket viktig händelse, nämligen den femte finsk-ugriska världskongressen där presidenter från fyra länder deltog - Ryssland, Ungern, Finland och Estland.
En femmannadelegation från Europaparlamentet var också närvarande vid kongressen. Vårt huvudsyfte var att rikta uppmärksamhet mot de små finsk-ugriska folken, varav 19 lever i Ryska federationen, och att uppmärksamma det faktum att dessa folks språk och kulturer riskerar att utplånas.
Förhoppningsvis kommer den överenskommelse som grundlades vid toppmötet mellan EU och Ryssland i Khanty-Mansiysk också att innebära att man kommer att uppmärksamma den tyvärr bedrövliga situationen för de mänskliga rättigheterna.
(SK) Jag välkomnar att temat för rådets junimötet mellan EU:s hälso- och sjukvårdsministrar var ett initiativ med rubriken ”European Antibiotic Awareness Day”.
Syftet är att göra medborgarna medvetna om att antibiotika måste användas på ett ansvarsfullt sätt och bara i indikerade fall.
Felaktig användning är på väg att bli ett allvarligt hot mot folkhälsan.
Bakterier blir alltmer resistenta vilket leder till att antibiotika kommer att kunna användas i mycket begränsad utsträckning i framtiden.
Kampanjen drivs av Europeiska centrumet för förebyggande och kontroll av sjukdomar (ECDC), EU:s institutioner och Världshälsoorganisationen.
Det ska kompletteras av nationella strategier.
En workshop om bakterieresistens kommer att hållas i Paris och det tjeckiska ordförandeskapet förbereder en konferens om ämnet.
En logo har också framställts för kampanjen.
(RO) Herr talman, kära kolleger! Jag välkomnar Europeiska kommissionens initiativ som innebar att direktivet om gränsöverskridande vårdtjänster antogs i förra veckan.
Fördelen med det här förslaget är att det skapar en tydlig lagstiftningsram genom vilken regler fastställs för hur europeiska medborgare kan utnyttja vårdtjänster inom EU-området, i en annan medlemsstat än den där de bidrar till hälso- och sjukvårdssystemet, och även hur patienterna ska få ersättning för sina utgifter.
Förslaget, som skulle ha lagts fram för antagande i Europaparlamentet och rådet för länge sedan, är efterlängtat och lägligt, i synnerhet som hälso- och sjukvård undantogs från direktivet om avreglering av kommersiella tjänster.
Fram tills i dag var europeiska medborgare tvungna att hänvisa till EG-domstolen som i samtliga fall fastställde att medborgarna hade rätt till medicinsk behandling och som tvingade medlemsstaterna att ersätta deras utgifter.
Jag är fast övertygad om att detta direktiv kommer att få positiva effekter. Det kommer att främja hälsotillståndet för de medborgare som av olika skäl inte kan begära sådana tjänster i sitt ursprungsland och det kommer att öka de medicinska förfarandenas kvalitet i EU-området.
(PL) Herr talman! Vi polska ledamöter av Europaparlamentet har blivit mycket oroade på grund av situationen i Vitryssland, ett land som gränsar till EU.
Vitrysslands parlament har nyligen antagit en mycket restriktiv rättsakt om yttrandefrihet som kan leda till ytterligare begränsningar av den redan hårt begränsade yttrandefriheten i Vitryssland.
För att rättsakten ska träda i kraft behövs bara diktatorn Alexander Lukashenkos underskrift, vilket är en ren formalitet.
Rättsaktens mycket repressiva karaktär kommer framför allt att påverka oberoende journalister och förläggare.
Den innebär helt klart att man sätter munkavle på de fria medierna i Vitryssland, på den oberoende allmänna opinionen och på det framväxande civila samhället.
Europaparlamentet måste med tanke på denna situation framföra en erinran om de grundläggande normer som gäller på vår kontinent där Vitryssland ingår.
Det faktum att parlamentet för tre år sedan gav Sacharovpriset till Vitrysslands journalistförbund är ännu en anledning till att vi bör agera.
(DE) Herr talman! Platsen för toppmötet mellan EU och Ryssland valdes inte av en slump.
Khanty-Mansiysk är centrum för Rysslands oljeutvinning.
I det nya partnerskaps- och samarbetsavtalet lägger Ryssland tonvikten på ekonomin.
Utifrån ett EU-perspektiv borde de mänskliga rättigheterna betonas i större utsträckning.
Under Dmitri Medvedevs regim befinner sig Alexander Lebedev och Michail Chodorovski fortfarande i fängelse.
Förra veckan hotades de båda av nya anklagelser som kan leda till fängelsestraff på upp till 20 år.
De ryska myndigheterna utnyttjar tiden tills Medvedev tydligt tar ställning.
Det är mycket angeläget att Moskva gör framsteg och ger bindande löften i denna fråga. Man måste också lösa de politiska morden och klargöra situationen när det gäller inskränkningarna i press- och yttrandefriheten.
I framtiden måste EU visa fram en enad front och tala med en röst till Moskva för att öka den politiska pressen på landet.
Det handlar om ingenting mindre än EU:s trovärdighet.
(BG) Herr talman! De senaste veckorna har det i pressen förekommit kommentarer om att Europeiska kommissionens inställning till de olika medlemsstaterna skulle ge uttryck för dubbelmoral.
Naturligtvis kommer varje ny utvidgning att leda till en allt strängare tillämpning av kriterierna.
Bulgarien och Rumänien till exempel är föremål för en hittills okänd mekanism för samarbete och kontroll när det gäller rättsliga och inrikes frågor.
Det finns utan tvivel problem och de två länderna måste i hög grad reformeras, men har Europeiska kommissionen samma inställning till alla?
Det finns länder där den organiserade brottsligheten har fått grundligt fotfäste och där konsekvenserna är uppenbara: missbruk av EU-medel, underutveckling, gatuvåld och främlingsfientlighet.
Men jag har inte hört en enda officiell kommentar eller något förslag till motsvarande åtgärder från kommissionens sida.
När man talar om korruption i maktens korridorer kan jag föreställa mig hur kommissionen skulle reagera om en bulgarisk premiärminister införde en lag som skulle skydda honom från att ställas inför rätta.
Sådana åtgärder låter man emellertid passera under tystnad när det handlar om det land som den tidigare kommissionsledamoten för rättsliga och inrikes frågor kommer ifrån.
Jag skulle kunna citera flera andra exempel.
För att tala i klartext: jag begär inte några kompromisser för Bulgariens och Rumäniens del, jag begär en rättvis och jämlik behandling av varje medlemsstat.
(SK) I mars 2003 när Castros regim orättfärdigt dömde och fängslade 75 kubanska dissidenter införde EU sanktioner mot Kuba.
Mer än 50 politiska fångar, vars familjer vi under lång tid stött genom en slags ”adoption”, hålls också fängslade under inhumana villkor i kubanska fängelser.
Vi är bekymrade över deras dåliga hälsotillstånd.
Har de ansvariga, innan EU:s sanktioner mot Kuba upphörde, frågat Sacharovpristagarna ”Kvinnor i vitt” om situationen för de mänskliga rättigheterna och medborgerliga friheterna på Kuba har förändrats efter Raul Castros tillträde?
Herr talman! Jag vill tacka er för ert personliga engagemang i frågan om frisläppandet av politiska fångar på Kuba, och jag vill om igen be er att på Europaparlamentets vägnar uppmana den kubanska presidenten att omedelbart släppa alla kubanska dissidenter.
(CS) Mina damer och herrar! Ett centralt gemensamt värde i EU är dess språkliga och kulturella mångfald.
En hel rad stater har antagit stadgan om minoritetsspråk vid sidan av den egna lagstiftningen till stöd för denna mångfald.
En av dessa stater är Tyskland.
Jag vill framhålla att enligt kraven i stadgan ska minoriteternas kulturella institutioner ges finansiellt stöd.
När det gäller Załožby za serbski lud (föreningen för det sorbiska folket) har anslagen gradvis skurits ned genom åren.
Detta är inget gott exempel på hur stadgan efterlevs.
Vi uppmanar den tyska regeringen att hålla sina löften.
Vi bör inte tillåta att ännu en nation försvinner från Europas karta.
(EN) Herr talman! I förra månaden kunde Mohammed Omer, en ung palestinsk journalist från Gaza som arbetar för försoning och fred med israelerna, med stöd från den nederländska regeringen resa till EU och motta ett pris för sin journalistiska gärning.
På återvägen blev han anhållen, förödmjukad, slagen och torterad av den israeliska underrättelsetjänsten.
Den nederländska regeringen har enligt vad jag hört uttryckt sin bestörtning, men detta uppträdande från Israels sida ingår i ett mönster.
Varför överväger vi att inleda närmare förbindelser med Israel när den israeliska regeringens agenter utför sådana våldshandlingar mot just de människor vars arbete för fred och försoning stöds av den stora majoriteten av ledamöterna här i parlamentet?
Varför stöder vi sådana initiativ när vi vet att Israels regering inte kommer att göra minsta ansträngning för att kritisera eller fördöma dessa handlingar?
(CS) Mina damer och herrar! Den fria rörligheten för människor inom Schengenområdet är förvisso ett positivt europeiskt värde.
Det innebär emellertid fri rörlighet för många och olika slags samhällsfiender.
Tack vare informationssystem och Europols och Interpols insatser fungerar jakten på kriminella och rymlingar ganska bra, men vi stöter regelbundet på problem när det gäller att verkställa de avhjälpande åtgärder i form av straff som domstolarna utdömer.
Jag tänker på åtgärder som förbud mot att bedriva viss verksamhet, obligatorisk psykiatrisk eller sexuell behandling och alla former av övervakning av människor som villkorligt frisläppts från fängelse.
Arbetet med ett europeiskt informationssystem bör utan tvivel påskyndas. Framför allt bör man se till att nationella institutioner blir skyldiga att inte bara bidra till ett sådant system utan också hämta lämpliga uppgifter från det.
(RO) Före Rumäniens anslutning till EU hördes många röster här i Europaparlamentet som hävdade att romerna diskrimineras i Rumänien.
Av den anledningen har flera icke-statliga organisationer publicerat olika undersökningar på detta område.
Rumänien har hela tiden hävdat att romerna är en angelägen fråga för myndigheterna, men man kan inte säga att diskriminering sker.
Rumänien har genomfört program för integrering av romerna i samhället, huvudsakligen i form av utbildning och till och med positiv särbehandling.
Efter 2007 har romerna, och inte bara romer från Rumänien utan även från andra östländer, spritts runt om i Europa av ekonomiska skäl, men främst på grund av sina nomadtraditioner.
Detta har inneburit ett tillfälle för dem som gav råd att tillämpa detta själva.
Tyvärr har EU inte lärt sig något av det som har hänt i Italien.
Det är oacceptabelt att ta fingeravtryck på EU-medborgare, särskilt barn, och det är inte normalt att sätta eld på läger, med myndigheternas tysta medgivande.
Jag anser att romernas situation är ett ämne för gemenskapen, och jag uppmanar alla ansvariga - EU:s institutioner, regeringar och icke-statliga organisationer - att vara med och utforma en gemensam, sammanhållen politik för romernas integrering som helt grundas på EU:s principer.
(EN) Herr talman! Jag vill demonstrera vår solidaritet med arbetarna på Fujitsu i Birmingham som hotas av friställning.
Det finns planer på att utlokalisera delar av Fujitsus verksamhet till Förenta staterna, och det kan innebära att upp till 140 personer förlorar sina jobb.
Den fackförening som är inblandad i fallet är kommunikationsarbetarnas fackförening, och den har varit beundransvärt flexibel i kontakterna med Fujitsus ledning.
Det enskiftssystem som de föreslog Fujitsu skulle ha räddat 60 jobb. Men i styrelsens slutliga beslut den 30 juni, som inte föregicks av något tecken från styrelsen på att ett beslut skulle fattas så snabbt, avvisades alternativa förslag utan vidare.
Jag vill be Fujitsu att överväga utlokaliseringen på nytt eller åtminstone se till att bara de som går frivilligt behöver sluta och att de som vill fortsätta jobba kan göra det.
I EU:s lagstiftning stadgas klart och tydligt att ett företag måste ha samråd med sin anställda, och ändå fortsätter arbetsgivarna att göra för lite och för sent för att följa denna lagstiftning.
(FR) Herr talman! Jag skulle vilja ställa en administrativ fråga som rör parlamentet.
I mer än två år har tjänsten som direktör för Europaparlamentets kontor i Luxemburg varit vakant.
Tjänsten har utannonserats en gång, för ett halvår sedan.
Kandidater valdes ut men inget beslut fattades sedan jag ställt frågor till förvaltningen. Ert sekretariat, herr talman, har inte heller kunnat ge mig något svar.
Jag vill veta om det finns några särskilda skäl till varför denna tjänst inte har besatts och varför de utvalda kandidaterna inte har förordnats.
(RO) Kommissionens arbetsprogram för 2008 omfattar, bland de strategiska initiativen, antagandet av ett paket för utvecklingen av miljövänligare transporter.
Under hösten kommer kommissionen att lägga fram ett lagförslag om översyn av Eurovinjettdirektivet 2006/38.
Syftet med översynen är att se till att transportinfrastrukturen används på ett mer effektivt sätt samt att minska de negativa effekterna för miljön av transporter, grundat på principen ”förorenaren betalar”.
Detta direktiv får allt större betydelse, med ökande bränslepriser.
En hållbar ekonomisk utveckling av unionen är också beroende av att man utvecklar mer miljövänliga och effektiva transporter i energihänseende.
Jag hemställer hos Europeiska kommissionen att internalisering av externa kostnader som uppkommit genom transporter ses i ett större sammanhang, genom att man också ser över de låga mervärdesskattesatser som tillämpas i unionen samt direktiv 2001/14 om beskattning och uttag av avgifter för utnyttjande av järnvägsinfrastruktur och direktiv 2003/96 om energibeskattning.
(NL) Herr talman! För tio dagar sedan inledde vi vår kampanj mot barnsexturism på www.sayno.eu.
Varje år reser tusentals män från Europa, Förenta staterna, Australien och Korea till fattiga länder i Sydostasien, Afrika och Latinamerika inom denna motbjudande form av turism, och de kommer nästan alltid undan utan straff.
Det budskap vi vill föra fram med detta medborgarinitiativ är att detta inte längre är acceptabelt.
EU kan heller inte längre blunda för detta, och vi måste bland annat stärka Europols roll.
Det gläder mig att kunna berätta att vi, på denna mycket korta tid, redan har samlat in 14 000 underskrifter.
Kampanjen fortsätter naturligtvis.
Jag vill också framföra ett tack för det breda stöd kampanjen har fått, också från ledamöter av Europaparlamentet.
Inte bara ledamöter från min egen grupp, gruppen Alliansen liberaler och demokrater för Europa, har skrivit på. Jag har också sett namn på ledamöter från gruppen för Europeiska folkpartiet (kristdemokraterna) och Europademokrater, den socialdemokratiska gruppen i Europaparlamentet, gruppen Europeiska enade vänstern/Nordisk grön vänster och andra på listan - vilket självfallet är högst välkommet.
Jag vill passa på när det franska ordförandeskapet är närvarande och tacka den franska regeringen för dess tidigare initiativ på detta område, oftast i opposition mot andra medlemsstater.
Jag hoppas att ni inte har blivit avskräckta av det utan kommer att utarbeta ytterligare initiativ under detta halvår också.
(PL) Herr talman! För flera månader sedan hade vi en debatt här i kammaren om situationen vid varvet i Gdansk.
Företrädare för alla grupper pekade på behovet av verklig konkurrens mellan europeiska varv och andra varv på världsmarknaden, särskilt den koreanska varvsindustrin.
De betonade att avvecklingen av två av tre stapelbäddar skulle omöjliggöra för varvet i Gdansk att konkurrera och innebära att dess chans att överleva försvann.
Vi sammanträder i Strasbourg, en stad som symboliserar den europeiska integrationen.
Att bibehålla denna symbol som Europaparlamentets säte kostar hundratals miljoner euro varje år, men vi har respekt för denna symbol.
Varvet i Gdansk är en symbol för kommunismens fall och integrationen mellan Västeuropa och Central- och Östeuropa.
Det skulle vara värdefullt att låta denna symbol förbli en levande ekonomisk verksamhet, en arbetsplats för tusentals anställda.
Detta var den vädjan som de demonstrerande varvsarbetarna i Bryssel nyligen riktade till Europeiska kommissionen.
(FR) Herr talman! Jag vill fästa er uppmärksamhet på de nyligen inträffade händelserna i Tunisien, i gruvområdet i Gafsa.
Under flera veckor har möten organiserats mot fattigdomen i detta område, som är rikt på fosfater.
Lokalbefolkningen får ingen del i vinsterna, och vi kan nu se ett mycket allvarligt förtryck av polis och militär, med trakasserier, fängslanden, arresteringar och städer som stängs - jag talar här om Redeyef.
Jag ber chefen för EU:s delegation - och jag framför min begäran genom er, för jag menar att det krävs att Europaparlamentet ingriper - att denna fråga tas upp till diskussion med de tunisiska myndigheterna.
(RO) Yttrandefriheten är en grundläggande princip i Europeiska unionens stadga om de grundläggande rättigheterna.
Varje land måste garantera yttrandefriheten och se till att det finns förutsättningar för oberoende medier.
Journalistförbundet i republiken Moldavien påtalar emellertid de mediefientliga åtgärder som skett 2001-2008 från regeringen Chisinau.
De ingrepp som journalisterna nämner, som regeringen använt sig av för att försöka få politisk kontroll över offentliga medier är följande: Censur av information, polisutredningar riktade mot journalister för spridande av åsikter som går emot statens politik, olika falska anklagelser, snedvridning av konkurrensen i pressen, maximala begränsningar av utrymmet för debatt i offentlig radio och tv.
Mot bakgrund av dessa åtgärder anser jag att EU borde övervaka respekten för yttrandefriheten i detta land mera noga.
(HU) Jag skulle vilja återge vad András Léderer, ordförande för det ungerska liberala partiet Ny generation, har sagt.
I lördags inleddes den ungerska demonstrationen för värdighet i Budapest.
Liksom tidigare år uppmärksammades kampen för att minska fördomar mot homosexuella, om så bara för en dag.
Efter angreppen med molotovcocktails de senaste veckorna deltog många hundra medborgare som sympatiserar med homosexuella i tåget.
Demonstrationståget möttes av ett våld utan motstycke.
Många civila, poliser och demonstranter skadades, även kanslichefen vid det ungerska liberala partiet, Gábor Horn, och en socialdemokratisk ledamot av Europaparlamentet, Katalin Lévai.
Sedan högerrörelsen Magyar Gárda bildades har flera nynazistiska extremhögerportaler fortlöpande organiserat aggressiva angrepp, dels mot ett judiskt biljettkontor, dels mot romska bosättningar. Nu senast drabbades homosexuella.
Regeringen är uppenbarligen svag och de rättsliga myndigheterna oförmögna att åstadkomma resultat. Tack så mycket.
Jag vill uppmärksamma er och det franska ordförandeskapet på frågan om Europaskolorna. De tjänar som riktmärke och modell för utbildningen i Europa men ändå tar man där ingen hänsyn till inlärningssvårigheter (dyslexi, stamning) som gör att många barn hindras från att nå framgång i skolan och efterföljande yrkesliv.
Vi har sett misslyckanden och elever som hoppar av skolan, vilket leder till stora problem för deras föräldrar - våra kolleger i parlamentet och EU-tjänstemän. De tvingas flytta så att deras barn kan gå i vanliga skolor i medlemsstaterna där man är lyhörd för särskilda behov hos barn med inlärningssvårigheter, såsom lagen och mänsklig värdighet kräver, särskilt mot bakgrund av barns skyddsbehov.
Parlamentet kommer att få ytterligare tillfällen att fundera över de problem som dessa barn ställs inför.
(EN) Herr talman! Det som händer i Zimbabwe är fruktansvärt sorgligt och avskyvärt.
Robert Mugabe, som fordom kämpade för frihet från kolonialväldets slaveri, har nu blivit en hänsynslös diktator och en barbarisk förtryckare av rättvisa och mänskliga rättigheter för miljoner landsmän.
Det internationella samfundet - inklusive EU - har uttömt sina krafter med retoriska uttalanden, fördömanden och i stort sett verkningslösa sanktioner.
Det har blivit dags för omval.
Robert Mugabe borde därför ställas inför en internationell brottmålsdomstol för brott mot mänskligheten.
Jag är övertygad om att en sådan åtgärd är helt och hållet motiverad och realistisk, och det kommer att ge den angelägna efterlängtade effekten, nämligen att hjälpa folket i Zimbabwe att bli av med det totalitära styre som för landet mot dess ruin.
Jag menar att EU måste gå före för att Robert Mugabe ska ställas inför rätta i den internationella domstolen.
(EL) Herr talman! Jag vill återigen här i Europaparlamentet ta upp en fråga som gäller fiskarna i mitt land, Medelhavsfiskarna och alla som bryr sig om miljön.
Grekerna, och europeiska fiskare i allmänhet, är föremål för strikta begränsningar - med rätta - när det gäller fiskemetoder, redskap, fiskeperioder etc.
Tredjeländer - de turkiska fiskarna är ett typiskt exempel - fiskar dock hur och när de vill, med de redskap de själva väljer, vilket leder till en minskning av fiskbestånden och att haven och miljön fördärvas.
Jag menar att vi bör ta initiativ i fråga om Turkiet, så att landet använder riktiga fiskemetoder.
Miljön är viktigast, och när jag talar om Turkiet syftar jag självfallet på alla tredjeländer som använder sig av icke standardiserade fiskemetoder.
(FR) Herr talman! Också jag gläds åt att välkomna det franska ordförandeskapet, med den franske ministern Jean-Pierre Jouyet här hos oss.
Det stämmer att det är ovanligt att ordförandeskapet är här på en måndag, även om det gäller dessa frågor.
Jag vill ta upp utposteringen av poliser, kravallpoliser, utanför parlamentet i dag.
När jag kom hit tidigare gick jag igenom två poliskedjor.
Jag undrade vad som kunde utgöra ett sådant hot mot parlamentet att en sådan ansamling av kravallpoliser skulle posteras ut.
Två gånger blev jag tvungen att intyga min identitet - jag blev tillfrågad vad jag gjorde på Europaparlamentets område.
Jag blev verkligen överraskad, herr Jouyet, för jag känner mig inte hotad här utan tvärtom känner jag mig ganska betryckt av alla dessa avspärrningar.
Jag vill påminna er om att det är ett märkligt sätt att inleda det franska ordförandeskapet, att omringa EU-folkets hus med kravallpoliser, och jag vill gärna framhålla att vi vill att detta ska fortsätta vara ett folkets hus, som är öppet för medborgarna.
(SK) Eftersom vi inte kommer att träffas på nytt förrän efter den 21 augusti, 40-årsdagen av Warszawapaktstruppernas ockupation av Tjeckoslovakien, känner jag att det är min plikt att uppmärksamma dessa dramatiska händelser.
Då framgick det tydligt att kommunistregimen innebar ett brott mot mänskligheten, precis som alla totalitära styren.
Efter augusti 1968 upplevde vi i mitt hemland ytterligare 20 år av olika former av kommunistiskt våld och terror från detta organiserade ondskans maskineri.
Vi bör visa respekt för dem som inte gav sig och som uppträdde med värdighet.
Tillåt mig parafrasera några ord av den slovakiske prästen Anton Srholec, ordförande i den slovakiska organisationen för politiska fångar: ”Vi får aldrig upphöra att vittna om att det finns hundratusentals hedervärda människor i Slovakien som gjorde insatser för att bevara friheten och de mänskliga rättigheterna.
Det är tack vare dem som vi återigen är på demokratins, frihetens och rättigheternas sida.”
(HU) Tack så mycket.
Det ryska toppmötet kommer att äga rum i staden Khanty-Mansiysk i den sibiriska provinsen Yugra, och om två dagar kommer den femte världskongressen för de finsk-ugriska folken att äga rum där.
EU ger också ekonomiskt stöd till de finsk-ugriska folken för deras kamp att bibehålla sin identitet.
I talen från den närvarande EU-delegationen och de fyra statsöverhuvudena, särskilt det ungerska statsöverhuvudet, har betonats hur viktigt det är att hotade folk inte bara har dansgrupper och körer utan också får utbildning i sitt modersmål och självbestämmande.
Denna kongress har två budskap till EU.
Det första är att Europeiska året för interkulturell dialog inte bara ska vara ett år för dialog mellan de stora folkens kulturer.
Det andra är att vi står inför obegripliga företeelser när ett parlament i ett europeiskt land vill rösta om att landet ska vara enspråkigt, när det i det landet finns 75 regionala språk.
Om EU och Ryssland anser att det är viktigt att bevara kulturer och modersmål för de folk som bor på deras territorier borde detta också vara ett exempel för EU-medlemsstaterna att följa.
Tack.
(PL) Fru talman! Några veckor före de olympiska spelen i Peking slutade den enda oberoende nyhetskanalen New Tang Dynasty Television att sända till Kina.
Denna situation har nu varat i flera veckor, och vi vet fortfarande inte vad som orsakade stoppet, som rapporterades av satellitoperatören Eutel Communications. Vi vet inte heller när det kommer att rättas till.
Men vi vet vem som tjänar på detta stopp, och vem som förlorar.
Miljoner kunder till oberoende tv-utsändningar utan vinstsyfte på kinesiska och engelska tvingas genomlida censur av information från de kinesiska myndigheterna, information om hur effektivt de kinesiska styrkorna handskas med tibetanska terrorister.
De vill inte höra om strejker, oroligheter och problem under anordnandet av spelen.
Vi medborgare och företrädare för EU behandlar Kina med den respekt som landet obestridligen förtjänar, som en stor nation som har gjort en stor insats för hela mänsklighetens kulturarv.
Det är synd att vi i gengäld behandlas så oerhört nonchalant av myndigheterna i Peking.
Efterlevnad av överenskommelser och respekt för samma principer är något vi måste kräva, både av oss själva och våra kinesiska partner.
(EL) Fru talman! Enligt en artikel i New York Times för några dagar sedan emotses en överenskommelse mellan den amerikanska regeringen och Europeiska kommissionen som kommer att möjliggöra för europeiska regeringar, banker och företag med säte i EU att lämna över information om EU-medborgare till amerikanska organ, såsom kreditkortstransaktioner, uppgifter om gjorda resor, e-postmeddelanden och besök på webbplatser - allt för att försöka bekämpa terrorismen.
Förhandlingar pågår om EU-medborgares möjligheter att väcka talan mot den amerikanska regeringen om de anser att deras personliga rättigheter kränks till följd av behandlingen av deras personuppgifter.
Jag uppmanar talmannen och ledamöterna i Europaparlamentet att titta närmare på frågan, och jag uppmanar Europeiska kommissionen att komma med klargöranden, så att parlamentet får information om innehållet i och arten av dessa samtal.
Det är Europaparlamentets plikt att skydda individens rättigheter och den personliga integriteten för EU-medborgare, om dessa kränks.
(EN) Fru talman! Jag vill ta upp frågan om de stigande oljepriserna, särskilt terminsmarknaden för olja.
Det finns många skäl till prisstegringen på oljemarknaderna.
En är efterfrågan, den andra är tillgången och de låga investeringarna i infrastrukturen för olja under många år.
Fackmän inom oljeindustrin och oljemarknaden tar hela tiden upp den löjligt låga initialsäkerheten för råoljeterminer, som ligger på mellan 5 och 7 procent.
Med andra ord, om man vill köpa oljeterminer till ett värde av 10 miljoner euro behöver man bara investera en halv miljon euro.
Trimtabs Investment Research, en ledande oberoende amerikansk forskningstjänst, har sagt att om initialsäkerheten höjdes med mellan 25 och 50 procent, vilket är vad de flesta som investerar på aktiemarknaden betalar, så skulle det få en avgörande inverkan för sjunkande oljepriser.
Den låga initialsäkerheten på marknaden innebär att marknaden går att manipulera - det råder inget tvivel om det.
För mig är det inget problem att folk investerar i terminer och råvaror, men detta är en löjligt låg initialsäkerhet.
Vi måste gå vidare i denna fråga.
Initialsäkerheten måste höjas, för konsekvenserna på världsnivå är enorma och vi måste göra allt som är möjligt för att få till stånd ett lägre världsoljepris.
(PL) Fru talman! Den polske presidenten har beslutat att inte skriva under ratificeringen av Lissabonfördraget, efter att ha förklarat fördraget för dött, i ett läge där irländarna har avvisat fördraget i en folkomröstning.
Den polske presidenten erinrade om den grundläggande principen för EU:s funktion, nämligen att fördrag träder i kraft först när alla EU- medlemsstater har ratificerat dem.
Hittills har tillämpningen av denna princip varit självklar, och den tillämpades efter att fransmännen och nederländarna hade avvisat konstitutionsfördraget.
När så skedde förklarades konstitutionsfördraget för dött, men ratificeringsprocessen för det fortsatte ändå i många länder.
Tyvärr hördes röster i EU, både efter folkomröstningsbeslutet på Irland och efter den polske presidentens beslut, även från framstående politiker, med krav på att Polen skulle ratificera fördraget, vilket är ett förnekande av den europeiska demokratins själva väsen.
Jag vill protestera å det starkaste mot dessa röster, de påtryckningar och den speciella typ av utpressning som de utövar.
Därmed är anförandena på en minut om frågor av politisk vikt avslutade.
Budgetkalender: se protokollet
4.
Ändring av förordning (EG) nr 881/2004 om inrättande av en europeisk järnvägsbyrå (
Röstförklaringar
Muntliga röstförklaringar
(LT) I dag har vi i Europaparlamentet antagit resolutionen om gemensamma regler för tillhandahållande av lufttrafik i gemenskapen vid andra behandlingen.
Vi ändrar den förordning som har varit i kraft sedan 1992, och jag skulle återigen vilja framhäva de ändringsförslag som är viktigast för våra medborgare och framför allt för flygplanspassagerare och besättningar.
Jag syftar på de föreliggande åtgärder som skulle göra det möjligt för oss att få insyn i flygpriser och att bli mer aktiva när det gäller att förbjuda vilseledande reklam och ohederlig konkurrens inom flygtrafiken.
De ändringsförslag som syftar till att garantera större efterlevnad av flygsäkerhetsnormerna samt de sociala bestämmelserna för flygplansbesättningar är viktiga.
Det ser ut som om alla meningsskiljaktigheter mellan kommissionen och rådet har lösts, så förordningen borde träda i kraft till årsslutet.
Jag hoppas att den ändrade förordningen kommer att genomföras på lämpligt sätt i alla EU:s medlemsstater.
(CS) Mina damer och herrar! Efter 16 år har vi i dag äntligen gett grönt ljus åt en förenkling, ett enande och samtidigt åt hårdare restriktioner när det gäller utfärdande och återkallelse av operativa licenser.
Jag hoppas att förordningen inte leder till att små sportflygarklubbar går i konkurs.
Jag röstade för förordningen. Jag tror uppriktigt sagt att den verkligen kommer att göra det möjligt att återkalla operativa licenser från företag som lurar kunderna genom att enbart ange priser utan skatter, avgifter eller bränsletillägg och därmed inte anger det totala priset för flygbiljetten.
Jag hoppas att kontrollorganet även kommer att fokusera på prisdiskriminering på grund av bostadsort.
Jag anser att den ändrade förordningen kommer att medföra ökad säkerhet för tillhandahållandet av lufttrafik, särskilt genom att man förenar de villkor som styr leasingen av flygplan med besättning från såväl EU som tredjeländer.
(HU) Tack så mycket herr talman! Som den socialdemokratiska gruppens ansvarige för denna fråga har jag ställt mig bakom Miroslav Ouzkýs kompromissförslag.
Jag ser det som en framgång för parlamentet och även för den socialdemokratiska gruppen att rådet även har accepterat att vi borde begränsa de två glykollösningsmedlen mer, för att på så sätt skydda våra medborgares hälsa.
Ämnet 2-(2-metoxietoxi)etanol är hälsofarligt när det tas upp via huden.
Det är väl känt att det begränsar reproduktionsförmågan och det är alltså en stor framgång att vi har förbjudit användandet av detta, inte bara i färger utan även i rengöringsmedel och golvvårdsprodukter.
Från början ville kommissionen endast förbjuda 2-(2-metoxietoxi)etanol i färger, men tack vare samarbetet med alla parter har vi även lyckats begränsa det i rengöringsmedel.
Det är skadligt för människors hälsa att andas in 2-(2-metoxietoxi)etanol.
Enligt kommissionens rapport skulle det bara ha förbjudits i sprutlackeringsfärger, men det har, återigen efter rekommendationer från den socialdemokratiska gruppen, även begränsats i rengöringsmedel med aerosol.
Eftersom vi inte hade någon debatt i kammaren ville jag bara nämna det viktigaste innehållet i kompromissförslaget.
(MT) Det är viktigt att Europaparlamentet känner till prissituationen för vatten och elektricitet i mitt land och närmare bestämt effekterna av dagens beslut när det gäller detta.
Det är därför jag avger en röstförklaring.
Ända sedan regeringen höjde oljepriset har den ökat konsumenternas kostnader genom att lägga på tilläggsavgifter.
Denna månad meddelade den att tilläggsavgifterna kommer att öka till 96 procent.
Detta kommer att medföra en ny fattigdom, en energifattigdom.
Regeringen kommer varken med kortsiktiga eller långsiktiga lösningar.
Trots att vi i vårt land har gott om sol och vind saknas det politik för alternativa energikällor, till och med när det gäller renare energikällor som gas, och regeringen har fortfarande inte ens börjat överväga detta.
Det var därför som jag röstade så här och det är därför som det vi har gjort i dag är viktigt, för att inte säga historiskt.
(CS) Herr talman, mina damer och herrar! Jag vill förklara varför jag röstade som jag gjorde om förslaget till Europaparlamentets och rådets direktiv om ändring av direktiv 2003/55/EG om gemensamma regler för den inre marknaden för naturgas.
Direktivets huvudsakliga del gäller utan tvekan förslaget till åtskillnad av ägandet, som uttryckligen skulle förhindra vertikalt integrerade företag från att ha både ett leverans- och ett överföringsintresse när det gäller gas.
Jag röstade för det ändrade kompromissförslaget därför att jag är övertygad om att man måste ta hänsyn till oron hos de länder som var emot en åtskillnad av ägandet.
Jag håller med kommissionen om att den europeiska marknaden för naturgas saknar investeringar i infrastruktur för energiöverföring och en bra samordning mellan enskilda systemansvariga för överföringssystemen.
Jag anser dock att vi måste ta hänsyn till naturgas- och elmarknadernas strukturella olikheter och därför göra en åtskillnad mellan dem.
Liberaliseringen av gasmarknaden måste ske gradvis och symmetriskt.
Fokus måste särskilt ligga på harmoniseringen av graden av öppenhet på de nationella marknaderna.
Jag lade ner min röst i den slutliga omröstningen och röstade mot förslaget till det så kallade ”tredje paketet” gällande åtskillnaden mellan leverantörer och nätföretag på gasmarknaden, eftersom vi har missat ett gyllene tillfälle att bekräfta principen om fri konkurrens på gasmarknaden. Vi borde ha följt med i det som har hänt på elmarknaden.
I det här tredje paketet ger man i stället praktiskt taget garantier för monopol och tidigare monopol i Europa. Våra nationella marknader kommer därför även i fortsättningen att vara ojämförbara, vilket gör att utsikterna för en verklig europeisk energimarknad blir ännu sämre.
Än värre är att detta tvetydiga tredje paket i praktiken innebär att de tidigare monopolen kommer att få ännu mer uppmuntran och hjälp att ingå avtal liknande dem med den ryska gasjätten Gazprom.
(DE) Herr talman! Som alla i kammaren vet har vi haft en EU-förordning om samordningen av de sociala trygghetssystemen sedan 2004, men tyvärr har vi inte haft någon tillämpningsförordning.
Med Europaparlamentets beslut får vi äntligen även tillämpningsbestämmelser, vilket innebär att vi har ett instrument som vi kan använda för att främja rörligheten i Europeiska unionen utan att man förlorar den sociala tryggheten.
Upprättandet av förbindelseorgan gör att vi även kan ge praktisk hjälp åt dem som arbetar utanför sitt hemland, till exempel genom att svara på frågor om var och hur de ska ansöka om pension.
Vi i Europaparlamentet har med andra ord sett till att människor kan få riktig hjälp i frågor som rör välfärden.
(NL) Jag avstod från att rösta om Bozkurtbetänkandet, även om jag i princip inte har något emot en begränsad form av samordning av EU-medlemsstaternas olika sociala trygghetssystem, i synnerhet inte om det fungerar till fördel för EU-medborgare som bor i en annan medlemsstat än sin egen.
Jag vill dock återigen varna för en harmonisering eller, ännu sämre, enhetlighet mellan de olika medlemsländernas sociala trygghetssystem.
Som flamländare har jag så att säga förmånen att se att ett enhetligt socialt trygghetssystem för enbart två befolkningsgrupper i Belgien, flamländare och valloner, är helt ogenomförbart och leder till ett oerhört omfattande missbruk.
Låt för guds skull varje medlemsstat organisera och finansiera sitt eget sociala trygghetssystem, annars kommer vi på ett eller annat sätt att få ett system som missbrukas och som är sämre, dyrare och mindre effektivt och som i slutändan leder till mindre i stället för mer solidaritet bland människorna i Europa.
(DE) Herr talman! Jag vill också förklara att jag röstade för det här betänkandet därför att det innehåller ett förslag till ny förordning i stället för den gamla och därmed en garanti för att våra sociala trygghetssystem nu kan samordnas mer effektivt, eftersom man har förenklat och ändrat de tillämpliga bestämmelserna.
Med Lambertbetänkandet blir det också möjligt för oss att uppnå våra mål för att bidra ytterligare till större rörlighet i EU och ge människor möjligheten att ta med sig sina sociala förmåner när de får anställning i ett annat medlemsland.
Detta bidrar till social trygghet i Europeiska unionen.
(NL) Tack, herr talman!
Då är vi i dag vid steg två av Richard Corbetts försök att uppfostra parlamentet ännu mer till de politiskt korrekta eurokraternas knähund.
I går beslutades det att vi parlamentsledamöter knappt får lägga fram parlamentsfrågor och att parlamentets talman kommer att bedriva självcensur.
I dag blir det svårare att bilda grupper, och föredraganden medger uttryckligen, och i viss mån ärligt, att denna åtgärd främst är riktad mot den EU-skeptiska högern i parlamentet.
Så det hela slutar där man började.
EU-skepsisen här i kammaren, i synnerhet hos den politiska högern, måste tystas ned.
Det EU-skeptiska resultatet av folkomröstningar i Irland, Nederländerna och Frankrike nonchaleras som vanligt som om de inte fanns.
Detta är en europeisk version av ”Mugabedemokrati”. Vilken demokrati!
Föredraganden Richard Corbett uttryckte faktiskt sina åsikter - på ett förolämpande sätt kan tilläggas - utanför utskottet för konstitutionella frågor angående den politiska familj som jag tillhör här parlamentet. Detta väcker naturligtvis stort tvivel när det gäller hans opartiskhet.
Betänkandet är mycket tvivelaktigt och innehållet försvagades drastiskt i utskottet. Det enda som fanns kvar var bestämmelserna för att säkra överlevnaden för politiskt korrekta grupper vars totala antal ledamöter skulle hamna under det minimiantal som krävs, och ett ändringsförslag har smugits in särskilt för att hindra vår politiska familj från att bilda en grupp.
De skäl som uppges stämmer inte alls överens med fakta. Det räcker att titta i bilagan till betänkandet så ser man att det inte finns något nationellt parlament där det minsta antalet ledamöter som krävs för att bilda en grupp är högre än 20.
Det råkar faktiskt vara så att antalet ofta är mycket lägre, till exempel 15, 10 eller 8, och i vissa fall räcker det med en person för att bilda en politisk grupp.
Corbettbetänkandet är därför ett angrepp mot demokratin och helt enkelt mot de grundläggande reglerna för rent spel.
. - (NL) Corbettbetänkandet syftar bara till en sak, bara en sak, nämligen att tysta ned de högerorienterade nationella rösterna i Europaparlamentet.
Richard Corbetts gruppordförande sticker inte under stol med detta.
När ITS-gruppen bildades i januari 2007 sa han helt öppet att förordningen skulle ändras särskilt i syfte att stoppa bildandet av högerorienterade grupper i framtiden.
Andra grupper kommer säkerligen att bli indirekt lidande till följd av detta, men Richard Corbett kommer inte att ligga sömnlös för det.
Hans förslag är förmodligen riktat mot en EU-skeptisk grupp.
Det är uppenbart att socialdemokraterna i parlamentet avskyr att grupper av alla politiska färger ska ha samma medel och politiska rättigheter.
Detta Mugabeliknande sätt att tänka utgör en väsentlig del av bristen på demokrati i Europa, på samma sätt som man på ett orubbligt sätt ignorerar de franska, nederländska och irländska väljarnas demokratiska röster.
Herr talman! Vi kommer att göra detta till en valfråga nästa år i Flandern, var så säker!
(EN) Herr talman! Det faktum att vi över huvud taget röstade om detta i dag tycker jag är ett brott mott parlamentets arbetsordning.
Utskottet röstade ned betänkandet därför att, som jag tror, utskottets ordförande hade missbedömt dem som var i rummet, varför han helt enkelt bara rev upp arbetsordningen och fortsatte med en ändrad version av det.
Varför har vi sträckt oss så långt?
Vad är det som är så viktigt att vi måste riva upp vår arbetsordning på detta sätt?
Ja, skälet är naturligtvis som vi vet - och föredraganden har varit tydlig med detta - att hindra EU-skeptiker från att bilda en grupp.
Men varför är ni så rädda?
Vad är det som gör er så nervösa?
Vi är bara 50, kanske högst 60 personer, av 785 parlamentsledamöter.
Kan det bero på att de personer ni egentligen bekymrar er över är era egna väljare och att ni överför och riktar det förakt och den rädsla ni känner för EU:s väljare, som röstar nej så fort de får chansen, mot oss och att ni tar ut det ni inte vågar säga om de människor som skickar tillbaka er hit på oss, som är deras synliga talesmän här i parlamentet.
Om jag har fel kan ni bevisa det genom att genomföra den folkomröstning ni en gång lovade.
Pactio Olisipiensis censenda est!
(PL) Herr talman! Jag röstade mot Corbettbetänkandet eftersom jag anser att det är ett uttryck för extrem diskriminering i Europaparlamentet, som påstår sig vara demokratiskt och som ändå försöker använda administrativa metoder för att göra det omöjligt att bilda politiska grupper som inte tänker eller agerar på det sätt som majoriteten anser vara politiskt korrekt.
Detta är en dubbel diskriminering eftersom man använder administrativa metoder för att hindra bildandet av grupper och därför att man samtidigt ger betydande ekonomiskt stöd i tillägg till organiserade politiska grupper, vilket innebär ytterligare fördelar för dessa.
Denna diskriminering strider mot Europeiska unionens grundvalar och de grunder som EU ska byggas på.
Jag protesterar högljutt mot detta och ni ska inte inbilla er att ni, även om ni lyckas driva igenom detta, kommer att kunna få igenom det i nationerna i Europa, som definitivt kommer att protestera.
. - (EN) Herr talman! Det är sällan jag hör sådant struntprat som jag precis hörde från Vlaams Blok, Front national och Dan Hannan.
Det här betänkandet förbjuder inte någon, och regeländringen skulle inte heller innebära att någon förlorade sin rösträtt eller sin rätt att tala och sin rätt att agera som ledamot av Europaparlamentet.
Det regeländringen handlar om är vilken tröskelnivå vi ska fastställa för det minsta antalet ledamöter som krävs för att bilda en grupp och därmed tilldelas extra skattepengar och extra resurser för att bedriva sin politiska verksamhet.
Alla nationella parlament med gruppsystem fastställer tröskelnivåer.
Vi har haft en väldigt låg tröskel - lägre än nästan alla nationella parlament procentuellt räknat.
Det är helt rätt att vi stannar upp och undersöker det.
Jag noterar att nästan alla grupper stödde kompromissförslaget i slutändan, såväl stora som små grupper.
Jag noterar att även talaren för gruppen Självständighet/Demokrati - den EU-skeptiska IND/DEM-gruppen - föreslog en alternativ nivå på 3 procent, det vill säga 22 ledamöter.
Så de inser själva att vi måste höja det nuvarande antalet, som för närvarande är för lågt.
Ärligt talat, är skillnaden mellan deras nivå på 22 och den nivå på 25 som har antagits verkligen ett angrepp mot demokratin?
Äh, försök inte!
(PL) Herr talman! Buzekbetänkandet innehåller en detaljerad utvärdering av alla strategiska åtgärder inom området energiteknik.
Tyvärr innebar bristen på finansiering till all den forskning som behövdes, i kombination med den plötsliga prisökningen på gas och olja, att vi blev tvungna att inrikta vår forskning på metoder för att minska användningen av dessa källor i energiförsörjningssyfte.
Denna prioritering kommer också att innebära minskade koldioxidutsläpp och borde inkluderas i strategin.
Jag tycker det är viktigt att främja forskning om uppbyggnaden av säkra, moderna kärnkraftverk och uppbyggnaden av de nyaste kraftverken som bygger på produktion av helium och vätgas, liksom om tredje generationens biobränslen som kan produceras lokalt så att man minskar överdrivna bränslekostnader.
Vid omröstningen röstade jag för de ändringsförslag där man tog upp dessa prioriteringar.
(PL) Mina damer och herrar! Vi har antagit det viktiga betänkande som professor Jerzy Buzek har utarbetat.
Europeiska unionens växande beroende av energiimport, som 2030 kommer att nå en nivå på 65 procent, har tvingat oss att vidta åtgärder för att garantera försörjningstrygghet när det gäller råvaror som används för kraftproduktion mot bakgrund av solidaritetsprincipen.
Det borde även skapas ytterligare instrument för att minska de risker för de enskilda medlemsstaternas energiförsörjningstrygghet som en fortsatt liberalisering av energisektorn medför.
För att nå EU:s mål för förnybara energikällor och minskade växthusgaser måste vi främja utvecklingen av nya tekniker, särskilt tekniker för avskiljning och lagring av koldioxid.
Det är viktigt att stödja ren kolteknik och att intensifiera vårt arbete när det gäller andra och tredje generationens biobränslen samt att utöka forskningen om kärnkraft.
Det har också blivit mycket viktigare att arbeta för förbättringar när det gäller energieffektivitet och energisparande.
Skriftliga förklaringar
skriftlig. - (IT) Herr talman! Jag röstar för denna resolution.
Jag är utvecklingsutskottets föredragande om Erasmus Mundus-programmet och mitt betänkande antogs nyligen enhälligt.
Jag hoppas att vi kommer att kunna godkänna den slutliga texten vid sammanträdesperioden i september, så att det nya programmet kan inledas i januari 2009.
Syftet är att sprida fördelarna med vårt utmärkta universitetssystem utanför unionens gränser och göra det möjligt för utländska studenter att komma och studera vid våra fakulteter - och att ge studenter från EU möjlighet att, genom stöd, samla på sig erfarenhet i ett land utanför EU.
Jag anser att Erasmus är ett centralt instrument för hållbar utveckling, eftersom syftet med det, vilket jag betonar i mitt betänkande, är att bidra till att studenterna kommer tillbaka till sina hemländer och därmed, med hjälp av de idéer, kunskaper och internationella kontakter de har samlat på sig, bidrar till sitt hemlands ekonomiska tillväxt.
En betydande andel av finansieringen när det gäller åtgärd 2 tas från de anslag som öronmärkts för utveckling.
Jag anser att vi måste se till att de ekonomiska anslagen för de årliga handlingsprogrammen för Brasilien och Argentina 2008, som är speciellt öronmärkta för främjandet av ekonomisk utveckling och välfärd, faktiskt används till både utbildning och konkreta åtgärder på området och att de bidrar till infrastruktur och produktionsmetoder anpassade till en hållbar utveckling.
skriftlig. - (PT) Eftersom det är omöjligt att ta upp alla viktiga punkter i det här betänkandet skulle jag vilja betona att Europaparlamentet, efter det irländska folkets bestämda NEJ till Lissabonfördraget, fortsätter att låtsas och agera som om ingenting hade hänt.
Men det har tvärtom hänt väldigt mycket, vilket man ser av det skamlösa syftet med det här betänkandet.
Majoriteten i Europaparlamentet anser bland annat att
varje lands ställning, det vill säga deras utrikespolitik, borde kopplas samman med en bindande politisk plattform som EU har upprättat,
EU borde överväga en omorganisering och utökning av sina kontor inom FN med anledning av ”de ökade befogenheter och ansvarsuppgifter som EU:s företrädare kommer att förväntas utöva med tanke på ratificeringen av Lissabonfördraget”,
rådet så snart som möjligt borde ”fastställa den operativa status som EU:s ”observatörer” ska ha i FN”,
medlemsstaterna borde enas om ”en mer samstämd ståndpunkt om reformeringen av FN:s säkerhetsråd - en ståndpunkt som, samtidigt som det slutliga målet med ett permanent mandat för Europeiska unionen inom ett reformerat FN kvarstår, under tiden syftar till att öka unionens inflytande”.
En målmedveten och tydlig federalism i stormakternas ledband, med Tyskland i täten ...
skriftlig. - (EN) Ledamöterna från Labour Party i Europaparlamentet välkomnar detta betänkande, i synnerhet den starka uppmaningen till EU:s medlemsstater om att fokusera och stärka sina åtaganden gentemot millennieutvecklingsmålen.
Vi håller helt med om att tyngdpunkten måste ligga på att uppfylla de avlagda löftena och trappa upp det befintliga arbetet.
Ledamöterna från Labour Party instämmer dock inte i rekommendationen om ett enda mandat i FN:s säkerhetsråd och kan inte stödja denna.
Vi anser inte att det skulle vara bra för Europas proportionerliga representation.
Enligt artikel 19 lägger inte EU-medlemmar i FN:s säkerhetsråd uttryckligen fram EU:s ståndpunkter i rådet.
Det står dessutom i FN:s stadga att så inte kan ske.
Men det pågår en sund informell samordningsprocess, såväl i New York som på ett större plan, och det är detta som bör uppmuntras.
skriftlig. - (IT) Gruppen De gröna/Europeiska fria alliansen har alltid ansett att Europeiska unionen borde ha ett permanent mandat i FN:s säkerhetsråd, vilket läggs fram i Lambsdorffbetänkandet.
Vår grupp godtar dock inte ”prioriteringen” av initiativet med en ”övergripande process”, som innebär att antalet permanenta nationella medlemmar skulle öka, och som vi anser bara måste ses som ett av flera möjliga alternativ.
skriftlig. - (EN) Jag gläds över Alexander Graf Lambsdorffs betänkande där man lägger fram EU:s prioriteringar för FN:s generalförsamlings 63:e session.
Jag stöder särskilt det som sägs om behovet av att fortsätta arbeta för ett målmedvetet engagemang för millennieutvecklingsmålen vid toppmötet.
EU:s agenda för millennieutvecklingsmålen borde utgöra ett globalt exempel och vi borde arbeta för att resten av världssamfundet följer detta exempel vid FN:s generalförsamling i september.
Jag röstade för betänkandet.
skriftlig. - (EN) I dag antogs Alexander Graf Lambsdorffs förslag till Europaparlamentets rekommendation till rådet om EU:s prioriteringar för FN:s generalförsamlings 63:e session utan omröstning i kammaren.
Detta förfaringssätt - som är möjligt genom ”artikel 90” - är inte bara väldigt tvivelaktigt. Det ger dessutom det falska intrycket av att hela Europaparlamentet håller med om innehållet i betänkandet, vilket verkligen inte är fallet.
Vi är starkt emot rekommendationen att Lissabonfördragets nuvarande ställning skulle nödvändiggöra en omorganisering och utökning av rådets ”kontor i New York och Genève med anledning av de ökade befogenheter och ansvarsuppgifter som EU:s företrädare kommer att förväntas utöva med tanke på ratificeringen av Lissabonfördraget”.
Detta är inte bara ett hån mot de irländska väljarna, som förkastade Lissabonfördraget med bred majoritet vid folkomröstningen. Det är dessutom ett försök att tolka Lissabonfördraget som att EU görs till en juridisk person och därmed till en överordnad stat.
skriftlig. - (IT) Lambsdorffbetänkandet (och den tillhörande rekommendationen) ger en klar politisk signal om att stärka Europeiska unionens profil inom FN.
Genom kommissionen och medlemsstaterna bidrar ju unionen totalt med över 40 procent av FN:s ekonomiska medel, men den har hittills inte fått något utbyte i form av politiskt inflytande eller förmåga att påverka.
En del av texten är emellertid vilseledande och till skada för den diskussion som har påbörjats i New York om reformen av FN:s säkerhetsråd.
Samtidigt som man betonar det grundläggande målet med ett permanent mandat för EU som sådant tar man i rekommendationen bland de olika förhandlingsinitiativen enbart upp den så kallade övergripande processen.
Denna drivs av de länder som endast stöder ett av de olika förslag som lagts fram, det vill säga förslaget om en utökning av antalet permanenta nationella medlemmar.
Detta förslag, som har fått stöd från mindre än en tredjedel av medlemmarna, verkade redan från början vara splittrande och obalanserat, vilket ordföranden för FN:s generalförsamling själv har påpekat.
Vi vill betona att vi varmt välkomnar den politiska uppmärksamhet som Europaparlamentet ägnar åt ett generellt stärkande av Europeiska unionens profil i FN, men vi anser samtidigt att våra reservationer och invändningar när det gäller rekommendationen om den ”övergripande processen” bör föras till protokollet.
skriftlig. - (IT) Herr talman! Jag vill säga något positivt om Lambsdorffbetänkandet, i vilket man återigen betonar Europaparlamentets engagemang för att stärka EU:s ställning i FN.
Jag vill dock understryka att man i betänkandet, när det gäller frågan om reformen av FN:s säkerhetsråd, lägger fram en värdering som inverkar negativt på de diskussioner som fortfarande pågår i New York.
Bland de olika reformalternativ som lagts fram tar man särskilt upp den ”övergripande processen” (punkt Q), som är ett förslag som innebär att man vill öka antalet permanenta medlemmar i FN:s säkerhetsråd.
Detta förslag har hittills fått stöd av mindre än en tredjedel av medlemmarna i FN:s generalförsamling.
Jag ber er därför att anteckna i protokollet att jag reserverar mig mot denna del av rekommendationen.
skriftlig. - (PT) Det är oroväckande att frågan om reformen av FN kommer på tal så ofta.
Behovet av en reform har varit känt under några år, men det har även det faktum att det är omöjligt att genomföra en sådan reform.
Detta dödläge är viktigt av två skäl.
För det första förvärrar det de faktorer som bidrar till organisationens misslyckanden, vilka är ganska många.
För det andra främjar det uppkomsten av en diskussion som stöds och rättfärdigas av behovet av alternativ.
Att stärka samarbetet mellan demokratier är helt klart en fin tanke att främja, även om det inte medför en omfattande anslutning till projektet demokratiernas förbund.
Men det vore även klokt att vara realistisk.
Det är därför som FN måste anpassa sig till maktens verklighet, inte så mycket på grund av rimligheten utan snarare på grund av genomförbarheten.
När det gäller Europeiska unionens roll måste vi inse att inget av de länder som har ett mandat i FN:s säkerhetsråd eller som kan få ett mandat där går med på att ersättas av ett enda EU-mandat.
Avslutningsvis har vi sett att FN:s nya råd för mänskliga rättigheter långt ifrån har övervunnit sin föregångares brister.
skriftlig. - (ES) Herr talman!
Med anledning av rekommendationen till FN:s generalförsamlings 63:e session i september i New York, fastställs det i artikel 90.4 i arbetsordningen att en rekommendation inom ramen för den gemensamma säkerhets- och utrikespolitiken, som gått till omröstning i ett utskott, ska anses antagen och föras upp på föredragningslistan för ett plenarsammanträde utan att parlamentet behöver godkänna texten och utan någon debatt eller något ändringsförfarande.
Därför, då vi är nöjda med praktiskt taget hela dokumentet med undantag för en punkt, skulle min grupp vilja uttrycka sin åsikt om denna punkt som gäller rätten till sexuell och reproduktiv hälsa.
Det konceptet, som är något tvetydigt, ger upphov till frågor som till stor del rör det individuella samvetet och moralen, och vi anser INTE att dessa bör utgöra ämnet för några av parlamentets uttalanden, i synnerhet inte med anledning av FN:s nya session.
Vår grupp begärde särskild omröstning i utskottet för utrikesfrågor och röstade emot på grund av ovannämnda skäl.
skriftlig. - (PL) Herr talman! Alexander Graf Lambsdorffs betänkande och rekommendation är politiskt sett mycket viktiga, eftersom syftet är att främja en förstärkning av EU inom FN.
Det kan vara bra att veta att även om kommissionen och medlemsstaterna står för mer än 40 procent av FN:s budget, är EU:s inflytande fortfarande mycket svagare än det borde vara.
Betänkandet innehåller dock ett missvisande stycke om de diskussioner som just nu förs i New York om reformen av säkerhetsrådet.
Samtidigt som det långsiktiga målet om ett permanent mandat för EU bekräftas, citerar man i rekommendationen endast ett av de förslag som lagts fram, nämligen den s.k. övergripande processen, trots att det finns många fler förslag.
Det är allmänt känt att detta förslag har visat sig vara högst splittrande och har godkänts av mindre än en tredjedel av FN:s medlemmar, vilket generalförsamlingens ordförande påpekat.
Samtidigt som vi vill uttrycka stor uppskattning för det huvudsakliga innehållet och strukturen hos denna rekommendation från Europaparlamentet, anser jag det därför nödvändigt att betona våra uttryckliga reservationer och protester mot det stycke där den ”övergripande processen” nämns.
skriftlig. - (IT) Herr talman! Lambsdorffbetänkandet ger en klar politisk signal om att stärka Europeiska unionens profil inom FN.
Genom kommissionen och medlemsstaterna bidrar ju unionen totalt med över 40 procent av FN:s ekonomiska medel, men den har hittills inte fått något utbyte i form av politiskt inflytande eller förmåga att påverka.
En del av texten är vilseledande och till skada för den diskussion som har påbörjats i New York om reformen av FN:s säkerhetsråd.
Samtidigt som man betonar det grundläggande målet med ett permanent mandat för EU som sådant tar man i rekommendationen bland de olika förhandlingsinitiativen enbart upp den så kallade övergripande processen, vilken stöds av länder som endast vill ha ett av de olika förslag som lagts fram, det vill säga förslaget om en ökning av antalet permanenta nationella medlemmar.
Detta förslag, som har fått stöd från mindre än en tredjedel av medlemmarna, verkade redan från början vara splittrande och obalanserat, vilket ordföranden för FN:s generalförsamling själv har påpekat.
Jag vill betona att jag varmt välkomnar den politiska uppmärksamhet som Europaparlamentet ägnar åt ett generellt stärkande av Europeiska unionens profil i FN, men jag anser samtidigt att min reservation och min invändning när det gäller rekommendationen om den ”övergripande processen” bör föras till protokollet.
skriftlig. - (PL) Herr talman! Det gläder mig att Europaparlamentet i dag har tänkt över frågan om EU-prioriteringar inför det kommande FN-mötet.
I föredragandens förslag nämns att FN vill se ”inrättandet av nya organ, en radikal översyn av andra organ, en omstrukturerad ledning för FN:s fältinsatser, en omorganisering av FN:s tillhandahållande av bistånd och en djupgående reform av dess sekretariat”.
Detta är oerhört viktigt.
Vi får dock inte glömma att all denna verksamhet bedrivs för människans skull och för de mänskliga rättigheter som människans värdighet medför.
Påven Johannes Paulus II talade om detta för ett par år sedan vid ett FN-möte, och sa att det första systematiska hotet mot de mänskliga rättigheterna har att göra med fördelningen av materiella tillgångar, som ofta är orättvis, att den andra sortens hot hade att göra med olika slags själsliga orättvisor, och att det är möjligt att skada en människas syn på sanningen, hennes medvetande och uppfattning av det vi kallar medborgerliga rättigheter, som alla har rätt till oavsett bakgrund, ras, kön, nationalitet, religion eller politiska åsikter.
Jag anser att hans ord bör vara vägledande i FN:s arbete.
skriftlig. - (PT) Herr talman! Det aktuella förslaget utgör en del av ett paket (tillsammans med förslagen till direktiv om driftskompatibilitet och inrättandet av en europeisk järnvägsbyrå) som syftar till att ”underlätta rörligheten för lokomotiv i gemenskapen”, som en del av liberaliseringen av järnvägstransporten inom EU.
Före alla andra överväganden, måste vi därför betona att huvudmålet för detta direktiv är att undanröja alla hinder för liberaliseringen av järnvägstransporten genom att harmonisera lagstiftningen om järnvägssäkerhet i medlemsländerna.
Det står klart att de mest avancerade normerna för järnvägssäkerhet i varje land måste antas och tillämpas.
Vi måste dock komma ihåg att liberaliseringen och privatiseringen av järnvägen ifrågasattes i vissa länder, till exempel i Storbritannien, efter en försämring av tjänster och andra allvarliga händelser som ledde till att man på nytt måste tänka igenom angreppet mot denna allmänna tjänst.
Jag betonar att harmonisering av lagstiftningen om järnvägssäkerhet på gemenskapsnivå aldrig får leda till att de mest avancerade lagarna på detta område hotas, och länderna får inte heller förbjudas att ha sådan lagstiftning.
skriftlig. - (EN) Herr talman! Jag röstade för Paolo Costas betänkande ”Säkerhet på gemenskapens järnvägar”.
Föredragandens rekommendation kommer att bidra till att rationalisera lagstiftningen och förenkla fri rörlighet för tåg i hela EU.
Med dessa rekommendationer kommer byråkratin att minskas och de bör ge utvecklingen av järnvägstransporten i EU ett uppsving.
skriftlig. - (PT) Herr talman! Det är helt och hållet nödvändigt att harmonisera de nationella säkerhetsförfarandena i medlemsstaterna.
Denna fråga är ännu ett exempel på hur viktigt det är att insistera på investeringar i järnvägstransport.
Om vi vill ha en hållbar utveckling av Europas transportsystem och om vi ska nå de mål och respektera de löften vi gett till medborgarna och på internationell nivå under de senaste åren, måste vi investera i järnvägen och garantera det europeiska järnvägssystemets driftskompatibilitet.
Förenklingsåtgärder och införandet av principen om ömsesidigt erkännande är de viktigaste punkterna i detta betänkande.
En annan väldigt viktig punkt är tillämpningen av strängare utbildnings- och certifieringsåtgärder för alla berörda och ansvariga aktörer på gemenskapens järnvägsmarknad, från järnvägsföretag till infrastrukturförvaltare.
Jag anser att detta betänkande är ännu ett positivt steg i vårt sökande efter multimodalitet som grund för den gemensamma transportpolitiken.
skriftlig. - (EN) Herr talman! Jag röstade för att de järnvägar som är kulturarv inte skulle omfattas av detta direktiv.
Detta speglar min uppskattning för dessa tågföretags speciella karaktär.
Om dessa företag hade tvingats att följa villkoren i direktivet, skulle det ha inneburit en mängd förödande kostnader för organisationer som till stor del finns kvar på grund av frivilliga och medlemmar.
Järnvägar såsom Romney, Hythe och Dymchurch Railway samt Kent och East Sussex Light Railway (där jag själv är medlem på livstid) är delar av den historiska turistindustrin i sydöstra England och i hela EU.
Det är skamligt att somliga här, som säger sig vara ”nationalistiska”, inte kunde stödja detta undantag.
skriftlig. - (PL) Herr talman! Skapandet av en gemensam järnvägsmarknad för transporttjänster kräver att vi förändrar de nuvarande reglerna.
Medlemsstaterna har utvecklat sin egen säkerhetsstandard, i första hand för inrikessträckor, baserade på nationella tekniska och operativa koncept.
Det börjar bli oerhört viktigt att skapa harmoniserade rättsliga strukturer i medlemsstaterna, gemensamma texter för säkerhetsregler, enhetliga säkerhetscertifikat för järnvägsföretag samt enhetligt ansvar och befogenheter för säkerhetsmyndigheter och för förfaranden vid utredning av järnvägsolyckor.
Varje medlemsstat bör ha ett oberoende organ för reglering och övervakning av järnvägssäkerheten.
För att säkra ett gott samarbete mellan dessa organ på EU nivå bör man fastställa minimiregler för arbetsuppgifter och skyldigheter som ska gälla för alla organ.
Skyddet av den allmänna säkerheten och ordningen, vilket omfattar uppehållande av ordningen vid allmänna järnvägskommunikationer, borde vara en av de grundläggande uppgifter som EU ansvarar för.
skriftlig. - (PT) Herr talman! Det aktuella förslaget är en del av ett åtgärdspaket (tillsammans med förslagen till direktiv om driftskompatibilitet och säkerhet) för att liberalisera järnvägstransporten inom EU, där ”byrån” tar på sig rollen som ”regleringsmyndighet”.
Denna politik kommer att leda till en gradvis försämring av järnvägstransporten som allmän tjänst, och de mer lönsamma sträckorna kommer att ges till privata företag genom privatisering (offentlig-privata samarbeten) på skattebetalarnas bekostnad och utan att ta hänsyn till de enskilda ländernas och befolkningarnas intressen och behov.
I Portugal har det visat sig att genomförandet av denna politik har lett till en försämring av de allmänna tjänsterna, begränsad rörlighet och ökade färdkostnader.
Det har resulterat i avstängning av hundratals kilometer järnvägssträcka, stängning av stationer, minskat passagerarantal och försämring av servicekvaliteten, minskat antal anställda inom järnvägssektorn samt en attack mot deras löne- och arbetsrättigheter.
Järnvägssektorn är strategisk för den socioekonomiska utvecklingen.
Vi behöver en politik som främjar utvecklingen och förbättringen av de offentliga järnvägstransportsystemen i våra länder.
skriftlig. - (DE) Herr talman!
Jag röstade för Paolo Costas betänkande om ändring av förordning (EG) nr 881/2004 om inrättande av en europeisk järnvägsbyrå.
Förbättrandet av den tekniska och lagstiftningsmässiga ramen för gemenskapens järnvägar som en del av det tredje järnvägspaketet är en viktig och välkommen utveckling som omfattar åtgärder för att förstärka den europeiska järnvägsbyrån.
Som centralt organ måste byrån garantera att en enhetlig strategi eftersträvas i hela EU.
Synnerligen viktig är den fortsatta utvecklingen av ERTMS-systemet (European Railway Traffic Management System). Dess driftskompatibilitet och kompatibilitet måste till varje pris garanteras.
Inrättandet av ett EG-kontrollförfarande är ett passande sätt att nå detta mål, men dess effektivitet kommer att vara beroende av en stabil och effektiv europeisk järnvägsbyrå.
Av denna anledning stöder jag en ytterligare utveckling av byrån såsom föredraganden föreslår.
skriftlig. - (EN) Herr talman! I Costabetänkandet om inrättande av en europeisk järnvägsbyrå stöder man uppenbarligen behovet av att införa ERTMS-systemet, vilket innebär högteknologisk järnvägssäkerhet.
Jag stöder detta initiativ som tillsammans med betänkandet om säkerhet på gemenskapens järnvägar kommer att ge utrymme för ett mer sammanhängande europeiskt järnvägssystem.
Jag röstade för betänkandet.
skriftlig. - (FR) Herr talman! Frågan om järnvägens driftskompatibilitet är oerhört viktig för de europeiska järnvägarnas utveckling och framgång.
Jag är därför väldigt glad att vi har kunnat nå en kompromiss om förbättringen av gemenskapens lagstiftning på det här området.
Trots att jag röstade för de förslag som föredraganden Paolo Costa lagt fram, är jag icke desto mindre medveten om kompromissens begränsningar.
Tio år för att få alla slags förflyttningar av rullande materiel godkända är en ansenlig tidsperiod.
När det gäller den europeiska järnvägsbyråns roll kunde den ha varit mer omfattande, i synnerhet gällande utvecklandet och införandet av ERTMS-systemet (European Rail Traffic Management System).
Medlemsstaterna beslutade annorlunda av rädsla att nyinrättade järnvägsbyråer och andra nationella organ skulle ses som föråldrade.
Vi står dock där vi står just nu på grund av att man 2004 inte vågade göra en ordentlig europeisk insats för järnvägen.
Det är så som den europeiska integrationen går vidare: sporadiskt och med små steg.
Men om vi agerar på detta försiktiga sätt kommer vi säkerligen att missa vissa chanser, och därför hoppas jag att medlemsstaterna kommer att agera genom att strängt tillämpa sina egna förslag.
skriftlig. - (PT) Herr talman! För att understryka vår kritik mot betänkandets huvudsakliga mål, avreglering av luftfarten som allmän tjänst inom EU, vill vi påminna er om vad vi påpekade för ett år sedan.
Här försöker man att
dölja det faktum att avregleringen har haft negativa konsekvenser för anställnings- och arbetsvillkoren, och man bör undersöka hur detta har påverkat säkerheten och underhållet vid större luftfartsföretag,
undvika att värna om full respekt för arbetstagarnas rättigheter, samt att låta bli att nämna att
a) kabinpersonalens anställningsavtal och arbetsvillkor kommer att regleras av det lands lagstiftning, kollektivavtal och närstående avtal i vilket arbetstagarna vanligtvis utför sitt arbete eller i vilket de påbörjar och återvänder till efter arbetet, även om de för en kort tid arbetar i ett annat land,
b) för arbetstagare vid ”gemenskapens” lufttransporter som tillhandahåller tjänster från en verksamhetsbas som befinner sig utanför medlemsstatens territorium gäller den sociala lagstiftning och de kollektivavtal som gäller i landet där operatören har sitt huvudkontor,
c) slippa ifrån kravet att representanter för arbetstagarnas organisationer garanterat kommer att delta i alla beslut som fattas inom lufttransportsektorn.
skriftlig. - (PL) Herr talman! I och med den förordning som har antagits av Europaparlamentet förändras den lagstiftning som styr tillhandahållandet av lufttrafik i EU, till förmån för både lufttrafikföretag och passagerare.
Förordningen är viktig för att den inre marknaden ska fungera ordentligt.
Den bidrar till att skapa en mer konkurrensinriktad miljö för de europeiska lufttrafiksföretagens verksamhet, vilket stärker dem gentemot internationella konkurrenter.
Genom förordningen kommer samma villkor att gälla för utfärdandet och återkallandet av operativa licenser, vilket bör undanröja den snedvridna konkurrens som just nu dominerar marknaden och som bl.a. beror på olika regler när det gäller villkor för operativa licenser, diskriminering av vissa EU-lufttrafikföretag på grund av deras nationalitet eller diskriminering när det gäller flygrutter till tredjeländer.
Den som vinner mest på förändringarna som presenterats kommer dock att vara konsumenten.
Att det blir obligatoriskt att inkludera skatt och pristillägg i biljettpriset kommer att ge en mer öppen prissättning och understödja principen om att pristillägg ska vara valfria.
Det kommer också att förhindra att konsumenter tvingas betala högre avgifter och gör det möjligt för konsumenterna att fatta välgrundade beslut.
Genom att eliminera flygbolag som är finansiellt osunda utsätts passagerarna dessutom inte för risken att deras lufttrafikföretag går i konkurs.
skriftlig. - (DE) Herr talman! Jag röstade för Arūnas Degutis betänkande om gemensamma regler för tillhandahållande av lufttrafik i gemenskapen.
Åtgärder som vidtas för att förstärka och förbättra de befintliga bestämmelserna bör uppmuntras, speciellt i fråga om öppen prissättning på flygresor.
Passagerarna har rätt till en detaljerad beskrivning av priset på deras flygbiljetter.
Detta nya instrument kommer att bidra till att prissättningen blir mer öppen och mer begriplig.
På så sätt vill EU bekämpa vilseledande reklam och skapa en marknad baserad på kvalitet och inte på de till synes attraktiva erbjudanden som man ofta kan hitta på Internet.
Åtgärderna för att garantera att skyddsnormerna efterlevs är ännu en förbättring som det nya instrumentet medför, och detta ger de anställda ett bättre skydd och mer enhetliga arbetsvillkor.
De gemensamma reglerna kommer att skydda konsumenternas och de anställdas rättigheter och garantera att gemenskapens lufttrafikföretag är öppna och inte döljer någon information.
skriftlig. - (PL) Herr talman! Jag röstar för föredragandens åsikt om antagandet av rådets gemensamma ståndpunkt utan några ändringar.
Jag anser även att vi med denna förordning kommer att förstärka och förbättra de befintliga lagbestämmelserna om övervakning av operativa licenser, leasing av luftfartyg, lufttrafikfördelning och öppen prissättning.
skriftlig. - (EN) Herr talman! I och med Arūnas Degutis betänkande om reglerna för tillhandahållandet av lufttrafik i gemenskapen kommer det att garanteras att det flygpris man ser är det pris man faktiskt kommer att betala.
Slutliga priser för flygresor måste nu inkludera flygpris, skatter, flygplatsavgifter och övriga tilläggskostnader.
Detta är ett steg framåt mot större öppenhet i luftfartssektorn och när det gäller konsumentskyddet.
Arbetstagarna i luftfartssektorn kommer också att få ett mer heltäckande socialt skydd i och med betänkandets förslag.
Jag röstade därför för rekommendationerna i betänkandet.
skriftlig. - (EN) Herr talman! Jag stöder helt och fullt detta betänkande som kommer att leda till att vi kan sätta stopp för vissa flygbolags oärliga taktik, där man anger flygpriser som inte inkluderar skatter, avgifter och ett stort antal andra tilläggskostnader.
I dagsläget är det möjligt för flygbolagen att ange vilseledande priser som helt enkelt visar sig vara felaktiga.
Resultatet av detta är en allvarlig brist på öppen prissättning när det gäller flygresor, vilket leder till att konkurrensen snedvrids och påverkar konsumentens förmåga att fatta välgrundade beslut.
Ofta får människor till slut betala mycket mer än vad de hade räknat med eftersom det angivna priset inte ens är i närheten av den slutliga kostnaden.
Kommissionen och parlamentet har arbetat tillsammans för att garantera denna förändring.
Detta betänkande kommer att medföra att flygpriset måste anges enkelt och tydligt samt inkludera alla skatter och tilläggskostnader.
EU:s nerslag på den här taktiken är goda nyheter för konsumenterna.
skriftlig. - (PL) Herr talman! Statistik används inom många områden, inte bara av företag eller institutioner på det ekonomiska området.
Den fyller en viktig funktion när det gäller att planera och följa marknadsutvecklingen.
Av denna anledning är det viktigt att de målindikatorer som används för att samla in statistiken är pålitliga och speglar verkligheten och marknadsförändringarna på ett korrekt sätt.
Befintliga målindikatorer bör ses över, men man bör även överväga nya områden för datainsamling.
Behovet av att modernisera vår statistik beror även på att det finns så många olika system och statistiska metoder i medlemsstaterna, vilket ofta gör det svårt att jämföra data inom EU.
Förändringarna på detta område får naturligtvis inte öka den administrativa bördan för företag, särskilt inte för de små och medelstora företagen.
Den avancerade metod som används i Meets-programmet bör bidra till både rationalisering och samordning av metoder för datainsamling från olika källor, och dessutom, vilket är mycket viktigt, medför den att företagen inte behöver vidarebefordra samma data till olika institutioner som är involverade i datainsamling.
Jag anser att Meets-programmet är ett steg i rätt riktning för att minska den administrativa bördan för företagen, vilket kommer att bidra till att nå det mål som kommissionen satt upp, att minska bördan med 25 procent till 2012.
skriftlig. - (EN) Herr talman! Jag stöder Christoph Konrads betänkande om programmet för modernisering av den europeiska företags- och handelsstatistiken.
Syftet med betänkandet är att tillhandahålla investeringar för att effektivisera statistikframställningen så att nya efterfrågningar kan mötas samtidigt som bördorna för företagen minskas.
Jag röstade för betänkandet.
skriftlig. - (PL) Herr talman!
Jag är för detta betänkande. Batterier och ackumulatorer som inte uppfyller kraven i direktiv 2006/66/EG bör dras in och inte få säljas.
Kommissionen har beslutat att batterier som uppfyller nuvarande krav och som har släppts ut på EU:s marknad före den 26 september 2008 inte ska dras in.
Detta anser jag vara en rimlig lösning.
Indragningen av batterier som inte uppfyller kraven kommer att leda till mer avfall.
Jag anser att det enklaste och bästa sättet att hantera denna situation är att märka dessa batterier och ackumulatorer för att ange att de inte uppfyller EU-kraven.
skriftlig. - (EN) Herr talman! I och med Miroslav Ouzkýs betänkande kommer användandet av de två ämnena 2-(2-metoxietoxi)etanol och 2-(2-butoxietoxi)etanol till stor del att begränsas och i vissa fall förbjudas i produkter som släpps ut på marknaden för försäljning till allmänheten.
Konsumentskyddet betonas särskilt i betänkandets rekommendationer och jag röstade för det.
skriftlig. - (PL) Herr talman! Giftiga ämnen som går att hitta i rengörings-, skölj- och desinficeringsprodukter, samt i färg och lösningsmedel, kan utgöra en risk för människors hälsa genom att irritera luftvägarna och orsaka allergier.
Att begränsa marknadstillträdet för produkter som inte uppfyller säkerhetskraven kan bidra betydligt till skyddet av vår hälsa och vår miljö.
Majoriteten av dessa produkter kan vara skadliga när de används och orsaka olika obehagliga symptom.
De kan även vara skadliga för miljön när de kommer in i ekosystemet.
När de förorenar mark eller vattenresurser är de ofta svårt att förutsäga vad följderna kommer att bli.
Att begränsa nivåerna av dessa ämnen i olika sorters tvättmedel och rengöringsprodukter är ett positivt steg och därför anser jag att EU bör anstränga engagera sig för att få bort dessa ohälsosamma ämnen från våra liv och från miljön.
skriftlig. - (PT) Herr talman! Vi röstade mot detta betänkande eftersom det utgör en del av avregleringspaketet för gasmarknaden och man uttryckligen stöder åtgärderna för att fullborda den inre marknaden så fort som möjligt, men generellt sett inte godkänner de instrument och bestämmelser som kommissionen har föreslagit.
Intressant kritik riktas mot förslagen till konsekvensbedömningar, att subsidiaritetsprincipen delvis inte beaktas och att det inte görs någon konsekvent uppdelning av behörigheten mellan EU-organen.
Vad man vill i betänkandet är dock att underlätta tillträdet till naturgasöverföringsnäten för företag, d.v.s. att underlätta privatiseringen av det som finns kvar av den offentliga sektorn och ställa den till förfogande för ekonomiska gruppers strategier, ekonomiska grupper som vill ta sig in på marknaden.
skriftlig. - (EN) Herr talman! Atanas Paparizovs betänkande om villkor för tillträde till naturgasöverföringsnäten kommer att bidra till att underlätta integreringen av EU:s inre gasmarknad.
I betänkandet behandlas gränsöverskridande frågor mellan medlemsstaterna och man vill öka tillsynen på EU-nivå.
Det är viktigt att EU arbetar för en inre gasmarknad och jag röstade för betänkandet.
skriftlig. - (PT) Detta betänkande förtjänar en röst från mig och från alla mina kolleger som ansåg att konsekvensen i det tredje energipaketet var beroende av en effektiv lagstiftning om handel med naturgas och inte bara en lagstiftning som ser bra ut på ytan.
Jag välkomnar viljan att skapa villkor för att öka investeringar i gasöverföringssystem.
Detta kan i sig leda till en potentiell ökad konkurrenskraft och konkurrens inom sektorn.
Jag välkomnar insatserna för en effektiv avreglering av nationella gasmarknader och tillträde till överföringssystemet, vilket ökar öppenheten.
Slutligen välkomnar jag den goda viljan i betänkandet att hörsamma EU-medborgarnas önskan om en öppnare och mindre monopoliserad energimarknad.
Det tredje energipaketet behöver vårt godkännande av detta betänkande, och det gör även EU-medborgarna.
skriftlig. - (EN) Herr talman! Min ståndpunkt avspeglar min åsikt om vikten av naturgas och att den finns tillgänglig för konsumenterna till lägsta möjliga pris.
En gasledning kommer att koppla samman Libyen och Sicilien.
Ledningarna kommer att dras i närheten av Malta, så att för att mitt land ska kunna dra fördel av detta måste det antingen ansluta sig till gasledningen eller, vilket har föreslagits, så måste en gasledning anläggas mellan Sicilien och Malta.
Mitt land har inte någon stor marknad och dess konsumtion varierar mellan 16 och 18 miljoner enheter per år.
Om användandet av naturgas skulle bli mer utbrett skulle detta säkerligen medföra en förändring av energipolitiken i både Malta och Gozo.
Detta är möjligt om gasen används i själva energiproduktionen.
Jag påpekade detta för den dåvarande nationalistiska regeringen och underströk vikten av att ha gasstationer för ungefär 15 år sedan.
Regeringen visade inget intresse och installerade till sist endast en liten gasstation.
Eftersom avstånden på Malta är små är det möjligt att använda gas som bränsle till privata och kommersiella fordon.
Omvandlingen av fordonens motorer utgör inget problem.
Naturgas är dessutom mycket billigare och renare än bensin eller diesel.
Regeringen och det statliga bolaget har dock inte tänkt över den infrastruktur som behövs i anknytning till distributionen av gasen.
Herr talman! Förslaget till ett direktiv om den inre gasmarknaden är en del av ”det tredje energipaketet” som fullbordar privatiseringen av tillhandahållet av naturgas.
Förslaget till ett direktiv och betänkandet syftar tillsammans till att eliminera den höga nivån av centralisering som fortfarande finns i vissa länder och att fullborda EU-monopolens intrång på marknaden. På så sätt snabbar man på genomförandet av avregleringen samtidigt som man inför sanktioner mot de medlemsstater som ännu inte har genomfört den helt och hållet.
Paketet har två nyckelpunkter: åtskillnad när det gäller ägandet mellan gasleveransverksamhet och gastransport och lagringsverksamhet, så att kapitalet effektivt kan dra nytta av denna offentliga infrastruktur för produktion, lagring och transport av gas som finns kvar i medlemsstaterna.
Bemyndigandet av till synes oberoende tillsynsorgan som syftar till att göra det omöjligt för medlemsstaterna att göra nationella förändringar eller statliga ingripanden, garanterar total immunitet för de företagsgrupper som är intresserade av gassektorn.
Denna EU-politik kommer att ge samma dåliga resultat för de anställda som privatiseringen av andra energisektorer: höjda priser och försämrad kvalitet på tjänsterna.
Kampen mot monopolintressena för att avskaffa denna politik är det enda sättet att tillgodose de behov som arbetarklassfamiljerna för närvarande har.
skriftlig. - (PT) Herr talman! Denna åtgärd visar tydligt på vår gemensamma vilja att nå målet att avreglera energimarknaden.
Jag röstar därför ja.
Jag anser att åtskillnad när det gäller ägandet av produkttillgångar och överföringsnät för naturgas är nödvändig för att nå detta mål, men det är inte nödvändigtvis det enda som behövs.
Därav viljan att skapa de villkor som är nödvändiga för att uppmuntra transnationella investeringar i nätinfrastrukturer.
Därav kravet på likabehandling för tredjeländer som planerar att investera i den europeiska energimarknaden.
Därav viljan att förbättra samordningen mellan nationella tillsynsorgan för energisektorn.
Med denna åtgärd kommer marknaden att bli konkurrenskraftig och den är därför viktig för konsumenterna som kommer att dra fördel av de nya reglerna på en sundare, friare och öppnare energimarknad.
skriftlig. - Jag röstar för detta betänkande, eftersom det kommer att underlätta för medborgare som flyttar och reser mellan medlemsländerna utan att makt förflyttas till EU.
skriftlig. - (RO) Herr talman! Jag röstade för Jean Lamberts betänkande eftersom det är lösningen på ett av medborgarnas problem.
Vi lever i en globaliserad värld där tusentals människor arbetar i ett annat land än sitt hemland, och vi behöver samordna de sociala trygghetssystemen för alla personer som utnyttjar sin rätt att arbeta i andra medlemsstater. Syftet är att garantera och främja rörligheten, som är en grundläggande rättighet inom EU.
Vi kan röra oss fritt inom EU, men det bör finnas större sociala rättigheter som inte upphör att gälla vid de nationella gränserna.
Med förhoppningen om att de europeiska medborgarna kommer att kunna dra fördel av likabehandling och icke-diskriminering när det gäller social trygghet, stöder jag initiativet för att underlätta arbetstagarnas fria rörlighet. Vi måste undanröja alla hinder för rörligheten.
skriftlig. - Jag röstar emot detta betänkande, eftersom det innehåller förslag till detaljerad reglering på EU-nivå av bl.a. utbetalning av svensk föräldrapenning, vilket kommer att försvåra för individuella bedömningar och ger EU för mycket makt.
skriftlig. - (PL) Herr talman! Syftet med detta dokument är att göra EU-reglerna om samordning av de sociala trygghetssystemen i de individuella medlemsstaterna bättre och mer effektiva.
Bestämmelserna i betänkandet kommer definitivt att förenkla livet för den genomsnittlige EU-medborgaren som kan röra sig fritt i hela EU.
Oavsett om man är anställd, tjänsteman inom administrationen, student, pensionär eller företagare kommer man att behålla sin rätt till sociala trygghetsförmåner efter att ha flyttat till ett annat land.
Jag stöder definitivt avlägsnandet av ännu ett hinder för människors fria rörlighet inom EU, och detta dokument är ett viktigt steg i denna process.
skriftlig. - (FR) Herr talman! Jag har två kommentarer till Jean Lamberts betänkande och ändringarna av den berörda förordningen.
1.
Trots att föredraganden förnekar detta förutsätts det i förslaget till förordning att tredjelandsmedborgare åtnjuter fri rörlighet, etableringsfrihet och fritt tillträde till arbetsmarknaden i hela EU.
Vi måste dock komma ihåg att ingen av dessa punkter har förverkligats ännu, tack och lov.
Vad man gör är att skala bort ännu en liten bit av medlemsstaternas befogenheter vad det gäller invandringspolitik, eller med andra ord deras suveräna rätt att välja vilka utlänningar som har tillåtelse att vistas på deras territorium och att kontrollera inträde, vistelse samt omfattningen av dessa utlänningars rättigheter.
2.
Det är viktigt att ge EU-medborgarna möjlighet att kunna dra fördel av en samordning av de sociala trygghetssystemen och att garantera att det sociala skydd som de har rätt att förvänta sig (beroende på deras arbete och berättigade förmåner) inte påverkas negativt av den ”internationella” rörlighet som de uppmuntras att delta i.
Att inom detta område göra allt för att garantera likabehandling av EU-medborgare och tredjelandsmedborgare, utan någon som helst tanke på att garantera någon motsvarande behandling, ökar bara invandringen, vilket våra enorma, icke-diskriminerande och alltför generösa sociala trygghetssystem redan gör.
skriftlig. - (DE) Herr talman! Människors tillit till EU beror till stor del på deras förtroende för EU:s sociala stabilitet, och det är ett av de områden som har förändrats mest under de senaste åren och årtiondena.
I praktiken har deltidsarbete och nya anställningsvillkor (”McJobs”) lett till att europeiska anställda i slutändan ofta inte tjänar särskilt mycket mer än vissa arbetslösa gör.
Baksidan av okontrollerad ekonomisk tillväxt och konstanta välfärdsbesparingar är en ökning av fattigdomen och den sociala utslagningen.
I EU, ett av de rikaste områdena i världen, levde år 2005 16 procent av befolkningen under fattigdomsgränsen.
Resultatet av de höjda olje- och livsmedelspriserna är att ännu fler människor nu har hamnat under fattigdomsgränsen eller lever på gränsen till fattigdom.
EU måste arbeta för att bekämpa fattigdom bland sina egna invånare och se detta som en brådskande angelägenhet, och välfärdssystemen måste finnas tillgängliga för EU-medborgarna i första hand.
skriftlig. - (FR) Herr talman! I dag röstade jag för betänkandet av Richard Corbett om ändringen av artikel 29 i Europaparlamentets arbetsordning om bildande av politiska grupper, dvs. kravet på att ledamöterna i en politisk grupp ska representera minst en fjärdedel av medlemsstaterna (i stället för det nuvarande kravet på en femtedel) och att det lägsta antalet ledamöter ska vara 25 (i stället för 20), och detta gjorde jag av flera anledningar.
För det första för att jag anser att denna reform är absolut nödvändig för att vår institution ska kunna fungera effektivt och för att förhindra att den blir ännu mer uppdelad, med regler som förblir oförändrade trots successiva utvidgningar och utökningen av vår församling sedan 2004.
Dessutom verkar den lösning som föreslagits av min kollega från den socialdemokratiska gruppen, vars outtröttliga ansträngningar lett till en kompromiss om de politiska gruppernas majoritet, väldigt rimlig jämfört med praxis på nationell nivå inom EU.
Med tanke på resurserna, både mänskliga och finansiella, som gjorts tillgängliga av parlamentet för de politiska grupperna, verkar tydlig representativitet vara nog för att rättfärdiga denna förändring.
Slutligen är syftet helt enkelt att främja en viss konsekvens bland de politiska krafterna på europeisk nivå. Allt detta kan bara göra vår demokrati starkare.
skriftlig. - (PL) Detta dokument utgör ännu ett försök av majoriteten att ta kontroll på bekostnad av minoriteten.
Arrogansen hos de största politiska grupperna i Europaparlamentet har nått nya höjder.
Målet med dokumentet är att höja minimiantalet ledamöter för att bilda en politisk grupp, från 21 till 30.
Små grupper som exempelvis gruppen Självständighet/Demokrati blir allvarligt hotade av sådana villkor.
Självfallet röstade jag nej till det här dokumentet.
skriftlig. - (EN) ALDE-gruppen röstade emot en ändring av artikel 29 av följande skäl:
Dagens sju grupper orsakar inga verkliga effektivitetsproblem.
Minoritetsuppfattningar har lika stor rätt att vara organiserade som majoritetsuppfattningar.
Europaparlamentet bör spegla den mångfald av politiska uppfattningar som finns i unionen på ett korrekt sätt: vi behöver inte exakt kopiera de nationella parlamenten, vars arbete det är att tillsätta en regering.
Att lägga ned mindre grupper tvingar antingen parlamentsledamöterna att motvilligt ansluta sig till större grupper, vilket minskar deras sammanhållning, eller att bli grupplösa, vilket ökar ineffektiviteten.
Parlamentets storlek ska ändå minskas från 785 till 751 (Lissabon) eller 736 ledamöter (Nice).
skriftlig. - (PT) Vi röstar mot detta betänkande och det åtagande som görs eftersom vi försvarar pluralism, demokrati och respekt för åsiktsskillnader.
Betänkandets ändrade bestämmelser om bildande av politiska grupper är oacceptabla, och fler hinder införs för att bilda politiska grupper i Europaparlamentet efter nästa val.
Hittills har det krävts minst 20 ledamöter från sex medlemsstater för att bilda en politisk grupp.
Enligt det förslag som nu har godkänts krävs det 25 ledamöter från sju medlemsstater för att bilda en politisk grupp.
Detta innebär att det kommer att bli svårare att bilda små politiska grupper i Europaparlamentet, vilket är ännu ett hinder för att hävda åsikter som skiljer sig från den dominerande ideologin i detta alltmer nyliberala, militaristiska och federalistiska EU.
En sista kommentar om de metoder som har använts av majoritetsgrupperna, PPE-DE-gruppen och PSE-gruppen.
De började med att lägga fram ett förslag om att det skulle krävas 30 ledamöter för att bilda en politisk grupp.
Sedan utpressade de några av de mindre grupperna för att vinna deras stöd för ett så kallat kompromissförslag, det som just har antagits.
Vi parlamentsledamöter från det portugisiska kommunistpartiet har ända från början konsekvent vidhållit att vi är mot införandet av fler hinder för att bilda politiska grupper.
skriftlig. - (ES) Jag lade ned min röst för det här betänkandet eftersom jag anser att även om praktiska regler för bildandet av parlamentsgrupper helt klart behövs, så är antalet föreslagna ledamöter och medlemsstater för högt.
Om parlamentet vill försvara pluralism och mångfald är det bättre att de berörda bildar en politisk grupp, hellre än att utvidga den grupplösa delen, som blir alltmer olikartad och ineffektiv.
skriftlig. - (FI) De större grupperna föreslog ursprungligen att 30 ledamöter från sju medlemsstater skulle krävas för att bilda en politisk grupp.
Lyckligtvis röstades planen ned av en knapp majoritet i utskottet för konstitutionella frågor i maj, då omröstningen slutade 15 mot 14.
Jag har också röstat emot de föreslagna ändringarna nu, eftersom de små grupperna ofta bara kommer att stå som åskådare när besluten fattas.
Det är fel att inskränka mångfalden av åsikter eller att försvåra de mindre gruppernas verksamhet jämfört med tidigare.
Det är också märkligt med tanke på att de största åsiktsskillnaderna ofta återfinns inom grupperna.
Den största gruppen, de konservativa, har splittrats i två eller till och med tre grupper i många viktiga frågor.
skriftlig. - (EN) De konservativa parlamentsledamöterna har röstat emot Richard Corbetts båda föreslagna ändringar för att höja ribban för bildandet av politiska grupper i Europaparlamentet.
Balansen mellan parlamentets effektiva verksamhet och behovet av att ta hänsyn till mångfalden av röster och åsikter inom parlamentet måste vägas med omsorg.
Detta uppnås bäst genom att behålla dagens tröskelvärden för bildandet av politiska grupper.
Även om vi erkänner att det finns skäl för att höja minimiantalet ledamöter för att bilda en grupp, så leder varje höjning av minimiantalet medlemsstater till att mindre grupper och delegationer missgynnas på ett orättvist och onödigt sätt.
Efter att ha studerat Richard Corbetts betänkande rekommenderade följaktligen utskottet för konstitutionella frågor att inte göra några ändringar av de tröskelvärden som fastställs i artikel 29.
De konservativa ledamöterna röstade emellertid ja till den ändring som ursprungligen lades fram av Timothy Kirkhope, och som har antagits av utskottet för konstitutionella frågor.
Med denna ändring införs ett mer praktiskt och förnuftigt tillvägagångssätt i fall där en politisk grupp hamnar under de nödvändiga tröskelvärdena.
skriftlig. - (EN) Jag stöder Richard Corbetts betänkande om att ändra arbetsordningen vad gäller bildandet av politiska grupper.
Med 27 medlemsstater behöver EU:s regler i den här frågan aktualiseras.
Europaparlamentet kan inte rättfärdiga att man använder miljontals euro av skattebetalarnas medel för att finansiera politiska grupper, särskilt fascister, som endast sätts samman för ekonomisk vinning.
Europaparlamentet har det lägsta tröskelvärdet för bildande av grupper av nästan alla parlament.
Det föreligger inget hot mot någon existerande grupp - inte heller är ändringen av arbetsordningen ett försök att krossa euroskeptikerna, som är fler än minimiantalet.
Således röstade jag för Richard Corbetts betänkande.
skriftlig. - (NL) De bägge största grupperna föredrar helt klart ett tvåpartisystem.
Det främsta kännetecknet på ett sådant system är att de båda partierna delar ett gemensamt intresse, nämligen att det andra, tredje och fjärde partiet inte får in en fot i det politiska beslutsfattandet och därmed förblir fullkomligt irrelevanta i väljarnas ögon.
Endast de största grupperna räknas. Protester och alternativ måste skjutas åt sidan.
Om undantagsvis några andra fortfarande lyckas ta sig in i parlamentet får de normalt de sämsta platserna, i egenskap av personer med begränsade rättigheter.
Vissa ledamöter i parlamentet hör inte till någon grupp.
Detta är vanligtvis en följd av påtryckningar från andra.
Sådana påtryckningar tvingar andra ledamöter att gå med i en grupp som har åsikter som de inte instämmer till fullo i.
På grund av egenintresse accepterar grupper ledamöter även då de vet att dessa ledamöters åsikter skiljer sig markant från partilinjen.
Skälet är att man inte kan bilda en grupp här om man inte har 20 likasinnade ledamöter eller fler.
Om alla åsiktsriktningar i samhället ska representeras demokratiskt är det bättre att slopa minimiantalet, i stället för att höja det till 25 eller 30 och införa stränga regler mot oliktänkande.
Jag är helt och hållet emot det.
skriftlig. - (DE) Enligt min mening finns det inget rimligt skäl till att höja minimiantalet ledamöter som krävs för bildandet av en politisk grupp.
Vid en närmare granskning håller inte föredragandens argument, särskilt inte hans påstående om högre tröskelvärden för bildande av politiska grupper i medlemsstaternas parlament.
Om en rättvis jämförelse ska kunna göras med Europaparlamentet bör man endast ta hänsyn till den direktvalda kammaren.
Den andra kammaren består i allmänhet av delegater från förbundsstater eller regioner, och av det skälet är de inte jämförbara.
Det genomsnittliga värde som används av direktvalda nationella parlament för bildandet av politiska grupper är praktiskt taget likadant som det tröskelvärde som används av Europaparlamentet.
Hur som helst är steget att höja gränsvärdet för bildandet av politiska grupper tydligt motiverat av ett annat hänsynstagande.
I utskottet hänvisade exempelvis föredraganden till bildandet av gruppen Identitet, tradition och självständighet (ITS) som en olycklig omständighet, och underströk behovet av att förhindra sådant i framtiden.
På grund av detta angrepp på demokratin och yttrandefriheten och på parlamentsledamöternas jämlikhet, som fastställs i fördraget och i Europaparlamentets arbetsordning, röstade jag självfallet nej till detta betänkande.
Betänkandet, i dess antagna form, kompletterar Europaparlamentets oacceptabla arbetsordning, som syftar till att kontrollera och undertrycka möjligheterna för dem som inte helt samtycker till EU.
Detta är ett nytt odemokratiskt och auktoritärt beslut, som ytterligare hindrar bildandet av politiska grupper.
Det politiska målet är uppenbart: de vill utesluta radikala krafter, i synnerhet kommunistiska, för att tysta alla motröster och alla yttrandeformer som utmanar EU och dess politik.
Detta odemokratiska förfarande åtföljdes tydligen av politisk utpressning från koalitionen gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater tillsammans med socialdemokratiska gruppen i Europaparlamentet, för att även tvinga andra att acceptera höjningen, eftersom de hotade med att rösta för ett förslag om en ännu större höjning av minimiantalet ledamöter, till 30, om motståndarna inte gav vika.
Omröstningen visar att den här matchen var uppgjord på förhand av krafterna bakom den europeiska enkelriktningen, som ett alibi för deras odemokratiska beslut.
Ledamöterna för Nea Dimokratia och Panellinio Socialistiko Kinima (PASOK) och ledamoten för Synaspismos har röstat ja till denna förkastliga ändring och beslutet i dess helhet, vilket bevisar att i nyckelfrågorna håller krafterna bakom den europeiska enkelriktningen samma kurs.
Vi, ledamöterna för Greklands kommunistparti, har röstat mot höjningen av antalet ledamöter till 25 och mot betänkandet i dess helhet, och därigenom fördömer vi odemokratiska intriger och politiskt spel.
skriftlig. - (PT) Att införa överdrivna begränsningar och skapa hinder för bildandet av politiska grupper kan aldrig vara bra för något parlament.
Förutom att det kan betraktas som en kränkning av de grundläggande rättigheterna blir följden av sådana åtgärder ofta det rakt motsatta mot vad förespråkarna hade i åtanke.
Detta är därför en dålig förändring.
Europaparlamentet måste göra sig gällande som en i grunden demokratisk referenspunkt, både i EU och i världen.
Detta kan inte uppnås om inte parlamentet visar en föredömlig inställning.
Jag håller inte med om att detta är den rätta riktningen.
Dessutom behöver EU mer än någonsin ständigt bevara förtroendet hos sina medborgare, alla medborgare, för sina institutioner.
Alla européer måste känna att de är representerade, oberoende av sina politiska ställningstaganden.
Därför är detta en dålig och oläglig reform, som jag röstar emot.
skriftlig. - Jag motsätter mig alla försök att minska demokrati och mångfald i åsikter i parlamentet genom att bland annat ändra antalet ledamöter och medlemsländer för att ha rätt att bilda politiska grupper.
Trots denna uppfattning, röstade jag för Corbettbetänkandets kompromissändringsförslag.
Skälet är pragmatiskt - det var det enda sättet att rösta för att inte riskera ett ur demokratisk synpunkt ännu sämre beslut som ytterligare skulle försvåra möjligheten att bilda en politisk grupp.
skriftlig. - (PL) I dag antog Europaparlamentet en ändring av arbetsordningen, som medför att riktlinjerna för bildandet av politiska grupper ändras.
Efter valet i juni 2009 måste de politiska grupperna i Europaparlamentet bestå av minst 25 ledamöter, som företräder minst sju medlemsstater.
Jag skulle vilja ge mitt fulla stöd åt denna höjning av tröskelvärdet för bildandet av politiska grupper i Europaparlamentet, eftersom detta kommer att bidra till att man undviker överdriven parlamentarisk splittring och göra parlamentets arbete mer effektivt.
Både sammanhållningen och effektiviteten i parlamentet har blivit lidande på grund av det överdrivna antalet små grupper i kammaren.
Små politiska grupper måste dock, för att stärka demokratin, skyddas mot tillfälliga minskningar i medlemsantal, om de hamnar under det nödvändiga tröskelvärdet.
skriftlig. - Vi röstade för betänkandet då ett bättre samarbete och mer öppenhet mellan nationella domstolar/domare och EG-domstolen är av yttersta vikt för ett fungerande europeiskt rättssystem.
Detta måste tydligt klargöras och sedermera verkställas genom förbättrad utbildning samt möjlighet till nätverkande och kunskapsutbyte.
Vi anser dock att diskussionen i punkterna 26 och 27 om EG-domstolens behörighet på vissa områden är en fördragsfråga som Europaparlamentet redan har yttrat sig om.
skriftlig. - (PT) Vi röstade emot det här betänkandet på grund av de påtryckningar som medlemsstaterna kommer att utsättas för, inklusive våra nationella domare, som utgör rättssystemets hörnsten i varje suverän stat.
I betänkandet tydliggörs syftet med den så kallade europeiska konstitutionen och det avsomnade Lissabonfördraget, som man försöker återuppliva på ett ytterst odemokratiskt sätt.
Betänkandet i sig bekräftar avsikten att införa en enhetlig europeisk rättsordning.
För att uppnå detta vill man ”i högre grad involvera de nationella domarna vid genomförandet av EG-rätten och ge dem ett större ansvar”.
Nationella domare spelar en väsentlig roll som garanter för rättssäkerheten, inklusive EG-rätten.
Men subsidiaritetsprincipen och konstitutionella frågor i varje enskild medlemsstat kan inte ifrågasättas med hänvisning till ”gemenskapsrättens företräde, direkt effekt, konsekvent tolkning och staternas ansvar för överträdelser av EG-rätten”, vilket åsyftas av kommissionen och en majoritet i Europaparlamentet.
Det är oacceptabelt att fortsätta med de här påtryckningarna, nu när fördraget har avslagits.
skriftlig. - (FR) Författaren till betänkandet är fullkomligt uppriktig.
Direkt i punkt 1 sätts målet upp: införandet av en enhetlig europeisk rättsordning.
I betänkandet, en sannskyldig stridsskrift för EG-rätten, försöker man verkligen i högre grad involvera de nationella domarna vid genomförandet av EG-rätten och ge dem ett större ansvar.
Följaktligen föreslås det att gemenskapslagstiftningen med tillhörande rättspraxis bör integreras i de nationella lagarna så snart som möjligt.
I betänkandet fortsätter man sedan med tanken att sammanföra de nationella rättsordningarna med EG-rätten, utan att överhuvudtaget ta upp frågan om överdrivna gemenskapsnormer, deras förvirrade ordalydelse och allmänna brist på konsekvens.
Detta steg mot en förenkling och kodifiering av gemenskapslagstiftningen är förvisso något positivt.
Detsamma gäller antagandet av förordningar för att se till att rättssäkerheten upprätthålls, jag tänker i synnerhet på dem som rör harmoniseringen av regelverket som styr lagkonflikter.
EG-domstolens rättspraxis visar sig emellertid ofta vara opålitlig för genomdrivandet av nationella lagar, vilka är underkastade domstolens bindande principer och dogmer även om de klart strider mot medlemsstaternas bästa rättstraditioner.
skriftlig. - (PT) ”Vänner, vänner, affärer åsido”...
Jag hänvisar till ytterligare en motsättning mellan EU och Förenta staterna, denna gång inom flygindustrin, där båda sidor, trots 1992 års avtal om statsstöd, försöker försvara sina intressen eftersom det är så kapitalistisk konkurrens fungerar.
Europaparlamentet klagar över att ”EU hela tiden har följt andan och bokstaven i 1992 års avtal och har regelbundet tillhandahållit styrkande handlingar” medan ”USA i stor utsträckning har åsidosatt sina förpliktelser”, ”ensidigt velat dra sig ur” avtalet och tog ”ett mål till Världshandelsorganisationen (WTO) mot EU med åberopande av europeisk återbetalningsskyldig finansiering som dock var helt förenlig med 1992 års avtal och som liknar den som Boeing åtnjuter”.
På samma gång försöker Europaparlamentet, som möts av ”bittra attacker” från Boeing och den amerikanska kongressen mot kontraktet som beviljats EADS tillsammans med Northrop Grumman Corporation för det amerikanska moderniseringsprogrammet för tankflygplan, gjuta olja på vågorna genom att framhålla behovet av ”att komma fram till en pragmatisk balans mellan EU:s civila stöd och USA:s militärindustriella system”.
Det verkar som om inte alla länder har rätt till suveränitet och ”frihandel”...
skriftlig. - (EN) Jag kommer att rösta ja till det här betänkandet, inte därför att jag finner nöje i WTO-tvister eller har paranoida föreställningar om Förenta staterna, utan därför att jag har fått nog av Förenta staternas protektionistiska politik under många år, särskilt inom civilflyget.
Amerikanerna har fulländat konsten att gnälla och klaga över andra länder och deras bristande frihandel, medan de själva har godkänt åtgärder som gör det möjligt för konkursmässiga flygbolag att fortsätta sin verksamhet, och har uppenbarligen slussat in miljontals dollar i understöd till Boeing.
Utskottet för internationell handel gör rätt i att stödja EU i dess process mot Förenta staterna i WTO.
Vad vi alla borde sträva efter i fråga om detta är en rättvis och öppen konkurrens mellan olika flygplanstillverkare, med frihet för flygbolagen att välja det bästa flygplanet som passar deras behov, till det bästa priset.
Det officiella valspråket för USA är ”Vi litar på Gud”.
Kanske det borde ändras till ”Gör inte som jag gör.
Gör som jag säger”.
skriftlig. - Vi svenska socialdemokrater har röstat för Buzeks betänkande om den europeiska strategiska planen för energiteknik.
Vi har ställt oss försiktigt positiva till avskiljning och lagring av koldioxid men ställer oss frågande till om det är nödvändigt att ge stöd till t.ex. gasifiering av kol för att vidareutveckla denna teknik.
Vi är även positiva till forskning och utveckling av nya energikällor med låga eller inga koldioxidutsläpp.
Vi stöder att unionen medfinansierar denna forskning, men anser inte att vi ska föregripa budgetarbetet genom att redan på förhand uppmana kommissionen att avsätta bestämda summor.
Vi har därför valt att lägga ned våra röster på dessa två punkter.
skriftlig. - (EN) Jag röstar nej till den andra delen av punkt 26, eftersom jag inte stöder tanken på att kärnkraften ska vara ett av de prioriterade initiativen.
Jag röstar ändå ja till betänkandet, eftersom dess mål är att snabba på utvecklingen av avancerad europeisk teknik för låga koldioxidutsläpp.
Det är centralt att EU har ett energiforskningsprogram för att stödja sin ambitiösa energipolitik och klimatförändringsmålen.
skriftlig. - (PL) Jag instämmer i Jerzy Buzeks åsikter om att vi behöver ny energiteknik för att bemöta de utmaningar EU står inför, dvs. miljöskyddet och behovet av att garantera en säker energiförsörjning och upprätthålla EU:s höga konkurrenskraft.
Jag håller även med föredraganden om att de resurser som anslås för ny energiteknik i EU:s nuvarande budgetram är otillräckliga.
Vi måste komma ihåg att det är genom offentlig-privata partnerskap som vi kan nå framgångar på området för ny energiteknik.
skriftlig. - (DE) Som vi vet av bitter erfarenhet har EU:s mål att snabbt öka den procentuella användningen av biobränslen haft ogynnsamma återverkningar.
Monokulturer, skövling av regnskogarna och konkurrens med säd för livsmedel och fodersäd, vilket har bidragit till dagens livsmedelskris, har uppenbarligen tvingat EU:s ministrar att tänka om och är ett slag mot deras mål att öka andelen förnybara energikällor i tillverkningen av motorbränslen till tio procent år 2020.
Vi bör välkomna att biobränslen inte längre kommer att tillverkas av säd för livsmedel och att det finns ett allmänt önskemål att invänta andra generationens biobränslen, såsom de som erhålls från avfallsprodukter, men detta får inte på något sätt leda till att EU:s insatser till förmån för förnybara energikällor mattas av.
Den oroande uppåtgående tendensen i oljepriserna gör det viktigare än någonsin att främja tillverkningen och användningen av energi från förnybara energikällor.
Alla de miljarder som spenderas på kärnkraft, med alla dess problem, måste i stället investeras i förnybara energikällor.
skriftlig. - (FR) De nationella placeringsfonderna, dessa statsägda fonder som investeras över hela världen, är de något bra eller dåligt?
Snarare något bra, om vi får tro resolutionen.
Det är dock sant att ett EU som stagnerar ekonomiskt på grund av sin egen ekonomiska politik och valutapolitik inte har råd att avfärda de tusentals miljarder euro i potentiella investeringar som de representerar.
Det är riktigt att de nationella placeringsfonderna för närvarande inte stör finansmarknaderna (de har till och med hjälpt det amerikanska banksystemet), och tenderar att vara inriktade på långsiktiga investeringar.
Detta kan dock förändras. Vi är alla medvetna om bristen på insyn i de flesta av dessa fonder när det gäller vidden av deras resurser, fördelningen av deras tillgångar, deras styrstrukturer och deras investeringsstrategier, som sträcker sig från etiska investeringar till att ägna sig åt investeringar med hög avkastning, skaffa sig maktpositioner och kanske potentialen att orsaka stor skada i framtiden.
De stater som innehar dessa fonder är inte alla vänligt sinnade mot EU, långt därifrån.
En av dem har redan gjort oss medvetna om hotet från dess ”finansiella kärnvapen”.
Vi lägger dock ned våra röster för denna text i stället för att rösta emot den. Skälet till detta är att kapitalets fria rörlighet i världen visserligen stöds i texten, men man efterlyser samtidigt en viss övervakning av och skydd mot dessa fonder.
skriftlig. - (EN) Resolutionen handlar om ett viktigt ämne.
Nationella investeringsfonder spelar en allt större roll för global handel och investering.
En del av detta är positivt, men så är inte alltid fallet, eftersom fondförvaltningar utan redovisningsskyldighet fattar beslut för att maximera kortsiktiga vinster på bekostnad av länder, samhällen och familjer.
Vi måste söka efter sätt att öka insynen i och ansvarigheten för dessa resurser, som ofta är större än de som är tillgängliga för nationalstaterna.
skriftlig. - (FI) Herr talman! Reinhard Racks betänkande om en ny kultur för rörlighet i städer, som vi har röstat ja till, är en viktig del av kommissionens nya övergripande tillvägagångssätt i dess energi- och klimatpaket: betydande utsläppsminskningar kan uppnås i Europa genom användning av en förnuftig och effektiv stads- och transportplanering.
Man måste dock ta hänsyn till att medlemsstaterna skiljer sig åt när det gäller geografiskt läge och levnadsförhållanden.
Just av det skälet röstade jag för de bägge ändringsförslagen från vår grupp.
Jag kommer från ett land med stora avstånd och jämförelsevis små städer.
Det står ganska klart att möjligheterna att minska privatbilismen är mycket mindre i exempelvis de glesbefolkade tätortssamhällena i Finland, i norr, än i de tätbefolkade områdena i Centraleuropa.
skriftlig. - (DE) Jag röstade för Reinhard Racks betänkande om en ny kultur för rörlighet i städer.
Förslaget till betänkande om grönboken är ett viktigt bidrag till frågan om stadsutveckling.
En tätorts eller stads ekonomiska utveckling och dess tillgänglighet är beroende av förbättrad rörlighet, men detta får inte uppnås på bekostnad av människors välbefinnande eller miljön.
Av det skälet borde man i betänkandet ta mer hänsyn till sociala faktorer och arbetsmarknadspolitik.
Vi måste också hålla i minnet att medlemsstaternas olikheter inte tillåter en enhetlig europeisk lösning, och att man därför bör fortsätta att strikt hålla sig till subsidiaritetsprincipen.
Jag är också av den åsikten att i de länder där en liberalisering redan har genomförts bör dess verkningar på sysselsättningen utvärderas.
Dessutom efterlyser jag ett certifieringssystem för anpassning av partikelfilter i bilar, transportfordon och terrängfordon i efterhand.
Medan man i grönboken pekar på de flesta problem som påverkar rörligheten i städer i dag, och även lägger fram ett par nya och innovativa idéer om hur man kan lösa dem, behandlas långt ifrån alla aspekter som skulle behöva tas upp och den kan därför endast betraktas som en utgångspunkt för diskussionen i denna fråga.
skriftlig. - (PL) Den viktigaste frågan som föredraganden tar upp handlar om att definiera de områden där EU bör delta när det gäller rörligheten i städer.
Föredraganden gör rätt i att framhålla att det finns liknande problem i hela EU vad gäller rörlighet i städer, men det är inte möjligt att utforma en enhetlig metod för att hantera dessa problem.
Föredragandens åsikter om att tätorten eller staden bör ha möjlighet att välja på vilket sätt den uppnår de fastställda målen är vettiga, och jag skulle vilja uttrycka mitt stöd för dessa åsikter.
skriftlig. - (NL) Tätorter och städer är tätbefolkade, med få öppna ytor och mycket trafik som färdas förhållandevis korta sträckor.
Genom att utrymmet är så värdefullt finns det helt enkelt ingen plats för tung fordonstrafik, och alltför höga buller- och luftföroreningar är ett ytterligare skäl till att vi måste försöka begränsa antalet bilar i städerna så mycket som möjligt.
Självfallet måste städerna vara tillgängliga för brandkåren, polisen, ambulanser, flyttbilar och fordon för personer med begränsad rörlighet, men de fåtaliga öppna ytorna bör i första hand reserveras för fotgängare, cyklister, spårvagnar, lekplatser och parker och trädgårdar.
Endast då blir staden beboelig.
I den text som vi röstar om i dag görs inte det tydliga ställningstagandet, utan man försöker bara sammanföra motsatta intressen och uppfattningar.
Lyckligtvis tillhör inte det här området EU:s behörighet.
Allt EU kan göra är att gynna bästa lösningar, goda erfarenheter som har vidareutvecklats och förbättrats.
Sådana förbättringar är viktiga inte bara för staden som har infört dem, utan även som ett föredöme för andra.
Bland föredömena återfinns Londons trängselskattsystem, det nya spårvägsnätet i Strasbourg och Bordeaux eller den sedan gammalt gällande begränsningen för trafik i centrum av Groningen.
Olyckligtvis bidrar EU knappast med någonting i och med det här betänkandet.
skriftlig. - (DE) Jag röstade emot det här betänkandet, eftersom EU inte är ansvarigt för dessa frågor.
Rättssäkerheten förbättras inte och man för inte EU närmare befolkningen när parlamentet producerar betänkanden i frågor som inte tillhör EU:s reglerande behörighet.
skriftlig. - Vi röstade för Olle Schmidts betänkande om ECB:s årsrapport.
Vi vill emellertid påpeka, med avseende på texten i betänkandets motiveringsdel där det talas om nödvändigheten av ett svenskt införande av euron, att vi respekterar det svenska folkomröstningsresultatet från 2003 då det beslutades att Sverige behåller kronan som valuta.
skriftlig. - (PT) Vi röstade emot det här betänkandet eftersom man återigen bekräftar stödet för Europeiska centralbankens arbete och inte anmärker på de gradvisa höjningarna av basräntan, trots att den redan har nått 4,25 procent, vilket är mycket högre än Federal Reserves basränta i Förenta staterna.
Vidare bortser man i betänkandet från att bankens åtgärder skadar arbetarna, befolkningen i allmänhet samt mikroföretag och små och medelstora företag.
Den tjänar endast de största ekonomiska gruppernas och finanskapitalets syften, trots att de orsakar problem för de bräckligare och mer beroende ekonomierna, såsom Portugals.
Till exempel i Portugal, där skuldnivån har nått 114 procent av BNP, utgör denna höjning, tillsammans med övervärderingen av euron, ytterligare en spik i kistan för mikroföretag och små och medelstora företag, förvärrar underskottet i handelsbalansen och förstärker landets beroendeställning.
Det kommer att bli svårare att hantera arbetslöshet, ökande användning av tillfällig arbetskraft, låga löner och den allmänna prishöjningen, med tanke på att skuldnivån för portugisiska familjer nu har nått 129 procent av deras disponibla inkomst.
Vi understryker därför åter behovet av att bryta med den här högerpolitiken och Europeiska centralbankens skenbara självstyre, vilket endast maskerar det faktum att den går i storkapitalets ledband.
skriftlig. - (FR) Olle Schmidts betänkande utgör parlamentets årliga klapp på axeln åt Europeiska centralbanken (ECB) för dess välvilja.
Som vanligt verkar man missa huvudproblemet: den fruktade minskningen av inkomstmarginalerna som krossar den europeiska befolkningens köpkraft och som ECB och EU delvis bär skulden för.
Ingen tror på att de officiella inflationssiffrorna (tre procent för 2008 enligt betänkandet), som bara är sammansatta index, speglar verklighetens stigande levnadskostnader för medborgarna, särskilt vad gäller basvaror, energi och boende.
Alla minns uttalandena av ECB, som varnade för löneökningarnas effekt på inflationen, som om lönerna för dessa EU-medborgare inte hela tiden pressas ned på grund av orättvis global konkurrens och den invandringspolitik som bedrivs av EU.
Vad gäller den kraftigt övervärderade eurokursen så är det sant att den besparar oss de värsta problemen i samband med de stigande oljepriserna.
Den hotar dock konkurrenskraften för många industrier, vilka i likhet med Airbus lockas att utlokalisera till dollarzonen.
Vi kan följaktligen inte stödja att man håller varandra om ryggen på det här sättet.
skriftlig. - (PL) I sitt betänkande om ECB:s årsrapport har föredraganden inriktat sig på de utmaningar Europeiska centralbanken står inför.
De senaste månaderna har det kommit en hel del oroande uppgifter om de europeiska ländernas ekonomi, och tyvärr är det mycket mer av den varan nu än under 2007.
Krisen på finansmarknaderna och de plötsliga prisökningarna på olja och livsmedel bromsar den ekonomiska tillväxten och driver upp inflationen, och det finns en oro för att arbetslösheten ska gå upp.
ECB kommer att vara en av de ledande institutioner som tvingas ta itu med dessa utmaningar.
Åtgärderna som vidtogs i augusti 2007 gav finansmarknaderna likviditet, men löste inte problemet.
Det sker också en ökning av antalet länder som ansluter sig till den gemensamma valutan.
Slovakien blir det första landet från Central- och Östeuropa som tar det steget.
Slovakien blir dock definitivt inte det sista landet.
Det verkar mest vara en tidsfråga när de andra nya medlemsstaterna går med i eurosamarbetet.
Slovakiens erfarenheter inom det området kommer säkerligen att studeras noga av andra länder i regionen som också planerar att ansluta sig till den gemensamma valutan.
Föredraganden konstaterar också med rätta att olika ekonomiska tillväxtnivåer, olika tillväxtindikatorer och olika grader av ekonomisk mognad i EU-länderna kan komma att skapa problem i ECB:s beslutsprocess.
Av det skälet anser jag att förslaget om att se över möjligheterna att göra förändringar i beslutsprocessen är förnuftigt.
En sådan översyn bör inte enbart omfatta eurozonens nuvarande medlemmar, utan även framtida och potentiella medlemmar.
skriftlig. - (EN) Jag välkomnar Olle Schmidts betänkande om ECB:s årsrapport.
Jag instämmer i föredragandens uppmaning till ECB om att fortsätta förbättra sina relationer till andra centralbanker och berörda institutioner.
Jag vill också upprepa Olle Schmidts rekommendation att man bör vara försiktig med fortsatta räntehöjningar för att inte skada den ekonomiska tillväxten.
Jag röstade för föredragandens bedömning.
I den resolution som vi ledamöter i Greklands kommunistparti har röstat emot försöker man på ett provocerande sätt att måla upp införandet av EMU och den gemensamma valutan för tio år sedan som en stor ”framgång”, samtidigt som arbetstagare och fattiga arbetarklassgrupper i EU-ländernas samhällen, däribland i Grekland, får känna av deras ödesdigra konsekvenser i form av bland annat höga priser, lönestopp och frysta pensioner, arbetslöshet, alltför hög beskattning av anställda och fattiga egenföretagare, slopade rättigheter för arbetstagare och slopade sociala och demokratiska rättigheter.
Den enda ”framgång” som uppnåtts handlar om de europeiska plutokraternas vinster och övervinster och går helt på tvärs mot arbetstagarnas och folkets intressen.
Europeiska centralbanken, ett renodlat verktyg för det europeiska kapitalet, ska nu spela en mer aktiv och effektiv roll i samma riktning via antifolkliga åtgärder som räntehöjningar och så vidare.
Genom resolutionens kommentarer om och oro för ”finanskrisen” och de ”sammanhållningsproblem” inom EU som kvarstår och faktiskt sprider sig, stärks vi i vår bedömning av de fortsatta och oundvikliga kriserna för det kapitalistiska systemet och dess orimliga tillväxt, liksom i vår övertygelse att detta system måste störtas och ersättas med ett folkligt planekonomiskt system där folket får makten, och att det är nödvändigt att kapa banden till det imperialistiska EU.
Inom EU finns det ingen väg till tillväxt som gynnar vanligt folk.
Inkomna dokument: se protokollet
Presentation av programmet för det franska ordförandeskapet (debatt)
Nästa punkt är rådets uttalande om presentationen av programmet för det franska ordförandeskapet.
President Sarkozy! Jag välkomnar er som rådsordförande till Europaparlamentet.
(Applåder)
Jag är medveten om att ni i dag besöker oss efter en lång resa från Japan.
Välkommen till Europaparlamentet, herr rådsordförande.
(Applåder)
Jag vill även välkomna Europeiska kommissionens ordförande José Manuel Durão Barroso, som i likhet med Europeiska rådets ordförande precis har återvänt från Japan.
Ni har en lång resa bakom er så jag ska inte ge några ytterligare kommentarer.
Herr rådsordförande! Härmed överlämnar jag ordet till er.
Herr talman, mina damer och herrar! Det är en stor ära för mig att få tala inför denna församling vid en sådan betydelsefull tidpunkt för Europa.
Jag är väl medveten om att ett tungt ansvar vilar på oss alla.
Naturligtvis har jag som rådsordförande ett stort ansvar, men alla vänner av Europa har samma ansvar.
Hur ska vi se till att Europa tar sig ur den kris det befinner sig i?
Hur förhindrar vi passivitet?
Hur gör vi för att överbrygga våra meningsskiljaktigheter och använda dem för att främja samma europeiska ideal?
Här står vi i hjärtat av den europeiska demokratin.
För var och en av er som har fått hedersuppdraget att vara parlamentsledamot har det varit ett måste att få era landsmäns stöd.
Det finns män och kvinnor från vänstern, från mitten och från högern. Det finns folkvalda representanter från 27 länder.
I dag måste vi emellertid förvandla våra meningsskiljaktigheter till en styrka för en plågad europeisk union.
Vi måste förvandla dessa meningsskiljaktigheter till en möjlighet att lugna de europeiska medborgare som är oroliga.
Vi måste hålla demokratin levande, vilket innebär att vi måste engagera oss i debatten samtidigt som vi visar att Europa inte accepterar passivitet.
Alla måste vara med i den europeiska familjen med dess 27 medlemsstater, ingen får lämnas på efterkälken.
Det återstår nu bara några månader till ett datum som är mycket viktigt för Europaparlamentet.
Det är rimligt att alla är medvetna om detta.
Samtidigt måste vi denna morgon visa att vi är ett Europa som arbetar för allas bästa.
Jag har upplevt enklare situationer än den som Europa nu befinner sig i.
Om jag får tala öppet, samtidigt som jag är medveten om att jag som rådsordförande måste tala på allas vägnar, så måste jag ta hänsyn till de frågor som är känsliga för de olika parterna samtidigt som jag kommer med de rätta svaren.
Min första iakttagelse är att vi har ett institutionellt problem.
Stats- och regeringscheferna har försökt att nå en kompromiss genom Lissabonfördraget.
Ingen har påstått att Lissabonfördraget kommer att lösa alla våra problem, men det har varit och fortsätter att vara ett uttryck för en kompromiss som är godtagbar för alla.
Som Frankrikes president har jag varit tvungen att ta mitt ansvar.
Frankrike röstade nej 2005 och det orsakade problem för Frankrike.
De frågor vi måste ta itu med är mycket svåra och komplicerade. Låt oss visa alla att vi arbetar med detta utan några baktankar eller fördomar.
Det är vad som förväntas av oss.
(Applåder)
Före valet erbjöd jag det franska folket parlamentsratificering av Lissabonfördraget.
Före valet sa jag att jag inte skulle hålla någon folkomröstning i Frankrike.
Jag sa detta till det franska folket i demokratisk anda. Det var ett val jag gjorde tre dagar innan jag valdes och det kunde ha fått stor betydelse.
Jag ångrar inte detta val.
Jag anser verkligen att beslut om institutionella frågor, det sätt vi hanterar saker och ting på i Europa, hellre bör fattas av parlamentsledamöterna än vid folkomröstningar.
Det är ett politiskt val som jag gör (applåder) och det är ett politiskt val som jag gjorde i mitt eget land före valet.
Därför är det helt demokratiskt.
Nu har vi ett problem i och med att irländarna röstade nej.
Det är inte min sak som fransman att sätta mig till doms när det gäller detta resultat, med tanke på att holländarna och fransmännen tidigare röstat nej.
Därför kommer jag den 21 juli att för första gången som rådsordförande resa till Irland för att lyssna, starta en dialog och försöka att hitta lösningar.
Det franska ordförandeskapet kommer att föreslå en metod och, förhoppningsvis, en lösning tillsammans med den irländska regeringen, i antingen oktober eller december.
Problemet är detta: vi måste både undvika att stressa våra irländska vänner och samtidigt fastställa på vilka villkor och med vilket fördrag vi ska organisera 2009 års val till Europaparlamentet.
Vi är skyldiga våra medmänniskor och medborgare detta.
Vi är skyldiga våra medmänniskor och medborgare att avgöra på vilken grund vi ska organisera valet till Europaparlamentet.
Grunden kommer att vara antingen Lissabonfördraget eller Nicefördraget.
Det kommer inte att hållas någon ny institutionell konferens.
Det kommer inte att upprättas något nytt fördrag.
Det är antingen Lissabon eller Nice.
Får jag även, bara för att vara helt tydlig, tillägga att jag - enligt min åsikt, men det innebär inte att det är sanningen - är en av dem som alltid har varit positivt inställd till den europeiska utvidgningen.
Utvidgningen 2004 var en framgång.
Familjen har återförenats, det bör vi inte beklaga.
Jag är emellertid även en av dem som alltid önskat att Europa hade varit tillräckligt klokt för att skapa nya institutioner före utvidgningen.
Detta var ett misstag som vi fortfarande betalar för.
Det skulle ha varit modigare att upprätta institutioner före utvidgningen.
Jag vill vara helt tydlig när det gäller detta.
Naturligtvis ångrar jag inte utvidgningen.
Familjen måste hålla ihop.
Det är dock min orubbliga ståndpunkt att vi inte får göra om samma misstag.
Om vi håller oss till Nice är det ett Europa med 27 länder.
Om vi vill ha en utvidgning - och jag personligen vill det - behöver vi nya institutioner före utvidgningen.
Vem skulle ha trott att EU med sina 27 medlemsstater skulle vara oförmöget att upprätta egna institutioner och att det inte skulle ha någon annan prioritering än att fortsätta utvidgas?
Förutsättningarna måste vara tydliga: om vi vill ha en utvidgning - och vi vill verkligen ha en utvidgning - behöver vi nya institutioner.
(Applåder)
Låt mig tillägga- och jag säger detta till Martin Schulz - att jag är för förslaget om att införliva Balkanstaterna, att våra kroatiska vänner precis som våra serbiska vänner utan tvekan är européer.
De länder som är mest positiva till utvidgningen kan emellertid inte säga ”vi vill inte ha Lissabon” och samtidigt säga ”vi vill ha en utvidgning”.
Vi ska ha Lissabon och vi ska ha utvidgning.
Det är inte utpressning eftersom vi i Europa inte sysslar med utpressning.
Det handlar om konsekvens, ärlighet och logik.
När det gäller Kroatien måste vi därför fortsätta med förhandlingarna, men alla bör ta sitt ansvar.
Om EU ska kunna växa, och det måste det, så måste det göra det med nya institutioner.
En annan punkt: då och då i de europeiska debatterna stöter jag på människor som säger ”det spelar ingen roll om vi har ett Europa i flera hastigheter”.
En dag kanske vi dessvärre är tvungna att ha ett Europa i flera hastigheter, men det bör endast vara en sista utväg.
Europa har betalat ett högt pris för att ha varit delat av en skammens mur.
Europa har betalat ett högt pris för den diktatur som 80 miljoner européer påtvingats.
Låt oss verkligen tänka efter innan vi låter någon hamna på efterkälken.
När vi förhandlade fram Lissabonfördraget i Bryssel stred Frankrike för att Polen skulle få inta sin plats i det fördraget.
Hur kan vi säga till 38 miljoner polacker att det är mycket lättare att göra sig av med oket från den diktatur de levde under och som de tack vare betydande personer som Lech Walesa och Johannes Paulus II själva befriade sig från, än att stanna kvar i ett fritt Europa?
Det finns 27 medlemmar i den här familjen.
Ingen får lämnas efter.
Vi måste få med oss alla i den europeiska familjen. Detta är åtminstone vad det franska ordförandeskapet kommer att arbeta för.
(Applåder)
När det gäller andra frågor, och jag tror att vi kan nå samförstånd om dem, skulle inget vara värre än att EU ger intryck av att vara passivt eftersom det går igenom ännu ett institutionellt drama.
Det vore en hemsk fälla för oss att hamna i.
Vi vill inte ha institutioner som dömer oss till passivitet, men samtidigt är européerna otåliga eftersom de tycker att vi är för passiva.
Trots det institutionella problemet, kanske till och med på grund av det institutionella problemet, har Europa en skyldighet att agera, och att agera nu.
Detta är det budskap som det franska ordförandeskapet vill förmedla till alla européer.
Vi arbetar med att lösa de institutionella problemen, men vi är inte dömda till passivitet.
Vilka är då våra prioriteringar?
Den första är att visa européerna att Europa kan skydda dem.
Jag skulle nu vilja säga något om ordet ”skydd”.
Sedan urminnes tider har människor valt en regering för att den ska skydda dem.
EU måste erbjuda skydd utan protektionism.
Protektionism leder oss ingenvart.
Att europeiska medborgare i dag tycker att EU, vars syfte är att skydda dem, är en källa till bekymmer snarare än skydd, är verkligen ett steg bakåt i utvecklingen.
Därför är det upp till oss att visa att EU kommer att skydda dem i konkreta frågor.
Den första frågan är energi- och klimatpaketet.
Om det finns ett område där våra nationer inte kan göra någonting på egen hand är det när det gäller att upprätthålla vår planets ekologiska balans.
När det gäller föroreningar, koldioxid och ozonskiktet är gränserna mellan våra länder irrelevanta.
Det är mycket som står på spel. Sedan mötet med IPCC:s experter har vi insett att vi är den sista generationen som kan förhindra en katastrof.
Den sista generationen!
Om vi inte gör något nu kanske de kommande generationerna kan begränsa skadorna, men de kommer inte att kunna stoppa dem.
Alla länder i världen säger: ”Jag är beredd att göra något om andra gör det först.”
Med denna typ av resonemang kommer våra barnbarns barnbarn aldrig att se några beslut fattas.
Om vi européer väntar på att andra ska göra något innan vi agerar kan vi få vänta länge.
Vi skapade EU för att föra ut vår civilisationsmodell i världen och försvara våra värden.
Bland dessa värden finns en förvissning om att världen är dömd till undergång om vi inte fattar ett beslut genast.
Europa måste föregå med gott exempel.
Europa måste leda vägen genom att föregå med gott exempel.
Vi har ett mål: konferensen 2009.
Vid denna konferens måste vi hantera och organisera fasen efter Kyoto.
EU måste komma enat till konferensen efter att ha beslutat sig för att anta energi- och klimatpaketet.
Om vi inte gör det kommer vi inte att ha något inflytande när det gäller att få kineserna, indierna, tillväxtekonomierna och amerikanerna att göra de ansträngningar vi har enats om.
Därför är det nödvändigt att vi under det franska ordförandeskapet antar det energi- och klimatpaket som lagts fram av kommissionen.
(Applåder)
Det är ett krävande paket, det är ett svårt paket, men jag vill vädja till allas ansvarskänsla.
Om varje land börjar vilja omförhandla frågor som rör deras egna orosmoment, de saker landet har problem med, kommer vi aldrig att nå en överenskommelse.
Det är därför det franska ordförandeskapet ber Europaparlamentet att gemensamt stödja oss så att vi kan anta energi- och klimatpaketet inom de kommande sex månaderna.
Det är en prioritering.
Det är inte en höger- eller vänsterprioritering, utan vanligt sunt förnuft.
Om vi ska inleda separata förhandlingar med varje medlemsstat har vi ingen chans att lyckas.
Nu finns det naturligtvis punkter där det krävs förtydliganden eller anpassningar.
Jag tänker framför allt på en mycket svår fråga, nämligen problemen för våra företag, för vilka vi med rätta kommer att införa bestämmelser för att upprätthålla planetens balans.
Bör vi i Europa införa nödvändiga lagar för våra företag samtidigt som vi fortsätter att importera produkter från länder som inte följer någon av de lagar vi förväntar oss att företagen i våra länder ska följa?
Det handlar inte om protektionism utan om rimlighet, rättvisa och en vägran att vara naiv.
Ett problem är att besluta om en mekanism för gränsöverskridande tillsyn.
Bör vi ha tullfria kvoter eller anpassningsmekanismer?
Jag vet inte, men vi måste under alla omständigheter diskutera detta.
(Applåder)
En andra fråga: Jag förstår att det för vissa länder krävs avsevärda ansträngningar - jag tänker framför allt på dem som blev EU-medlemmar 2004, som till stor del är beroende av fossila bränslen för att få energi.
Dessa länder säger: ”Vi har haft tillväxt i 10 år, snälla ta inte det ifrån oss”.
Det finns utan tvekan ett sätt att få med alla, och tillsammans med kommissionens ordförande måste vi arbeta för detta så att alla inser att de inte döms till lågkonjunktur, elände, fattigdom och arbetslöshet.
Detta energi- och klimatpaket är en absolut prioritering för oss.
Världen kan inte vänta.
Europa måste visa vägen.
Den andra punkten. Av de 27 länderna ingår nu 24 i Schengenområdet, dvs. 24 länder av 27.
23 säger ni?
Okej, 23 då, men det är fortfarande inget dåligt resultat.
Här ingår inte länder som står utanför Europeiska unionen men - och det är därför vi ofta har debatter - ingår i Schengenområdet.
Så vad innebär detta?
Det innebär att vi har beslutat att fullständigt fri rörlighet ska råda mellan länderna i Schengenområdet.
Till ledarna för de politiska grupperna och parlamentsledamöterna vill jag säga att vi i Frankrike, med Bernard Kouchner och Jean-Pierre Jouyet, har fattat ett beslut som inte var enkelt.
Sedan den 1 juli har det inte längre funnits några hinder för tillträde till den franska arbetsmarknaden eftersom jag har meddelat att jag kommer att avskaffa alla restriktioner som mina företrädare förhandlat fram.
Alla arbetstagare från alla EU-länder kan komma och arbeta i Frankrike.
(Applåder)
Det var inte enkelt, det var inte lätt.
Hur som helst, och de franska parlamentsledamöterna kommer att rätta mig om jag har fel, fick jag höra att det vore en katastrof om jag tillkännagav detta beslut.
Som vanligt fattade vi beslutet och ingen katastrof uppstod.
Jag var inte glad över kontroversen med den ökände polske rörmokaren, som inte gav vare sig mitt land eller för den delen Europa något särskilt gott rykte.
Det är inte därför vi alla har byggt upp Europeiska unionen.
(Applåder)
När vi nu inte längre har några gränser mellan oss, är det då rättvist och rimligt att var och en av oss får bestämma över sin egen invandringspolitik utan att behöva ta hänsyn till de andra ländernas restriktioner?
Den europeiska pakten för invandring och asyl är ett nödvändigt dokument för det franska ordförandeskapet, av två orsaker.
Den första av dessa - och får jag vända mig till den vänstra sidan av kammaren först - är att om vi alla, om alla europeiska länder, har en europeisk invandringspolitik, försvinner invandringsfrågan från nationella debatter där extremister utnyttjar fattigdom och rädsla för att främja värderingar som vi inte stöder.
Det enda sättet att ha en ansvarsfull debatt om invandringen är att göra den till en europeisk politik.
Inga fler partipolitiska baktankar som tvingar länder som har olika ömma punkter att samarbeta.
Det som Brice Hortefeux föreslog, som godkändes av alla ministrar och ska diskuteras av Ständiga representanternas kommitté och av Europeiska rådet, ser jag som en prioritering.
Det kommer att visa att Europa inte vill vara en fästning, att Europa inte vägrar att ta emot människor, att Europa behöver migrerande arbetstagare, men att Europa inte kan ta emot alla som vill komma hit.
Låt mig tillägga att när det handlar om politisk asyl så är det inte logiskt att en individ ska kunna skicka 27 ansökningar till 27 demokratiska länder och inte få samma svar varje gång på samma fråga.
Låt mig tillägga att när det gäller utvecklingen för Afrika kommer vi att bli starkare om vi samarbetar. Detta är det franska ordförandeskapets andra prioritering.
Den tredje prioriteringen: vi vill främja ett koncept som det ofta talas om i Europa, men där utvecklingen går långsamt, nämligen ett europeiskt försvar.
Jag är väl medveten om att det råder stor oenighet i denna fråga, men låt mig berätta vad jag anser.
Hur tror ni att Europa ska kunna bli en politisk makt och göra sin röst hörd om det inte kan försvara sig och utveckla resurser till stöd för sin politik?
Ta exemplet Kosovo, som enligt min mening är en framgångssaga för Europeiska unionen.
Detta är ett europeiskt problem, som måste lösas av européer.
Hur kan européer fortsätta att göra det om de inte skaffar de militära och mänskliga resurser som krävs för att driva igenom de beslut vi fattat tillsammans?
Hur tror ni att Europa ska kunna bli det mest blomstrande ekonomiska området i världen om vi inte kan försvara oss?
Ja, vi har Nato.
Det skulle inte falla någon in, minst av alla mig, att ifrågasätta nyttan med Nato.
Det handlar inte om att välja mellan en europeisk försvarspolitik eller Nato, utan om att ha Nato - alliansen med amerikanerna - och en självständig europeisk säkerhetspolitik.
Det handlar om att ha båda dessa tillsammans och inte det ena i stället för det andra.
Låt mig tillägga att vi inte kan fortsätta att garantera Europas säkerhet om endast fyra eller fem länder bidrar, medan de andra förlitar sig på insatserna från dessa fyra eller fem länder.
Medlemsstaterna kan inte fortsätta att bygga upp sin egen luftfart, och ha vapenindustrier som tävlar mot varandra så att de går under och medlemsstaterna i slutändan försvagas, bara för att de inte är tillräckligt starka för att ha en europeisk försvarspolitik.
Den fjärde prioriteringen: den ytterst svåra frågan om den gemensamma jordbrukspolitiken.
Jag närmar mig nu min slutsats som är kopplad till denna fråga.
Det är just för att den är så svår att tala om som vi måste tala om den.
Jag är väl medveten om att vi bland oss har jordbruksländer som kraftfullt försvarar sina jordbrukare och samtidigt medlemsstater som tycker att denna politik kostar för mycket.
Jag vill vädja till ert sunda förnuft.
År 2050 kommer världen att ha 9 miljarder invånare.
Redan nu dör 800 miljoner människor av svält.
Ett barn svälter ihjäl var trettionde sekund.
Är det rimligt att begära att Europa ska minska sin jordbruksproduktion vid en tidpunkt då världen har ett så starkt behov av livsmedel?
Jag tycker inte detta är rimligt.
Det handlar inte om franskt jordbruk utan om sunt förnuft.
(Applåder)
Låt mig lägga till en andra punkt: oavsett om ert land är ett jordbruksland eller inte så är livsmedelssäkerhet en fråga som berör alla.
Är det rimligt att våra uppfödare och jordbrukare ska omfattas av bestämmelser om spårbarhet och säkerhet samtidigt som vi fortsätter att importera kött till Europa från andra länder som inte följer de bestämmelser som vi kräver att våra jordbrukare ska följa?
(Applåder)
Den tredje punkten: jordbrukskostnaderna har aldrig varit så höga som nu.
Det är verkligen rätt tidpunkt att tala om kostnader, subventioner och gemenskapens preferenssystem.
Jag tror också att vi mellan den gemensamma jordbrukspolitikens hälsokontroll och ekonomiska förlikning kan enas om vissa begrepp såsom livsmedelsoberoende och livsmedelstrygghet för Europa.
Det finns en rad andra frågor. Den sociala dimensionen är ett exempel på en viktig fråga.
Låt mig påpeka något.
Ibland upplever jag en viss inkonsekvens. Ibland förekommer en ensidig åsikt som går ut på att EU inte bör blanda sig i allt utan endast bör ingripa på områden som det direkt berörs av.
Samma människor som anklagar EU för att lägga näsan i blöt överallt är de första som höjer rösten om vi inte talar om den sociala dimensionen.
Fram till nu har medlemsstaterna alltid velat att socialpolitiken först och främst ska omfattas av nationell behörighet, eftersom pensioner och hälso- och sjukvård främst är nationella frågor.
Det finns en rad sociala direktiv som ordförande Barroso gjort rätt i att sätta upp på dagordningen.
Jag tänker på dem som gäller företagsråd, tillfälligt arbete och ett antal grundläggande bestämmelser som alla i Europa måste följa.
Det franska ordförandeskapet kommer att prioritera detta.
Andra ämnen bör också sättas upp på det franska ordförandeskapets dagordning, även om de inte tillhör EU:s ansvarsområde.
Låt mig ge ett exempel på något som påverkar oss alla: Alzheimers sjukdom.
(Daniel Cohn-Bendit kommenterar utan mikrofon: ”Inte än”).
Herr Cohn-Bendit! Det skulle aldrig falla mig in att någon som är så ung som ni redan skulle ha drabbats av en sjukdom som även om den inte drabbat er, drabbar miljontals européer.
Dessa miljontals européer är lika viktiga för mig som er hälsa.
(Applåder)
Naturligtvis innebär subsidiaritetsprincipen att detta inte faller under europeisk behörighet.
Jag skulle ändå vilja att det franska ordförandeskapet anordnar ett möte för alla specialister från alla europeiska länder, så att vi kan utbyta bra metoder, så att våra forskare kan förena sina kunskaper för att få veta mer om denna sjukdom och så att vi tillsammans kan hitta en lösning.
Föreställ er bara vad européerna i så fall skulle säga om EU: att det är ett sätt att bota dessa hemska sjukdomar.
Det som jag sa om Alzheimers skulle även kunna gälla cancer, som splittrar familjer.
Det finns ingen anledning till att alla ska arbeta var för sig för att hitta sätt att bota cancer, när vi tillsammans har mer resurser och är starkare.
(Applåder)
Låt mig avslutningsvis säga att när det gäller kultur och idrott så är det ett stort misstag att inte prata om de frågor som påverkar européernas vardag.
Det finns ett europeiskt kulturellt undantag.
Vi måste göra kulturen till en del av den dagliga debatten i Europa.
Världen behöver inte underkasta sig ett språk och en kultur.
Vi måste helt klart ta itu med frågan om mervärdesskatt på videofilmer och cd-skivor, precis som mervärdesskatt på böcker, som ni har löst.
När det gäller idrott, som överbryggar politiska klyftor, så låt mig bara säga att jag skulle vilja att det fanns ett undantag för idrott i Europa, precis som det finns ett kulturellt undantag.
Jag är för den fria rörligheten för personer och varor, men jag accepterar inte förslaget om att vi ska tvinga våra fotbollsklubbar att betala, och undergräva den investering som många klubbar gör i tonårspojkar, som måste stanna i klubben av träningsskäl.
Ett undantag för idrott, som skulle innebära att idrotten inte står i tacksamhetsskuld till marknadsekonomin, borde stödjas av alla parlamentsledamöter.
(Applåder)
Jag vill avsluta med en sista iakttagelse - och jag ber om ursäkt för att jag utan tvekan talat för länge.
Jag är medveten om var jag gör denna iakttagelse: på den plats där den europeiska demokratins hjärta slår.
Europa har genomlidit mycket.
Det har först och främst drabbats av fegheten hos vissa av oss som varit nöjda med att låta Europa betala för sådant som i själva verket varit de politiska ledarnas ansvar, men som de varit ovilliga att offentligt fatta beslut om och vägrat att försvara i Bryssel.
(Applåder)
Detta är fel.
Till Europaparlamentets talman och kommissionens ordförande vill jag säga att ordförandeskapet kommer att arbeta sida vid sida med er.
Om någon medlemsstat har något emot detta kan den göra sin röst hörd.
Som jag sa till den polske presidenten, som själv förhandlat fram Lissabonfördraget, har han gett sitt löfte och ett löfte måste hållas.
Det handlar inte om politik utan om moral.
(Applåder)
Europa har emellertid drabbats av något annat också.
Europa har drabbats av avsaknaden av en debatt.
Jag vill avsluta med detta eftersom det är väldigt viktigt för mig.
Våra institutioner är oberoende, men oberoende är inte samma sak som likgiltighet.
Om vi, de politiska ledarna, inte har modet att debattera, vem ska då ha det?
Vad är det som ska debatteras?
Vilken är den rätta ekonomiska strategin?
Vilken är den rätta monetära strategin?
Vilken är den rätta växelkursstrategin?
Vilken är den rätta räntestrategin?
Naturligtvis har alla rätt till sina egna övertygelser, och det säger jag framför allt till våra tyska vänner.
Ingen har emellertid rätt att förhindra en debatt, en konstruktiv debatt.
Naturligtvis vill alla ha ett avtal som det handelsavtal som håller på att förhandlas fram.
Ingen får emellertid vara rädd för att säga att EU inte får vara naivt.
Vi måste diskutera fördelarna med frihandel, men vi måste även berätta för tillväxtekonomier att de inte har något skäl att kräva samma rättigheter utan att även omfattas av samma skyldigheter.
Vi får inte vara rädda för att ha en europeisk debatt.
Vi måste engagera oss i en värdig europeisk debatt, men vi får inte vara rädda för att försvara våra övertygelser.
Vi ifrågasätter inte Europeiska centralbankens oberoende när vi frågar om det är rimligt att höja räntesatserna till 4,25 procent när de amerikanska räntesatserna är 2 procent.
Vi har en debatt.
En fredlig debatt, där ingen har monopol på sanningen.
Jag har det sannerligen inte, och inte heller experterna, som måste bevisa effektiviteten i sina beslut.
Det är i denna anda som jag tillsammans med de franska ministrarna avser att ta mitt ansvar.
Jag vet att det är svårt.
Jag vet att man som rådsordförande inte försvarar sitt eget lands intresse utan unionens intresse.
Jag vet, herr talman och herr ordförande, att vi måste samarbeta i de 27 länderna i EU:s intresse och jag hoppas att alla om sex månader kommer att kunna säga: ”EU har gjort framsteg tack vare ert deltagande och stöd”.
(Livliga applåder)
Herr rådsordförande! Tack för ert anförande.
Vi önskar er fortsatt mod, beslutsamhet och framför allt framgång under ert ordförandeskap - eftersom er framgång är en framgång för Europeiska unionen och därmed för Europaparlamentet.
Ni kan vara säker på att Europaparlamentet finns vid er sida när ni med fasthet bidrar till att föra Europeiska unionen framåt mot en bra framtid.
Europaparlamentet kommer att stödja er i detta arbete.
Jag vill även välkomna de ministrar som är här med er i dag: Bernard Kouchner, Brice Hortefeux, tidigare parlamentsledamot, och framför allt er unge EU-minister, Jean-Pierre Jouyet, som nästan alltid är här i parlamentet.
Jag välkomnar er alla varmt till Europaparlamentet.
(Applåder)
kommissionens ordförande. - (FR) Herr talman, herr rådsordförande, mina damer och herrar! Jag är glad över att vara här med er i Europaparlamentet i dag för presentationen av Frankrikes sex månader långa ordförandeskap för Europeiska unionen.
Jag tror att det kommer att bli ett ordförandeskap fullt av drivkraft och beslutsamhet och rikt på konkreta resultat som vi alla kommer att bidra till.
Ni ville att Frankrike skulle återvända till Europa, herr rådsordförande, och detta är utan tvekan fantastiska nyheter för oss alla.
De europeiska medborgarna och Europaparlamentet som samlats här i dag förväntar sig stora saker av det franska ordförandeskapet.
Som jag sa vid vårt möte i Paris den 1 juli kommer kommissionen helhjärtat att stödja det franska ordförandeskapet för att se till att Europeiska unionen blir framgångsrik under dessa sex månader.
Det kommer inte att saknas utmaningar.
Globaliseringen har kommit för att stanna och den internationella konkurrensen blir allt hårdare.
Världen står inför nya utmaningar, såsom bristen på fossila bränslen och klimatförändringarna.
Vi måste agera nu för att hitta gemensamma lösningar på dessa utmaningar.
Alla dessa faktorer innebär att EU måste reformera sin ekonomi för att bli mer konkurrenskraftigt, modernisera sina sociala modeller och investera i utbildning, forskning och innovation.
EU har många ess i rockärmen, framför allt som en av världens ledande handelsmakter.
Det måste emellertid ha modet att anpassa sig.
Om vi vill erbjuda skydd måste vi anpassa oss.
Det är avgörande.
Det är ingen mening att förneka att EU genomgår en svår period: det irländska folkets nej i folkomröstningen och det globala ekonomiska klimatet, de ständigt ökande priserna på olja och handelsvaror, de kraftigt stigande livsmedelspriserna och inflationstrycket, som är köpkraftens största fiende.
Inflationen är även den sociala rättvisans största fiende eftersom de som drabbas mest vid en kraftig inflation är de som har låga löner eller lever på pension.
Alla dessa faktorer kastar en skugga över våra ekonomier och tvingar våra politiker på både EU-nivå och nationell nivå att fatta svåra beslut.
Vi måste möta denna verklighet utan omsvep och hantera den med realism och beslutsamhet.
Vi har precis återkommit från G8-mötet i Japan, där jag tydligt kunde se att det inflytande Europeiska unionen har och de förväntningar och den respekt den framkallar runt om i världen, står i bjärt kontrast till den förstämning som ofta uttrycks inom EU.
Jag kan informera er om att Europeiska unionen nu mer än någonsin tidigare av länderna utanför Europa betraktas som en positiv och bestämd aktör, en aktör med ett enormt inflytande på världsscenen.
Låt oss ta upp två konkreta ämnen som var centrala på G8-mötet: klimatförändringarna och utvecklingen - två frågor där Europa har tagit initiativet på global nivå.
Förenta staterna har nu förenat sig med oss i kampen mot klimatförändringarna genom att till stor del ansluta sig till våra åsikter.
Förra året i Heiligendamm - president Sarkozy var där - minns jag att vi hade stora svårigheter när det gällde att övertyga amerikanerna och ryssarna om att acceptera principen om obligatoriska mål för 2050.
Nu har vi uppnått detta.
Det var möjligt tack vare vår roll som europeisk ledare. Som ordförande för en europeisk institution är jag stolt över detta.
Det är en framgång som vi återigen har den europeiska enigheten att tacka för.
Det andra exemplet är utvecklingen, och framför allt de stigande livsmedelspriserna, som hotar alla millennieutvecklingsmålen.
Vi kunde fungera som katalysator även på detta område tack vare slutsatserna från förra månadens möte med Europeiska rådet som, jag citerar, välkomnade ”kommissionens planer på att lägga fram ett förslag till en ny fond för att stödja jordbruket i utvecklingsländerna”.
Europeiska kommissionen kommer att anta detta förslag nästa vecka.
Jag räknar med helhjärtat stöd från budgetmyndighetens båda grenar så att Europa snabbt kan förse jordbrukarna, framför allt dem i Afrika, med nödvändigt bistånd, i nära samarbete med behöriga multilaterala organisationer.
Detta stöd är nödvändigt för att garantera ”den gröna revolution” som krävs för att Afrika ska uppnå stabilitet och välfärd, vilket som ni alla vet, även ligger i Europas intresse.
Som Europeiska rådet efterfrågade kommer vårt förslag att ligga inom gränserna för den aktuella budgetramen.
Vår strategi går ut på att låta de besparingar som EU, som ett led i politiken för jordbruksstöd, kunnat genomföra tack vare ökningen av de internationella priserna gå till dem som drabbas hårdast av denna ökning.
Det inträffar nöd- och katastrofsituationer över hela världen.
Om ni hade hört vad ordföranden för Världsbanken sa, om ni hade hört några av ledarna för afrikanska länder och andra länder som var företrädda vid utökade möten tala om den hunger och svält som nu utgör ett verkligt hot mot så många människor i världen, skulle ni förstå hur nödvändigt och oumbärligt EU:s bistånd är.
(Applåder)
Det är därför jag tror att vi återigen kan föregå med gott exempel när det gäller solidaritet mellan europeiska och afrikanska jordbrukare, och illustrera det faktum att den gemensamma jordbrukspolitiken (GJP) och utvecklingspolitiken kan och måste fungera sida vid sida eftersom livsmedelstrygghet, precis som president Nicolas Sarkozy just sa, är en global fråga som vi behöver ta itu med gemensamt.
Inte var för sig utan tillsammans.
Därför är det sant att det finns orosmoment, men det är också sant att Europeiska unionen mer än någonsin tidigare har en central roll när det gäller att ta itu med dem.
Låt oss i stället för att vältra oss i vad jag ibland kallar ”kriskultur” - det förekommer till och med tal om en permanent tillbakagång i Europa - framhäva värdet av EU:s konkreta och positiva åtgärder.
Hur som helst är detta det bästa sättet att lösa de internationella problem som orsakats av att Irland inte ratificerat Lissabonfördraget.
Vi måste ta itu med detta eftersom Lissabonfördraget skulle kunna göra det möjligt för oss att arbeta mer effektivt, mer demokratiskt, men vi får inte använda det som en ursäkt för att underlåta att omedelbart svara på våra medborgares behov.
De europeiska medborgarna förväntar sig svar av oss.
Det bästa svaret vi kan ge dem är att tala uppriktigt med dem och visa att vi har politiskt mod.
Det franska ordförandeskapet har båda dessa kvaliteter i överflöd.
I ett hårt prövat EU måste vi bevisa att unionen fungerar.
Vi måste fokusera på politik som för EU närmare medborgarna och förändrar deras vardag.
Mer än någonsin tidigare planerar vi för ett EU baserat på resultat.
Personligen känner jag tillförsikt.
Genom ert ordförandeskaps prioriteringar blir det möjligt för Europa att möta de stora utmaningar det står inför, och samtidigt förbereda sig inför kommande problem.
Jag välkomnar det franska ordförandeskapets prioritering när det gäller en integrerad politik för energi och klimatförändringar.
Som ni sa, herr rådsordförande, är detta den viktigaste prioriteringen för ert ordförandeskap, och vi vet hur bestämd ni är när det gäller att slutföra detta strategiska avtal före årsskiftet, så att EU får en bra utgångspunkt för att inleda Köpenhamnsförhandlingarna om ett år.
Kommissionen kommer helhjärtat att stödja detta så att vi kan nå ett ambitiöst och balanserat avtal med Europaparlamentet och medlemsstaterna.
Jag har gjort detta till en prioritering för min institution, och jag vill återigen tacka rådsordföranden för hans outtröttliga stöd för det energi- och klimatpaket som presenterats av Europeiska kommissionen.
Vi måste också röra oss mot en politik för kontrollerad invandring i Europa.
Vi måste först hantera den invandring som ett åldrande Europa behöver i vissa viktiga ekonomiska sektorer och som måste vara förenad med en riktig integration, så att vi i vårt humanistiska Europa kan vara stolta över den integration vi erbjuder dem som verkligen vill komma hit för att arbeta.
Införande av blåkortet under det franska ordförandeskapet vore ett viktigt steg i denna riktning.
Vi måste emellertid även ta itu med den olagliga invandringen och den exploatering som den ofta ger upphov till, framför allt genom att stödja förslaget om påföljder för dem som anställer svart arbetskraft.
Det är här vi faktiskt måste göra den största insatsen. Vi ska inte hota de stackars arbetstagare som bara vill arbeta i Europa, utan straffa dem som vill exploatera dem.
Dessa tvivelaktiga metoder är en skam för Europa.
Det får inte råda något tvivel om att vi kommer att hantera invandringsfrågan på ett realistiskt sätt.
Jag är övertygad om att vår oförmåga att hantera denna fråga seriöst och ansvarsfullt är ett av de största hoten mot Europa.
Vi löser inte invandringsfrågan genom att vara släpphänta på alla fronter.
Det vore en perfekt ursäkt för extremistiska och främlingsfientliga krafter.
Vi måste vara hårda när det gäller olaglig invandring och samtidigt visa att vi är generösa och enade när det gäller att integrera invandrargrupper som vill bidra till Europas tillväxt och utveckling.
Jag anser att vi måste vara tydliga på den här punkten - vi måste vara hårda när det gäller brott och samtidigt fortsätta att respektera de mänskliga rättigheterna, som är kännetecknande för den europeiska civilisationen och våra planer för den europeiska integrationen.
Detta är naturligtvis känsliga frågor som kan ge upphov till polemik och missförstånd.
Det var därför kommissionen ville lägga fram ett balanserat förslag och skisserade 10 huvudprinciper, så att vi kan röra oss framåt tillsammans.
Det gladde mig verkligen att det franska ordförandeskapet och de franska justitie- och inrikesministrarna stödde denna integrerade strategi vid sitt informella möte i Cannes denna vecka.
Jag vill påpeka att det vore absurt att fortsätta med 27 olika typer av invandringspolitik i Europa och Schengenområdet, där fri rörlighet är en realitet.
Det vi behöver är en europeisk invandringspolitik.
Vår sociala agenda är också under planering.
Utan riktiga sociala investeringar som förhindrar risken för fattigdom, utanförskap och marginalisering kan det inte finnas någon dynamisk och konkurrenskraftig ekonomisk modell.
Frankrike har gjort den nya sociala agenda som Europeiska kommissionen presenterade för några dagar sedan till en av sina prioriteringar.
Jag välkomnar detta.
För att förbereda européerna inför framtiden måste vi erbjuda dem möjligheter, tillgång till kvalitetstjänster, utbildning, hälso- och sjukvård och fortsatt solidaritet.
Ingen i Europa får slås ut.
Möjligheter och solidaritet är vad EU handlar om.
Många andra projekt kommer att dras i gång de kommande sex månaderna.
Jag kan inte beskriva dem alla här, men om jag får ge en kortfattad översikt över två av dem skulle jag vilja berömma projekten för europeiskt försvar och unionen för Medelhavsområdet, som kommer att presenteras nästa söndag i Paris.
Jag ser dessa projekt som två möjligheter för EU att bekräfta sin roll i världen.
Även här är det upp till oss att omvandla denna ambition till konkreta åtgärder.
Jag önskar det franska ordförandeskapet all lycka och garanterar kommissionens helhjärtade stöd under de kommande sex månaderna, som ser ut att bli spännande.
Politikernas första plikt är att möta utmaningarna och intensifiera insatserna för att kunna ta itu med dem på ett framgångsrikt sätt.
Vi kan göra mycket tillsammans.
Jag vill hylla de insatser som den franska regeringen genomfört på högsta nivå under de senaste månaderna för att ha ett nära samarbete med de europeiska institutionerna.
Institutionerna, ordförandeskapet och medlemsstaterna måste alla arbeta sida vid sida.
Detta är avgörande för att nå den gemensamma framgång som vi är skyldiga Europas medborgare, och jag vill hylla det engagemang som rådsordföranden i dag återigen ger uttryck för, för att rådet, parlamentet och kommissionen tillsammans ska kunna hitta konkreta lösningar på de konkreta problem som våra medborgare möter varje dag.
Herr talman, herr rådsordförande, herr kommissionsordförande, mina damer och herrar! Frankrike har beslutat att dess ordförandeskap ska vara synonymt med politiskt engagemang.
Vi behöver politiskt engagemang för att besegra de svårigheter som den europeiska integrationen står inför.
Den största av dessa är utan tvekan det irländska folkets nej i folkomröstningen som vi diskuterat här denna morgon.
Vi måste engagera våra medborgare i Europa.
Det finns många orsaker till att de känner tvivel, bland annat rädsla för globaliseringen, de ökade priserna och förändringarna av traditionella familjevärden och sociala värden.
Om vi inte kan övertyga alla om att det endast är på EU-nivå som det går att förhandla effektivt om viktiga frågor som säkerhet, klimatförändringar, energi och migration kan vi inte räkna med att få en fredlig framtid - och när det gäller världens större regioner måste EU även vara tillräckligt starkt för att övertyga USA, Indien, Kina och Brasilien.
Det franska ordförandeskapet kommer också att behöva politiskt engagemang för att övertyga sina samarbetspartner om att Lissabonfördraget kommer att hjälpa oss att fatta beslut på ett mer effektivt och demokratiskt sätt när det gäller alla dessa gemensamma frågor.
De ledamöter av min grupp som tillhör Europeiska folkpartiet vill att alla medlemsstater som inte redan har ratificerat fördraget ska göra det under det franska ordförandeskapet.
Efter en period av reflektion och med all respekt ser vi precis som vi gjorde i fråga om Frankrike och Nederländerna fram emot att Irland ska erbjuda landets 26 samarbetspartner en lösning på dödläget.
Vi ber varje medlemsstat att avstå från att försöka platta till andra och agera ansvarsfullt.
Vår grupp vill se ett slut på denna institutionella debatt och vi är övertygade om att det franska ordförandeskapet kommer att arbeta mot detta mål.
Samtidigt som vi försöker förse oss med ett bättre verktyg för att fatta beslut ökar våra problem.
Detta stjäl energi som skulle behövas för att skapa sysselsättning, försvara våra intressen och främja vår sociala modell och Europa i allmänhet.
Som jag sagt kommer vi definitivt att behöva politiskt engagemang.
Vi bör även se till att vi har det engagemang som krävs för att ta itu med de prioriteringar som rådsordföranden just har presenterat.
Vi måste agera skyndsamt för att ta itu med klimatförändringar, energi, migration, livsmedelstrygghet och försvar.
När det gäller klimatförändringar och energi är alternativet tydligt: antingen är våra medlemsstater övertygade om att de måste gå vidare och föregå med gott exempel inför toppmötet i Köpenhamn, och i så fall måste vi fatta tydliga beslut före december för att garantera ömsesidighet från våra internationella samarbetspartner, eller så har de beslutat att det trots de försämrade klimatvillkoren och beroendet av energin inte finns något behov av att vidta brådskande åtgärder.
Jag behöver knappast säga åt vilket håll min politiska grupp lutar.
Även när det gäller migration vill vi ha ett slut på detta hyckleri.
Även om flera länder runt om i världen redan har antagit en invandringspolitik med relativt tillfredsställande resultat har de flesta av våra länder skjutit upp dessa val.
Det är dags för en debatt och ett beslut i frågan, som måste vara positivt, humant och ansvarsfullt.
Förslaget till en europeisk pakt för invandring och asyl, som kommer att debatteras i oktober, är ett steg i rätt riktning och jag gratulerar EU:s ministrar till deras svar på det förslag som utarbetats av Brice Hortefeux.
Ni har vårt stöd, herr Hortefeux.
Avslutningsvis vill jag nämna två ämnen som ligger mig mycket varmt om hjärtat och som är ytterst viktiga för framtiden och för vårt oberoende: livsmedelstrygghet och försvar.
Jag vill att vi ska tänka på dem som har det sämst ställt, både runt om i världen och i våra egna länder, dem som de ökande livsmedelspriserna verkligen är ett problem för.
Jag vill att EU och det franska ordförandeskapet gör en ansträngning för att hjälpa dem i dessa svåra tider.
När det gäller försvar vill jag bara ställa en fråga: Hur kan EU vara trovärdigt utan ett försvar värt namnet?
Vi behöver ett försvar för att garantera fred i Europa och för att hjälpa dem som har det sämst ställt i världen.
Vår grupp stöder det franska ordförandeskapets engagemang att leda vägen genom att komma med modiga förslag till sina samarbetspartner på dessa två strategiska områden.
Den europeiska integrationen är i högsta grad en politisk fråga.
Jag hyser inga tvivel om att våra medborgare återigen kommer att känna sympati för EU om vi är tillräckligt modiga för att fatta tydliga politiska beslut.
Jag har fullt förtroende för att det nya ordförandeskapet kommer att uppmuntra oss i detta, och vi har allt att vinna på att få våra medborgares tillit innan 2009 års val till Europaparlamentet.
Herr talman, mina damer och herrar!
Det finns aspekter av era åsikter som vi delar, herr Sarkozy, och jag vill först av allt gå närmare in på några av dessa.
Det gläder mig att ni har återvänt välbehållen från Japan.
Vi har nu återigen hört om de kommande åtagandena när det gäller klimatförändringarna och det är hög tid att vi genomför dessa.
Ni har rätt i att klimatpaketet är en prioritering. Vår grupp delar denna åsikt med er.
Ni har även rätt när ni säger att enskilda länder inte kan uppnå detta på egen hand - inte ens tyskarna eller fransmännen genom att nå egna överenskommelser i Straubing.
Det är 25 andra länder som ingår i detta och framför allt är det Europaparlamentet som fattar det slutgiltiga beslutet.
Vi kommer att göra det tillsammans med er, genom att samarbeta, men ta inga initiativ vid sidan om - inte ens med Angela Merkel, oavsett hur bra denna idé verkar.
Eftersom ni nämner idrott vill jag påpeka att jag tittade i de franska dagstidningarna i morse eftersom jag undrade vad de skulle skriva om president Nicolas Sarkozys besök i Europaparlamentet i dag.
Ingenting!
De skriver mycket om Tour de France, där det för närvarande är en tysk som har den gula tröjan.
(Häcklande)
Jag lyssnade noggrant på er, herr rådsordförande, och de punkter ni tog upp om klimatförändringarna och framför allt om Lissabonfördraget.
Om vi ska kunna uppnå resultat behöver vi verkligen instrument och detta försätter oss i ett dilemma.
Medborgarna vill att vi ska bli mer effektiva, mer öppna, mer demokratiska och de vill att de nationella parlamenten ska bli mer demokratiska och få mer inflytande.
Allt detta är rätt, men varje gång vi vill uppnå resultat rycks det instrument vi behöver - ett reviderat fördrag - bort från oss.
Ni har rätt, detta innebär att vi behöver en ny taktik, och en ny start.
Vi måste se till att detta fördrag träder i kraft.
Jag tycker att det är fantastiskt att ni ska åka till Irland och arbeta konstruktivt med det irländska folket.
Om jag får ge er ett personligt tips tycker jag att ni ska lämna kvar Bernard Kouchner i Paris denna gång.
Jag fick intrycket att hans tidigare bidrag inte direkt hjälpte oss att övertyga irländarna.
(Applåder, häcklande)
Jag talar emellertid om en fråga där vår uppfattning är raka motsatsen till er.
Ni talar om fyra prioriteringar för ert ordförandeskap och jag väntade för att se om det fanns en femte.
Sedan nämnde ni flera andra saker som ni sa var viktiga - inte prioriteringar, bara andra saker.
Dessa ”andra saker” var bland annat ett socialt Europa, som ni tyckte var ett ärende för nationalstaterna.
Jag anser att detta är ett allvarligt misstag.
(Applåder)
Jag vill säga er att vi förväntar oss en annan taktik från det franska ordförandeskapet.
Ett socialt Europa innebär inte att vi vill upprätta ett socialförsäkringskontor i Europa eller att vi vill göra barnbidrag till en EU-fråga.
Ett socialt Europa handlar om något annat: under en lång tid har människor trott - med rätta - att Europa kan göra ekonomiska framsteg möjliga.
Vi har ägnat 50 år åt att arbeta för att se till att ekonomiska framsteg i Europa leder till ökad tillväxt och fler arbetstillfällen och alltid till en garanti för ökad social trygghet.
Allt fler människor anser nu att det motsatta är sant - att Europas ekonomiska framsteg gynnar några få stora konglomerat, vissa försäkringsbolag, hedgefonder och stora företag, men inte folket.
Det är Europeiska unionens uppgift att återupprätta känslan hos dem att tillväxten i Europa och de ekonomiska framstegen på denna kontinent inte gynnar bankerna och de stora konglomeraten utan varje enskild medborgare.
Om nationalstaterna ska garantera detta är dessutom ni som ordförande för Europeiska rådet skyldig att meddela era stats- och regeringschefskolleger att de måste se till att social rättvisa snarare än frimarknadsradikalism blir dominerande i deras nationalstater.
(Applåder)
Jag vill tillägga att vi har en EG-domstol som utfärdar domar varje dag, och dess domar kan ändra graden av social välfärd i de enskilda medlemsstaterna, även om medlemsstaterna inte har några instrument att motsätta sig detta med.
Därför behöver vi ett socialt Europa, herr rådsordförande, och därför förväntar jag mig att ni ändrar åsikt i denna fråga före december.
Annars kommer den socialdemokratiska gruppen i Europaparlamentet inte att kunna stödja er.
Herr rådsordförande! Rädslan för social utestängning leder till en farlig utveckling, bland annat till att regeringar som intar en försvarsställning tror att de kan få människor att glömma denna rädsla för social utestängning genom att förfölja minoriteter.
För närvarande ser vi detta i en EU-medlemsstat.
Jag vet inte hur många procent av den italienska befolkningen som består av romska barn, men jag vet att när en regering säger ”de kommer att registreras på samma sätt som i polisregister, de måste lämna fingeravtryck”, under förevändning att ge dem socialt skydd, är detta ett grovt brott mot EU:s grundläggande rättigheter.
Ert land Frankrike gav den europeiska gemenskapen dess första stadga om de grundläggande rättigheterna.
Den första förklaringen om de mänskliga rättigheterna kom från ert land.
Som president för denna republik är ni en del av ert lands tradition.
Jag vill be er att i er funktion som ordförande för Europeiska rådet påverka Silvio Berlusconis regering och informera den om att EU är en gemenskap grundad på rättsstatsprincipen och inte en union som bygger på nyckfullhet.
(Livliga applåder)
Europeiska unionen står inför många stora utmaningar, men om vi inte garanterar social välfärd i Europa kommer människor att vända sig bort från EU, och när de vänder sig bort kommer vi inte att ha någon användning för Lissabonfördraget. Hela projektet kommer att misslyckas.
Därför måste vi ha mod.
Jag vet att ni är en modig man.
Vi stöder era prioriteringar och vill nu be er stödja våra - ett socialt Europa samt klimatförändringar, institutionell reform och mänskliga rättigheter.
Då kommer ert ordförandeskap att bli framgångsikt.
(Applåder från vänster)
för ALDE-gruppen. - (EN) Herr talman! Jag vill till rådets ordförande säga att det faktum att Irland röstade nej till fördraget har gjort hans noggrant förberedda ordförandeskap mer problematiskt.
Det innebär också att behovet av ett EU som kan handla praktiskt och lösa problem har blivit större än någonsin.
Energi- och klimatpaketen blir mer angelägna för varje dag som går.
Att sätta ett tak för momsen ger kortvarig tröst: EU måste minska sitt beroende av olja och gas.
Vi behöver investera mycket mer i förnybar energi: småskaliga satsningar, avsedda att minska hushållens kostnader, och storskaliga, som att använda oss av unionen för Medelhavsområdet för att investera i produktion av högspänningsel med hjälp av Nordafrikansk solkraft.
G8-länderna - som genererar nästan två tredjedelar av världens koldioxid - godkände i tisdags ett mål om att minska utsläppen med 50 procent.
Men tillväxtekonomierna har rätt i att målet borde vara högre satt - till kanske 80 procent - och innefatta delmål.
För att stabilisera livsmedelspriserna behöver vi goda idéer - som kommissionsledamot Mariann Fischer Boels nyligen genomförda reformer av den gemensamma jordbrukspolitiken - inte protektionism, i vilken form den än visar sig.
Sanningen är den att människor bryr sig mer om priset på bensin och bröd än om gemenskapens storslagna mål.
Numera ska ingen säga ”Qu'ils mangent de la brioche” (”Låt dem äta bakelser”).
Rådsordföranden gör rätt i att sätta fokus på migrationsfrågan.
Men vi kan inte hantera migrationen förrän vi lärt oss hantera den hopplösa situation som får så många att riskera så mycket för att komma hit.
Det behövs lagliga migrationsvägar, kraftåtgärder mot människosmuggling och reformer av jordbrukspolitiken i syfte att få fart på tillväxten i ursprungsländerna.
Det kan tyckas optimistiskt att be ett franskt ordförandeskap att liberalisera marknaderna.
Men för att skapa trygghet inom våra gränser måste vi skapa möjligheter bortom dem.
Det franska ordförandeskapet kan bryta ny mark på ytterligare ett sätt.
Frankrike gav oss mänskliga rättigheter - nu måste Frankrike gå i spetsen för deras försvar.
Hemmavid, genom att driva på arbetet med antidiskrimineringsdirektivet.
Utomlands, genom at förankra fred på Balkan i en gemensam europeisk framtid, genom att utnyttja unionen för Medelhavsområdet för att förbättra de mänskliga rättigheterna i Nordafrika, genom att stå enade i våra förbindelser med Ryssland samt genom att fördöma Kinas övergrepp på oliktänkande.
(FR) Herr rådsordförande! Res inte till Peking.
Var en lagspelare!
(Applåder)
Det var Voltaire som sa att alla människor föds jämlika - det är deras handlingar som skiljer dem åt.
(EN) Och genom att ta initiativet kan EU visa prov på handlingsförmåga och kräva ett erkännande av varje människas värde.
Herr rådsordförande! För att lyckas måste ni söka samförstånd.
Ni måste få parlamentet, rådet och kommissionen att arbeta tillsammans enligt en gemensam dagordning som fastställs av 27 medlemsstater och parlamentet.
Om vi måste tvista ska det vara om denna dagordning, inte om dess budbärare.
Ni har gått i polemik med ECB:s ordförande och med två kommissionsledamöter, men de representerar vår gemenskap och den politik vi enats om.
Det är inte Europas stil att söndra och härska.
Vi måste hålla på våra principer men också arbeta tillsammans för att nå våra gemensamma mål.
(FR) Herr talman! Jag ska snart avsluta, men var snäll och ge mig ”soixante petites secondes pour ma dernière minute” med Carla Brunis make.
(Skratt)
Herr rådsordförande! Om ni håller på era principer och verkligen låter oss arbeta tillsammans för att uppnå gemensamma mål, då kommer vi liberaler och demokrater att samarbeta med er.
(Applåder)
Herr talman, mina damer och herrar!
Som jag sa i Europeiska konventet om det nya fördraget så är det, för att minska avståndet mellan EU och medborgarna, nödvändigt att ge Europa en själ. En själ som respekterar olika språk och identiteter, och som bekräftar våra gemensamma rötter och värderingar - den själ som ni försökt ge uttryck för här i dag, herr rådsordförande.
Strasbourg är en symbol för förnyad fred, och i dag vajar EU-flaggan tillsammans med nationsflaggorna. Den bör vara en synlig symbol för alla medborgare som förenas i vårt gemensamma projekt för försvar, säkerhet och kulturell och ekonomisk tillväxt, och för insyn i centralbanken - kanske saknas det fortfarande i det nya fördraget.
Politikerna måste ge våra ungdomar klara mål.
Den framtida ekonomin kräver att vi respekterar miljön, och respekten för rättigheter kräver att vi erkänner de därmed sammanhängande skyldigheterna.
Vi hoppas att det franska ordförandeskapet i sina mål inkluderar den europeiska stadgan om skyldigheter.
Demokrati och frihet grundas på tillämpning av regler.
Internet får inte utnyttjas för terrorism och barnhandel eller som incitament för våldshandlingar.
Vi måste harmonisera våra länders lagar - från invandring till skydd av minderåriga, från energi till hållbar utveckling.
Ett nytt EU för en ny relation till Afrika.
En relation som inte bara handlar om gröna certifikat och handel utan också om ömsesidig tillväxt i och med samarbetsprojektet mellan Europa och Medelhavsområdet - vi måste vara medvetna om terroristgrupperna i Mogadishu och våldet i Zimbabwe som förhindrar demokratins utveckling.
Man tvekar för mycket inom EU: vi uppmanar rådet att godkänna ”made in”, så att den internationella handeln får tydligare regler.
Kampen mot förfalskning och kriminalitet innebär inte bara en påfrestning på ekonomin utan också på våra medborgares hälsa, och små och medelstora företag har kulturella värden som måste försvaras.
Vi erbjuder det franska ordförandeskapet vårt lojala stöd så att hoppet kan bli verklighet för alla medborgare och vi kanske, genom att bidra till den vetenskapliga utvecklingen i kampen mot sällsynta sjukdomar, också kan bekämpa den endemiska motvilja som vår skarpsinnige vän Martin Schulz känner för premiärminister Silvio Berlusconi.
Herr talman! Denna europeiska voluntarism, dessa höga ambitioner för Europa är en utmaning som vi i gruppen De gröna/Europeiska fria alliansen delar.
Man skulle faktiskt kunna säga, för att parafrasera en sång som ni känner till, ”it is a drug we are all hooked on”.
Det finns dock en sak jag skulle vilja säga.
Om vi den ena stunden ambitiöst säger att vi måste acceptera klimatpaketet som det är, och den andra knäböjer för den tyska bilindustrins lobbyister - då har vi förlorat, eftersom alla andra kommer att kräva liknande behandling.
Häri ligger problemet.
Vi kan inte klaga på att bensinen är för dyr och samtidigt tillåta bilindustrin att tillverka bensinslukande fordon.
Vi har i 15 år vetat hur man tillverkar energisnåla bilar, men eftersom det saknas regler som tvingar tillverkarna att göra det så får nu bilägarna betala det pris bensinen kostar.
Detta är sanningen, det är så det ligger till.
(Applåder från mitten och från vänster)
Ni nämner den europeiska pakten för invandring och asyl.
Så låt oss då bilda en europeisk pakt för invandring och asyl.
Starta en dialog: låt Europarlamentet delta enligt medbeslutandeförfarandet när det gäller laglig invandring - då får vi en genuin politisk debatt, en genuin demokratisk debatt.
Jag har fått nog. Varenda gång vi pratar om utvandring tar det bara 15 sekunder innan vi börjar prata om illegal invandring, om invandring som något hotfullt.
Först och främst: det är tack vare de män och kvinnor som har byggt upp Europa tillsammans med oss som Europa är vad det är i dag.
Detta är sanningen.
(Applåder från mitten och från vänster)
Snälla ni, jag är ingen ängel, men vi har byggt ett hus utan dörrar.
Människor tar sig in via fönstren.
Jag säger så här: låt oss öppna dörrarna så att människor kan komma in i Europa och sedan kan vi besluta vad vi ska göra med dem som tar sig in olagligt.
Ni säger att vi behöver kvalificerad arbetskraft, men samtidigt skickar Europa varje år hem tiotusentals studenter som har kommit hit för att studera.
Låt dem stanna - om de har studerat här är de inte illegala invandrare.
Nu går jag tillbaka till det ni sa om att den sociala dimensionen inte tillhör EU:s ansvarsområde.
Herr rådsordförande! Ni kan inte skydda EU-medborgarna om vi inte tillsammans arbetar för att bekämpa social och skattemässig dumpning.
Nu måste européerna ta sig an det här problemet.
Vi måste få ett slut på det och i detta arbete stöder vi er.
Behöver vi diskutera saken med centralbanken?
Så låt oss då diskutera.
Behöver vi diskutera saken med irländarna?
Så låt oss då diskutera.
Vi måste sluta hävda att den sociala dimensionen inte tillhör EU:s ansvarsområde.
Så kan det inte fortgå.
(Applåder från mitten och från vänster)
Nu skulle jag vilja ta upp de frågor där vi är djupt oeniga.
Ni ska resa till Kina för att tillsammans med den kinesiske presidenten närvara vid invigningen av de olympiska spelen.
Ha det så trevligt!
Själv kommer jag att tänka på alla de fångar som ruttnar bort i kinesiska fängelser.
Jag kommer att tänka på alla dem som har gripits.
Jag kommer att tänka på alla dem som misshandlas i Tibet.
Ni hade ett gyllene tillfälle att försvara europeiska värden som demokrati och frihet genom att säga: ”Jag kommer inte att närvara vid de olympiska spelens invigningsceremoni - denna maskerad som Kinas kommunistiska parti har iscensatt.”
Det är det vi vill höra.
(Applåder från mitten och från vänster)
Jag ska säga er att den dagen ni sitter och skriver era memoarer, då kommer ni att ångra er.
Ni kommer att ångra er därför att de som en gång låste in dessa oskyldiga medborgare kommer att säga till dem: ”Som ni ser kan vi göra vad vi vill - västvärlden är ändå bara ute efter den kinesiska marknaden. ”Det är skamligt och patetiskt att närvara vid de olympiska spelens invigningsceremoni.
(Applåder från mitten och från vänster)
Jag skulle vilja inrikta mitt anförande på att det franska ordförandeskapet är splittrat. Det uppvisar en utan tvekan stark sida och en bara alltför tydlig svag sida.
Ordförandeskapets starka sida är att det, till skillnad från hur det brukar låta i EU-sammanhang, inte hävdar att det går bra för Europa och att vi bör fortsätta på den inslagna vägen, trots att allt fler européer anser att det går dåligt för Europa och vill se en förändring.
Gott och väl - men sedan, då?
Det är just frågan.
Herr rådsordförande!
Vilka slutsatser föranleder denna klarsynthet om unionens nuvarande legitimitetskris, särskilt beträffande dess ekonomiska modell och funktionssätt?
Ni hävdar att ni vill förstå den oro som unionen utlöser hos européerna, och att ni respekterar den. Ändå sätter ni press på irländarna att upphäva sitt beslut, fast de inte gjort något annat än att, i likhet med fransmän och holländare, ge uttryck för tvivel som delas av miljoner européer.
Ni kritiserar med all rätt Europeiska centralbanken för hur den från sitt elfenbenstorn hanterar euron. Men ni aktar er för att ompröva den stadga som ger banken dess enorma befogenheter, bland annat just denna uppgift!
Angående invandringen säger ni att ni vill ”tjäna våra värderingar”. Ändå stödde ni det avskyvärda direktiv som fördömdes av FN:s högkommissarie för mänskliga rättigheter, av samtliga människorättsorganisationer och av de europeiska kyrkorna, just för att det kränker grundläggande mänskliga värden.
Ni struntar i den sociala frågan med argumentet att den är en angelägenhet enbart för medlemsstaterna. Sedan tiger ni när Europeiska gemenskapernas domstol tar artikel 43 och artikel 49 i fördraget till intäkt för att i dom efter dom låta medlemsstaternas olika sociala modeller konkurrera med varandra.
Ni sa att ni ogillade kampanjen om den ”polske rörmokaren”.
Det gjorde jag också.
Det var ett uttryck som högerpopulisterna hittade på och som blev välkänt genom Frits Bolkesteins uttalanden i tv.
För min del välkomnar jag arbetare från alla länder, på jämställda villkor och inom alla yrkesområden.
(Applåder från vänster)
Det är just detta som EU:s lagstiftning i dag förbjuder.
Jag vill påminna er om att det enligt kommissionen går för sig att en arbetare från en annan medlemsstat får hälften av den minimilön som gäller för en tysk arbetare, trots att båda utför samma uppgifter på samma byggarbetsplats i Niedersachsen.
Så vill vi inte ha det.
Europeiska fackliga samorganisationens generalsekreterare John Monks kan knappast beskyllas för att vara populist, och vet ni vad han anser?
Han anser att dessa domar är ”mycket problematiska”, eftersom de enligt hans bedömning föreskriver ”att de ekonomiska friheterna ges företräde framför de grundläggande rättigheterna och respekten för arbetsrätten”.
Hur vill ni svara på det?
Ni hävdar att ni vill bygga ett ”skyddande Europa”, men vi hör er aldrig kritisera de strukturåtgärder som utsätter européerna för risker, till exempel att allmännyttig verksamhet ska konkurrensutsättas, att stabilitetspakten pressar ned löneutveckling och sociala utgifter och de talrika ”riktlinjer” som kommissionen upprättar och rådet antar och som ni tillämpar energiskt i ert hemland.
Jag skulle kunna nämna riktlinje nr 2 om reform av pensions-, socialförsäkrings- och hälso- och sjukvårdssystemen, riktlinje nr 5 om flexibilitet på arbetsmarknaden och riktlinje nr 13 om att undanröja lagstiftningshinder, handelshinder och övriga otillbörliga konkurrenshinder.
Och då har jag inte nämnt dem alla.
Frankrikes och Italiens kovändningar har gjort det möjligt för rådet att gå längre än sina självpåtagna uppgifter. Det har enats om ett förslag till direktiv som tillåter en arbetsvecka på 65 timmar.
Det gör Charles Dickens till Europas nya skyddshelgon!
Nu i helgen talade ni inför era europeiska gäster, med parlamentets talman, kommissionens ordförande och 2 000 franska näringslivsdirektörer från högerkanten som åhörare. Ni avslutade då ert anförande med några ord som fackföreningsrörelsen såg som en tydlig och mycket oklok provokation.
Ni sa att när strejker i dag genomförs i Frankrike lägger invånarna inte ens märke till dem. Dagen efter denna högtidliga tilldragelse förklarade er utbildningsminister att detta var ert sätt att ”lugna våra europeiska partner i ett sammanhang där deras främsta företrädare närvarade”.
Om ni bara kan lugna Europas ledare genom att förolämpa fackföreningarna är det definitivt hög tid för förändring i Europa.
(Applåder från vänster)
Herr president! Tyvärr tvingas Europas invånare att varje dag leva med de katastrofala följderna av den politik som förs av de europeiska myndigheterna i Bryssel och Frankfurt.
Varje dag ser européerna hur alltmer av deras självbestämmande glider dem ur händerna och hur de steg för steg berövas sin frihet, oavsett om det handlar om köpkraften, den höga eurokursen, genmodifierade organismer, skatter, fiskeripolitiken, bristen på handelsskydd, invandringen eller till och med fotbollen, som ni själv nämnde för en liten stund sedan.
Allting glider dem ur händerna. Även er glider allting ur händerna.
Ni säger det ju själv, ni lyfter fram det som något som förtjänar att kritiseras.
Nu är det hög tid för er att handla, att omsätta era uttalanden i handling.
För en stund sedan kritiserade ni med all rätt att gemenskapens inhemska arbetssökande inte ges företräde.
Men låt mig påminna er om att gemenskapsföreträdet upphävdes genom Marrakeshavtalet, som ni godkände, och inte finns med i Lissabonfördraget, som ni upprättade.
Ni beklagar centralbankens oansvarighet och efterlyser en debatt.
För vår del efterlyser vi beslut.
Låt mig påminna er om att centralbankens oberoende, som utgör den oansvarighet vars följder vi kan observera dagligen, infördes och formaliserades genom Maastrichtfördraget.
Ni ångrar att ni fick Bryssel att gå med på att sänka skattesatsen för olja, men det är helt enkelt följden av Nice- och Amsterdamfördragen, som ni lät parlamenten ratificera.
Ni beklagar er alltså dag efter dag över följderna av något som ni ständigt uppmuntrar, det vill säga att statsmakten berövas sin auktoritet till förmån för postdemokratiska organ som utgörs av tjänstemän, bankirer och domare.
EU-ordförandeskapet ger er en historisk chans att få EU på rätt kurs igen, ett EU som grundar sig på nationellt självbestämmande och respekt för demokratin.
Det är därför vi uppmanar er att respektera irländarnas folkomröstning och dödförklara Lissabonfördraget.
Det är inte européerna som ska försonas med Bryssel, utan Bryssel som ska försonas med européerna!
(Applåder från talarens grupp)
(FR) Herr rådsordförande! De närmaste sex månaderna är det ni som ikläder er det rullande och kortvariga ämbetet som Europeiska rådets ordförande.
Ni har, till skillnad från en majoritet av den franska valmanskåren, framträtt som en hängiven Europavän. Ni gick till och med så långt att ni än en gång, nu i form av det föga förändrade Lissabonfördraget, lade fram den konstitution som de holländska och franska medborgarna avvisade 2005.
Nu har era planer tråkigt nog stött på patrull i form av det irländska folkets vilja.
Lissabonfördraget är därmed överspelat, trots alla storslagna planer som det skulle ha tvingat på européerna, och trots de härskande euro-globalistiska potentaternas vilja.
Som ung parlamentsledamot röstade jag 1957 mot Romfördraget, som enligt sina förespråkare Monnet, Coudenhove-Kalergi med flera utgjorde det första steget mot ett Europas förenta stater. Detta Babels torn kan bara uppföras på spillrorna av nationalstaterna.
Det gäller framför allt mitt eget hemland Frankrike. Jag har med kraft bekämpat denna idé ända sedan dess.
Man intalar oss att globaliseringen medför grundläggande förändringar överallt, som vi bara har att finna oss i. Men i själva verket växer sig nationalstaterna i hela världen allt starkare, drivna av en brinnande patriotism.
Det är bara i en region, nämligen Europa, som nationer och hemländer offras, monteras ned och förödmjukas för att främja ett projekt som saknar såväl styrka som identitet. Samtidigt sköljer utländska invandrare in i våg efter våg, och genom att öppna våra ekonomiska gränser utsätter vi oss för stenhård konkurrens från omvärlden.
Många löften har utfärdats till Europas invånare för att de skulle finna sig i att mista sitt oberoende, sitt självbestämmande, sin identitet och sin kultur. Inget av dem har hållits.
Vi har vare sig fått tillväxt, full sysselsättning, välstånd eller säkerhet. Allra mest känner vi oro när vi står vid randen till systemets förestående energi-, livsmedels- och finanskriser.
I går fotbolls-EM och tennis på Roland Garros, i morgon olympiska spelen i Peking. Och i dag den häpnadsväckande historien om Ingrid, kultfiguren som skrattar, gråter, ber och kommer och går, stödd på er broderliga arm!
Er lust att leka befriare fick er att förhandla med terroristerna i FARC, men det var varken ni eller Hugo Chávez som befriade den kolombianska senatorn Ingrid Betancourt.
Det var president Álvaro Uribe som genom sin uthållighet, och stick i stäv med de allmänna progressiva strömningarna i världen, vann en avgörande seger mot dessa brottslingar och terrorister.
Gång på gång gjorde ni misslyckade försök och gick till och med så långt att ni inbjöd ångerfulla kommunistiska FARC-terrorister att resa till Frankrike och söka asyl där. Vem ville ni skydda dem från?
President Uribe - en demokrat?
Varför inte ta steget fullt ut och bjuda in talibanerna, Hizbollah eller de tamilska tigrarna?
Ni är precis som den där tvehövdade draken som Césaire var så förtjust i.
Men en sak ska ni veta, herr rådsordförande: inte ens hela er fallenhet för att domptera medierna räcker för att avvärja de faror som förestår och som ni ställs inför innan året är till ända.
Vårt Europa är ett fartyg som hamnat ur kurs, som misshandlas av vind och våg. Det är den enda region i världen som med berått mod har monterat ned sina politiska och moraliska strukturer, som inte har några gränser och som steg för steg översköljs av en massinvandring som bara är början!
Europa har ruinerats ekonomiskt av ohämmat marknadstänkande, är socialt utfattigt, demografiskt försvagat och saknar vitalitet och försvarsmakt. I bästa fall är Europa dömt att bli ett amerikanskt protektorat, i värsta fall till ett slaveri som liknar dhimmins.
Det är hög tid att vi överger våra ödesdigra illusioner om federalism och bygger ett nationalstaternas Europa, som förenas av mer konkreta allianser - för all del blygsammare, men också mer verksamma.
Att såväl konstitutionen som fördraget gick i stöpet borde kunna tjäna som en varning.
Européerna vill inte ha något att göra med dessa planer, och kommer inte att underkasta sig dem frivilligt, eftersom de inte vill dö.
(Talmannen avbröt talaren)
Mina damer och herrar! Tack för era anföranden.
Låt mig först tacka Joseph Daul, ordförande för gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater, för stödet från honom och hans grupp, som är ovärderligt för det franska ordförandeskapet.
Jag instämmer i era analyser och är säker på att ni förstår om jag inte återkommer till varje enskild punkt i dem, även om ert försvarspolitiska engagemang definitivt är välbehövligt.
Herr Schulz! Låt mig få uttrycka min uppskattning för den ansvarsfulla inställning som ni gav uttryck för i ert anförande.
Vi har träffats, diskuterat och har inga hemligheter för varandra - precis som fallet är med Joseph Daul.
Demokratin får inte bli ett skuggspel.
Den ska låta oss jämföra varandras idéer och sträva efter en kompromiss.
Och precis som i Joseph Dauls fall kan ni vara förvissad om att det franska ordförandeskapet uppskattar stödet från den socialdemokratiska gruppen i Europaparlamentet, och ert stöd i frågan om enhällighet.
Och jag kan inte inse varför detta stöd skulle vara mindre värt för mig därför att det kommer från en gruppordförande som är socialdemokrat - eller varför ni försöker provocera fram konflikter med ordförandeskapet under förevändning att vi har olika politiska uppfattningar?
Låt mig beträffande energi- och klimatpaketet säga att parlamentet självfallet har sista ordet - nu riktar jag även ordet till Joseph Daul. Men bättre upp, det är inte bara en fråga om att få sista ordet.
Det handlar om att mobilisera parlamentet för att sätta press på medlemsstater som inte har samma ambitioner som parlamentet, kommissionen och ordförandeskapet.
Jag skulle inte vilja säga att ni, herr Schulz, får sista ordet, utan att ert engagemang är helt avgörande.
Till Daniel Cohn-Bendit skulle jag vilja säga att det inte handlar om att falla på knä inför någon, särskilt inte inför biltillverkarna, vare sig de nu är franska, italienska eller tyska.
Varför skulle det bara gälla tyska företag?
I detta fall måste rådsordföranden beakta samtliga medlemsstaters legitima intressen.
Vi behöver stå emot branschlobbyn samtidigt som vi ger branschen rimliga arbetsförhållanden och tydligt talar om att vi inte är naiva bara för att vi försvarar energi- och klimatpaketet.
Herr Cohn-Bendit! Jag skulle med andra ord inte vilja anklagas för att främja omlokaliseringar när vår strävan är att uppnå global balans.
Det handlar inte om att respektera miljön och finna sig i omlokaliseringar, utan om att respektera miljön och säga nej till omlokaliseringar.
Att resonera annorlunda är självmordstaktik.
Om ni uppmanar medlemsstaterna att välja mellan miljö och tillväxt hamnar vi i en återvändsgränd.
Hållbar utveckling och respekt för miljön är faktorer som främjar ekonomisk tillväxt.
Och därför tar ni säkert inte illa upp om jag för en gångs skull föredrar Martin Schulz och Joseph Dauls analyser framför er egen.
Herr Schulz! Nu till den punkt där ni anser att vi är oeniga.
Med förlov sagt: jag håller inte med.
Jag vill också tala om för er att det inte är EU:s fel att våra vänner tyskarna inte har lyckats komma överens om en minimilön.
Skyll inte brister i samhället på EU när de beror på den politiska debatten i ett medlemsland!
Här ankommer det inte på mig som rådsordförande att döma någon.
Jag skulle helt enkelt vilja säga: ”Herr Schulz!
Låt mig tillägga att vi fransmän anser att minimilönen är en mycket viktig samhällsfråga.
Vad skulle social harmonisering innebära?
Ni tyskar har avvisat en minimilön.
Vi fransmän vill behålla vår minimilön.
Social harmonisering skulle innebära att vi tvingas avskaffa vår minimilön eftersom tyskarna inte har någon.
Denna sociala tillbakagång vill jag inte ha, inte ens om man vädjar till mina europeiska ideal.
Tack, herr Schulz, för att ni gett mig möjlighet att förtydliga mitt sociala engagemang.
Jag skulle dock vilja tillägga att ni har helt rätt i att vi behöver höja den moraliska ribban för kapitalismen på finansmarknaden och skärpa bestämmelserna för kreditvärderingsföretag. Det är riktigt att vissa finansinstitut handlat på ett sätt som är fullständigt förkastligt.
När vi nu ser hur det har gått för ett antal stora privatbanker vill jag hävda att de som mästrade oss kastade sten i glashus, och nu får räkna med att själva bli måltavlor. Herr Schulz!
Låt mig inför Graham Watsons vakande öga tillägga att jag är emot protektionism och för frihet.
Men vi kan inte fortsätta att leva i en värld utan regler, där kreditvärderingsföretagen gör som de behagar och där ett antal finansinstitut vill tjäna miljardtals euro genom några sekunders aktivitet på börsgolven.
Det Europa som vi eftersträvar - och herr Schulz, det franska ordförandeskapet kommer att lägga fram förslag om det här, förslag till skärpta bestämmelser som höjer den moraliska ribban för kapitalismen på finansmarknaden. Vi inser ju nu att orsaken till att tillväxten i världen har avstannat det senaste året är subprimekrisen och förtroendekrisen för finansinstituten.
De har gjort vad som helst, när som helst, har lånat ut pengar till vem som helst, till vilka villkor som helst. Ett omdömesgillt EU måste avskaffa djungelns lag och någorlunda återställa ordningen.
Jag vill säga till Martin Schulz att jag helt håller med honom.
Beträffande den europeiska pakten för invandring skulle jag vilja svara Martin Schulz och Daniel Cohn-Bendit att det franska ordförandeskapet avser att rådgöra med Europaparlamentet.
Det är bästa sättet att undvika överdrifter.
Herr Schulz, ni nämnde överdrifter i ett land som det inte ankommer på mig att nämna. Om vi alla enas om ett golv för kostnaderna kommer de överdrifter som ni syftade på att upphöra.
Jag är säker på att Joseph Daul håller med mig - varför skulle inte Europaparlamentet vilja medverka till detta? Jag är inte säker på att det går rent institutionellt.
(Inpass av Daniel Cohn-Bendit utan mikrofon)
Herr Cohn-Bendit!
Jag vet att ni är en frikostig person som i regel gärna delar med sig av goda råd, särskilt till mig.
Det här rådet skulle jag inte behöva ens om jag vore lika blygsam som ni.
Jag visste att beslutet erfordrar enhällighet, men det krävs ändå ingen enhällighet för att jag ska kunna säga till Europaparlamentet att invandringsfrågan är tillräckligt viktig för att diskuteras politiskt, och för att parlamentet ska delta i diskussionen, även innan vi har ett Lissabonfördrag eller har ändrat det.
Detta är en politisk utfästelse från min sida. Jag, Bernard Kouchner och Brice Hortefeux kommer att presentera pakten för er och överlägga om den med er.
Vi ska diskutera era önskemål om hur detta bör genomföras med parlamentets talman och kanske med talmanskonferensen.
Herr Watson! I varje svårighet ligger en möjlighet.
Om man väljer att bli ett lands president, och att axla ordförandeskapet i Europeiska rådet under sex månader, och tycker att det är jobbigt med problem eller svårigheter - ja, då är det givetvis bättre att avstå från att vara europé och politiskt aktiv.
För egen del ser jag en möjlighet i dessa svårigheter.
Förstår ni varför?
Därför att de utgör en möjlighet för oss att övervinna vår nationella egoism och våra partipolitiska fördomar.
Med förlov sagt: om allting vore frid och fröjd skulle mitt framträdande inför Europaparlamentet inte nödvändigtvis ha fått ett varmare välkomnande.
Jag tror att det stora flertalet ledamöter av Europaparlamentet i stort sett är medvetna om hur allvarlig situationen är.
Alla måste dra sitt strå till stacken.
Jag är inte så säker på att Martin Schulz eller Daniel Cohn-Bendit hade varit mer vänligt sinnade till det franska ordförandeskapet om läget hade varit ljusare.
Själv ser jag en möjlighet i dessa svårigheter.
Herr Watson! I ett avseende hade jag definitivt fel.
Jag borde ha utvecklat resonemanget om den europeiska energipolitiken.
Ett antal personer här bär särskilda t-tröjor för att signalera att de är emot en viss energiform.
Jag respekterar er, men andra har en annan uppfattning.
Men på en punkt borde vi kunna vara överens, nämligen om att vi behöver en europeisk energipolitik, där vi är öppna med vår lagerhållning och lägger ihop våra resurser i form av solkraft, solceller, energi från biomassa och vattenkraft.
Jag ber om ursäkt för att jag inte sa detta under mitt inledningsanförande, men det franska ordförandeskapet kommer att prioritera utarbetandet av energipolitiken, oavsett våra meningsskiljaktigheter om kärnkraften.
Jag tror inte att kommissionsordförande José Manuel Barroso har något att invända mot detta, eftersom han instämmer i denna prioritering.
Vi har inte råd att dra benen efter oss i den här frågan.
Jag skulle också vilja framhålla för Graham Watson att jag varken är, har varit eller kommer att bli en protektionist.
Men det finns en sak som även liberalerna bör begrunda. Vi har öppnat gränserna och det har gagnat oss.
Men övriga parter kan inte uppmana oss att göra här vad de inte vill att vi gör där.
De stora tillväxtländerna Kina, Indien, Brasilien och Mexiko kan inte komma och säga: ”Öppna era gränser och minska era subventioner, medan vi gör som vi vill.”
Det är inte frihandel och skulle inte heller gagna dem.
Att älska sitt land är inte nationalism, och att eftersträva ömsesidighet och skydd är inte protektionism.
Man kan förespråka frihandel och ändå vilja eftersträva balans i denna frihandel.
Herr Watson, vi kommer att ha mer att diskutera.
Somliga ibland oss betonar skydd, andra betonar frihet.
Vi kanske kan mötas halvvägs.
Slutligen vill jag gratulera er eftersom det verkar som om vi har samma musiksmak.
(Skratt)
Jag ska vidarebefordra era vänliga ord till den person de gäller. Hon kommer utan tvekan att signera sin senaste cd åt er.
Jag hoppas att ni inte tar illa upp.
(Skratt)
Herr Cohn-Bendit! Jag har redan besvarat många av era frågor.
Jag skulle vilja ta upp två saker.
För det första den mycket viktiga utbildningsfrågan.
Givetvis behöver Europa öppna sig för att utbilda eliter från hela världen.
Jag har till och med en längre tid funderat på om inte utbildning av eliter från hela världen innebär att vi bör hälsa dem välkomna till våra universitet och samtidigt ge dem en chans att förvärva sina första yrkeserfarenheter.
Här menar jag särskilt läkare.
Men, herr Cohn-Bendit, vi måste se till att vi inte plundrar utvecklingsländerna på deras eliter.
Ni bör begrunda följande: I Frankrike arbetar fler läkare från Benin än det finns läkare i Benin.
Jag anser att Benin behöver sina eliter.
Att inte vilja plundra utvecklingsländerna på deras eliter är inte detsamma som att stoppa invandring.
Den här diskussionen går inte att slutföra på några få minuter.
Jag uppskattar ert sätt att ta upp det här temat, men ni måste inse att debatten behöver nyanseras och inte kan reduceras till karikatyrer.
Det här handlar inte om att vissa människor är frikostiga medan andra är hjärtlösa.
Vi är politiker som försöker hitta den bästa lösningen.
Tillåt mig att säga en sak om Kina, som är en mycket allvarlig och komplicerad fråga. Herr Cohn-Bendit!
Låt mig säga att jag, i likhet med alla andra här, hörde att ni talade känsloladdat, vilket hedrar er. Låt mig säga att jag delar era känslor.
Ni uppmanade mig att visa samarbetsvilja, och jag skulle vilja påstå att det är precis vad jag har gjort. Som rådsordförande samrådde jag med samtliga medlemsstater för att ta reda på vad de tyckte och om någon invände mot att jag deltog.
Än så länge talar jag om formen, jag återkommer till innehållet om ett ögonblick. Låt mig säga att samtliga medlemsstater höll med om att jag borde delta vid olympiska spelens invigningsceremoni.
Som ni vet så är detta en känslig fråga, och vi bör gå mycket varsamt fram eftersom vi inte har råd att hoppa i galen tunna.
Men Graham Watson uppmanade mig alltså att vara en ”lagspelare”.
Ni ska veta att jag diskuterade saken med samtliga medlemsstater.
Ingen invände mot att jag medverkade. För närvarande ser det ut som om tretton medlemsstater sänder företrädare till invigningsceremonin.
Detta är ju ingen motivering, herr Watson, utan jag bemöter helt enkelt er kritik när det gäller mitt lagspel.
Låt oss nu övergå till själva sakfrågan.
Jag förstår dem som hävdar att européer inte bör närvara vid olympiska spelens invigningsceremoni i Peking.
Var och en har rätt till sin egen uppfattning om hur de mänskliga rättigheterna bäst försvaras, och jag kan bara respektera dem som hävdar att vi bör bojkotta ceremonin.
Men min egen personliga uppfattning är att vi inte kan driva frågan om mänskliga rättigheter vidare genom att förödmjuka Kina, utan bara genom öppen och rak dialog. Detta är en anständig åsikt, och jag hävdar att den bör respekteras.
Jag skulle till och med vilja gå så långt som att säga att vi knappast kan bojkotta en fjärdedel av mänskligheten.
Rådsordföranden har ett ansvarsfullt ämbete men handlar varken klokt eller ansvarsfullt om han säger till en fjärdedel av mänskligheten: ”Vi stannar hemma.
Jag vill resa dit, och jag vill tala med dem.
I huvudfrågan, om försvaret av mänskliga rättigheter, är vi överens.
När det gäller hur dessa mänskliga rättigheter bäst försvaras bör ni finna er i att dessa frågor kan diskuteras och att denna diskussion inte tar slut med de olympiska spelen.
Jag vill därför resa dit för att diskutera och försvara de mänskliga rättigheterna.
Jag kan till och med gå ännu längre, herr Cohn-Bendit.
Vissa saker kommer jag inte att säga till Kina, eftersom Kina förtjänar att bemötas med respekt. Andra saker bör Kina inte säga till de europeiska länderna, och särskilt inte till Frankrike, eftersom Frankrike och länderna i Europa ska respekteras på samma sätt som Kina.
Det är inte kineserna som kontrollerar min kalender eller mitt mötesschema.
På motsvarande sätt är det inte jag som kontrollerar den kinesiske presidentens kalender eller mötesschema.
Jag kommer därför att försvara de mänskliga rättigheterna, samtidigt som jag, som statschef, behöver tänka på en sak.
Vi talar alltid om överenskommelser.
Här har jag invändningar, eftersom det är helt rimligt att en demokratiskt vald statschef försvarar sina medborgares ekonomiska intressen och arbeten.
Jag vill tala om något annat.
Kina är permanent medlem av säkerhetsrådet.
Vi behöver Kinas hjälp för att stoppa skandalen i Darfur, eftersom Kina har stort inflytande i Sudan.
Vi behöver Kina för att kunna isolera Iran, och förhindra att Iran - eller vilka andra aktörer som helst som säger att de tänker få bort Israel från kartan - får tillgång till kärnvapen.
Hur kan vi uppmana Kina att hjälpa oss att åstadkomma fred och stabilitet i världen, om vi bojkottar landet när det står värd för ett arrangemang av oerhörd betydelse för sina 1,3 miljarder invånare?
Det vore varken rimligt eller ansvarsfullt. Det vore inte värdigt en statsmans självrespekt.
(Applåder)
Efter att ha uttryckt min respekt för Daniel Cohn-Bendits uppfattningar och känslor, liksom för alla andra ledamöter som resonerar på samma sätt, skulle jag vilja lägga till följande: Inför resan har jag rådfrågat Graham Watson och den socialdemokratiska gruppens ordförande Martin Schulz.
Vad honom beträffar vågar jag påstå att han helt och hållet håller med om att vi inte bör bojkotta Kina.
Han är socialist - det är inte jag.
Jag rådfrågade Joseph Daul som instämde fullständigt.
Jag skulle vilja avsluta med en annan punkt.
Se hur pragmatiskt Kina har varit beträffande Hongkong.
Detta var ändå en väldigt besvärlig fråga.
För femton år sedan ägde demonstrationer rum i Hongkong, men Kina agerade pragmatiskt för att lösa Hongkongfrågan.
Eller se på Macao: Kina har löst Macaofrågan genom att medverka i överläggningar.
Jag ska gå ännu längre: se på Taiwanfrågan i dag, där president Hu Jintao har gjort stora framsteg.
För fem år sedan trodde alla att en konfrontation mellan Taiwan och Kina var oundviklig. Men så är det inte.
Påverkar vi Kina bäst genom uppriktig, modig och direkt dialog, eller genom förödmjukelser?
Jag väljer dialog, uppriktighet och mod.
(Applåder)
Herr talman! Bara en minut till, som en artighetsgest gentemot Francis Wurtz.
Låt mig lugna honom. Jag förolämpar inte alls fackföreningarna, utan tackar honom för att han understryker att det går att förändra Frankrike utan att förlama det - vilket är vad som sker nu.
Den som hävdar att fackföreningarnas enda funktion är att förlama samhället förolämpar dem.
Fackföreningarna har, precis som politikerna, en roll i den sociala demokratin, varken mer eller mindre.
Vad jag menar här är att ingen har rätt att ta användarna som gisslan.
Jag är säker på att en så belevad person som ni, herr Wurtz, som aldrig har blockerat något ärende, förstår vad jag menar.
Herr Wurtz! I övrigt tycker vi olika, men det hindrar mig inte från att varmt uppskatta det sätt som ni uttrycker er avvikande åsikt på.
Herr de Villiers! Jag önskar att jag hade ännu större förståelse för ert resonemang, med tanke på att ni utan tvekan företräder en politisk maktfaktor såväl i vårt land som i EU.
För att inte rentav säga så här: för min del anser jag att ni inte argumenterar mot EU, utan för att vi ska bygga EU på ett annat sätt.
Jag vill inte ställa förespråkare mot nejsägare, utan försöka finna en plats för alla i ett annat EU som bygger på demokrati, fred och tillväxt.
Jag har tagit till mig era förbehåll, är medveten om dem och ska försöka att reagera på dem med praktiska åtgärder snarare än med ord.
Och vad er beträffar, herr Le Pen: när jag hörde er tala sa jag till mig själv att Frankrike tyvärr i åratal hade Europas mäktigaste extremhöger.
När jag lyssnar till er blir jag väldigt glad över att det är slut på detta nu.
(Livliga applåder)
(EN) Herr talman! Låt mig hälsa rådsordföranden välkommen.
Låt mig först, för den brittiska konservativa delegationens räkning, tacka för er gästfrihet i förra veckan och tillägga att vi ser mycket fram emot att samarbeta med er för att göra ert ordförandeskap framgångsrikt.
Vi är övertygade om att ni är en energisk, engagerad människa, och efter att nyligen ha läst en bra bok är vi också övertygade om att ni är en visionär.
Här syftar jag förstås på er bok Témoignage.
Jag rekommenderar de kollegor som inte haft förmånen att läsa denna intressanta bok att göra det, och särskilt att slå upp sidan 146.
Där beskriver ni 35-timmarsveckans vanvett och alternativets fördelar - ”travailler plus pour gagner plus”, för att citera UMP:s slagord.
Vidare skriver ni: ”Jag tror inte att våra medborgare önskar sig en stelbent 35-timmarsvecka för alla, eller att pensionsgiljotinen avslutar deras arbetsliv när de fyller 60 år.
Där fick ni till det.
Ett sådant Europa är verkligt socialt.
Det är inte regeringarnas sak att tvinga på människor längre eller kortare arbetstid. Regeringarnas uppgift är att skapa förutsättningar för dem som vill arbeta mer att göra det.
Ledstjärnan för ert parti är frihet och valfrihet. Det är också det brittiska konservativa partiets ledstjärna.
Om dessa principer vägleder ert ordförandeskap kommer vi att vara era trogna bundsförvanter.
När arbetstidsdirektivet ses över ska vi kämpa för frihet och valfrihet. Och när direktivet om arbetsvillkor för personal som hyrs ut av bemanningsföretag ses över ska vi också kämpa för frihet och valfrihet.
Låt mig avslutningsvis säga att våra partiers politik inte enbart bör syfta till att öka valfriheten, utan också handla om att respektera invånarnas vilja när dessa väl har gjort sitt fria val.
Jag uppmanar er därför att respektera det irländska folkets vilja, så som den uttrycktes i folkomröstningen nyligen.
Jag uppmanar er att inte se beslutet som ett problem som behöver lösas, utan som en möjlighet för EU att återknyta banden till sina medborgare.
Detta kommer givetvis att kräva en stor arbetsinsats av er och era kollegor i rådet.
Men, som ni själv säger: travailler plus pour gagner plus.
(FR) Herr rådsordförande! Jag är socialist, fransman och europé.
Det betyder att jag inte är en av era anhängare i Paris. Men i Strasbourg räknar jag mig inte helt och hållet till era motståndare, särskilt inte när jag ser två socialdemokrater flankera er.
Min president kanske har fel i vårt hemland, men han förblir ändå min president.
Jag vill därför önska det franska ordförandeskapet, och därmed Europeiska rådets ordförandeskap, lycka till.
Jag har kunnat luta mig tillbaka sedan ni började ert anförande - jag förstår nämligen att ni vill vara i det franska parlamentet.
Jag ser naturligtvis en statschef, men också en ganska frispråkig premiärminister.
När det gäller socialpolitiken och era prioriteringar anser jag att man måste skilja på två saker.
Vissa saker måste förbli nationella uppgifter, exempelvis pensionssystem.
Men när det gäller sådant som den inre marknaden, en gemensam valuta och fri rörlighet, det vill säga alla frågor som påverkar sysselsättningen, måste vårt mål vara att genomföra en harmonisering i linje med bästa praxis.
Vi behöver alltså skilja på dessa saker.
Låt mig tillägga att jag i samband med detta kapitel gärna hade sett att ni gjorde en ordentlig insats för att få till stånd ett ramdirektiv om allmännyttiga tjänster.
Ni gjorde detta för restaurangsektorn, och samma sak behövs också för allmännyttiga tjänster.
Slutligen tror jag inte att EU:s kris enbart är socialt eller demokratiskt betingad.
Den är också, tror jag, en identitetskris.
När freden väl uppnåtts, friheten erövrats och demokratin segrat har omständigheterna i världen gjort det svårt för många av våra medborgare att ta till sig och förstå vad unionens historia egentligen innebär.
Därför är frågor som kultur, utbildning, rörlighet för konstnärer, ungdomar och studenter och vänkontakter av grundläggande betydelse. Vi kan inte längre ta ett europeiskt medvetande för givet.
Men det kommer att växa fram, och jag anser att dessa frågor bör genomsyra det franska ordförandeskapet.
Och avslutningsvis: ni kommer givetvis att dömas efter vad ni har uppnått under era sex månader.
Det har vi fransmän ingenting emot - i Frankrike är, som ni vet, sex månader en lång tid.
I december står resultatet klart.
En sak som vi definitivt kan utgå från är att fördraget inte kommer att ha ratificerats.
Ni vill förenkla fördraget, och situationen är komplicerad. Ni måste ta er ur den!
Låt mig avsluta med några ord som jag lånat av en polsk författare. Låt mig citera: ”Att vara fransman är att se något mer än Frankrike.”
Sådant är vårt rykte, och delvis kanske också ert, herr rådsordförande.
Jag skulle vilja be Cristiana Muscardini uppriktigt om ursäkt. Mitt i den entusiasm som Bernard Poignant var vänlig nog att uppmärksamma glömde jag alldeles bort att svara er och tala om hur mycket vi kommer att behöva er grupp.
Jag vet vilka som ingår i den, och jag vet att ni kan räknas till dem som älskar Europa, och att det finns parlamentsledamöter som älskar sina nationer lika mycket.
Fru Muscardini! Ni kan vara förvissad om att jag kommer att beakta era synpunkter helt och fullt, och att jag de närmaste sex månaderna ska försöka att, tillsammans med de europeiska institutionerna, bygga ett EU som tar hänsyn till era farhågor.
Ni har visat att jag glömmer bort hur överskattad jag är - vilket ger Bernard Poignant rätt.
(FR) Herr talman! För några veckor sedan röstade Irland nej, och jag tror att detta, som vi alla vet, är ett tecken på en växande klyfta mellan medborgarna i Europa.
Vi får naturligtvis inte underskatta detta nej. Tvärtom anser jag att det bör tvinga samtliga ledande politiker att beakta människors förväntningar och oro och försöka hitta ett svar på dem, oavsett vilket fördrag som är i kraft.
Om Lissabonfördraget trädde i kraft i morgon skulle ju inte för den skull alla problem försvinna som genom ett trollslag.
Det franska ordförandeskapet har valt att inrikta sig på fyra områden. Det är naturligtvis konstruktivt, särskilt som ett av dem är klimatförändringen.
Men när krisen nu fördjupas så att vi har en finanskris och en livsmedelskris medan råvarupriserna exploderar och oljan blir allt dyrare och knappare - då tror jag att människorna inte bara förväntar sig problemlösning, utan också visioner. Människorna önskar sig framtidsutsikter.
Det finns tre områden där vi, anser jag, har anledning till eftertanke.
För det första den grundläggande, väsentliga frågan om vår identitet.
Jag anser - jag är övertygad om - att det finns en europeisk modell, ett europeiskt sätt att inrätta samhället.
Den europeiska modellen är ekonomisk, hållbar och social.
Den europeiska modellen försöker exempelvis att göra något åt de växande klyftorna.
Det finns därför en europeisk modell som vi borde vara stolta över, hävda, lyfta fram, föra vidare, försvara och värna.
Detta är det första området.
Så till det andra området för eftertanke.
Jag tror att vi behöver en ny vision för hur vi ska organisera världen.
Här syftar jag framför allt på Afrika.
Jag syftar även på jordbruksprodukterna. Vi bör sluta subventionera exporten av våra jordbruksprodukter och i stället sikta på att Afrika ska bli självförsörjande på livsmedel och energi.
Detta är den nya revolution som behövs för att göra världen rättvisare i framtiden.
(Applåder)
Det handlar om demokrati och mänskliga rättigheter, och det är värden som är lika giltiga för oss i EU som de blir i framtiden i unionen för Medelhavsområdet. Där kommer det inte att handla om att göra affärer och samtidigt bortse från mänskliga rättigheter.
De mänskliga rättigheterna är av grundläggande betydelse de närmaste årtiondena. De utgör Europas innersta väsen, som förtjänar att försvaras.
Detta är några av de utmaningar som jag anser att vi ställs inför. De handlar om grundläggande frågor, det vill säga om vilken vision vi har för Europa och vilken djupare innebörd som vi bör och vill ge Europa.
Detta är inte bara politik, utan samvetsfrågor.
(EN) Herr talman! Jag välkomnar än en gång president Sarkozy till Strasbourg och gläder mig åt att han vill kommunicera med parlamentet och vara uppriktig beträffande sina idéer, även om han var väl medveten om att idéerna inte skulle få medhåll av hela parlamentet.
Alltför länge har gått i de gamla misslyckade ideologiernas fälla, oförmögna att blicka framåt mot de nya gränser som ligger framför oss och möta framtidens utmaningar med öppna ögon.
Vi har spelat säkert genom att bekvämt hålla oss till gamla imperialistiska ideal eller post-fascistiska budord eller till och med - om jag vågar säga det - idéer i fråga om människoliv och mänskliga rättigheter som härrör från början av 1900-talet.
Världen i dag är ju komplex på ett helt annat sätt och så mycket mer varierad än vad en enda ideologi eller en enda plan kan erbjuda.
Ni nämner också med rätta vikten av att kommunicera med andra regeringar runtom i världen: med Kina för att lösa problemen i Tchad och Sudan och se till att problemen med Afrika och utvecklingsländerna hanteras direkt.
Vi hedrar redan i dag minnet av de sju fredsbevarare i Sudan som miste livet under ett FN-uppdrag enbart på grund av att regeringarna inte har klarat av att ingripa på ett riktigt sätt och sätta press på myndigheterna i Tchad och i Sudan för att skydda flyktingars och asylsökandes liv.
Det är ju bra att tala stora ord här i parlamentet om vikten av invandring och fri rörlighet för personer.
Det skulle vara bättre om vi gjorde det möjligt för folk att stanna hemma.
Jag kommer från Irland, en nation som tvingades exportera 12 miljoner av sin befolkning under en tidsrymd på 100 år.
Ingen av dessa ville lämna Irland.
De tvingades lämna landet.
Om vi ger människor möjlighet att stanna i sina hemländer, ger dem stöd genom de politiska mekanismer vi har inrättat, antingen genom handel eller på andra områden, då kan vi göra det.
Slutligen, herr rådsordförande, så talade ni tidigare om att ni kände att legitimiteten i er position när ni lade fram ratificeringen av Lissabonfördraget för parlamentet var det enda sättet att göra det på.
Jag håller med er.
Det är rätt för Frankrike.
Men rätten att hålla en folkomröstning är lika legitim, och den rätten ska alltid värnas.
Det handlar inte om antingen eller.
Det finns problem och svårigheter med resultatet i Irland, men problemen handlar inte bara om Irlands förhållande till EU.
Det återspeglar en allvarligare kris för folket och för EU.
(FR) Herr rådsordförande! Jag vill ta tillfället i akt och fråga vad det franska ordförandeskapet har för inställning i fråga om den språkliga mångfalden.
Mångfald är en av unionens grundprinciper.
Alla världens språk är en del av människans arv och det är de offentliga institutionernas skyldighet att vidta åtgärder för att skydda dem.
(ES) Herr rådsordförande! I rådets slutsatser av den 22 maj om flerspråkighet uppmanades kommissionen att utarbeta förslag till en övergripande ram för en flerspråkighetspolitik, vilket kommissionen har uppgett att den kommer att göra till hösten.
Vilka blir det franska ordförandeskapets ståndpunkter och åtgärder i fråga om flerspråkighetspolitiken?
Vad har ordförandeskapet för inställning och vilken roll kommer det att ge de inofficiella EU-språken, också kallade regionala språk eller minoritetsspråk?
I väntan på omröstningen i den franska senaten nästa vecka är nämligen Frankrike ett riktigt dåligt exempel för alla oss som anser att den språkliga mångfalden är alla européers gemensamma arv.
(Talaren fortsatte sitt anförande på baskiska.)
(EN) Herr talman! Jag vill svara Nicolas Sarkozy.
Ni är en mycket god talare, herr Sarkozy, men jag är inte säker på att ni är en lika god lyssnare.
Det program för ordförandeskapet som ni lade fram i morse visar att ni vill ha en Europeisk union som kontrollerar bokstavligen varje aspekt av våra liv. Här finns allt från en gemensam invandringspolitik till hur vi ska styra våra sjukhus och fotbollsklubbar.
Av era kommentarer framgick också att ni vill isolera oss från resten av världen, att vi inte ska handla med folk som inte har samma standard som vi.
Värst av allt är dock er arrogans när ni påstår att ni vet bäst när det gäller det europeiska projektet.
Ni visar förakt inte bara för det irländska folket, utan också för själva det demokratiska koncept som ni påstår er vara mästare på.
Ni säger att Polens president måste hålla sitt ord, att han måste ratificera fördraget eftersom han gått med på detta.
Nåväl, det irländska folket har talat.
Kommer ni att respektera den irländska folkomröstningen?
Kommer ni att hålla er del av avtalet, som innebär att fördraget är dött?
Jag tror faktiskt inte att ni har förstått.
Europas folk vill inte ha en djupare politisk integration.
Det är därför som fransmännen sa nej, och holländarna sa nej och irländarna sa nej och om vi hade haft en folkomröstning i Storbritannien hade en överväldigande majoritet av oss också sagt nej.
Demokrati till vilket pris, herr Sarkozy? Ni ska till Dublin den 21 juli.
Var snäll och försök inte göra som ni gjorde i Frankrike för att undvika en andra folkomröstning, få dem att ändra reglerna och ratificera fördraget bakvägen.
Det vore att visa ett ytterligt förakt för demokratin.
Var snäll och låt bli.
(FR) Herr talman, herr rådsordförande! För att tillgodose våra och övriga medborgares förväntningar måste rådet, som ni nu är ordförande för, och parlamentet visa en klar, tydlig och konkret politisk vilja.
Ert ordförandeskap är redan det en garant för beslutsamhet.
I detta avseende har vi alla sett, här i Strasbourg och i Bryssel, kvaliteten på förberedelserna inför dessa sex månaders ordförandeskap och hur tillgängliga den franska regeringens medlemmar har visat sig.
De prioriteringar ni lagt fram är de rätta för att bemöta EU-medborgarnas farhågor.
På samma sätt är de övriga utmaningar som ni tog upp, bland annat den ekonomiska styrningen av euroområdet för att hantera den explosionsartade prisökningen på råvaror och kolväteprodukter, eller upprättandet av ett område med stabilitet och välfärd kring Medelhavet, mycket representativa för ert engagemang för en Europeisk union som är mer reaktiv inför problem och mer lyhörd gentemot befolkningen.
När den allmänna opinionen tvivlar och folk ibland ger efter för frestelsen att gå tillbaka till den nationella nivån för att lösa problemen, är det viktigare än någonsin att påpeka att vår kontinent förfogar över stora tillgångar och fortfarande är ett av de sällsynta stabila områdena i en värld som blir alltmer oförutsägbar.
Europeiska unionen bör försöka visa att den inte låter sig globaliseras utan att skydda sitt folk, och jag välkomnar er beslutsamhet att visa detta.
Slutligen hoppas vi att det franska ordförandeskapet, nu när unionen genomgår en betydande förtroendekris, ska kunna få ett slut på de ansträngningar som nu pågått i över femton år för att reformera den utvidgade unionens sätt att fungera.
Lissabonfördraget måste träda i kraft så snart som möjligt, vilket ni också har bekräftat.
Vi förlitar oss alla på att ni ska förhandla med våra irländska vänner och övertyga de få medlemsstater som fortfarande tvekar att ratificera fördraget en gång för alla.
Förra helgen talade ni om att ni inte var beredd att stoppa tillbaka EU-flaggan i fickan, och vi har också sett att ni har hissat den under triumfbågen bredvid den franska.
Vi tolkar denna symboliska gest som bevis för er beslutsamhet att handla i gemenskapens tjänst, och det tackar vi er för.
(EN) Herr talman! Jag vänder mig till rådsordföranden och vill bara påpeka att jag är Rasmussen I, inte att förväxla med Rasmussen II, men jag vill försäkra er om en sak.
Ni talar klokt om det nya Lissabonfördraget, och jag ska säga Nigel Farage att han har glömt fallet Danmark.
Vi röstade nej till Maastricht, men vi röstade ja till Edinburghavtalet och vi skulle aldrig drömma om att säga att vi ska blockera resten av Europa eftersom vi röstade nej i första omgången.
Det skulle vi aldrig säga.
Nigel Farage har fel - det är inte demokrati.
Jag vill bara försäkra er och Frankrike om att vi har hittat lösningen för Danmarks del, och vi kommer att hitta en för det irländska folket också.
Min andra punkt är en vädjan till er från det europeiska socialdemokratiska partiet och alla mina kolleger och ledare och min politiska familj.
Min vädjan är att ni ska lägga till ytterligare en prioritering till era fyra prioriteringar.
Min prioritering - som jag hoppas ni delar, som jag vet att ni delar - gäller jobben, tillväxten, hållbarheten.
Ni sa att vi behöver en bättre reglering av finansmarknaderna, och det gladde mig så att höra.
Jag håller fullständigt med er.
Vi arbetar faktiskt just nu här i parlamentet med ett betänkande och jag hoppas att vi snart kan lägga fram ett klokt betänkande om bättre lagstiftning för det franska ordförandeskapet - här vädjar jag till mina kolleger i PPE-DE-gruppen och ALDE-gruppen.
Jag talar om öppenhet.
Jag talar om bättre lagstiftning i fråga om rättvisa, bonusar och aktieoptioner och allt annat ni talade så klokt om.
Jag talar om ansvarsskyldighet, ansvarstagande, att se till att finansmarknaden är en långsiktig, tålmodig finansieringskraft för våra långsiktiga investeringsbehov för mer och bättre sysselsättning.
I det sammanhanget har jag en annan idé jag vill nämna för er.
Ni har rätt i att vi just nu tappar i tillväxt och sysselsättning, särskilt i Storbritannien och Spanien, men också i Frankrike.
Varför lanserar vi inte ett nytt initiativ för tillväxt, en ny samordnad investeringsåtgärd?
Tänk er följande scenario: om vi investerar bara en procent mer i utbildning, i struktur, i alla relevanta frågor, så kommer vi inom de närmaste fyra åren att få minst 10 miljoner fler jobb än vad vi nu har.
Tänk vad vi skulle kunna göra tillsammans.
Ni sa att idrott är mer än bara marknadsekonomi.
Jag håller med, och vill tillägga att det gäller hela EU.
Europa är mer än bara marknadsekonomi.
Det är arbete och människor.
Låt oss ta hand om dem.
Jag önskar det franska ordförandeskapet all lycka och framgång.
(FR) Herr rådsordförande! Ni sa att Frankrike inte kan döma om irländarnas nej.
(DE) Det håller jag med om.
Irlands nej måste respekteras.
Irländarna är i sin fulla rätt att rösta som de gjort.
Alla EU:s övriga länder är dock i sin fulla rätt att fortsätta på vägen mot ett mer demokratiskt, öppnare och mer handlingskraftigt EU.
Lissabonfördraget är ett steg i den riktningen.
Jag välkomnar därför att ratificeringen fortsätter.
Jag anser emellertid också - och här delar jag inte er ståndpunkt, utan tvärtom - att det vore bra att tala öppet om att vi redan har ett Europa i flera hastigheter.
Tänk på euron, Schengenavtalet, stadgan om de grundläggande rättigheterna och många andra områden.
EU-medlemsstaternas hjärtefrågor och önskemål avspeglas i deras val av olika hastigheter för de projekt de genomför tillsammans.
Europa i flera hastigheter gör det möjligt för de länder som vill göra mer tillsammans att göra det, för det är viktigt att vi slår vakt om principen om frivillighet i Europa.
Det är viktigt att de länder som vill göra saker tillsammans gör det frivilligt och att alla länder har möjlighet att ansluta sig när de vill.
Inget land ska tvingas in i större solidaritet än det önskar.
Europa i flera hastigheter gör det också lättare att fortsätta anslutningsförhandlingarna.
Jag tycker det vore fel att straffa Kroatien och Turkiet för att majoriteten av det irländska folket röstade nej.
Ni är med rätta stolt över att ert land är de mänskliga rättigheternas hemland.
Mänskliga rättigheter är tidlösa, de är universella. Olympiska spelen är ett idrottsevenemang, inte ett politiskt evenemang.
Jag tycker därför det är fel av er att vilja åka till Kina för öppningsceremonin, och jag är glad att Europaparlamentets talman Hans-Gert Pöttering inte kommer att åka till Kina.
Låt mig avslutningsvis nämna att ni på er plats fann en hälsning från många av mina kvinnliga kolleger - en ros och ett brev.
I brevet uppmanas ni att göra ert för att fler kvinnor ska nå toppen i Europeiska unionen.
Kvinnorna fäster sitt hopp vid er som en ”kvinnornas man”.
Låt mig tillägga ytterligare en uppmaning: som demokratiskt vald företrädare hoppas jag att ni kommer att ge oss ert stöd för att se till att detta parlament kan fatta ett självständigt beslut om var det ska vara baserat.
(PL) Herr talman, herr rådsordförande! Jag vill börja med att uppriktigt gratulera er till ordförandeskapet för Europeiska unionen.
Detta blir inte något lätt ordförandeskap.
Det sammanfaller med en svår period, men jag önskar er naturligtvis all framgång.
Irland har förkastat Lissabonfördraget.
Vi kan inte utesluta möjligheten att Irland kommer att ändra sig i framtiden, men det är definitivt inte acceptabelt att försöka påverka irländarna med hot, precis som varken fransmännen eller nederländarna hotades när de avvisade fördraget för tre år sedan och startade dagens problem.
EU-länderna får inte delas upp i bättre och sämre.
Jag vill därför tacka er för era ord att ingen av de 27 medlemsstaterna kan uteslutas från EU-familjen, vilket damen som talade före mig, Silvana Koch-Mehrin, kanske hade velat göra.
Jag vill också ta tillfället i akt och tacka er för att ni nyligen öppnat den franska arbetsmarknaden för bland andra polacker.
Vi har väntat länge på detta - mycket längre än i andra länder, men bättre sent än aldrig.
En sak jag saknade i dagens anförande var någon hänvisning till vår största granne i Europa, Ukraina.
Jag hoppas ändå att det toppmöte som är planerat till den 9 september 2008 i Evian kommer att föra oss betydligt närmare undertecknandet av ett associeringsavtal med Ukraina.
När allt kommer omkring vore en tydlig signal från oss just nu mycket viktig för våra ukrainska vänner, med tanke på det ökande hotet från Ryssland.
På alla de miljontals européers vägnar som för närvarande drabbas av de ständigt ökande priserna vill jag slutligen tacka er, herr rådsordförande, för era ansträngningar att minska mervärdesskatten på bränsle.
Jag hoppas att ni under det franska ordförandeskapet kommer att lyckas vinna över de andra stats- och regeringscheferna för denna tanke, särskilt premiärministern i mitt land Polen.
(DE) Herr talman, mina damer och herrar! Jag vill lyckönska rådets ordförande.
Detta är det 29:e rådsordförandeskapet som jag är med om, och jag kan helt ärligt och förbehållslöst säga att jag aldrig har sett en så övertygande programpresentation och en så europeisk tanke som denna.
(Applåder)
Bara en tidigare rådsordförande har fått ett ännu varmare mottagande, men det var bara vid inledandet.
I slutet av perioden hade han inte levererat någonting på agendan.
Det var den brittiske premiärministern Tony Blair.
Vi är säkra på att ni, president Sarkozy, kommer att avsluta ert ordförandeskap om sex månader med goda resultat.
Ert sätt att förklara allting i dag - ert sätt att svara våra ledamöter, det faktum att ni satt er in i ärendena och att ni inte lägger fram en ”önskelista” utan en rad prioriteringar som backas upp av bra resonemang - allt detta ger mig hopp om att ni faktiskt är kapabel att genomföra ert ambitiösa program.
När det gäller att samarbeta med er för att slutföra klimatpaketet kan ni räkna med parlamentet.
Tyvärr är jag rädd att det är troligare att det blir nya svårigheter med rådet, svårigheter med rådets de enskilda medlemsstaternas ansvar - att de kvoter som planeras inte kommer att godtas där.
Vi håller också med om att kärnenergin måste vara med i klimatpaketet.
Här i parlamentet finns en klar majoritet för civilt utnyttjande av kärnenergi.
Låt er inte förvirras av t-tröjorna.
När det gäller Tysklands och Frankrikes önskan att tillsammans ta över ledarskapet för Europeiska unionen i fråga om innehållet - inte för större deklarationer av världspolitisk art - står vi på er sida.
Jag måste säga att Silvana Koch-Mehrin uppenbarligen inte lyssnade när ni förklarade skälen till ert ställningstagande om Kina.
Det var en lektion i utrikespolitik för parlamentet och jag kan bara uppmana er att förbli lika konsekvent och orubblig i dessa frågor.
(FR) Herr talman, herr rådsordförande, herr kommissionsordförande! Tio nationer producerar 60 procent av de globala koldioxidutsläppen.
Bland dessa tio länder återfinns endast ett europeiskt land - Tyskland.
De 27 EU-medlemsstaterna står för endast 14 procent av de globala utsläppen.
USA står för 17 procent, medan Brasiliens, Rysslands, Indiens och Kinas sammanlagda utsläpp utgör drygt en tredjedel av världens totala koldioxidutsläpp.
Allt detta visar att europeiska initiativ för att bekämpa klimatförändringen fortsätter att vara meningslösa så länge inte motsvarande insatser görs av USA, Kina och övriga industrialiserade länder.
Medan vi väntar på en överenskommelse i denna fråga måste Europa bekämpa koldioxidläckaget.
För närvarande finns det ingen stor industrikoncern som investerar i Europa.
Arcelor Mittal stänger ner i Frankrike, men investerar i Brasilien, Ryssland, Turkiet, Indien och Kina.
Thyssen Krupp investerar i Brasilien, österrikiska Vöest Group investerar i Indien.
I Nordafrika byggs för närvarande tio fabriker som ska producera flytglas för den europeiska marknaden.
Med tanke på att det saknas specifika åtaganden från övriga industriländer måste Europa visa att man är fast besluten att försvara sin industriella struktur, sitt industriella know-how.
Att kräva uppoffringar av EU-medborgarna är meningslöst så länge övriga världen inte gör likadant.
(Applåder)
(FR) Herr talman, herr rådsordförande! Precis som Europaparlamentets talman, precis som många andra parlamentskolleger är jag ett barn av Andra världskrigets ruiner, och jag uppskattar storligen det engagemang som ni på grund av detta visar prov på i ert anförande, som är så befriat från all misstro.
För mig är misstro något som hör ihop med München-andan, och misstro är som en syra som fräter på den europeiska viljan.
Det är därför som jag så starkt uppskattade den energi som ni lade in i ert anförande, som vi, i likhet med vad Astrid Lulling sa i TV nyss, tycker var tydligt och precist, och utan vidare åtbörder vill jag även säga att det var övertygande.
En annan sak jag vill framföra, herr rådsordförande, är att naturligtvis har ni rätt och att detta måste sägas här.
Visst var det främst under Europas uppbyggande under 1950-talet som farhågorna och hoten mot Europa var som störst, men en hel del av dem finns förstås kvar än i dag, även om de har ändrat karaktär.
Det är därför som det behövs en fullkomligt entydig reaktion.
Jag är mycket nöjd med prioriteringarna. Jag säger detta rakt ut, för de är förankrade i verkligheten, i synnerhet den invandringspolitik som er minister Brice Hortefeux, vår f.d. parlamentskollega, har för avsikt att föra.
För två år sedan hade jag äran att företräda Europaparlamentet vid den euroafrikanska konferensen i Rabat.
Där samlades för första gången länder med samma ansvar i invandringsfrågan, oavsett om det var i egenskap av ursprungsland, transitland eller mottagarland, och i likhet med vad Graham Watson sa för en stund sedan anser jag att det är mycket viktigt med en generös närhets- och övervakningspolitik, i synnerhet - ja, varför inte? - via den struktur som unionen för Medelhavsområdet utgör.
Glöm inte att anledningen till Europas unika inflytande världen över är att Europa är en kulturens vagga. För det är i kulturen som våra skillnader befästs.
Kulturen utgör plattformen för våra politiska system, och det är därför som man ser på oss på ett speciellt sätt. Er energi kommer antagligen också att behövas om det ska bli något engagemang även på detta kulturområde.
Först och främst vill jag uttrycka min tillfredsställelse med att Frankrike den 1 juli öppnade sin arbetsmarknad för nya medlemsstater och därigenom undanröjde ett av de sista hindren mellan de gamla och de nya medlemsstaterna.
Jag hoppas bara att förbundskansler Angela Merkel kommer att följa detta exempel.
Frankrike, Tjeckien och Sverige har tillsammans utarbetat ett 18 månader långt rådsordförandeprogram, och jag ser positivt på att man i detta program prioriterar energifrågan, en absolut nyckelfråga, och även reformen av den gemensamma jordbrukspolitiken, eftersom detta rör budgetramen efter 2013 och därmed hur mycket pengar vi kommer att ha tillgång till i framtiden.
Jag förstår att Frankrike vill nå en lösning på dessa aktuella frågor och problem, eftersom det är detta som oroar och intresserar människor.
När det gäller institutionella frågor uttalar jag mig inte i egenskap av medlem av PPE-gruppen, utan som medlem i DE-gruppen, så det kommer förmodligen inte som någon överraskning att vi inte kommer att vara helt överens här.
Vi kan inte bete oss inför Lissabonfördraget likt en hare som får panik i strålkastarljuset.
Det är inte världens undergång, och vi vill inte skapa en krisstämning, så situationen måste lösas lugnt och sansat, utan något politiskt tryck, utan något juridiskt trixande och i enlighet med de regler som vi själva satt upp. Enligt dessa regler kan inget fördrag träda i kraft utan att man först enhälligt har nått en överenskommelse, och någon sådan överenskommelse har vi inte för närvarande.
Jag anser inte att det är omöjligt med en fortsatt utvidgning även utan Lissabonfördraget. Enligt min mening kan åtminstone Kroatien beviljas inträde i EU utan Lissabonfördraget.
På samma sätt anser jag inte att vi måste välja antingen Nice eller Lissabon. Vi har naturligtvis fler alternativ, och vi måste kunna titta på dem lugnt och sansat utan hysteri för att nå fram till en lösning på situationen.
I vilket fall som helst, herr rådsordförande, önskar jag er lycka till när ni nu ska leda Europeiska unionen.
(IT) Herr talman, mina damer och herrar! Vi har följt initiativet Union för Medelhavsområdet, som toppmötet nästa söndag i Paris kommer att fokusera på, och vi hoppas att detta initiativ blir en framgång.
Jag vill dock komma med ett par förtydliganden.
Detta initiativ syftar till att stärka den multilaterala dimensionen i Europa-Medelhavssamarbetet.
Jag anser att detta är rätt, och att det är i denna riktning vi bör gå.
Om det finns en politik som är i behov av en kritisk granskning så är det just relationerna med de sydligare länderna, eftersom grannskapspolitiken snarast skapar konkurrens mellan länder som är mycket splittrade.
Vi måste arbeta för att integrera dessa länder med varandra och för att integrera dem med Europa, och även kanalisera resurser dit.
Jag säger detta rakt ut, herr rådsordförande: Vi uppskattade verkligen inte - och detta säger jag även till kommissionsordförande José Barroso - att ni satte stopp för finansieringen av programmet Euromed Audiovisuel, som utgjorde det enda samproduktionsinstrumentet på kulturområdet.
Ni har sagt att det finns ett europeiskt ”kulturellt undantag”, men jag skulle vilja tillägga, herr rådsordförande, att det finns ett kulturellt undantag även för Europa-Medelhavsområdet.
Av världens tjugo främsta intellektuella kommer flera av de tio främsta av dessa från den muslimska kulturen och ännu fler från Europa-Medelhavsområdet.
Låt oss därför hjälpas åt att vidta effektiva åtgärder så att vi kan förändra livet för många människor i dessa länder, särskilt ungdomar och kvinnor, som sätter sitt hopp till Europa.
Det är inte goda lärjungar vi behöver, utan vi behöver förändra den verklighet som finns bakom denna relation, och parlamentet är redo att samarbeta med ert ordförandeskap om ni väljer att gå framåt i denna riktning.
(ES) Herr talman! Det franska EU-ordförandeskapet har ställt upp realistiska prioriteringar som enligt min mening mycket väl svarar mot det som kommissionens ordförande José Durão Barroso framfört angående kritiken om att EU är kraftlöst och inte klarar av att lösa de dagliga problem som medborgarna ställs inför, dvs. det konstitutionella problemet, livsmedels- och energipriserna, Försvarseuropa och invandringen.
En flykting hittas död i en kylcontainerbil i tunneln under Engelska kanalen, en flykting kastas överbord från en liten öppen båt med kurs på Kanarieöarna - detta hände för bara några timmar sedan, och händelser av detta slag är en av de största tragedierna i vår tid.
Det är ett allvarligt och akut problem, och EU måste agera adekvat.
Ordföranden i gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater, Joseph Daul, talade om behovet av en mobilisering av den politiska viljan, och enligt min mening visar detta rådsordförandeskap ingen som helst brist på politisk vilja.
Men, herr talman, även om det behövs politisk vilja räcker det inte med det: de rådande omständigheterna är också en viktig faktor, och även om de är övergående, kortvariga eller tillfälliga påverkar och begränsar de oss medan de varar, och jag ser positivt på att president Nicolas Sarkozy säger att vi måste se till att omvandla omständigheter till möjligheter.
Jag beklagar att inte Martin Schulz är här just nu, för när han talade om sport kom jag att tänka på en viss speciell omständighet.
Jag önskar att Spanien fick ha den gula tröjan än en gång, precis som i första etappen av Tour de France.
Ni har dock rätt i, herr rådsordförande, att det behövs en europeisk dimension i sportsammanhang, och flera parlamentsledamöter har bett mig framföra en förfrågan till er om ni kunde överväga om de franska idrottare som ska delta i OS (som har varit en diskussionspunkt här i dag) skulle kunna ha EU-emblemet bredvid nationsflaggan på sina dräkter. Sedan kunde övriga medlemsstater själva välja om de också vill delta i ett sådant initiativ.
Herr rådsordförande! Vi hoppas att det franska ordförandeskapet kommer att lyckas mobilisera alla krafter och nå samförståndslösningar, så att, som ni själv uttryckte det, EU kan gå framåt med beslutsamhet under ert ordförandeskap.
(FR) Herr talman, herr rådsordförande! Ni önskade att ledmotivet för ert ordförandeskap skulle vara ”EU som värnar”, och jag tror att förväntningarna nu verkligen är höga bland EU:s medborgare.
Men just därför finns det en motsägelse här - och ni har förstått huvudbudskapet från den socialdemokratiska gruppen i Europaparlamentet - med tanke på att den sociala dimensionen i den europeiska integrationsprocessen inte har getts status som en av ert ordförandeskaps fyra huvudprioriteringar.
Vid de senaste folkomröstningarna tillfrågades människor om EU:s institutioner och fördrag, men svaren de gav baserades på hur framgångsrik den europeiska integrationsprocessen och EU:s politik varit.
Jag tror att det är denna obalans som har uppstått under de senaste åren mellan å ena sidan framstegen i den ekonomiska integrationen - som i sig är något positivt - och stagnationen när det gäller den sociala dimensionen å den andra som också ligger bakom denna besvikelse, detta missnöje gentemot EU-institutionerna som människor inom EU känner.
Problemet är således inte att EU måste vara involverat i alla sociala frågor, utan snarare att så snart det finns en gemensam inre marknad, inklusive en gemensam inre arbetsmarknad, kommer det att behövas gemensamma regler för att bekämpa de skillnader som finns, skillnader som annars leder till social dumpning, och för att se till att konvergenselementen drar oss uppåt, dvs. i riktning mot de bästa förebilderna, istället för att den sociala situationen dras nedåt.
Kommissionen har nyligen offentliggjort en social agenda, men reaktionen på behovet av skydd kommer att utebli om inte rådet tar sig an ett antal konkreta frågor - ni talade ju om ett konkret EU - för att stärka de europeiska företagsrådens befogenheter, skydda tillfälligt anställda arbetstagare, förbättra direktivet om utstationering av arbetstagare så att - och detta måste tilläggas - det finns ett direktiv om skydd av offentliga tjänster och allmännyttiga sociala tjänster.
En av era prioriteringar är invandringspolitiken, som dock inte får reduceras till en ren utvisningspolitik.
Det är därför vi även måste ha en integrationspakt, något som vi talade med Brice Hortefeux om - och en utvecklingspakt.
Ni har just kommit från G8-mötet.
EU och vissa medlemsstater, däribland Frankrike, anklagades för att inte ha uppfyllt sina åtaganden när det gäller offentligt utvecklingsstöd.
Se till att åtagandet att vi ska närma oss 0,7 procent av BNP uppfylls under ert ordförandeskap, ett åtagande som kommer att vara effektivare än det skamliga ”återvändandedirektivet” när det gäller att bidra till en effektivare hantering av den internationella invandringen.
(PL) Herr talman, herr rådsordförande, herr kommissionsordförande!
Jag håller med rådsordförande Nicolas Sarkozy: Det är en svår tid för Europa.
Var och en av oss känner av detta personligen, även jag.
När jag var ansvarig för förhandlingarna i samband med mitt lands anslutning till Europeiska unionen gjorde jag allt som stod i min makt för att säkerställa att det europeiska samarbetet skulle fungera bra i framtiden.
Jag vill även betona att i dag, som tur är, finns det inga problem när det gäller Polens stöd för EU och fördraget.
En betydande majoritet i det polska parlamentet röstade för fördraget, och nästan 80 procent av det polska folket är för EU-medlemskapet.
Jag stöder rådsordförandens bedömning.
Vi måste agera för våra medborgare och på deras vägnar.
Vi politiker måste prioritera energi- och klimatpaketet, men vi måste göra allt vi kan för att se till att genomförandet av detta paket inte slår tillbaka på EU-medborgarna med stora prisökningar och förlorad konkurrenskraft för vår ekonomi.
Detta paket måste antas relativt omgående, men det vore inte bra om man satte snabbhet före ett genomtänkt förslag.
Vårt paket blir beviset på vårt ledarskap i kampen mot den globala uppvärmningen.
Jag håller med om att det är detta vi behöver, först i Poznañ och senare i Köpenhamn, men detta paket kommer inte att fungera som ett föredöme för någon, ingen kommer att följa vårt exempel om den europeiska ekonomin drabbas negativt vid genomförandet.
Jag är därför glad att ni ser dessa risker, herr rådsordförande, och att ni menar att principerna om handel med utsläppsrätter - för det är ju främst det som detta rör sig om - kommer att ses över i en positiv anda.
Erfarenhet har vi.
Reach-förordningen ändrades avsevärt i parlamentet, under medverkan av rådet och kommissionen, till fördel för oss alla.
Den vägen kan vi gå igen.
Herr rådsordförande! Jag vill gratulera till att det nu är ni som håller i tyglarna i EU.
Jag önskar er framgång i de två viktigaste frågorna under de kommande sex månaderna: Fördraget och energi- och klimatpaketet.
(FR) Herr talman, herr rådsordförande! Ni kommer att få ta tjuren vid hornen när det gäller misstron mot Lissabonfördraget.
Frankrike har redan en hel del erfarenhet av konsten att ibland föra den europeiska integrationen framåt, ibland bakåt.
Jag ber er finna en lösning på problemet för Irland, samtidigt som respekten måste upprätthållas för åsikterna hos en överväldigande majoritet européer, eftersom de ju också räknas.
När det gäller sociala frågor vill jag även påpeka att stadgan om de grundläggande rättigheterna och den europeiska sociala modellen ingår i Lissabonfördraget.
Så har t.ex. mer än en miljon underskrifter redan samlats in från funktionshindrade i EU, som utgör vart fjärde hushåll och som är för fördraget eftersom det eliminerar sekulär diskriminering.
Ni har därför stöd för att gå framåt och integrera den sociala modellen.
När det gäller invandringen talade ni till vänstersidan, men ni bör vara medveten om att det är olika vänsterregeringar som för fram idéer som har gjort det möjligt för er att arbeta fram ett mindre slutet och mer progressivt paket, som enligt min mening parlamentet kan förbättra ytterligare, men vi måste fortsätta arbeta ihärdigt med denna fråga.
Dessutom, herr rådsordförande - och detta är direkt kopplat till invandringen: Ni talade om den gemensamma jordbrukspolitiken, men ni nämnde inte Doha.
(IT) Herr talman, herr rådsordförande, mina damer och herrar! I egenskap av ordförande för gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater vill jag uttrycka min tillfredsställelse över att ni har tagit över rodret i Europa, och jag ser positivt på det ni har framfört här.
Ni utstrålar entusiasm och stolthet.
Ni tror själv och får andra att tro på institutionen EU, en institution med många problem och som verkligen är i behov av kloka, upplysta och medvetna ledare, och en sådan har ni visat att ni är.
Italien och Frankrike har alltid haft starka kulturella och sociala band sinsemellan. Båda våra länder har gjort stora uppoffringar för att grunda och bygga Europa, som det nu är alla medlemmars plikt att vidareutveckla.
Var och en av oss som arbetar inom denna institution vet hur många svårigheter vi kan komma att stöta på när vi för utvecklings- och integrationsprocessen framåt, med tanke på att denna process byggs mellan folk med olika historia, kultur, social status och traditioner.
De politiskt sett opportunistiska åsikter som Martin Schulz nyss framförde om den nuvarande mycket populära italienska regeringen hjälper föga.
Men processen måste föras vidare trots de besvikelser som den ibland ger upphov till.
Lissabonfördraget, som är ett utmärkt fördrag, har satts på sparlåga, och det kommer att krävas stor viljekraft för att gjuta nytt liv i det, om vi inte vill stöta bort dem som inte har förstått fördragets innebörd.
Jag håller dock med om det ni sa om att innan det kan bli fråga om någon fortsatt utvidgning måste vi utarbeta nya regler, utan att Irland för den skull lämnas utanför.
Vågen av invandrare som kommer till Europa, särskilt till vissa medlemsstater, och framför allt till mitt hemland och övriga Medelhavsländer, måste regleras och ses som ett gemensamt problem snarare än som en anledning att särskilja eller att rent ut utnyttja situationen genom att straffa de länder som redan fått göra så många uppoffringar.
Vi måste värna om invånarna i våra länder och basera integrationen på en rimlig grund.
Herr rådsordförande! Italiens regering och folk följer ert ordförandeskap med stor uppmärksamhet och tillförsikt, i visshet om att den historia och det sociala anseende som ni representerar här i dag kommer att ingjuta hopp och leda till utveckling i Europa.
(HU) Tre saker - som enda talare från den östra sidan av Berlinmuren.
Jag är besviken över att lika möjligheter inte fanns med i presidentens tal.
Som tur är, herr rådsordförande, har vi kvinnor från de sju politiska partierna noggrant beskrivit vad vi vill i ett brev: det är blomman, det är vår blomma till er, herr president.
För det första välkomnar jag det franska ordförandeskapets insatser på EU-nivå för att skapa social jämställdhet mellan könen. Samtidigt förefaller det motsägelsefullt att de lokala institutioner som arbetar med lika möjligheter läggs ned.
Rekommenderas det någon annan politik på EU-nivå än den som Frankrike tillämpar?
För det andra har presidenten informerat de franska medborgarna om att det kommer att inrättas 350 000 förskoleplatser de närmaste fem åren.
Det är en viktig åtgärd eftersom den ger män och kvinnor lika möjligheter på arbetsmarknaden och en möjlighet att kombinera arbete och familj.
Här är det oerhört viktigt med en förskola av god kvalitet som alla har råd med och tillgång till eftersom det är ett verktyg för lika möjligheter och integration.
När det gäller familjelivet undrar jag om han menar att kvinnor kommer att kunna kombinera arbete och familj om de arbetar 65 timmar i veckan?
Kvinnor är mer utsatta på arbetsplatsen och är i allmänhet inte medlemmar i fackliga organisationer.
Ja, vi behöver en gemensam europeisk invandringspolitik men den måste innehålla en diskussion om medborgarnas och invandrarnas rättigheter och skyldigheter.
Migrationspolitiken måste kompletteras med mottagarlandets integrationspolitik.
Tack så mycket.
(EL) Herr talman! Jag skulle vilja vända mig till rådets ordförande och säga: Jag såg fram emot ert tal i dag med särskilt intresse.
Er ståndpunkt i dag har övertygat mig om att ni kommer att få saker och ting att hända under de sex månader som ni innehar ordförandeskapet.
Hela världen står inför en av de allvarligaste ekonomiska kriserna de senaste årtiondena men EU står också inför sina egna kriser.
Det är uppenbart att EU27 i dag inte kan verka enligt de regler som gällde för EU15.
Det här är den institutionella kris som EU går igenom.
Det är också uppenbart att vissa medlemsstater i dag inte vill ha någon politisk enighet i Europa och inte vill att våra föregångares visioner ska förverkligas.
Det här är en identitetskris.
Den institutionella krisen kommer att lösas men hur ska vi lösa identitetskrisen?
Jag är rädd att det endast finns en lösning. De medlemsstater som vill ha politisk harmonisering bör gå i förväg och de medlemsstater som bara ser EU som en ekonomisk union bör komma efter.
Jag är faktiskt rädd att om vi inte går vidare med den här lösningen kommer EU till slut att upphöra att vara en spelare på det internationella schackbrädet.
Kriser kan leda till stora framsteg men endast om det finns erforderligt mod.
Jag tror att ni har både visioner och mod.
Var modig!
(DE) Herr talman, herr rådsordförande! Er huvudsakliga inriktning har mitt fulla stöd.
Jag tror att ni är rätt rådsordförande vid denna oerhört känsliga tidpunkt, och att ni har den lyhördhet för människors oro och den beslutsamhet att leda och förlika som behövs.
När ni besvarade frågorna vältrade ni inte över ansvaret på någon annan och ni talade rent ut.
Ni vek inte undan utan tog itu med saker och ting.
Jag vill särskilt framhäva ert starka engagemang för parlamentarisk demokrati.
Detta engagemang är särskilt viktigt i dessa tider. I åtskilliga medlemsstater - inklusive mitt hemland, Österrike - har vi upplevt en kamp mellan direkt demokrati och parlamentarisk demokrati, vilket har lett till att parlamenten i parlamentariska demokratier har förlorat mark i EU-frågor.
Låt oss tillsammans stå upp för den parlamentariska demokratin och förhindra att den sätts ur spel.
(Applåder)
Jag tycker också att det är viktigt att ni direkt har tagit upp många regeringars och regeringsmedlemmars feghet eller, det skulle kunna hävdas, dubbelmoral, när det gäller deras gemensamma europeiska ansvar. Denna dubbelmoral är nämligen ett av de främsta skälen till den brist på förtroende och det ömsesidiga fingerpekande som vi måste sätta stopp för.
Vi kräver inte att alla måste bli djärvare men vi kräver att alla är ärliga och principfasta.
Jag skulle vilja gå in på ytterligare tre frågor.
Den första är er ståndpunkt om fördraget.
Ni är inte rädd eller handlingsförlamad, ni väntar inte på Irland utan ni fortsätter ratificeringen samtidigt som ni försöker påverka Irland.
Jag är helt övertygad om att vi inte kommer att hitta en överenskommelse med Irland förrän alla de andra 26 medlemsstaterna har ratificerat fördraget.
Vi får emellertid inte lämna Kroatien åt sitt öde.
Jag välkomnar ert åtagande att inleda förhandlingar om samtliga kapitel före årets slut.
Vi behöver även en tidsplan för Makedonien.
Jag vill be rådet att också fatta ett beslut om en Small Business Act vid toppmötet i december eftersom huvudansvaret ligger hos medlemsstaterna.
Vi behöver juridiskt bindande åtaganden och inte bara ytterligare ett offentligt politiskt uttalande.
(PL) Herr talman! Jag har lite goda nyheter från Polen.
I dag hålls det en debatt i det polska parlamentet som kommer att mynna ut i en resolution som innehåller en uppmaning till den polska presidenten att leva upp till sin konstitutionella skyldighet och underteckna Lissabonfördraget.
Det är det polska folkets vilja. 80 procent av folket stöder EU och är mycket glada över att vara medlem.
Visa mig en annan stat där stödet för EU är så högt.
Det här är en signal om att Polen kommer att fullgöra sina skyldigheter i fråga om fördraget.
Över till någonting annat.
Jag har en uppmaning till er, herr president. Kan ni sätta barnens situation i EU på dagordningen och tillsätta en ombudsman, en advokat i barnfrågor, i stil med Europeiska ombudsmannen för mänskliga rättigheter?
Vi skulle vilja se att rådet kommer överens och godkänner denna institution som EU har ett så stort behov av.
(DE) Herr talman, mina damer och herrar! Om jag skulle summera förmiddagens debatt så skulle jag säga att det är bra att Frankrike innehar ordförandeskapet vid den här tidpunkten och att det är bra att ni, president Nicolas Sarkozy, innehar befattningen som rådets ordförande.
Det har varit en bra dag för EU och för parlamentet. För första gången på länge har vi åter en person framför oss som talar för EU med passion, inte bara med goda argument.
Kanske är det just det som vi behöver för att övertyga irländarna och återfå våra medborgares förtroende: passion och gott omdöme, och gott omdöme innebär också att EU håller sig inom vissa gränser.
Jag skulle vilja ge er receptet på framgång: Vi behöver inte bara fördraget på Irland utan även en ny subsidiaritetskultur.
Vi behöver gränser för EU i förhållande till resten av världen men vi behöver också gränser inom EU.
En ny subsidiaritetskultur kommer att skapa en ny acceptans för EU. Jag håller helt med ordförande José Manuel Barroso om det.
Lycka till, president Nicolas Sarkozy.
(EN) Herr talman! Jag hälsar president Nicolas Sarkozy välkommen till Europaparlamentet.
Jag uppskattade verkligen hans väl övervägda och välformulerade anförande.
Som irländsk ledamot kommer jag också att välkomna honom när han besöker Irland som EU:s ordförande, som en ordförande som vidtar praktiska åtgärder för att förbättra medborgarnas liv.
Det framgick tydligt av hans prioriteringar.
Jag uppskattar även hans synpunkter om livsmedelstrygghet och om att hitta en balans när det gäller att införa förordningar och restriktioner för våra företag och jordbrukare.
Som han själv sa, skydd utan protektionism.
Jag kunde höra hans engagemang för Europa i hans presentation och i hans röst.
Jag och väldigt många irländare delar detta engagemang.
Han talade om att övervinna våra svårigheter.
Det kommer att ta tid och det kommer att krävas en kompromissvilja från alla parter.
Det kan inte sättas några tidsfrister.
Som en person som värvade röster på ja-sidan vet jag att han kommer att hålla med mig när jag säger att ett irländskt nej är precis lika legitimt som ett franskt, nederländskt eller danskt nej.
Det måste behandlas med samma respekt. Sedan kan vi gå vidare.
Vi kan göra framsteg.
Jag ser fram emot det och jag önskar honom lycka till med sitt ordförandeskap.
(FR) Herr talman, herr rådsordförande! Det franska ordförandeskapet har precis presenterat sina mål och jag önskar det all framgång.
Det viktigaste mål som ni har framför er är att stärka EU och dess handlingsförmåga.
Med detta i åtanke vore det en försutten möjlighet att inte ratificera Lissabonfördraget.
EU behöver Frankrike, särskilt i denna svåra tid.
EU behöver det Frankrike som omvändes, av er president Nicolas Sarkozy, efter den franska folkomröstningen.
Det är tyvärr inte Polen som för EU framåt i dag, men en dag kommer det att vara så och jag tror att det kommer att ske snart.
Jag hoppas att det franska ordförandeskapet, med sin politik för europeisk integration, för önskvärd invandring, för utvidgning på Balkan, och inte nödvändigtvis Turkiet, kommer att få européerna att återfå förtroendet och smaken för EU.
(EN) Herr talman! Det tog Irland 700 år att få ut britterna ur Republiken Irland och jag måste sitta här gång på gång och höra de människor som vi slängde ut berätta för oss vad vi bör göra på Irland.
Jag tycker att det är lite väl magstarkt.
Låt det beslut som fattas i Republiken Irland fattas av folket i Republiken Irland.
För det andra vill jag säga följande till Frankrikes president: Om ni vill förändra det irländska folkets åsikt kan ni ju ta Jean-Marie Le Pen med er.
Det skulle räcka för att få det irländska folket att ändra åsikt.
Jag var valgeneral för Fine Gael-partiet, som är en del av Europeiska folkpartiet, i fyra folkomröstningar om EU-frågor: europeiska enhetsakten, Maastrichtfördraget, Amsterdamfördraget och Lissabonfördraget.
Regeringen har suttit vid makten sedan 1994. Politikerna inställer sig i undersökningsdomstolar.
Regeringen och oppositionspartierna - det politiska etablissemanget - ville att det skulle gå igenom. Det fanns en rädsla när det gäller försvar och värnplikt, abort och eutanasi - åtföljt av sprutor som delades ut av ledamöter av parlamentet - skatter, sysselsättning, invandring.
Mycket av detta leddes av höger- och vänsterextremister.
Jag vill bara säga följande till rådets ordförande: Förbered er inför ert besök på Irland.
Om det är viktigt att ni bidrar till att förändra situationen på Irland bör ni vara förberedd när ni kommer och vara beredd att lyssna.
Ni kommer att vara mycket välkommen men det är komplicerat och det kommer att ta tid att lösa denna svåra situation.
(FR) Herr talman! Européerna sätter stora förhoppningar till det franska ordförandeskapet och dessa förhoppningar måste förvaltas väl.
Ordförandeskapet måste undvika att underblåsa orealistiska drömmar och orimlig rädsla, bland annat i grannländerna och kandidatländerna.
När det gäller Lissabonfördraget finns det inte tillräckligt med diplomatisk uppmuntran för en ratificering.
Ordförandeskapet måste hjälpa oss att utarbeta en nödlösning eller säkerhetsstrategi för om saker och ting går fel.
För att undvika det värsta måste vi från början visa att vi är beredda på det värsta.
Jag vill avsluta med ett par ord om det farliga fenomenet med åternationalisering i EU.
Nationalpopulism är det mest oroväckande uttrycket för detta fenomen och det ligger också bakom propagandan för det irländska nejet, den rasistiska främlingsfientligheten i Italien men också retoriken om socialpolitikens nationella karaktär.
Antingen blir EU socialt eller också kommer det att gå under.
Jag hoppas att det franska ordförandeskapet kommer att vara lyhört för den sidan av saken.
Jag är ledsen men jag kan inte ta några fler talare.
Vi har redan dragit långt över tiden.
Jag är mycket tacksam för att president Nicolas Sarkozy och naturligtvis även ordförande José Manuel Barroso har tagit sig tid för oss i dag.
Jag vill därför avsluta med att ge ordet först till ordförande José Manuel Barroso och därefter till president Nicolas Sarkozy.
Jag vill börja med att mycket kort stämma in i de gratulationer som har uttryckts av de allra flesta parlamentsledamöter som har haft ordet. Jag gratulerar till den övertygelse, entusiasm, energi och politiska vilja som president Nicolas Sarkozy har uttryckt här i dag och som jag är övertygad om att han och hans ministrar och kolleger kommer att visa under hela det franska ordförandeskapet.
Jag skulle vilja säga att det här inte alls kommer som någon överraskning för mig.
Jag var fullkomligt övertygad om att det var mycket positivt att Frankrike fick överta ansvaret för ordförandeskapet i rådet under denna särskilt svåra period.
Naturligtvis skulle både vi och president Nicolas Sarkozy ha föredragit om framtiden såg ljusare ut ur institutionell synvinkel. Jag tror emellertid att det är just i dessa svåra tider som vi kan se den politiska handlingskraften och den fulla betydelsen av en stark politisk vilja.
Jag är för den här demokratiska politiska debatten.
Jag har många gånger sagt att vi politiskt behöver erkänna att det finns skillnader och många olika perspektiv, till exempel här i parlamentet.
Vi behöver veta hur vi ska uttrycka dessa skillnader med tanke på att EU skiljer sig från ett nationellt politiskt system.
I våra demokratiska nationella system ifrågasätter vi inte statens legitimitet varje gång vi har en politisk diskussion, inte ens om den ibland är väldigt polariserad. I EU är det emellertid ofta så att när vi som är för EU framför dessa invändningar måste vi konfrontera dem som är emot EU och som försöker ta till all möjlig slags populism för att skada våra institutioner och äventyra det enastående freds- och solidaritetsprojekt som EU-projektet är.
(Applåder)
Därför behöver vi verkligen kunna uttrycka alla dessa åsikter, samtidigt som vi stärker EU-förespråkarna i denna särskilt svåra tid.
Vi ska ha klart för oss att vi har Europaparlamentsvalet i juni 2009.
Om de olika europeiska politiska krafterna och institutionerna inte samarbetar och har en konstruktiv ståndpunkt kommer vi att ge argument åt dem som i sin mest extrema form vill utnyttja populism, främlingsfientlighet och nationalism genom att skapa ett samband mellan nationalism och hemland, vilket är fel.
Vidare citerar jag ofta en stor fransk författare som sa att patriotism är kärlek till det egna folket, nationalism är att hata andra.
Vi kan älska vårt hemland och samtidigt försvara EU-projektet med övertygelse, som president Nicolas Sarkozy precis sa.
Jag hoppas därför att den debatt som kommer att föras under de kommande sex månaderna kommer att stärka EU:s institutioner och vårt projekt för EU:s framtid.
Jag vill gärna besvara en specifik fråga.
Det är den enda specifika fråga som ställdes och jag kommer naturligtvis att lämna resten till president Nicolas Sarkozy som är bättre lämpad att ta itu med dem än jag.
Denna specifika fråga kom från Pasqualina Napoletano angående Euromeds kulturprogram.
Det gläder mig att kunna informera er om att det nuvarande programmet, Euromeds kulturprogram, fortfarande har 15 miljoner euro i anslag för i år.
Det stämmer att ingenting är beslutat ännu för 2009-2010. Det finns dock ett ganska hårt tryck på externa utgifter och det som händer i det fallet är, uppriktigt sagt, att berörda tredjeländer tenderar att prioritera bilateralt samarbete, vilket går ut över de regionala budgetarna.
Det är därför en fråga som bör diskuteras med Euromedländerna.
En av de intressanta aspekterna av det franska initiativet för att skapa en union för Medelhavsområdet - som jag för den delen stod bakom från allra första början - är att det innebär ett ökat regionalt samarbete.
Ibland undrar människor vad unionen för Medelhavsområdet tillför Barcelonaprocessen.
Den tillför naturligtvis ökat politiskt inflytande, och även en uppvärdering av politiken, särskilt tack vare det toppmöte som hålls vartannat år.
Den tillför emellertid också den dimension som tillkommit genom specifika regionala projekt och jag hoppas också genom mycket specifika projekt där vi kan låta den privata sektorn spela en mer framträdande roll, eftersom vi fortfarande behöver mer resurser.
Det här är alltså det specifika område som vi arbetar med. Avslutningsvis vill jag bara säga följande: ”Lycka till Frankrike, och lycka till min käre vän, president Nicolas Sarkozy!”.
(Applåder)
Jag vill tacka ordförande José Manuel Barroso och vice ordförande Jacques Barrot för att de har varit här i tre timmar utan avbrott.
Jag vill börja med att säga att jag tycker att det är naturligt när man har äran att vara rådets ordförande att vara i parlamentet under så många timmar som parlamentet önskar, inte bara under ordförandeskapets första dag. Jag vill snarare säga er, herr talman för Europaparlamentet, liksom alla gruppordförandena och talmanskonferensen, att jag står till ert förfogande om ni vill att jag ska komma vid vissa tillfällen under ordförandeskapet.
Man måste spela EU-institutionernas spel.
Europaparlamentet är hjärtat i den parlamentariska demokratin.
Det är inte en fråga om tillgänglighet. Det är en fråga om prioritering.
Ordförandeskapet behöver Europaparlamentet och står därför till dess förfogande.
(Applåder)
Om talarna ursäktar vill jag säga ett par ord till var och en av dem.
Först av allt vill jag säga till Philip Bushill-Matthews att jag hör till dem som anser att EU behöver Storbritannien.
Jag har aldrig hört till de européer eller fransmän som har tyckt att vi borde vara på vår vakt mot våra brittiska vänner.
Storbritannien kan tillföra mycket mer till EU än det tror att det kan.
Storbritannien är nyckeln till den anglosaxiska världen. Det representerar det ledande språket i världen och det har en dynamisk ekonomi, vilket har visat sig på senare år.
Jag vill säga följande till våra brittiska konservativa vänner: ”Ni måste tro på att EU behöver er, på att ni har en plats där, och på att EU skulle bli svagare om britterna hade en fot i och en fot utanför EU”.
Storbritannien är en storslagen nation.
Den har ingenting att frukta av EU och EU har en hel del att förvänta sig av Storbritannien.
Till Bernard Poignant, som såg djupt in i mig och därför förstod att jag älskade politik och att parlamentet var lite som min trädgård, vill jag säga att ja, parlamentet är demokratins kärna och jag respekterar och förstår inte de politiska ledare som inte skulle vilja uttrycka och försvara sina idéer i den parlamentariska demokratins vagga.
Jag hoppas att det i er kommentar fanns ett uns av beklagande, snarare än en ytterlig åsikt om harmoniseringen av arbetsmarknaden.
Detsamma gäller även Harlem Désir. Jag håller med er helt och hållet.
Jag är emot en fullständig harmonisering eftersom folket skulle förkasta det. Det är emellertid helt naturligt att ha minimiregler på en arbetsmarknad, på en inre ekonomisk marknad.
Vi bör alla vara medvetna om svårigheterna.
Ta till exempel Österrike, som har en socialdemokratisk förbundskansler och regering. De kommer att säga er att pensionsåldern är 65 år och att avgiftsperioden är 45 år.
Ni vet vilka problem jag stötte på när jag försökte införa en avgiftsperiod på 40 år och jag fick inte något omedelbart stöd från det franska socialdemokratiska partiet.
Så förklara för mig hur det kommer sig att jag, när jag stötte på så stora problem när jag införde en avgiftsperiod på 40 år i Frankrike, bara behöver vara EU:s ordförande i sex månader för att helst åstadkomma en avgiftsperiod på mellan 45 år i Österrike och 40 år i Frankrike.
Hur ska det gå till?
Det är långt mellan dröm och verklighet men det är kanske det som är skillnaden mellan det franska socialdemokratiska partiet och Europeiska socialdemokratiska partiet.
Ibland känner jag att jag till och med står närmare Europeiska socialdemokratiska partiet än det franska socialdemokratiska partiet.
Jag medger denna brist och ber om ursäkt för den.
(Martin Schulz avbröt talaren utan mikrofon)
Det fungerar inte så.
Det är inte upp till er att avgöra vem som talar.
Talartiden kan inte delas mellan den socialdemokratiska gruppen i Europaparlamentet och rådets ordförande.
President Nicolas Sarkozy! Är ni beredd att låta Martin Schulz ställa en fråga?
Om ni är det så ska jag ge honom ordet.
rådets ordförande. - (FR) Herr talman! Ja, förutsatt att jag inte hamnar mitt i korselden i en heltysk debatt.
(DE) Tack så mycket, herr talman, det var mycket vänligt av er.
President Nicolas Sarkozy! Det är trevligt att ni vill närma er socialdemokratin på det här sättet.
Efter att ni i ert tal alldeles nyss ställt er bakom de tyska socialdemokraternas ståndpunkt och därmed distanserat er från förbundskansler Angela Merkel föreslår jag att ni gör enligt följande.
Om ni känner er så bekväm inom den europeiska socialdemokratiska församlingen tycker jag att ni först ska ansluta er till den tyska socialdemokratin så ska vi gradvis föra er närmare den franska socialdemokratin och så kommer ni att bli en riktigt god kamrat till slut.
Herr Schulz! Det här har inte så mycket att göra med vänlighet som med att följa reglerna - någonting som vi i EU när allt kommer omkring vill göra.
rådets ordförande. - (FR) Herr talman! Som ni kommer att märka har jag redan en socialdemokrat till höger om mig men det finns plats för en socialdemokrat till vänster om mig.
(Applåder)
Mina damer och herrar! Som ni vet tycker jag inte att vi slösar bort någon tid eftersom jag anser att demokrati på EU-nivå kan vara fri från det våld som ibland finns på nationell nivå.
På EU-nivån kan alla ta ett steg tillbaka från valförfarandet, som är brutalt, ofta orättvist och alltid svårt.
Slutligen kan man i ett forum som ert tala och samtidigt le och respektera varandra, vilket kanske också är någonting som kommer att få människor att bli vänligare inställda till det europeiska idealet och göra det till sitt eget.
I vilket fall som helst ser jag det inte som slöseri med tid och jag vill försäkra Bernard Poignant och Martin Schulz om detta.
Mariell De Sarnez har helt rätt.
Vi måste ändra vår utvecklingspolitik och prioritera livsmedel och jordbruk.
Det är absolut nödvändigt. De afrikanska länderna måste ha resurser för att bli självförsörjande på livsmedel och delar av de pengar som vi har anslagit för att utveckla stora infrastrukturer måste säkerligen investeras i mikroprojekt inom jordbruket.
På den punkten delar jag er åsikt helt och hållet.
Ni uppmanade mig också att försvara en vision om Europa.
Jag delar den ambitionen.
Jag hoppas att ni kommer att vara generös nog att vägleda mig om vad denna vision ska innehålla.
Som ni mycket väl vet är vårt problem återigen att någonstans mellan det något avknoppade stora idealet och alla tekniska problem i vardagen ständigt behöva avgöra vad vi ska göra med de stora idéerna, som ibland är mycket större än de dagliga svårigheter som våra medborgare möter i sin vardag, och vad vi ska göra för att lösa de tekniska problem som påverkar deras vardag.
Det är inte så enkelt men jag ska i alla fall göra ett försök.
För att svara er, herr Crowley, så stämmer det att vi behöver utveckling för att undvika olaglig invandring.
Vidare är alla medvetna om att utveckling är det bästa sättet att ta itu med invandringsfrågan.
Det finns 475 miljoner unga afrikaner under 17 år och det är 12 km av Gibraltar sund som skiljer Europa och Afrika åt.
Afrikas katastrofer kommer att bli Europas katastrofer och det finns inga hinder eller gränser som kommer att kunna stå emot det.
Vi behöver därför verkligen en utvecklingspolitik.
Återigen är det mycket svårt att välja mellan multilateralism och bilateralism.
Det här är en viktig fråga och jag avser att ägna en hel del uppmärksamhet åt den.
Mikel Irujo Amezaga talade om den språkliga mångfalden.
Jag håller med honom fullständigt, bland annat när det gäller de officiella språken - och jag förstår att ni inte tycker om uttrycket ”regionalt språk”.
Ni förstår att jag hör till dem som anser att vi skulle hjälpa alla rörelserna för självständighet och oberoende om vi gav dem monopol på att försvara de regionala språken och det vore ett mycket allvarligt misstag.
Jag talar om Korsika i Republiken Frankrike, där det finns människor som är korsikaner, som älskar Korsika och som talar korsikanska i byarna, men det utgör inte något hot mot den nationella enigheten.
Därför är den språkliga mångfalden i mina ögon precis lika viktig som den kulturella mångfalden och det kommer i vilket fall som helst inte att bli någon kulturell mångfald om det bara finns ett språk.
Herr Farage! Jag tyckte mycket om ert anförande men jag ska säga er en sak: Britterna var glada över att jag lade ned Sangatte, för det var faktiskt jag som lade ned Sangatte, och det var ni som bad mig att göra det.
Även om man är britt och älskar sitt land kan man inte lösa landets alla invandringsproblem och jag måste säga er att Frankrike inte tänker bli Storbritanniens gränsvakt.
Låt mig säga att det är en sak att säga att ”i mitt land vill jag inte ha id-kort eller en gemensam invandringspolitik”. Det hindrar er dock inte från att vara glad över att invandrare som inte har sina papper i ordning stoppas i Frankrike så att ni inte behöver ha dem i Storbritannien.
Precis som Frankrike kan Storbritannien inte klara det på egen hand.
Jag vill tillägga att jag respekterar polackerna. Ni stod dock inte på mitt kontor och förhandlade om Lissabonfördraget med ett antal kolleger.
Vi var i Bryssel och vem var på mitt kontor?
Inte premiärminister Donald Tusk, för premiärministern vid den tiden var Jarosław Kaczynskis bror.
President Lech Aleksander Kaczynski var där och jag ska säga en sak. Det är en man som jag litar på och det är en man som jag respekterar.
Om man undertecknar någonting i Europa och börjar med att inte respektera det finns det emellertid inte något Europa kvar, ingenting alls, inga förhandlingar.
När någon av oss gör åtaganden för sitt lands räkning i Bryssel måste denne göra åtaganden även på hemmaplan.
Det var det jag sa, varken mer eller mindre.
(Applåder)
Detta är med full respekt för Polen. Herr Farage!
Jag anser att jag försvarade Polen. Ordförande José Manuel Barroso kommer att kunna säga detta bättre än någon annan.
Vi behöver Polen men vi måste även ha respekt för en persons ord.
Fru Sudre! Tack för ert stöd.
Jag håller helt och hållet med om er analys och jag tackar er uppriktigt för den.
Herr Rasmussen, som jag förstod var Rasmussen I, och jag är nästan på det klara med vem Rasmussen II är! Jag vill säga att Danmark är ett bra exempel på ett land som har lyckats göra framsteg och det innebär att jag kan svara alla talare om Irland.
Vi bör naturligtvis inte tvinga irländarna och vi måste respektera dem men vi måste ha modet att säga till våra irländska vänner: ”Ni måste också respektera de andra länderna som har ratificerat fördraget.
Vi läxar inte upp er men tänk på att andra också har en åsikt och att vi någon gång måste hitta en gemensam väg.
EU vill inte fortsätta utan er men EU kan inte stanna av bara på grund av er.”
Jag säger det med alla den respekt jag har för ett land som har röstat nej.
Vi, fransmännen, har ställt till med stora problem och svårigheter för er. Någonstans måste vi dock ta oss ur den här situationen, där alla tittar på varandra och väntar på att någon annan ska ta initiativet.
Det franska ordförandeskapet, tillsammans med ordförandeskapet för kommissionen och Europaparlamentet måste ta initiativet. Därefter kommer vissa att säga ja och andra säga nej.
Personligen tror jag att det finns en lösning.
Den handlar dock verkligen inte om att låta saker och ting vara som de är eller om att säga att ”vi får vänta och låta tiden göra sitt”.
Personligen tycker jag att vi har tiden emot oss, att EU har väntat i åratal och att det inte är någon idé att vänta längre.
Jag är övertygad om att vi kommer att hitta en lösning, precis som danskarna gjorde.
Fru Koch-Mehrin! Jag blev mycket rörd över er bedömning av mig som en ”fruntimmerskarl”.
Jag kommer att låta er stå för innebörden. Jag vet ärligt talat inte exakt vad det innebär och jag kommer att vara noga med att inte att ge mig in på det spåret eftersom jag inte vill att ni ska missförstå mig.
Jag vet att vi har ett Europa i flera hastigheter.
Vi är inte alla med i eurosamarbetet och vi är inte alla med i Schengen.
I slutändan vill jag dock att vi, innan vi bygger ett institutionellt Europa i flera hastigheter, försöker att göra det hela tillsammans.
Kritisera inte ordförandeskapet för sin ambition att få alla med sig. Om vi innan vi ens hade börjat hade sagt ”det spelar ändå ingen roll, vi låter det vara” så skulle vi ena dagen förhandla om ett socialt undantag för britterna, nästa dag förhandla om ett institutionellt undantag för irländarna och nästa dag förhandla om ett undantag för polackerna.
Då är jag rädd att vi kommer att hamna i en situation där alla länderna, med rätta, kommer att be om ett undantag och vad kommer det att bli av EU då?
Var kommer det projekt som grundarna lanserade vara då?
Det är det jag menar.
Kanske kommer vi att hamna där ändå. Jag vill dock att vi hamnar där efter att ha försökt att få med oss hela familjen.
Jag vill också säga till dem som är oroade över Kroatien att jag naturligtvis är för fortsatta förhandlingar. Jag anser att det vore ett allvarligt misstag att stänga EU:s dörr mot Balkan, eftersom Balkan behöver den fred och demokrati som EU kan ge dem.
Jag skulle vilja säga till Adam Bielan att jag inte vill hota Irland. Dessutom skulle jag inte kunna göra det och det skulle inte heller falla mig in att göra det.
Samtidigt måste alla inse att i opinionsmätningarna säger 80 procent av folket att de är för EU. Vi kan ändå arbeta med dem utan att hota dem.
Momsen på bränsle är ett franskt förslag. Jag vill inte tvinga det på någon.
Jag vill bara göra er uppmärksamma på att jag är övertygad om att priset på olja kommer att fortsätta att öka.
Vi måste ha modet att säga det till våra medborgare.
Oljeproduktionen minskar med 3 procent varje år på grund att tillgångarna sinar. Samtidigt ökar oljeförbrukningen med 2-3 procent på grund av tillväxten i de framväxande ekonomierna.
Jag menar helt enkelt att momsen är en skatt som står i proportion till priset.
Om oljan imorgon kostar 175 dollar per fat kommer vi, utan att säga någonting, att kunna fortsätta att ta ut 20 procent skatt på kraftigt stigande oljepriser?
Det är den frågan som jag vill ställa.
Vi kommer tillsammans med kommissionens ordförande att rapportera om detta i oktober.
Jag kommer att försöka styra det hela enligt min övertygelse och så får vi se vad resultatet blir.
När det gäller Ukraina kommer det att hållas ett toppmöte och vi kommer att göra framsteg.
Vi behöver uppmuntra Ukraina att gå mot demokrati och vi behöver föra landet närmare EU.
Ukraina är inte betydelselöst. Det har 42 miljoner invånare.
Det är inte något litet beslut.
Just nu står vi inför en associering men alla som promenerar genom Kievs gator kan se att det är en europeisk huvudstad.
Herr Langen! Jag vill tacka er för era komplimanger, som verkligen berörde mig.
Jag gillade faktiskt hänvisningen till Tony Blair.
Jag vet inte om det är därför som ni gjorde hänvisningen men jag tycker att Tony Blair är en av de statsmän som har gjort en hel del för EU och en hel del för sitt land. Uppriktigt sagt vet jag inte om han skulle ha någonting emot att jag säger det men på många områden tycker jag att han har återskapat tilltron och styrkan i den brittiska politiska debatten och i den europeiska politiska debatten.
Jag tycker att vi i Europa behöver ledare och att Tony Blair under sin tid obestridligen var en sådan ledare.
Det här kommer att ge er intrycket av att jag är mer vänsterinriktad, även om jag har lagt märke till att Tony Blair inte alltid får komplimanger från den sidan av det politiska spektrumet.
Herr Goebbels! Ja, andra måste göra en insats, och det är precis den fråga som kommer att tas upp under förhandlingarna om klimatförändringen, men Europa måste föregå med gott exempel.
Jag är inte naiv för att jag säger det.
Jag tycker att vi har mer trovärdighet när vi lever som vi lär.
Vissa kanske säger att det är bättre att vänta.
Jag tycker personligen att vi måste ta risken att handla.
Herr Goebbels! I grund och botten är min politiska filosofi att det inte finns någonting värre än passivitet.
Den värsta risken är att inte ta några risker.
Herr Cavada! Ni har helt rätt.
Vi behöver ta itu med denna rädsla. Tack för ert stöd.
När det gäller unionen för Medelhavsområdet skulle jag, för att ta vid efter ordförande José Manuel Barroso, vilja säga att jag inte har någon kritik mot Barcelonaprocessen.
Jag vill trots det säga en sak.
Barcelona var en mycket god idé men det fanns ett problem vid toppmötet i Barcelona.
Så vitt jag minns så var det bara en arabisk statschef där, premiärminister Abu Mazen.
Hur tror ni att vi ska kunna skapa en union för Medelhavsområdet, som går ut på att föra nord- och sydkusten närmare varandra, om sydkusten in kommer?
Vid toppmötet i Paris tror jag, även om Bernard Kouchner kanske kommer att rätta mig senare, att samtliga arabiska statschefer kommer att närvara.
Det kanske inte spelar så stor roll men för mig är det helt avgörande.
Jag vill också säga till Jan Zahradil att det inte är en fråga om att skapa en kris om Lissabon men att vi inte heller bör agera som om ingenting har hänt.
Vi bör inte vara överdramatiska men samtidigt är det ändå oroande att de senaste tre folkomröstningarna i EU slutade med ett nej. Det berodde visserligen på andra saker men faktum kvarstår att det åtminstone inte är ett särskilt uppmuntrande tecken.
Jag tänker inte svara er, fru Napoletano, eftersom ordförande José Manuel Barroso gav er ett bra svar.
Herr Sánchez-Neyra! Ja, idrotten behöver en europeisk dimension och jag tycker att det bara vore bra om OS-statistiken räknades nation för nation men att det fanns en särskild kolumn för europeiska medaljer.
Det vore ett sätt att visa att vi även finns i idrottens Europa.
Herr Désir! Jag svarade er när det gäller standarderna på arbetsmarknaden.
När det gäller socialpolitiken har vi en berömd debatt.
35 timmars arbetsvecka är inte tillräckligt för att vinna valet, eller för att få en ordentlig socialpolitik.
Jag skulle vilja tillägga att skälet till varför jag gjorde mig så mycket besvär för att övervinna de automatiska, stela reglerna för 35 timmars arbetsvecka i Frankrike var just för den europeiska harmoniseringens skull, för att inget annat land hade följt efter er i den frågan.
Inget.
Inte ett enda.
Inte ens i de europeiska socialdemokratiska regeringarna.
Därför är jag som ni förstår glad över att vi uppmanar till social harmonisering. Jag skulle dock vilja säga till våra franska socialdemokratiska vänner att social harmonisering handlar om att inte förespråka idéer i Frankrike som ingen annan förespråkar i Europa, för det är ett undantag och vårt land drabbas därför av det.
Jag vill tacka Jerzy Buzek för Polens engagemang i EU.
Jag har aldrig någonsin tvivlat på Polens engagemang i EU.
Polen är ett av de sex befolkningsrikaste länderna i Europa och det är just därför som jag säger till president Lech Aleksander Kaczynskis att vi behöver hans underskrift, för Polen är inte vilket europeiskt land som helst.
Det är oerhört viktigt, det är en symbol, och naturligtvis måste vi minska den institutionella krisen till att bara handla om Irland.
Herr Barón Crespo! Doha, ja jag sa det till ordförande José Manuel Barroso, jag sa det till Gordon Brown, men kort sagt, Doha, dock inte till vilket pris som helst.
Jag skulle vilja försvara två idéer som ligger mig varmt om hjärtat.
För det första sägs det att utan överenskommelse blir det ingen tillväxt.
Ursäkta mig, men det har inte funnits någon överenskommelse på sju år, och i sex år har världen haft en exempellös tillväxt.
WTO-överenskommelsen är att föredra framför att inte ha någon överenskommelse. Därmed inte sagt att det inte kan bli någon tillväxt utan överenskommelse.
Vi har haft tillväxt i sex år.
För det andra säger ordförande José Manuel Barroso, den kanadensiska premiärministern och till och med Angela Merkel för närvarande att det inte är bra nog.
Brasilien gör inte någon insats för att sänka tullhindren i industrin. Det gör inte några insatser när det gäller tjänster.
Vad kan man säga om stängningen av den kinesiska marknaden?
Det finns inte något franskt undantag ur det perspektivet.
För det första måste jag, som rådets ordförande, lojalt försvara unionens ståndpunkt.
När det gäller unionens ståndpunkt har jag emellertid inte hört någon, inte ens den brittiska regeringen, säga att överenskommelsen borde undertecknas i det nuvarande skedet i förhandlingarna.
Vi är därför helt överens i Europa, även om det inte är av samma skäl, när vi säger att det inte är bra nog som saker och ting ser ut.
Europa har gjort hela jobbet och kan inte fortsätta göra insatser om de andra stora regionerna i världen inte är engagerade i att göra framsteg.
Ur det perspektivet tror jag att vi alla är överens.
Jag skulle vilja säga till Stefano Zappala' att jag tackar honom för hans stöd för den europeiska invandringspolitiken. Till Zita Gurmai vill jag säga att jag tycker att jämställdheten mellan män och kvinnor är mycket viktig men jag vet inte om hennes kommentar även var riktad mot mig.
I vilket fall som helst är det faktum att hon är från Ungern redan en obestridlig tillgång.
Jag skulle vilja säga till Ioannis Varvitsiotis att jag är väl medveten om att det finns en europeisk identitetskris och kanske också att Europaparlamentet skulle kunna hjälpa alla institutionerna med den frågan.
Varför inte tänka sig en ordentlig debatt, talman Pöttering, om vad den europeiska identiteten är?
Frågan om den europeiska identiteten är ett ämne för debatt i Europaparlamentet snarare än en fråga för stats- eller regeringschefer.
Kanske skulle Europaparlamentet till och med kunna anordna debatter i den här frågan och i så fall kommer vi att komma och säga vår åsikt.
Personligen tycker jag att det är parlamentets uppgift att definiera den europeiska identiteten snarare än regeringarnas, som naturligtvis har hand om den dagliga förvaltningen i sina länder.
Om den europeiska identiteten bör definieras någonstans så tror och hoppas jag att ordförande José Manuel Barroso kommer att hålla med om att det inte är i Europeiska rådet, eller i kommissionen, utan först och främst i Europaparlamentet.
Jag skulle vilja svara Othmar Karas, som sa att jag måste vara diplomatisk.
Ja, uppfattat, jag ska försöka att vara diplomatisk.
Jag hoppas att han å sin sida inte ifrågasatte huruvida mitt temperament skulle hindra mig från att vara diplomatisk.
Det är inte bara en fråga om att vara svag men smart, eller om att vara dynamisk men klumpig.
Kanske är det till och med möjligt att vara både dynamisk och skicklig. Jag vill i vilket fall som helst tacka er för att ni gav mig möjlighet att visa detta.
(Livliga applåder)
Tack president Sarkozy!
Jag har varit ledamot av Europaparlamentet i 29 år och jag kan inte minnas någon rådsordförande som stannat i tre och en halv timme för att diskutera med oss och svara på varje anförande.
Vi ser fram emot ert nästa besök.
Punkten är härmed avslutad.
Skriftliga förklaringar (artikel 142)
skriftlig. - (RO) Frankrike har tagit över ordförandeskapet i Europeiska unionen vid ett avgörande ögonblick, då EU letar efter tillfredsställande lösningar på flera utmaningar av strategisk karaktär.
Frankrike har fått uppgiften att garantera den fortsatta ratificeringen av Lissabonfördraget, fokusera på energiområdet och konsolidera Europeiska unionens säkerhets- och försvarspolitik.
Jag stöder det franska ordförandeskapets prioriteringar och hoppas att de genomförs framgångsrikt.
Som ledamot av utrikesutskottet och föredragande för samarbetet i Svartahavsområdet vill jag fokusera på en viktig aspekt som bör främjas i EU:s utrikespolitik.
Jag välkomnar Frankrikes initiativ att konsolidera den europeiska grannskapspolitiken men jag insisterar på att den östliga dimensionen ska få lika mycket uppmärksamhet och engagemang som Medelhavsdimensionen.
Denna målsättning bör gälla både de bilaterala förbindelserna, i samband med förhandlingar om EU:s framtida avtalsförbindelser, och multilaterala förbindelser inom Svartahavssynergin.
Frankrike tar nu över ordförandeskapet i EU under Europeiska året för interkulturell dialog och bör framgångsrikt kunna fortsätta med åtgärderna på det området.
Jag vill först och främst välkomna det europeiska engagemanget från rådets ordförande Nicolas Sarkozy och hans klarsynthet när det gäller de utmaningar som EU står inför.
Jag stöder det politiska uttalandet om att nya institutioner baserade på Lissabonfördraget är nödvändiga och att det utan dem skulle vara oansvarigt att planera ytterligare anslutningar.
Ett resultatinriktat EU måste beakta medborgarnas förväntningar och visa att vi är en lösning och inte ett problem.
Jag stöder idén om en mekanism vid gränserna som ska se till att konkurrensen är rättvis och inte snedvriden, med beaktande av miljöåtgärdernas inverkan i samband med energi- och klimatfrågorna.
Prioriteringen av en EU-politik för laglig invandring är också en mänsklig, ekonomisk och social nödvändighet.
Jag vill gratulera Brice Hortefeux till hans utmärkta arbete med den europeiska pakten för invandring och asyl.
När det gäller EU:s försvar kommer presidentens modiga ståndpunkter att ge oss möjlighet att gå framåt i denna svåra fråga, särskilt genom att inkludera soldater från samtliga länders befolkningar och stödja utvecklingen av en europeisk försvarsindustri.
Presidenten gör rätt i att försvara den gemensamma jordbrukspolitiken. Den har aldrig varit mer nödvändig.
Avslutningsvis vill jag betona behovet av en bättre politisk dialog med Europeiska centralbanken för att få en europeisk ekonomisk styrning som ligger i linje med dagens globala krav.
Herr talman!
Jag vill lyckönska president Nicolas Sarkozy till hans arbete när han nu övertar ansvaret för rådet under de kommande sex månaderna.
Tyvärr samlas nu orosmolnen över EU:s framtid.
Vi måste hitta styrkan och kompetensen för att återlansera en europeisk väg som kan entusiasmera medborgarna, som fortfarande uppfattar EU som någonting avlägset och rätt svårbegripligt.
Jag vill även ta tillfället i akt och utmana rådets ordförande: för att föra medborgarna närmare EU måste konkreta signaler skickas ut.
Låt oss koncentrera all vår verksamhet till Bryssel och undvika den månatliga flytten till Strasbourg (där lokalerna i stället kunde användas till annat, exempelvis ett centrum för teknisk kvalitet). Denna ”resa” varje månad innebär faktiskt ett enormt och omotiverat slöseri med ekonomiska resurser och energiresurser.
Det franska ordförandeskapet har prioriterat rätt och satsar på till exempel klimat, invandring och försvar. Men jag vill fokusera på en aspekt som fått mindre uppmärksamhet men likväl är extremt viktig för våra ungdomar och hela idrottssektorn i EU.
Det franska ordförandeskapet stöder ”sex-plus-fem”-regeln inom idrotten, det vill säga en begränsning av antalet utländska spelare.
Målsättningarna är goda: att tvinga klubbarna att investera mer i sin egen utbildning för ungdomar och därmed till viss del bidra till att återupprätta jämvikten i konkurrensen.
Parlamentet stöder detta till hundra procent.
Därmed stöder vi också regeln om ”inhemsk skörd”, som - om än mer blygsamt - har likadana målsättningar.
Frågan är om sex-plus-fem-regeln är möjlig på EU-nivå.
Den strider mot den fria rörligheten för arbetstagare och kan endast tillämpas om det görs en avvikelse från EU-fördraget, och vi befinner oss långt bort från detta handlingssätt.
Det är tveksamt om EG-domstolen någonsin skulle acceptera någonting sådant, trots den nya artikeln om idrott i Lissabonfördraget.
Europaparlamentet vill hjälpa till att hitta en lösning som främjar den europeiska fotbollen.
Vi uppmanar helt enkelt till en stabil lösning, en lösning som inte gör att fotbollen kastas in i ett kaostillstånd.
Ingen vill ha en Bosman del 2.
President Nicolas Sarkozy använde ungefär en tredjedel av sitt anförande till att försvara Lissabonfördraget och fortsätta sätta press på och utöva utpressning mot Irland. Han glömmer vad som står i EU:s regelverk om ikraftträdandet av ett nytt fördrag - det ska ratificeras av alla medlemsstater.
Om en majoritet av den irländska befolkningen förkastade det så är fördraget stendött.
Ratificeringsprocessen bör inte fortsätta.
Att insistera på en ratificering av fördraget är en odemokratisk hållning.
En annan prioritering är att skärpa invandringspolitiken, där återvändandedirektivet, även känt som det skamliga direktivet, utmärker sig på grund av att det åsidosätter grundläggande mänskliga rättigheter och behandlar illegala invandrare som brottslingar istället för som människor som har flytt undan svält i sina egna hemländer på jakt efter en bättre framtid för sig själva och sina familjer.
Det sociala området nonchalerades helt.
Han känner till det motstånd som finns mot förslaget om att ändra arbetstidsdirektivet och de förslag som rådet godkände och skickade till Europaparlamentet, som syftar till att försvaga arbetstagares rättigheter, öppna möjligheten till en längre genomsnittlig vecka med upp till 60 eller 65 timmar, avreglering av sysselsättning och lägre löner.
skriftlig. - (PL) Jag vill uttrycka min förhoppning om att de sex månaderna med det franska ordförandeskapet kommer att kännetecknas av ett givande och effektivt arbete som ska gynna samtliga EU-medborgare.
Jag vill dock betona jordbrukets stora betydelse inom EU.
I till exempel Polen arbetade 2005 över 17 procent av landets anställda inom jordbruket.
Jordbruksfrågan är av indirekt betydelse för medlemsstaterna - här tänker jag främst på problemet med livsmedelstrygghet i samband med stigande livsmedelspriser på världsmarknaderna.
Jag hoppas att det franska ordförandeskapet kommer fram till en lösning i flera omtvistade frågor med anknytning till EU:s jordbruksmodell.
EU har inte tillräckligt bra klimat eller jordbruksförhållanden för att kunna avstå helt från sitt stöd till jordbrukarna.
Kostnaden för att producera kött, mjölk eller spannmål kommer alltid att vara högre på vår kontinent än i Sydamerika, Förenta staterna eller Australien.
Vi måste komma ihåg att dessa länder också stöder sina jordbrukare.
Jag anser att högre priser på jordbruksprodukter skapar en utvecklingsmöjlighet för EU:s jordbruk.
Det finns dock en fara att extrainkomsten snappas upp av mellanled. Med andra ord skapar ökade livsmedelspriser en oproportionerlig ökning av kostnaderna för jordbrukets produktionsmetod.
Resultatet blir att överskottet absorberas av mellanled.
Jordbruket är fortfarande en viktig ekonomisk sektor.
Villkoren för dess funktion har ändrats men huvudprioriteringarna - att garantera en anständig inkomstnivå för jordbrukarna och livsmedelstrygghet - finns fortfarande kvar.
Efter att Nicolas Sarkozy slagit blå dunster i ögonen på det franska folket genom att säga att han skulle respektera resultatet från den omröstning som hölls 2005 - varigenom den ”europeiska konstitutionen” förkastades - samtidigt som han körde vidare med ”minifördraget”, som i stort sett var en omstuvning av innehållet i det nedröstade fördraget, genom att presentera det i en annan form och undvika ytterligare en folkomröstning, ansvarar han nu för den process som sattes i gång av Angela Merkel. Man försöker alltså ännu en gång tvinga igenom detta federalistiska, nyliberala och militaristiska fördrag som redan har röstats ned tre gånger.
Mot bakgrund av den fördjupade krisen för kapitalismen, storfinansen och EU:s långtgående befogenheter visar särskilt Frankrike och Tyskland ”vägen ut” genom att pressa fram sin federalistiska, nyliberala och militaristiska politik och detta förslag till fördrag, som ett försök att stärka grunden för en ”superstat” för att bygga upp mekanismerna för imperialistiska ingripanden i tätt samarbete med Förenta staterna och Nato.
För att lyckas har det utövats påtryckningar och utpressning (utvidgning, ett EU med två hastigheter, etc.).
Döv, stum och blind för irländarnas uttryckta vilja konspirerar unionen mot den senare för att få dem att hålla ytterligare en folkomröstning 2009, till och med före valet till Europaparlamentet.
skriftlig. - (HU) En av de viktigaste uppgifterna för det franska ordförandeskapet kommer att vara samordningen av medlemsstaternas skyldigheter när det gäller klimatförändringar.
Det är mycket viktigt att vi minskar utsläppen av växthusgaser på EU-nivå.
Detta kan ske om vi tar Kyotoprotokollet på allvar och fortsätter att minska utsläppen betydligt i jämförelse med basåret 1990, i enlighet med dess bestämmelser.
Det skulle vara skandalöst om de medlemsstater som inte minskade utan snarare ökade sina utsläpp mellan 1990 och 2005 nu skulle belönas av Europeiska unionen och få behålla sin fördel, som är oförenlig med Kyotoprotokollet.
Det skulle vara ännu mer upprörande om de medlemsstater som tar Kyotoprotokollet på allvar och ärligt minskar sina utsläpp - inklusive Ungern - skulle bestraffas med ännu fler restriktioner.
Jag hoppas att det franska ordförandeskapet aldrig kommer att acceptera ett sådant hån mot Kyotoprotokollet och den negativa särbehandlingen av de nya medlemsstaterna, inklusive mitt hemland.
skriftlig. - (PL) Jag vill tacka den franske presidenten för hans anförande, där flera av EU:s grundläggande problem tas upp.
Det stämmer att vi måste överväga hur vi ska lösa krisen inom EU.
Det är en klen tröst att praktiskt taget hela världen befinner sig i en situation som är mer eller mindre kritisk.
Detta har en viktig ekonomisk och social dimension.
Jag talar om svälthotet i flera områden i världen, eftersom livsmedelpriserna stiger snabbt, om energitrygghet och även om miljöns status.
Världens ekonomiska system blir alltmer instabilt.
Varför betonar jag detta?
Därför att det inte är läge att vara självrättfärdiga.
De cirka 500 miljoner EU-medborgarna utgör för närvarande mindre än 8 procent av världens befolkning, och om 40 år kommer denna del knappt att nå upp till tröskelnivån för valbarhet - 5 procent.
Vår europeiska utgångspunkt får därför inte förbise högre stående värden som är förenade med upprätthållandet av den euroatlantiska civilisationen.
Detta har också en etisk dimension.
I varje EU-land behöver vi därför visa vederbörlig omsorg om familjen, som även om den är en mycket liten gemenskap samtidigt utgör en av hörnstenarna i hela den europeiska gemenskapen.
Vi får inte glömma detta.
Om vi gör det kommer vi att tappa greppet, som vi håller på att göra nu, genom att missbruka begreppet ”äktenskap” och använda det om förbindelser som inte är äktenskap.
Det stämmer att vi behöver nya rättsliga ramar men de måste vara sådana som människor kan förstå.
EU-medborgare är föremål för åtgärder som vidtagits av Europaparlamentet, rådet och kommissionen.
Vi tillhandahåller bara en tjänst.
Det är just precis ur den aspekten vi måste se på Irland.
skriftlig. - (PL) Som väntat har en av det franska ordförandeskapets prioriteringar blivit frågan om ratificering av Lissabonfördraget.
Oväntat för de flesta observatörer var dock att huvudrollen i början av det franska ordförandeskapet spelades av Polen eller för att vara mer exakt den polske presidenten Lech Kaczyński.
Jag förstår inte de argument som Polens president anför för att låta bli att underteckna Lissabonfördragets ratificeringsdokument.
Fördraget ratificerades av sejmen och av senaten.
Inget har hänt som kan försena presidentens undertecknande.
Fördraget har till exempel inte hänskjutits till författningsdomstolen.
Detta liknar respektlöshet för Europaparlamentet och brott mot en överenskommelse med premiärministern Donald Tusk.
Jag håller med rådets ordförande om att detta inte är av politisk utan etisk karaktär.
Polen förhandlade sig till fördraget, undertecknade det och är enligt internationell rätt skyldigt att slutföra ratificeringsprocessen.
Jag hoppas också innerligt att situationen när det gäller ratificeringen av fördraget kommer att förändras snart och att hållningen kommer att vara avsevärt bättre när det franska ordförandeskapet går mot sitt slut än vad den är nu för tillfället.
skriftlig. - (FI) Herr talman! Jag respekterar den tydliga önskan från rådets ordförande Nicolas Sarkozy om att inta en ambitiös hållning i fråga om EU:s energi- och klimatpaket och att nå en överenskommelse i frågan under det franska ordförandeskapet.
Jag hoppas att detta framför allt innebär att utmaningarna med klimatförändringarna till sist befinner sig i politikens centrum.
Jag vill dock påminna rådets ordförande om uppgiftens allvar - handel med utsläppsrätter är ett väldigt viktigt marknadsverktyg och påverkar så många människor att vi inte har råd att sträva efter det slags politiska tidtabell som tillämpas på bekostnad av miljön och en hållbar utveckling.
Annars kan det sluta med att Frankrike får stå där med skammen, något som landet knappast kan känna stolthet över.
Förra månaden organiserade jag ett seminarium där miljöorganisationer, forskningsorgan och organ som påverkas av handeln med utsläppsrätter kunde uttrycka sina åsikter om de ekonomiska effekterna. Budskapet jag fick var tydligt.
Kommissionens förslag kommer att innebära mycket högre kostnader utan att det leder till jämförbara miljöfördelar.
Jag syftar på McKinseys oroväckande analys av frågan.
Handeln med utsläppsrätter måste förbättras.
Situationen är allvarlig.
Vi kommer inte att kunna använda den europeiska industrin, som har hanterat sin egen verksamhet bra, som försökskanin igen såvida inte systemet hanteras vårdslöst.
Det är bättre att misslyckas med att uträtta något än att lyckas med att misslyckas.
Jag anser att vi kan leverera ett gott resultat med tiden men det krävs vissa väsentliga justeringar.
Utsläppen av koldioxid förebyggs inte med fromma förhoppningar och löften, såvida de inte blir en del av själva direktivet.
Vi måste behålla vår beslutsamhet när det gäller att dra ned på skyldigheterna, men förfarandet är i högsta grad öppet för diskussion.
I Europaparlamentet har vi uppvisat en bred front mot kommissionens sätt att närma sig de föreliggande alternativen.
Jag vill be rådets ordförande att bekanta sig med den.
skriftlig. - (RO) Herr talman! Ni har presenterat ett mycket ambitiöst program, som jag hoppas att ni kommer att slutföra med framgång.
Den europeiska pakten för invandring och asyl är en nödvändig prioritering för att minska den illegala invandringen och skapa en enhetlig politik för laglig invandring.
Likväl vill jag betona en aspekt som ni bör beakta innan ni påbörjar de planerade åtgärderna. Pakten bör omfatta ett antal åtgärder som tar hänsyn till de restriktioner på den europeiska arbetsmarknaden som vissa nya medlemsstater påtvingat arbetstagarna.
Det är inte normalt att den ekonomiska migrationen från tredjeländer är större än den fria rörligheten mellan länder inom EU.
Det finns medlemsstater som har övergångsbestämmelser som reglerar tillträdet till arbetsmarknaden för EU:s arbetstagare.
När väl politiken för laglig invandring börjat gälla finns det en risk för att EU:s medborgare missgynnas jämfört med tredjelandsmedborgare.
I detta avseende vill jag gratulera Frankrike till att ha tagit det första steget i denna riktning den 1 juli när landet öppnade sin arbetsmarknad för medborgare från de länder som anslöt sig till EU 2004.
Jag hoppas att Rumänien och Bulgarien behandlas på samma sätt så fort som möjligt och jag uppmuntrar de andra medlemsstaterna att följa Frankrikes exempel.
Frankrike har tagit på sig ansvaret att leda den europeiska agendan i sex månader i ett mycket svårt läge, som uppstått efter Irlands förkastande av Lissabonfördraget.
Det franska ordförandeskapets program är ambitiöst men man ska även vara medveten om EU-medborgarnas förväntningar.
Den senaste Eurobarometerundersökningen visar att endast 52 procent av EU-medborgarna anser att medlemskapet gynnar deras hemland.
Det behövs en strategi för att få EU:s medborgare att förstå att våra gemensamma intressen är mycket viktigare från ekonomisk och politisk synvinkel än de saker som skiljer oss åt.
Självklart är det franska ordförandeskapets prioritering att hitta en metod att sluta den irländska sprickan, eftersom EU-processen måste fortsätta med tanke på att Nicefördraget blockerar en utvidgning.
När det gäller det franska ordförandeskapets andra prioritering - den gemensamma jordbrukspolitiken och dess förberedelse inför framtida utmaningar - bör det nämnas att upprätthållandet av ett system med samlat gårdsstöd är tillämpligt i Rumänien från och med 2013.
Även som mottagare av stöd från den gemensamma jordbrukspolitiken kommer Rumänien att ta emot 735 miljoner euro i år i europeiskt direktstöd till rumänska jordbrukare.
Jag vill ta upp följande två punkter:
För det första är det helt omöjligt att söka asyl i 27 länder.
Vi har Dublin II-förordningen, som reglerar frågan om mottagarländernas ansvar.
Det finns dock fortfarande skillnader mellan medlemsstaterna när det gäller att inse behovet av internationellt skydd och det är ett stort problem.
För det andra vill jag nämna mänsklighetens grundläggande problem i dagens värld.
Hur kan vi alla leva tillsammans i en globaliserad värld?
Vi måste ta itu med de underliggande orsaker som driver vissa desperata människor att lämna sina hemländer. Den europeiska pakten för invandring och asyl anser jag inte uppnår den rätta jämvikten mellan att bekämpa människosmugglare, främja laglig invandring och upprätta en ambitiös gemensam utvecklingspolitik.
skriftlig. - (ET) I år har EU möjlighet att se sig självt i spegeln och se om de beslut som vi tog förra året burit frukt.
Förra året inleddes handlingsplanen för miljö och energi för att minska utsläppen av växthusgaser och bekämpa den globala uppvärmningen.
Vi har diskuterat en gemensam invandringspolitik för Europeiska unionen, och för en stund sedan fick vi höra uppgifter om den illegala invandringens enorma ökning.
Vi har också gett oss i kast med skyddsfrågor: gemensamma europeiska styrkor har utfört militära operationer ute i världen, och sedan 2004 har vi skapat EU:s stridsgrupper och enheter för nödinsatser.
Det nya ordförandeskapet under den franske presidenten Nicolas Sarkozy har gett EU-politiken fräschör och nytt liv. Det har gett oss tanken på en miniöverenskommelse och en ny inställning till de nya medlemsstaterna.
Det finns många exempel på detta.
Tack vare sin egen drivkraft och företagsamhet kommer han säkert att kunna starta eller påskynda många utmanande projekt.
Med tanke på det vill jag understryka att det land som innehar ordförandeskapet inte ska driva EU-frågor separat, även om det har rätt att föreslå vissa punkter på arbetsplanen.
Det är av grundläggande betydelse att ordförandeskapet inte är ansvarigt för beslut som fattas i Europeiska rådet, och det är något som landet bör fokusera sitt ordförandeskap på, i stället för att pryda det med tomma löften.
Framför allt hoppas jag väldigt mycket på att det franska ordförandeskapet ska kunna ge nytt hopp till EU-medborgarna i fråga om specifika projekt.
skriftlig. - (EN) Herr rådsordförande! Vid det senaste EU-toppmötet i Bryssel diskuterades inrättandet av en union för Medelhavsområdet - ett viktigt initiativ för hela Medelhavsregionen och en prioritering för det franska ordförandeskapet.
Men jag hoppas innerligt att Östersjöregionen och Östersjöstrategin inte kommer att försummas när ordförandeskapet betonar unionen för Medelhavsområdet.
Östersjön har i stort sett blivit en EU-sjö, omringad av åtta medlemsstater sedan 2004.
EU-strategin för Östersjön innefattar områden som miljö, ekonomi, kultur och utbildning samt säkerhet. Den utgör en hållbar plan för utvecklingen av denna region.
Det skulle glädja mig om det franska ordförandeskapet tog sig tid att uppmärksamma frågorna beträffande Östersjön och att prioriteringen av Medelhavet inte drar undan mattan för Östersjöregionen.
Med tanke på det nästkommande svenska ordförandeskapet skulle det vara förnuftigt att börja inrikta sig på Östersjöstrategin för att garantera en bättre överensstämmelse mellan ordförandeskapen.
skriftlig. - (RO) Under de kommande sex månaderna kommer det franska ordförandeskapet att ha ett stort ansvar för EU:s framtid.
EU behöver Lissabonfördraget.
Den befintliga institutionella ramen, där det krävs enhällighet för vissa beslut, väger tungt.
Genom Lissabonfördraget ökar dessutom demokratiseringsgraden och de nationella parlamentens befogenheter, och medbeslutandeförfarandet införs på de flesta områden.
Det franska ordförandeskapet bör även stödja den gemensamma jordbrukspolitiken, som gör det möjligt för EU:s jordbrukare att producera mer.
Tillsammans med de andra medlemsstaterna bör det franska ordförandeskapet försöka hitta lösningar på EU:s dödläge efter den irländska folkomröstningen.
Det franska ordförandeskapet tillkännagav sina prioriteringar inför den kommande perioden: klimatförändring, invandring, den gemensamma jordbrukspolitiken, EU:s försvars och säkerhet.
I Köpenhamn nästa höst ska EU delta i slutandet av ett internationellt avtal efter Kyoto.
EU bör ge exempel på handlingskraft i kampen mot klimatförändringen, och av det skälet bör EU:s antagande av paketet för energi och klimatförändring vara ett av målen för det franska ordförandeskapet.
skriftlig. - (EN) Ingen kan förklara anledningen till resultatet i den irländska folkomröstningen.
En norm blir en lag efter ett allmänt godkännande av folket.
Dess innebörd bör motsvara allas övertygelse.
En landsman till er, en tänkare som vilar i Pantheon, Rousseau, skrev att ”varje lag som folket inte själva har ratificerat är utan verkan, det är inte någon lag”.
Det är därför som människorna ska kontrollera sina regeringar, som annars riskerar att åsidosätta deras rättigheter.
Men hur ska människorna kunna ta kontrollen med hjälp av ett verktyg som de inte förstår sig på, vars struktur är lika komplicerad och otydlig som i det senaste fördraget?
Jag tvivlar inte på att ni i detta Europaparlamentets ”tempel” vill framstå som - för att parafrasera Dominique de Villepin -- en ”väktare av ett ideal och ett samvete”.
Jag räknar dock med att ni kommer att vara mer intresserad av att förmedla information om plattformarna för ett gemensamt förverkligande av europeiska intressen till den allmänna opinionen, vilket i sin tur gör att medierna håller sig borta från ert privatliv och i stället fokuserar på er politik.
(Sammanträdet avbröts kl. 13.40 och återupptogs kl. 15.00.)
1.
Gemenskapsstatistik över utrikeshandeln med tredjeländer (
Datum för nästa sammanträdesperiod: se protokollet
Meddelande om rådets gemensamma ståndpunkter: se protokollet
Parlamentets sammansättning: se protokollet
Inkomna dokument: se protokollet
Återupptagande av sessionen
Jag förklarar Europaparlamentets session återupptagen efter avbrottet torsdagen den 4 december 2008.
Omröstning
Nästa punkt är omröstningen.
(För omröstningsresultat och andra uppgifter som rör omröstningen: se protokollet.)
Situationen i Mellanöstern/Gaza (debatt)
Nästa punkt är rådets och kommissionens uttalanden om situationen i Mellanöstern/Gaza.
Det gläder mig särskilt att välkomna rådets tjänstgörande ordförande, den tjeckiske utrikesministern Karel Schwarzenberg, som måste resa vidare till Sydafrika i dag.
Tidigare ordförandeskap har ordnat det så att en ställföreträdare har kommit i stället för deras utrikesminister, så vi uppskattar särskilt att ni är här i dag, herr Schwarzenberg.
Ni är varmt välkommen!
Det gläder oss naturligtvis också att den ansvariga kommissionsledamoten, Benita Ferrero-Waldner, är närvarande - som hon nästan alltid är.
Som ni vet känner kommissionsledamoten också mycket väl till problemen i Mellanösternkonflikten och hon har, i likhet med Karel Schwarzenberg, besökt området.
Också ni är varmt välkommen, fru kommissionsledamot!
rådets ordförande. - (EN) Herr talman! Tack så mycket för att ni ger mig ordet i denna mycket lägliga debatt om den dramatiska situationen i Mellanöstern.
Situationen har försämrats snabbt på alla nivåer sedan Israel inledde sin militära offensiv i Gazaremsan den 27 december.
De humanitära konsekvenserna av denna operation är dramatiska för befolkningen i Gaza.
Sedan operationen inleddes har över 900 palestinier omkommit, varav cirka 30 procent var kvinnor och barn.
Vi är ytterst oroade över förlusten av människoliv, vilket vi vid upprepade tillfällen har gett uttryck för i ordförandeskapets uttalanden.
Europeiska unionen beklagar djupt de pågående fientligheterna, som har lett till så många civila dödsoffer, och vi vill förmedla våra uppriktiga kondoleanser till offrens familjer.
Vi är särskilt oroade över incidenter som attacken mot FN-skolan i Jebaliya och beskjutningen mot humanitära hjälpkonvojer, då humanitär biståndspersonal dödades.
Över 4 200 palestinier har skadats enligt FN:s kontor för samordning av humanitära frågor (OCHA).
Enligt detta FN-organs beräkningar har 28 000 personer blivit internflyktingar sedan fientligheterna började.
Många av internflyktingarna söker sin tillflykt till läger, resten av dem vistas hos släktingar.
De största humanitära behoven rör det stora antalet skadade och de överbelastade sjukhusen, medan internflyktingarna och deras värdfamiljer behöver särskild hjälp som livsmedel, husrum, vatten och nödvändighetsartiklar.
Eftersom vattenförsörjningssystemet skadades allvarligt och är i behov av en snabb reparation, har Gazas befolkning knappt tillgång till rent vatten.
Att tillhandahålla dricksvatten är därför av yttersta vikt.
Det råder också en omfattande livsmedelsbrist bland hela befolkningen.
Utländska icke-statliga organisationer har inte fått komma in i Gaza för att leverera och övervaka det humanitära biståndet på lämpligt sätt sedan den 4 november förra året.
Det antal lastbilar som kommer in i Gaza har ökat sedan operationerna inleddes.
Men det nuvarande dagliga genomsnittet på 55 lastbilar är fortfarande skriande otillräckligt med tanke på att det krävs minst 300 lastbilar per dag för att täcka behoven hos 80 procent av befolkningen, som har blivit biståndsberoende.
EU har nära följt de tragiska händelserna ända från början.
Tre dagar efter det att operationen inleddes möttes utrikesministrarna för ett extra sammanträde i Paris för att diskutera situationen.
De var överens om behovet av en omedelbar och permanent vapenvila och brådskande humanitära åtgärder för att påskynda fredsprocessen.
Syftet med mötet var främst att diskutera hur man kan bidra till att få slut på våldet och mildra den humanitära krisen.
Ordförandeskapet ledde ett diplomatiskt uppdrag i Mellanöstern och EU:s ministertrojka besökte regionen den 4-6 januari för möten i Egypten, Israel, med den palestinska myndigheten och i Jordanien.
Den höga representanten besökte även Syrien, Libanon och Turkiet.
Grunddragen för en lösning på krisen börjar skönjas.
Först och främst måste Hamas ovillkorligen upphöra med sina raketattacker mot Israel, och Israel måste upphöra med sina militära aktioner för att möjliggöra oavbrutna leveranser av humanitärt bistånd och återupptagandet av de offentliga tjänster och den sjukvård som Gaza är i så stort behov av.
Den sex månader långa vapenvilan, som löpte ut den 19 december, var långt ifrån perfekt.
Israel led sig genom regelbundna raketbeskjutningar, i vetskapen om att de hade större eldkraft än sin fiende.
Gaza uthärdade verkligt pressande ekonomisk blockad, som fullständigt raserade dess ekonomiska utveckling.
För att nå en hållbar vapenvila måste vi finna en förnuftig kompromiss som omfattar ett slut på raketuppskjutningarna och återöppnande av gränsövergångarna.
För att lösningen ska vara genomförbar måste man ta itu med tunnlarna över gränserna, särskilt längs Philadelphiarutten, för att förhindra vapensmuggling.
Lösningen måste också leda till ett systematiskt och kontrollerat öppnande av alla gränsövergångar för att ge Gazas ekonomi möjlighet att utvecklas.
Vi anser att utplacering av internationella uppdrag för att övervaka genomförandet av vapenvilan och agera som en kontaktpunkt mellan de två sidorna skulle kunna vara en användbar lösning i detta avseende.
EU är redo att skicka tillbaka sina observatörer till Rafah-gränsövergången och förlänga mandatet för EU:s gränsuppdrag i omfattning och innehåll.
Vi vet att Israel har gått med på ett dagligt uppehåll för att livsmedel, bränsle och läkemedel, som det finns ett så trängande behov av, ska kunna komma in i Gaza.
Endast en fullständig och omedelbar vapenvila skulle emellertid möjliggöra leverans och distribution av de stora kvantiteter bistånd som Gaza så desperat behöver och återupptagandet av grundläggande tjänster.
Israel måste garantera obehindrat och säkert tillträde för det humanitära biståndet och andra nödvändiga varor, inklusive livsmedel, läkemedel och bränsle till den palestinska civilbefolkningen i Gazaremsan, samt en säker passage för civila och humanitär personal, in i och ut från Gazaremsan.
En varaktig och allomfattande lösning i Gaza kommer dock inte att vara tillräcklig för att skapa fred i regionen.
Det finns mer allmänna och komplicerade utmaningar som vi måste hantera.
Vi behöver en ny och integrerande strategi för att komma till rätta med den palestinska politiska situationen och återuppta fredsförhandlingarna, som har ställts in till följd av Gazakrisen.
Försoning i Palestina och en regering som avspeglar det palestinska folkets ambitioner är mer nödvändigt än någonsin.
Vi stöder därför de medlingsinsatser som genomförts av Egypten i enlighet med Arabförbundets resolutioner av den 26 november 2008.
Som det påpekas i rådets (allmänna frågor och yttre förbindelser) slutsatser från december 2008 är EU berett att stödja en stabil palestinsk regering som för en politik och vidtar åtgärder som avspeglar kvartettens principer.
EU betonar behovet av att uppnå en rättvis, varaktig och allomfattande fred i Mellanöstern och efterlyser ett återupptagande av förhandlingarna mellan Palestina och Israel, samt att alla kvarstående frågor i den israelisk-palestinska konflikten, inklusive alla grundfrågor, kan lösas.
En varaktig och allomfattande lösning kommer slutligen att vara beroende av att det görs verkliga framsteg i fredsprocessen i Mellanöstern.
Det kommer att krävas snabba och omfattande insatser från parterna för att nå en heltäckande fred, som grundas på visionen av en region där två demokratiska stater, Israel och Palestina, existerar sida vid sida inom säkra och erkända gränser.
Det senaste våldsutbrottet i Mellanöstern kanske inte bara leder till ett bakslag när det gäller utsikterna till en fredlig lösning på konflikten mellan Israel och Palestina.
Den politiska skada som striderna orsakar, både när det gäller regional polarisering och radikalisering, och det försämrade anseendet för de mer moderata krafterna får inte heller nonchaleras.
Endast en livskraftig palestinsk stat kommer att skapa säkerhet i denna region, som redan har lidit alltför länge.
Detta ligger särskilt i Israels och dess grannars intresse.
Därför måste kraftfulla åtgärder omedelbart vidtas för att motverka den skada som de militära aktionerna har orsakat för att blåsa nytt liv i förhoppningen om ett rättvist och förhandlat resultat.
(Applåder)
ledamot av kommissionen. - (EN) Herr talman! Jag tror att vi alla hade hoppats på en bättre inledning på 2009.
Tyvärr står vi inför en fruktansvärd och skrämmande konflikt i Gaza, som nu är inne på tredje veckan.
Detta skapar mycket stor oro.
Vi diskuterade frågan i går vid ett möte med utskottet för utrikesfrågor, utskottet för utveckling och de parlamentsledamöter som besökte Gaza under helgen.
Rådsordföranden har redan tagit upp den ohyggliga statistiken över döda och skadade, som förvärras varje dag.
Det dyker upp allt fler exempel på offer som drabbats av extrema brännskador och hjälporganisationerna rapporterar att befolkningen lider akut brist på mat, bränsle och medicin. Dessutom är byggnaderna och infrastrukturen förstörda.
Israel har dock också drabbats av förluster och har träffats av hundratals raketer som Hamas avfyrat in på landets territorium, med civila israeler som mål.
Krig skapar tyvärr alltid stort mänskligt lidande och det här kriget är inget undantag.
Konflikten har inte bara förödande effekter, utan fördröjer också möjligheterna till fred, undergräver det arabiska fredsinitiativet och kan få en mycket negativ inverkan på stabiliteten i hela regionen.
Jag vill bara snabbt beskriva den diplomatiska aktivitet som vi tillsammans bedrivit i syfte att få slut på den här konflikten och sedan titta på vilka utmaningar som finns på medellång och lång sikt.
Vi har varit aktiva redan från början, vilket jag menar är viktigt.
Vi vet att vi inte är någon huvudaktör i Mellanöstern, men vi har varit, och är, en viktig aktör.
Det extrainsatta mötet mellan EU-ländernas utrikesministrar som hölls i Paris den 30 december 2008 med anledning av krisens utbrott var därför mycket viktigt för att kunna ta fram förslag redan från början - Parisdeklarationen - i syfte att få slut på den här konflikten. Detta använde vi sedan i vår delegation och vid besöket i Mellanöstern.
Deklarationen kan delas in i tre delar.
Först och främst efterlyser vi ett omedelbart eldupphör av humanitära skäl, vilket skulle innebära att både Hamas raketattacker mot Israel och Israels militära angrepp måste upphöra.
Vi vill också att ett eldupphör ska åtföljas av ett permanent och normalt öppnande av alla gränsövergångar, i enlighet med avtalet om rörlighet och tillträde från 2005.
Vi uttryckte vår beredskap att på nytt skicka ut Europeiska unionens gränsövervakningsuppdrag (BAM) till gränsövergången i Rafah så att den kan öppnas på nytt, och vi indikerade också att vi är beredda att undersöka möjligheten att skicka hjälp till andra gränsövergångar, förutsatt att våra säkerhetskrav uppfylls.
För det andra betonade vi det omedelbara behovet av humanitärt bistånd, som måste uppfyllas.
Här efterlyste vi att gränsövergångarna omedelbart ska öppnas för att medicinsk hjälp, bränsle och livsmedel snarast ska kunna levereras till Gazaremsan och för att hjälparbetare ska kunna nå fram och sårade evakueras.
För det tredje upprepade vi vår ståndpunkt att det inte finns någon militär lösning på konflikten mellan Israel och Palestina, att fredsprocessen är den enda vägen framåt samt att insatserna måste intensifieras så snart som det finns ett varaktigt eldupphör.
Som ni vet genomfördes vår delegationsresa samtidigt som president Sarkozy var på besök. Han hade sedan tidigare planerat en resa till Syrien och Libanon och beslutade nu att även besöka Egypten och Israel för att ge extra stöd för de här insatserna, med utgångspunkt från vår deklaration från den 30 december 2008.
Frankrike leder för närvarande FN:s säkerhetsråd och det var därför ett viktigt initiativ.
Besöken samordnades noggrant och inkluderade ett gemensamt möte i Ramallah, där president Sarkozy beskrev sin plan för eldupphör, som vi - trojkan - i viss mån hade berett väg för genom våra samtal med viktiga intressenter, framför allt Egypten och Jerusalem.
De här insatserna förstärkte varandra och sände ett kraftfullt, samordnat budskap från EU. Trojkan förmedlade inte bara EU:s hållning i frågan, utan manifesterade också vår närvaro.
Jag anser att det var viktigt att också president Sarkozy reste till Syrien och att Javier Solana följde med honom till Syrien och Libanon och även hade överläggningar med Turkiet.
Jag menar att allt detta var nödvändigt.
Jag betonade, som redan nämnts, den humanitära situationen och jag efterlyste framför allt att gränsövergångarna måste öppnas och en möjlighet till åtminstone några timmars eldupphör ges så att de internationella organisationerna kan genomföra sitt arbete.
Israel tog till sig en del av de här punkterna och i förhandlingarna med den israeliska regeringen utverkade jag också att en representant för ECHO kan placeras hos den israeliska förvarsmakten för att samordna distributionen av humanitärt bistånd med de israeliska styrkorna, på samma sätt som gjordes under kriget i Libanon, då det var ett kraftfullt verktyg för ökad samordning.
Jag vill utnyttja det här tillfället till att tacka alla de modiga kolleger som fortfarande arbetar i Gaza, representanter för UNWRA och ICRC, som vi arbetar med och som tar emot en stor del av vårt ekonomiska stöd, men också många andra.
(Applåder)
Jag vill också säga att mina tankar går till familjerna till de hjälparbetare som redan har blivit offer för dessa tragiska händelser.
Kommissionen har också fört över stora medel till humanitära fonder och vi är beredda att göra mer i framtiden.
Vad har vi uppnått med de här förhandlingarna?
Som rådsordföranden nämnde omfattade förhandlingarna också de viktigaste delarna i säkerhetsrådets senaste resolution, som antogs ett par dagar efter förhandlingarna, då USA lade ner sin röst.
Ett omedelbart eldupphör, egyptiska garantier för att smugglingen genom tunnlarna ska stoppas, öppnande av gränsövergångarna för humanitärt bistånd, inklusive utpostering av en styrka - eventuellt med internationellt deltagande och/eller den palestinska myndighetens säkerhetsstyrkor - som bevakar den 15 km långa Philadelphia-korridoren mellan Gaza och Egypten.
Vår uppfattning är att den palestinska myndigheten har accepterat det här förslaget och att Israel och Hamas nu studerar det.
Vi menar att det är mycket viktigt att man mycket snart kan få någonting som fungerar.
De senaste uppgifterna jag har är att alla arbetar med detta och att vi om ett par dagar faktiskt kommer att ha ett eldupphör.
Jag hoppas att så kommer att vara fallet.
När det gäller utsikterna på medellång sikt har beklagligtvis både Israel och Hamas inledningsvis avvisat FN:s säkerhetsråds resolution, men genom den dagliga kontakten hoppas jag att ett avtal snart kan komma till stånd.
Det är viktigt att påpeka och vara medveten om att Egypten har spelat en ledande roll när det gäller direktkontakter med Hamas och att president Sarkozys besök i Syrien och de turkiska insatserna har varit mycket viktiga i det här avseendet.
Det verkar också som om arabländernas toppmöte kommer att hållas i Qatar i slutet av veckan.
Som denna intensiva diplomatiska aktivitet visar har vi som mål att stödja alla relevanta aktörer som kan påverka Hamas och som kan hjälpa till att leverera en hållbar lösning i enlighet med FN:s säkerhetsråds resolution 1860.
Så snart som man kommit överens om eldupphör måste vi fundera över - förmodligen i form av en konferens - hur vi ska kunna formulera mer konkreta åtgärder för att uppfylla de humanitära behoven hos den palestinska befolkningen i Gaza.
Vi måste dock vara tydliga med att påpeka att oavsett vad vi gör får det inte bidra till en oändlig cykel av förstörelse och återuppbyggnad utan fred.
När omständigheterna är de rätta kommer jag eventuellt tillbaka till er för att söka er hjälp att på ett meningsfullt sätt bidra till konstruktiva insatser, på samma sätt som jag tidigare gjort.
Som ni känner till reser FN:s generalsekreterare Ban Ki-moon runt i regionen och förhoppningsvis kan också han bidra till den slutliga framgång som är absolut nödvändig för att få till stånd detta varaktiga eldupphör.
I ett långsiktigt perspektiv måste vi konstatera att den nuvarande offensiven tveklöst bidrar till att försvaga förtroendet mellan palestinierna och israelerna.
Militära operationer kan aldrig leda till en varaktig fred. Det kan endast ett politiskt avtal göra.
Dialogen måste därför återupptas mellan både israelerna och palestinierna och bland palestinierna själva.
När angreppen upphört tror jag att det kommer att vara viktigt att återuppta samtal som syftar till en omfattande fred så snart som möjligt.
Här måste vi arbeta med den nya amerikanska administrationen för att se till att den kan ställa sig bakom bilaterala förhandlingar från början.
Utifrån det perspektivet välkomnar jag den blivande utrikesministern Hillary Clintons ställningstaganden vid utfrågningen i senaten i går.
Vi kommer att insistera på att parterna förhandlar om innehåll, och inte bara om process, och att Anapolis-processen kan avslutas på ett framgångsrikt sätt.
Krisen visar att detta är mer brådskande än någonsin tidigare.
Frågan om försoning mellan palestinierna kommer också att vara central.
Hamas kommer sannolikt inte att utplånas genom det här angreppet.
Möjligen kommer organisationen att försvagas militärt, men stärkas politiskt.
Hamas ståndpunkt att president Abbas mandat går ut den 9 januari är en annan fråga som har nära koppling till reformeringen av PLO och Fatah.
För att få till stånd en varaktig fred är det tydligt att en stark palestinsk myndighet måste kunna tala för alla palestinier och att den måste ta ställning för en tvåstatslösning genom fredliga metoder.
Konflikten i Gaza har tyvärr också negativa återverkningar när det gäller det regionala stödet för fredsprocessen.
Flera fredsförespråkande arabregimers bild av Israel har solkats av det stora lidande som drabbat civilbefolkningen i Gaza.
Israeliska ledare och Israels befolkning bör vara medvetna om hur negativt detta är för deras ambitioner att leva i fred.
Vi är deras vänner och måste berätta för dem hur det ligger till.
Israel har därför ont om tid om de vill uppnå fred.
Detta är min första, korta - eller kanske inte så korta - analys och vi måste försöka arbeta för att få till stånd ett varaktigt eldupphör för att sedan kunna få i gång fredsförhandlingarna med den nya amerikanska administrationen.
Herr talman! Sjutton dagars strider i Gaza efterlämnar endast djup smärta.
Det allra värsta, som inte går att reparera, är att människor fått sätta livet till, bland dem oskyldiga civila och barn. Men vi kan också se förstörelse, kaos, hat och hämnd.
Radikalerna blir allt starkare på moderaternas bekostnad. Och fredsprocessen har spårat ut fullständigt.
Som talmannen betonade så beror detta på att man kan vinna ett krigs alla strider, men det viktigaste slaget kan fortfarande gå förlorat - kampen för fred.
Hellre än att försöka utmäta ansvar eller lägga skulden på den ena eller båda sidorna, är den viktigaste frågan - som kommissionsledamoten precis nämnde - att få till stånd ett eldupphör, enligt FN:s resolution 1860.
Som FN:s generalsekretare precis påminde oss om måste bägge sidor efterleva resolutionen.
Det är också mycket viktigt att lindra den hemska humanitära och ekonomiska situation som råder i Gazaremsan, som ”styrs” - inom citationstecken - av Hamas, som är en organisation som finns med på EU:s lista över terroristorganisationer.
Men vi måste komma ihåg att Hamas inte bara utgör orsaken till konflikten, utan Hamas är också konsekvensen av hemska förhållanden.
Min politiska grupp stöder och vill erkänna de ansträngningar som alla politiska grupper i parlamentet gör för att stödja förslaget till resolution som vi antar i morgon.
Vi vill också hylla de ledamöter som deltog i förhandlingarna, i synnerhet Elmar Brok som representerade min grupp och hade en mycket svår uppgift.
Min grupp stöder kommissionens och rådets ansträngningar för att få ett eldupphör så fort som möjligt, i samarbete med de arabiska länderna - i synnerhet Egypten - och andra medlemmar i Mellanösternkvartetten.
Vi är förhoppningsfulla efter den nya utrikesministern Hillary Clintons uttalande i går inför den amerikanska senatens utrikesutskott, om erbjudandet av pragmatisk och effektiv diplomati grundad på dialog.
Slutligen kommer jag till det allra viktigaste: Europeiska unionen är en union med värderingar och sätter freden på första plats.
Jag anser att Europeiska unionen måste göra alla ansträngningar och använda all sin politiska kraft i denna saks intresse, utan att vi låter våra tankar besudlas eller vårt hjärta förhärdas av konflikten.
(Applåder)
för PSE-gruppen. - (DE) Herr talman, mina damer och herrar! Debatter som den som vi för i dag är svåra för oss alla.
Anledningen till att de är svåra är att Israel är en vän, och många av oss - och det är sant särskilt för mig - är bundna till landet genom djup vänskap.
Det är särskilt viktigt att diskutera kontroversiella frågor öppet med vänner.
Fram till i dag har konflikten skördat 1 000 liv under 17 dagar.
Det är en blodig konflikt, och kvinnor och barn lider alldeles särskilt.
Det finns en FN-resolution som utgör grunden för att utropa ett omedelbart eldupphör och inleda förhandlingar.
Det är kristallklart att konflikten endast kan lösas utifrån internationell lagstiftning, och att internationell lagstiftning och internationell humanitär lagstiftning måste respekteras bör vara självklart för ett demokratiskt land som grundas på rättsstatsprincipen.
Det är faktiskt skamligt att vi måste diskutera det här.
Allt vi kan göra för att övervinna den humanitära krisen är att vädja om omedelbart eldupphör.
Det vi menar i vår resolution är inte vad som helst, utan något som är mycket viktigt för att få ett direkt och omedelbart slut på dödandet, hungern och lidandet.
Det är alldeles klart att staten Israel har rätt att försvara sig.
Staten har rätt att försvara sig mot folk som har som mål att förstöra den.
Men ett demokratiskt land som grundas på rättsstatsprincipen måste ändå fråga sig självt om de medel som används i det syftet är proportionella.
Enligt min åsikt - och jag tror de flesta ledamöterna i kammaren anser detsamma - är medlen inte proportionella.
(Applåder från vänster)
Vi måste säga till våra vänner i Israel, oavsett deras politiska ställning, att vi är medvetna om att Hamas inte är någon fredsrörelse.
Vi vet att organisationen leds av människor som inte delar våra grundläggande värderingar, och varje raket som avfyras mot Israel är ett angrepp som staten har rätt att försvara sig emot - men trots allt är det ett misstag att vägra inleda en dialog.
Om dialog utgör det grundläggande villkoret för en fredlig utveckling, då innebär en vägran att inleda en sådan dialog en fortsatt väpnad konflikt.
Därför krävs en grundläggande anpassning.
En dialog med Hamas måste komma till stånd.
Om Israel inte kan inleda dialogen direkt - jag kan förstå israeliska politikers inställning när de säger att de inte kan tala med Hamas, även om många medborgare anser att de borde - och om ledamöter av parlamentet och medlemmar i regeringen säger att de inte vill, finns det tillräckligt många möjligheter till internationell medling.
Det finns till exempel Mellanösternkvartetten, och en av Europeiska unionens uppgifter inom kvartetten är att få till stånd en medling om dialog.
Det är fundamentalt fel att tro att det i slutändan kan bli en militär lösning på Mellanösternkonflikten.
Jag anser att det är ett fundamentalt fel oavsett vilken sida som tror det.
Terrorattacker leder inte till någon lösning och konventionella militära strider leder inte till någon lösning.
Den enda lösningen är en dialog mellan konfliktens bägge parter, med hjälp av internationell medling.
Det krävs ett omedelbart eldupphör.
Det måste det internationella samfundets system se till, om så med hjälp av en multinationell styrka där arabiska och i synnerhet muslimska stater ingår.
Det vore en väg för att få till stånd ett eldupphör och en förbättring.
När jag var en ung grabb och började med politik fick jag lära mig att man inte talar med terrorister.
Vid den tiden var Yasser Arafat den störste terroristen.
Ett par år senare såg jag bilder på tv när den här terroristen fick Nobels fredspris tillsammans med israeliska politiker.
Det som var möjligt då kan också bli möjligt i framtiden.
Frågan är därför om tillräckliga framsteg görs så att de system som finns kan få till stånd den nödvändiga dialogen.
På min grupps vägnar vill jag tacka alla dem, också från andra grupper, som har arbetat med vår resolution.
Om resolutionen, som alla grupper i kammaren stöder - jag anser att det är ett gott tecken - kan bidra till en förbättrad atmosfär, har vi bidragit, om än i liten utsträckning, till att få slut på ett dödande som ingen kan acceptera.
(Applåder från vänster)
för ALDE-gruppen. - (FR) Herr talman, fru kommissionsledamot! Den dagen kommer då vi måste skilja det goda från det onda, men jag anser att det i dag är mer brådskande att vi ställer följande krav: en omedelbar vapenvila, upphörande av raketanfallen mot Israel och israeliska operationer i Gaza, humanitärt bistånd, en hållbar vapenvila, upphörande av smuggling av vapen och ammunition, effektiv övervakning av gränsen mellan Egypten och Gaza, tillbakadragande av israeliska trupper och återöppnande av gränsövergångar; och slutligen, upphävande av embargot - allt detta, samtidigt.
Det blir en mycket omfattande fas, som utan tvekan eller högst sannolikt kommer att kräva närvaron av en internationell styrka, och jag tror att unionen bör förbereda sig för att ingå i den.
Jag skulle vilja göra två tillägg.
För att nå resultat måste Europeiska unionen tala och agera tydligt och organiserat.
Det är väldigt bra att ha goda avsikter, men det är viktigare att vara effektiv.
Förenta staterna måste också ta på sig en uppgift, liksom Arabförbundet och dess medlemsstater.
Slutligen vill jag tillägga att, för att erbjuda ett verkligt alternativ till situationen i Gaza måste Israel i hög grad förbättra situationen på Västbanken: 634 gränsövergångar, avskärningen av vägnätet, 8 meter höga murar och otaliga kränkningar av palestinierna innebär inte ett tillräckligt attraktivt alternativ för invånarna i Gaza för att få dem att vända ryggen mot Hamas.
Sammanfattningsvis skulle jag vilja säga att den dagen kommer onekligen då alla måste tala med varandra.
(Applåder)
Herr talman, mina damer och herrar! Precis som alla andra är vi tydligt involverade i och upprörda över situationen, men jag anser att det är en plikt, åtminstone för mig, att förkasta allt hyckleri.
Problemet har mycket djupa rötter. Palestiniernas legitima och heliga rätt till en fri stat är förknippad med Israels lika heliga rätt till erkännande, och vi vet att Israel har raderats från kartan i många länder.
Vi vet att Frankrike, Italien, Spanien och Tyskland absolut inte skulle ha accepterat att bli utraderade från kartan. De skulle inte ha accepterat att betraktas som icke-befintliga.
Vi vet att det inte var Israel som startade det här femtioelfte kriget och att terrorism fortfarande utgör ett av huvudproblemen.
Jag anser därför, om vi lämnar hyckleriet därhän, att vi är skyldiga att börja tänka på ett annat sätt.
Vi kan inte tro att en dialog med terrorister kan motiveras med att så många civila har omkommit, för det skulle medföra en anledning för alla terrorister att i framtiden använda våld, tvång och död för att nå politisk legitimitet.
Jag anser att vi inom Europeiska unionen till slut bör agera mer konsekvent och finna förmågan att hantera problemet med ekonomiska relationer med länder som inte erkänner Israel och tillhandahålla humanitära korridorer så att civila, både palestinier och israeler, kan känna sig trygga.
I det här fallet lider palestinierna mer, och med det vill jag säga att jag anser att det också vore riktigt att se över stödet som vi har gett och som vi ger för närvarande, men som vi inte har någon kontroll över.
Herr talman, mina damer och herrar! Situationen är så man kan gråta.
Hoppet om fred och säkerhet för dem som är berörda gick upp i rök i Gaza och försvann under liken, under barnens, kvinnornas, männens och de skadades kroppar.
Vi står längre än någonsin från hoppet om säkerhet.
Alla som tror att kriget, enligt israelernas logiska argument, är ett krig som motiveras av ett raketanfall mot Israel och att palestinierna måste lära sig läxan, har inte förstått något alls.
De har inte förstått något alls, för att lära någon läxan är ett sorgligt sätt att utbilda dem och det har aldrig fungerat.
Sedan Clausewitz tid vet vi att den som startar ett krig måste kunna avsluta det, måste veta vad syftet är.
Nåväl, syftet med kriget är ökad säkerhet för Israel.
I dag kan vi säga att krigets syfte aldrig kommer att nås genom det här kriget och det sätt som det utkämpas på.
Ju fler civila som dödas, ju fler palestinier som dödas, desto mindre säkerhet i regionen!
Där är dramat, tragedin som för närvarande utspelas i regionen.
Och därför måste vi vara väldigt tydliga.
Martin Schulz har rätt. Israel måste skyddas mot sig självt!
Israel måste räddas från frestelsen i en lösning som innebär krig och väpnad styrka.
Palestinierna måste skyddas mot Hamas.
Palestinska civila måste skyddas mot Hamas.
Det är vår uppgift.
Det är inte lätt, men vi måste vara tydliga.
Jag uppmanar rådet att sluta tänka i termer av uppgraderade, djupare, förbättrade relationer med Israel samtidigt som situationen förblir som den är.
Det är en klen lösning, det är inte den rätta lösningen!
(Applåder)
Jag uppmanar alla som förespråkar en dialog, en diskussion med Hamas, att inte vara naiva, att komma ihåg att en diskussion måste äga rum med Hamas för att förbättra situationen i Gaza, eftersom de har makten, men samtidigt vara medvetna om att Hamas strategi kräver förluster.
Israel har fallit i Hamas fälla: ju fler döda i Gaza, desto bättre för Hamas.
Det är en av de sanningar som vi också måste säga till Hamas.
Vi vägrar acceptera Hamas självmordsstrategi som går ut på att skapa offer och martyrer i syfte att utlösa attacker mot Israel.
Vi måste tala om detta för Hamas också.
Slutligen vill jag säga något till er. De enda som kan lösa problemet med Hamas är palestinierna.
Så länge Israel fortsätter att ockupera Västbanken, så länge Israel misslyckas med att erbjuda en positiv lösning till palestinierna på Västbanken, så kommer allt fler palestinier att vända sig till Hamas.
Om vi ger palestinierna på Västbanken ett hopp om liv så kommer de att resa sig mot Hamas och de kommer att befria oss från Hamas.
Befria palestinierna från Israels ockupation av Västbanken och palestinierna kommer att befria sig själva från Hamas.
(Applåder)
för GUE/NGL-gruppen. - (IT) Herr talman, mina damer och herrar! Rahed är 50 år gammal, han har förlorat sitt hem, sina tre barn, sin hustru och två svägerskor.
Rahed är förtvivlad och befinner sig i det center som vi besökte.
Han sa i djup förtvivlan att Hamas kommer att säga att de har vunnit när anfallet är över, och Israel kommer att säga att de har vunnit, men i verkligheten är det vi civila som är döda. Jag skulle vilja säga en sak till.
Med liken av kvinnor och barn som vi såg och med över 4 000 skadade på sjukhus utan behandling, är det faktiskt rättvisan som håller på att dö. Drömmen om ett Europa som strävar efter mänskliga rättigheter för alla håller på att dö, och det är en tragedi!
Vi är ineffektiva.
Fru Ferrero-Waldner! Ni vet att jag har stor respekt för er och jag vet att ni vidtar åtgärder och arbetar med andra för att nå resultat.
Jag anser att vi tydligt och klart måste förstå att det militära kriget, militarismen från Israels sida, inte leder till Israels räddning, utan till landets undergång, inklusive dess moraliska undergång.
Det är det som David Grossmann säger, dessutom, när han firar minnet av Yitzhak Rabin som dödades av en judisk fundamentalist, inte en islamisk fundamentalist, för att han ville uppnå fred.
Se till att det blir eldupphör!
Se till att det blir eldupphör!
Det är vad den norske läkaren sa till mig, han som opererar varje dag och arbetar dygnet runt (vi skickar läkare till Gaza).
Ett eldupphör är vad vi vill ha!
Säkerhetsrådet måste börja omvandla sina ord till konkreta handlingar.
Vi är överens om diplomati, men vi kan inte bara använda diplomati, utan vi måste använda alla instrument som vi har.
Ett instrument som vi har i förhållande till Israel är uppgraderingen, och jag är glad över att höra att Europeiska kommissionens representant i Tel Aviv i dag sa, till exempel, att tiden inte är inne att tänka på uppgradering.
Vi bör göra ett uppehåll, för vad vi verkligen måste få till stånd är ett eldupphör.
Det är oerhört viktigt.
Jag anser att det är viktigt, och det är ett starkt budskap.
Ni talade om beskydd och internationellt beskydd.
Jag anser att det är fel att bara tänka på Gaza och Rafah.
Beskydd av civilbefolkningen kommer norrifrån, det kommer från de israeliska attackerna som kommer från Herez.
Gränskontroll är kontroll av de viktigaste gränserna, Rafah och Herez, för under lång tid, sedan 1992, sedan Osloavtalet, som ni väl vet, har palestinierna inte haft möjlighet att ta sig ut genom Herez. Inte ens sjuka kan ta sig ut den vägen.
Vi måste därför tänka inte bara i termer av tunnlar och vapen med vilka Hamas kan beväpna sig, utan i termer av absolut alla förbud som finns för palestinierna.
Vi behöver ett eldupphör och öppnandet av inte enbart humanitära korridorer, utan öppnandet av alla gränsövergångar, för om folket inte har mat att äta, om folket inte kan handla, vad kan då göras?
Det skulle vara en riktigt allvarlig påtryckning på Hamas att upphöra med sin existens och att upphöra med sina anfall som skadar den israeliska befolkningen.
Men Israel bör veta att det är Västbanken som är militärt ockuperat och Israel bör verkligen söka fred i stället för att bygga nya bosättningar.
(Applåder)
Tack så mycket, fru Morgantini.
Jag vill uttrycka all min respekt till er och övriga ledamöter som tog initiativet och nyligen reste till Gazaremsan.
för IND/DEM-gruppen. - (NL) Herr talman! Palestina är islamiskt territorium, det kan inte ifrågasättas.
Sedan den islamiska rörelsen Hamas inrättades 1987 har den stått fast vid den grundprincipen.
I detta avseende får den fullt stöd av den islamiska republiken Iran.
Den ideologiska ståndpunkten lämnar absolut inget utrymme för den judiska staten Israel i Mellanöstern, och de skadliga konsekvenserna av muslimsk totalitarism märks på ett grymt sätt i Gazaremsan.
Typiskt för Hamas filosofi är att använda moskéerna i Gaza för militära ändamål, med alla tragiska följder det innebär.
Jag skulle här vilja referera till den klarsynta rapporten i förra måndagens Frankfurter Allgemeine.
Om Europa verkligen värdesätter en fortsatt existens för den judiska staten Israel, lutar det åt en konfrontation mellan Hamas och dess allierade Hizbollah i Iran.
Är vi redo att samla oss inför dessa bistra, om än realistiska, utsikter?
När allt kommer omkring är ett eldupphör eller en tillfällig vapenvila för Hamas och kompani endast en andningspaus i jihad mot Israel.
(IT) Herr talman, mina damer och herrar! Jag måste säga att jag tror att den stora majoriteten av oss i kammaren delar önskemålen om fred och den oro som många av oss här hittills har uttryckt.
Jag tror också att vi kan skriva under det som rådet sa, och jag skulle vilja säga att kommissionen hittills har följt en väg som kan gynna dialog: öppnandet av humanitära korridorer och bilateralt eldupphör kan förebåda ett åtagande att inrätta en internationell säkerhetszon.
Här har kanske Luisa Morgantini rätt när hon efterfrågar att zonen inte bara ska relatera till Gaza, utan bör utvidgas till alla palestinska territorier.
I grunden har jag intrycket att önskemålen och Benita Ferrero-Waldners diplomatiska aktivitet åtminstone i visst avseende kan ses som att hon intar samma hållning i frågan som påven.
I all ödmjukhet önskar jag dela denna typ av hållning: efter alla dessa år måste vi fortfarande söka efter en lösning för två folk och två stater - det är en punkt som vi inte får glömma - och vi måste slutligen sträva efter att följa internationell lagstiftning.
Det finns ingen militär lösning och det kommer aldrig att finnas någon - Martin Schulz sa det också - emellanåt måste jag hänvisa även till honom - och jag måste säga att problemet i det heliga landet utan tvekan aldrig kommer att lösas militärt.
På den punkten tror jag att Europeiska unionen har verktygen för att stödja vilka diplomatiska ansträngningar som än görs här.
Jag är övertygad om att Martin Schulz kommer att bli nöjd med att höra att ni nämner hans namn i samband med den helige Fadern!
(DE) Herr talman, fru kommissionsledamot, herr rådsordförande! Jag skulle vilja beskriva min utgångspunkt.
Hamas motsätter sig en tvåstatslösning, förkastar statens Israels rätt att existera, har kommit till makten genom en brutal kupp mot sitt eget folk, avfyrar raketer mot civila och använder civila, skolor och moskéer som mänskliga sköldar.
När man försöker skydda sin egen civilbefolkning, hur är det möjligt att reagera proportionellt om den andra sidan använder sin egen civilbefolkning som mänskliga sköldar?
Principen att jämföra antal och proportionalitet är därför inte tillämplig i en situation som denna.
I en krigssituation finns ingen proportionalitet - varje krig och varje skadad är ett eller en för mycket och det är omöjligt att svänga sig med siffror för den ena sidan eller mot den andra.
För mig förefaller detta vara utgångspunkten.
Vi ska därför inte ägna oss åt den här typen av fingervisning som vi har sett, utan i stället försöka få till stånd ett eldupphör och se till att hjälpa till i det avseendet.
Jag tror att rådets tjänstgörande ordförande Karel Schwarzenberg och hans delegation, och även kommissionsledamot Benita Ferrero-Waldner, med hjälp av andra nationella delegationer har gjort mer än någon annan part, och det vill jag uppriktigt tacka dem för - jag har inte sett några tecken från Förenta staterna, knappt något tecken från FN och inget tecken från övriga medlemmar i kvartetten.
Vi måste se till att eldupphöret omfattar två aspekter: Israels attack måste upphöra och Hamas måste hindras från att lägga vantarna på nya raketer från Korea och Iran, som skulle sätta Tel Aviv inom räckhåll.
Av den här anledningen måste man inte bara se till att eldgivningen upphör utan också, genom internationella avtal som omfattar kvartetten och arabförbundet, med Egypten i nyckelpositionen, se till att den 15 kilometer långa gränsen patrulleras i en omfattning så att inga fler skott kan nå Gaza.
Samtidigt måste den israeliska attacken stoppas.
Jag skulle vilja göra en sista kommentar.
Det här är bara ett första litet steg.
Om Israel önskar förhandla med moderata palestinier i framtiden - vilket skulle innebära en tvåstatslösning - då, när allt det här är över, måste man se till att moderata palestinier som stödjer president Abbas äntligen kan uppvisa resultat för sitt eget folk, vilket betyder ett stopp för bosättningspolitiken och många andra saker.
När allt kommer omkring kommer radikalerna att segra om de moderata krafterna inte har några framgångsrika resultat att visa sitt folk.
Det här måste bli utgångspunkten för en ny israelisk politik.
(IT) Herr talman, mina damer och herrar! Inför denna ofantliga tragedi är våra ord troligen otillräckliga.
En armé som dödar hundratals civila, kvinnor och barn placerar sig själv på samma nivå som den terrorism den hävdar att den bekämpar.
Å andra sidan så vet alla som känner till Gaza, även om man bara sett området på en karta, att ingen militär operation kan planeras utan att man medger att följden troligen blir en massaker på civila.
Kan Israel säga att landet i dag är säkrare, efter att ha åstadkommit så mycket hat och förtvivlan?
Om inte med Hamas, direkt eller indirekt, så med vem ska man söka en väg bort från det blinda våldet?
I vår resolution stärker vi den uppmaning till eldupphör som Förenta nationernas säkerhetsråd tidigare uttryckt.
Vi uppmanar parterna att följa den och vi uppmanar Europa att vidta åtgärder så att det blir möjligt.
Risken, herr Brok, är att massakern, långt ifrån att besegra Hamas, kommer att försvaga den palestinska myndigheten ytterligare och också de i den palestinska världen som har satsat allt på förhandlingar med Israel.
Vi måste fråga oss själva ärligt vad de hittills har vunnit?
Ingenting.
Det är svaret som vi måste ge om vi verkligen vill börja utrota hatet och våldet.
- (FR) Herr talman! Vi är alla delvis ansvariga för vad som händer i dag i Mellanöstern.
Vi i Europa och vi i det internationella samfundet har tillåtit situationen att förvärras. Vi gjorde ingenting när Israels säkerhet hotades och vi gjorde ingenting när blockaden gjorde livet i Gaza fullständigt omöjligt.
I dag är det krigets nittonde dag; 995 människor har dödats, varav 292 barn, och tusentals har skadats, varav några fortfarande väntar på att evakueras.
Det finns tio tusentals flyktingar som inte har något hem längre och inte vet vart de ska ta vägen.
Den humanitära situationen förvärras allt mer: 700 000 invånare i Gaza har inte längre någon elektricitet, en tredjedel av dem har inte längre vatten eller gas, och snart är det tre veckor sedan denna situation började, tre veckor under vilka folket har levt eller snarare gjort sitt bästa för att överleva.
Det finns för mycket lidande, för många prövningar, och det måste få ett slut, det måste sluta nu!
Vårt ansvar gentemot oss själva, som européer, är inte att tillmötesgå någon.
Vårt ansvar gentemot oss själva, som européer, är att sätta press på bägge parter så att de till slut går med på förhandlingar.
Det är en fråga om dagar, kanske rentav timmar, innan det inte finns någon väg tillbaka, när det blir en landoffensiv, i synnerhet i Gaza stad.
Israels säkerhet måste garanteras och befolkningen i Gaza måste garanteras ett framtida liv i fred.
Gränserna måste övervakas och blockaden måste hävas.
Vi vet alla att en förutsättning för att nå det avtalet kanske är att Europa, Förenta staterna och arabstaterna - som träffas i övermorgon - agerar samfällt.
Innan jag slutar skulle jag vilja uttrycka min starka övertygelse. Det är inte kriget som måste vinnas, utan freden.
(Applåder)
(IT) Herr talman, mina damer och herrar! Jag välkomnar verkligen kommissionsledamotens och Hans-Gert Pötterings kommentarer, som i tydliga ordalag fördömer och lägger ett tungt ansvar på Hamas för att ha brutit vapenvilan, men som också tydligt fördömer Israels oproportionerliga reaktion.
Men bakom orden kvarstår krisen och tusentals människor - den civila befolkningen och barn - som är i desperat behov av humanitärt bistånd.
I vårt samvete och utan hyckleri borde vi kanske ställa oss några frågor.
Hur många barn dog i Gaza medan våra barn firade jul?
Två eller tre hundra. Och hur många israeliska civila?
Skulle det internationella samfundet ha kunnat göra mer?
Jag anser att svaret är ja.
Mer borde ha gjorts.
Vi måste ta vårt fulla ansvar.
Det räcker inte att tv-sända åsikter om Hamas, om Israel, om det ursprungliga ansvaret eller om vem som bär skulden.
Utöver krissituationen är Europa tyvärr fortfarande otillräckligt.
Jag anser att det är en allvarlig svaghet. En oförmåga att bygga upp en verklig, strategisk och hållbar fredspolitik.
I dag måste vi utfärda en tydlig begäran om eldupphör, men det räcker inte.
Vi måste lägga fram stränga villkor för freds- och utvecklingsprocessen i Mellanöstern.
Slutligen skulle jag vilja hänvisa till påvens ord, nämligen att vi måste ge specifika svar till de allmänna förhoppningar, som många i dessa länder har, att få leva i fred, trygghet och dignitet, så som Luisa Morgantini också betonade.
Jag avslutar nu.
Våld, hat och misstro utgör olika former av fattigdom - kanske de värsta att bekämpa.
- (FR) Herr talman! I Gaza har vi sett krig och död, men vi har också sett människor, levande människor som har rätt att leva och som det är vår uppgift att skydda.
Att skydda civilbefolkningen är det som är det viktigaste.
Det finns inga ursäkter för det faktum att vi inte har gjort allt för att skydda befolkningen och jag vill fråga er, herr rådsordförande, om ni i dag anser att ni har gjort allt ni kan för att se till att de israeliska myndigheterna omedelbart upphör med denna urskillningslösa och oproportionerliga militära operation?
Svaret är med säkerhet nej.
När rykten om operationen florerade på ambassaderna bekräftade rådet på nytt, mot parlamentets önskan, sin beslutsamhet att intensifiera förbindelserna.
Detta var ett tragiskt misstag!
När icke-statliga organisationer uppmanar säkerhetsrådet att låta internationella brottmålsdomstolen utreda påstådda krigsförbrytelser är rådet oförmöget att åberopa klausulen om mänskliga rättigheter i avtalet med Israel.
Jag är trött på att höra att vi inte kan göra något mer, att vi har gjort allt vi kan.
Det största misslyckandet är i själva verket dödläget i er i grund och botten humanitära politik för att lindra den skada som den militära ockupationen och kriget orsakat.
Hur långt ska vi låta det gå när det gäller brott mot internationell rätt innan vi ser till att klausulen om mänskliga rättigheter tillämpas?
Om vi inte i dag kan ställa frågor om räckvidden för effektiva mekanismer när det gäller utövande av påtryckningar och genomförande vet jag sannerligen inte vilken slags situation som skulle kunna rättfärdiga att vi äntligen vidtar åtgärder.
Jag säger det rent ut: Om strategin att låta allt fortsätta som vanligt fortsätter att vara del av våra förbindelser med Israel kommer ni, genom de 1000 dödsfallen i Gaza, att begrava artikel 11 i fördraget samtidigt som ni begraver unionens politik för mänskliga rättigheter och det europeiska projektet!
(Applåder)
(EN) Herr talman! Efter att ha återkommit från Gazaremsan, där jag sett massakern på framför allt civila, känner jag att jag måste uttrycka min helhjärtade solidaritet med det palestinska folket.
I 17 dagar har de ställts inför den enorma israeliska krigsmaskinen, som på ett flagrant sätt bryter mot internationell rätt.
Jag vill också uttrycka mitt stöd för fredsrörelsen i Israel som vill ha ett slut på kriget.
Efter en lång avstängning och belägring, som förvandlade Gaza till det största öppna fängelset i världen, byggandet av den skamliga muren runt Västbanken, den fortsatta utvidgningen av bosättningarna och den effektiva uppdelningen av palestinsk mark har de ockuperande styrkorna övergått till en våldsam militär operation.
I det här sammanhanget användes raketattackerna mot södra Israel - och jag vill betona att jag är emot alla attacker från båda sidor mot civila - som en förevändning.
Att eldupphöret bröts mot bakgrund av maktspelet i samband med det israeliska valet är en förolämpning mot hela landet.
FN:s säkerhetsråd har antagit en resolution.
Israel är en stat, inte någon organisation - landet är medlem av Förenta nationerna.
Landet har ett ansvar gentemot det internationella samfundet och måste följa denna och andra resolutioner som antagits av Förenta nationerna.
Den internationella rätten måste respekteras.
Straffrihet ska inte längre tillåtas.
En fullständig internationell undersökning måste genomföras.
Det internationella samfundet kräver ett omedelbart eldupphör, att de militära styrkorna omedelbart dras tillbaka, tillgång till humanitärt bistånd och rörelsefrihet för befolkningen.
Låt UNWRA genomföra sitt uppdrag.
EU har vidtagit åtgärder, men bara på humanitär nivå.
EU måste visa handlingskraft på politisk nivå.
Använd klausulerna i associeringsavtalen.
Sluta uppgradera relationerna med Israel.
Stoppa vapenexporten till Israel.
Det kan bara finnas en politisk lösning på den här konflikten.
En fullständig återgång till internationell rätt måste genomföras, vilket innebär att den 42 år långa ockupationen av Palestina måste upphöra och en självständig och livskraftig palestinsk stat etableras. På så sätt kan en fredlig framtid byggas upp för såväl palestinska som israeliska barn.
För att rädda framtida generationer måste vi stoppa kriget nu.
- (FR) Herr talman! För flera tusen år sedan konfronterade David Goliat för att få klarhet i huruvida landet var avsett för moabiterna, filistéerna eller hebréerna.
Just nu utspelas samma drama i detta land som är källan till en av vår civilisations tre pelare.
I dag är det angeläget, rätt, berättigat och nödvändigt att garantera säkerhet för och erkännande av staten Israel.
För att lyckas med detta krävs det en lösning, nämligen att garantera att en suverän palestinsk stat upprättas.
Här, precis som på andra områden, finns det en gräns för multikulturalismen.
Där det finns två befolkningar måste det finnas två stater.
Om Europeiska unionens bistånd ska vara effektivt måste det fokuseras på ett mål: att garantera att denna palestinska konstitutionella stat utvecklas och att rättssäkerheten fungerar som ett skydd för de svaga och en hjälp för de starka.
Detta brådskar eftersom extremisterna på alla sidor är mäktiga och orättfärdiga, medan barnen är offer.
Lösningen när det gäller att distansera sig från kravet ”öga för öga” är vare sig moralisk eller militär utan politisk.
Så det är dags att sätta i gång med arbetet!
(EN) Herr talman! Jag avskyr terrorism.
Jag avskyr terrorismens propaganda.
Jag är kanske mer medveten om detta eftersom jag kommer från Nordirland och när jag hör Hamas utgjuta sig över de nödvändiga vedergällningarna för åratal av urskillningslösa raketregn över oskyldiga medborgare i Israel blir jag inte berörd, eftersom jag vet att Hamas, i likhet med IRA i mitt land, är mästare i de besläktade konstarterna terrorism och propaganda.
Situationen är mycket tydlig.
Israel accepterar en tvåstatslösning.
Hamas kan inte ens tolerera Israels rätt att existera och genomför därför oupphörliga, obarmhärtiga terroristattacker på landets territorium.
Och när Israel, efter att ha visat stor fördragsamhet, slår tillbaka menar Hamas att det är de som är offret.
Tyvärr: det är de som är gärningsmännen och om de vill ha fred ligger svaret i deras egna händer.
Sluta bomba Israel.
(EL) Herr talman! Vi inser alla att situationen i Gaza är tragisk.
Vi står på tröskeln till en humanitär katastrof som kräver omedelbara åtgärder.
Jag vill gratulera Europeiska kommissionen till att ha ökat sina insatser, ordförandeskapet till dess initiativ och till att ha samordnat de nationella åtgärder som vidtas och Egypten till den viktiga och lyhörda roll landet spelar.
Behovet av eldupphör och av att fientligheterna på båda sidor upphör, av korridorer från det israeliska territoriet, av att Egypten tar itu med de humanitära behoven och av gränskontroller för att sätta stopp för den olagliga förflyttningen av vapen och människor är brådskande.
Som kommissionsledamoten sa är det uppmuntrande att det finns tecken på en plan för vapenvila och jag hoppas att den kommer att godkännas omedelbart och respekteras i praktiken.
Så hur ska vi agera härnäst?
Både kommissionsledamoten och rådets ordförande har redan sagt att vi måste främja våra mål för en genomförbar fred och skapandet av en palestinsk stat som existerar i fred och respekt bredvid Israel.
De är inte nya.
Vi har tillkännagivit dem och vi har försökt främja dem utan resultat.
Den onda cirkeln av våld fortsätter med negativa konsekvenser, inte bara för människorna i Israel och för palestinierna, utan för alla människor i området och för det internationella samfundets säkerhet.
Nu måste vi granska våra åtgärder, våra politiska val och våra metoder och vidta andra modigare åtgärder.
Det är angeläget att vi självkritiskt inleder en ärlig, ingående dialog på bilateral nivå med Israel inom ramen för våra vänskapliga förbindelser och vårt partnerskap och att vi identifierar de misstag som gjorts i främjandet av ömsesidig tillit mellan dessa båda folkgrupper.
Vi måste även stärka dialogen med alla palestinier, för att få dem att förstå vikten av fred, sammanhang, mänskligt liv och enighet mellan dem.
(DE) Herr talman! Efter premiärminister Topoláneks skämtsamma kommentarer i dag vill jag säga att jag som österrikisk parlamentsledamot är nöjd med att både kommissionen och det tjeckiska ordförandeskapet representeras av österrikare.
Ni är varmt välkommen!
Herr rådsordförande! Jag inser naturligtvis att er lojalitet finns hos Tjeckien.
När jag en kort tid före Israels ensidiga tillbakadragande från Gazaremsan reste till landet, som medlem av en delegation där Martin Schulz var ordförande, sa den dåvarande biträdande premiärministern: ”Lägg er inte i, det här kommer att fungera bra”.
Andra, däribland den tidigare utrikesministern Josip Elin, sa: ”Detta kommer att leda till kaos”.
Det finns ingen mening med ett ensidigt tillbakadragande, utan förhandlingar och utan att ha en förhandlingspartner.
Det var emellertid inte heller särskilt klokt av oss att besluta oss för att inte inleda en dialog ens med sansade företrädare för Hamas. Dessa kanske inte ens tillhörde Hamas, men Hamas hade nominerat dem till den gemensamma regeringen.
Genom att inta denna ståndpunkt bidrog vi till att denna gemensamma regering upplöstes.
Jag vet att det fanns vissa här som ville genomföra samtal, men som inte tilläts göra det - även detta var ett misstag.
Vi behöver en dialog!
Jag tycker inte om Hamas. För det första eftersom det är en terroristorganisation och för det andra på grund av dess fundamentalistiska åsikter, men detta handlar inte om att tycka om eller att tycka illa om något - det handlar om att hitta lösningar.
Därför måste vi återgå till dialog och samtal, precis som många av våra parlamentskolleger redan har sagt i dag.
Dessutom måste människorna i Gaza få chansen att leva ett någorlunda anständigt liv.
Varför röstar de på Hamas?
Svaret är att de ser dem som sin enda chans, sin sista chans, att ens överleva - och detta måste förändras.
Vi måste även erbjuda dessa människor ett ekonomiskt underlag så att de kan överleva. Vi måste häva bojkotten och se till att deras isolation upphör.
Detta är det enda riktiga kravet.
Elmar Brok, som jag hyser stor aktning för, sa att proportionalitetsprincipen inte var tillämplig - men detta är inte sant.
Proportionalitetsprincipen kan tillämpas på såväl privat som internationell rätt.
Den som bryter mot den bryter även mot internationell rätt - och det är något som parlamentet verkligen inte kan acceptera.
(Applåder)
(EN) Herr talman!
En vän som vet att jag var i Gaza för bara tre dagar sedan ställde en fråga till mig. ”Har du aldrig sett bilderna av femåriga judiska barn som står framför nazisternas gevär med händerna i luften?”, skrev hon. ”Det är fruktansvärda bilder.”
Hennes ord illustrerar varför vi gör eftergifter för Israel som vi inte skulle göra för något annat land.
Det förklarar dock inte varför ett folk som har lidit så mycket under 1900-talet nu utsätter andra människor för så mycket lidande under det här århundradet. Israel har gjort Gaza till ett helvete: marken skakar av explosioner, också under ett eldupphör.
Åsnekärror kör på gatorna och F-16-plan flyger i luften ovanför, 2000-talets dödsmaskiner som släpper ner bomber. 300 barn har redan dödats, ytterligare hundratals har slitits sönder i bitar.
Detta är inte ett proportionerligt svar från en civiliserad stat.
Det är ren ondska.
Det är ren ondska.
Ja, Hamas raketbeskjutning måste upphöra.
Det har jag själv sagt till Hamas representanter i Gaza tidigare, men låt oss slippa det skenheliga talet från israeliska företrädare om behovet av att bekämpa terrorismen. Palestinierna som bombas skulle också kunna peka ut terrorister och de namn de skulle nämna är Olmert, Livni och Barak.
Vi har ett visst ansvar för Israels handlingar.
EU har aldrig, i varje fall inte som jag kan minnas, backat upp sin kritik av israelernas behandling av palestinierna med någon form av handling.
Vi ger Israel grönt ljus att fortsätta som de vill och vi förstärker detta genom att strunta i det man kan lära av historien.
Man kan inte uppnå fred utan att tala med fienden, ändå vägrar vi att tala med de folkvalda företrädarna för det palestinska folket.
Nu slutförhandlar vi med Israel om ett utökat samarbetsavtal.
Vi har inga planer på att fördöma Israel: vi tänker belöna landet.
De som vill ha fred i Mellanöstern, de som vill se rättvisa för båda sidor, måste inse att det är dags att tänka om.
- (GA) Herr talman! Kriget i Gaza är skrämmande och skandalöst.
Alla vet att en militär lösning inte kommer att fungera i Mellanöstern.
En politisk lösning är det enda sättet att återupprätta fred och försoning i detta område.
För att detta ska kunna ske måste våldet upphöra omedelbart.
Jag stöder skapandet av en självständig och bärkraftig palestinsk stat, men detta kräver en tillräckligt god ekonomi och en ordentlig politisk plan.
Det bör vara vår målsättning att se till att dessa båda stater kan existera i regionen och att de respekterar varandra.
Israel har rätt att skydda sig självt, men landet har gått för långt med dessa attacker.
Attackerna är omoraliska och det internationella samfundet kan inte acceptera dem.
Fredsprocessen i Mellanöstern måste genomföras omedelbart.
Jag hoppas att USA:s nyvalde president, Barack Obama, kommer att arbeta med detta.
Vi önskar honom lycka till med denna viktiga uppgift och med den utmaning han har framför sig.
(ES) Herr talman! Även jag var i Gaza för några dagar sedan och det var en mycket intensiv upplevelse.
Vi reste även till Egypten.
Jag anser att vi befinner oss i slutet av en era, Bush-eran, och att de sista av president Bushs kval har visat sig vara särskilt blodiga och smärtsamma.
Vi har nått en vändpunkt där vi kan anta en annan Mellanösternpolitik och där vill jag att Europeiska unionen ska ta initiativet.
President Obama ger uttryck för samma ståndpunkt när han säger att kan kommer att tala med Iran.
Ja, president Obama kommer att tala med Iran och vi måste tala med alla, inklusive Hamas, i Mellanöstern.
Den nya Mellanösternpolitiken måste vara en samarbetsinriktad politik som överensstämmer med våra värderingar och med internationell rätt.
De hundratals barn vi såg i Gaza, som klängde sig fast vid våra armar och såg på oss med ögon fulla av hopp, förtjänar ett svar, precis som barnen i Israel.
Detta kräver konkreta åtgärder, det kräver åtgärder på plats, för att ge hopp till de sansade.
Den mest beklagliga aspekten är att premiärminister Fayad, president Abbas, president Mubarak och kung Abdullah nu anklagas för förräderi på gatorna i arabvärlden.
När jag under en taxiresa gjorde ett uppehåll i Sinaiöknen för att dricka kaffe var Khaled Meshaal det enda jag såg på de stora skärmarna.
Detta är resultatet och de oavsiktliga skadorna av attacken mot Gaza.
Den kommer inte att leda till fred för Israel eller till den trygghet vi vill ha, än mindre till någonting bra för oss.
Om vi inte sätter stopp för denna konflikt kommer den att leda till att hatet sprids till Europas egna gator.
(PT) Ettusen är dagens siffra, ettusen dödsfall som ger oss en dyster lärdom.
Ursäkta min rättframhet, men hur många fler liv kommer det att krävas för att välja Tzipi Livni och Ehud Barak i valet i februari?
Vi är här i dag för att kräva eldupphör och ett slut på slakten av civila.
Resolutionen väcker emellertid även frågor om vårt eget ansvar.
Den påminner oss om att rådet beslutade att uppgradera de diplomatiska förbindelserna med Israel, i strid med parlamentets åsikt.
Detta var delaktighet genom föregripande.
I dag hör jag: ”Det är nödvändigt att tala med Hamas”.
Vi kunde ha sparat år om vi hade respekterat valen i Palestina.
Europas roll handlar inte om att stödja politikerna och den ödeläggelse som den starkare sidan orsakar.
Den handlar om att lyssna på de protester som gatorna och torgen i våra städer fylls av.
Vi kräver ett eldupphör nu, men vi måste inse att ockupationen måste upphöra för att fred ska kunna uppnås.
Detta ord har missbrukats, men det måste tas bort från listan över förbjudna ord där mäktiga politiker placerat det.
(EN) Herr talman! Det som händer i Gaza är hjärtskärande.
Att förödelsen vidmakthålls av en förment västerländsk nation är ofattbart.
Jag håller helt och hållet med om att israelerna har rätt att leva utan hotet om raketattacker.
Men det som händer i Gaza är inte rättvisa: det är slakt.
Det finns ingen ursäkt. Det går inte att rättfärdiga.
Det mest skamliga för oss inom EU är att det genomförs av en av våra främsta handelspartner.
Under 2007 uppgick värdet av handeln mellan EU och Israel till 25,7 miljarder euro.
Med tanke på den stora mängd pengar vi bidrar med till Israels ekonomi har vi ett tungt ansvar när dessa pengar också bidrar till att civila och barn dör.
Om vi inte agerar kommer blodet från människorna i Gaza att fläcka även våra händer.
Jag vill uppmana parlamentet och alla EU-organ att omedelbart införa handelssanktioner mot Israel och att behålla dem till dess att ett verkligt eldupphör kommit till stånd.
Om vi inte gör vårt allra yttersta för att stoppa detta dödande blir vi medskyldiga till slakten.
- (FR) Herr talman! Återigen är det vapnen som talar i Mellanöstern.
Återigen är de huvudsakliga offren kvinnor, barn, varav tusentals har skadats och hundratals dödats.
Återigen upprepar sig historien med all dess ohygglighet på tröskeln till Europa.
Vi konstaterar dock att Europa, trots dess initiativ, inte bidrar på ett effektivt sätt i denna stora konflikt, trots att den äger rum i ett område som Europa har inflytande över.
En överväldigande majoritet av allmänheten upplever att detta är svårt att förstå och de vägrar i allt större utsträckning att acceptera sådan maktlöshet.
Fru kommissionsledamot! Vi måste kraftfullt och myndigt ta på oss ledarskapet för att skapa fred.
Unionen för Medelhavet måste spela en viktig roll, liksom den parlamentariska församlingen för Europa-Medelhavsområdet.
I enlighet med detta måste Europaparlamentet stödja den fransk-egyptiska fredsplanen för ett omedelbart eldupphör, skydd av gränserna mellan Israel och Gazaremsan, öppnande av gränsövergångsställena och framför allt upphävande av blockaden mot Gaza.
Vi måste även kräva en omedelbar tillämpning av FN-resolutionen.
När detta första skede är över måste vi gå vidare genom att föreslå en militär styrka, inte en multinationell styrka utan en styrka från Europa-Medelhavsområdet.
Genom denna gest skulle vi bekräfta vår politiska vilja att uppnå en ”europeisk fred”, något som alla människor i Medelhavsområdet har väntat så länge på.
Jag vill även uppmärksamma er på en ny situation.
Genom konflikten i Mellanöstern går vi steg för steg in på ett mycket farligt område, nämligen sammandrabbningar mellan civilisationer.
Ända sedan konflikten mellan israeler och palestinier tog sin början har det funnits underströmmar av en allmän arabisk opinion.
I dag är det en muslimsk allmän opinion som sträcker sig långt bortom Arabländernas gränser.
Detta tyder på en radikal förändring av konfliktens karaktär.
Europa har ett historiskt ansvar som handlar om att enträget stärka dialogen mellan civilisationer.
Jag har här i parlamentet så många gånger sagt att vi bör utnyttja varje möjlighet till fred, hur liten den än är, och att vi trots allt som hänt bör tala med Hamas, eftersom de vann valet. Jag vill därför inte återkomma till denna fråga.
Jag är utom mig av sorg och ilska och samtidigt som jag i dag inte vill tillåta mig själv att överväldigas av känslor när jag ställs inför denna massaker, denna krigspropaganda som jag hör runt omkring mig, denna förvirring och denna våg av hat och antisemitism som börjar sprida sig på våra gator, har jag något jag vill säga: Europa måste börja om från början och för mig är dessa fakta självklara, men ibland är det bra att poängtera dem.
För det första är en palestiniers liv lika mycket värt som en israels liv, men inte bara hans liv utan även hans framtid och frihet.
För det andra måste internationell rätt respekteras och internationell rätt innebär naturligtvis ett omedelbart eldupphör.
Det finns många FN-resolutioner och Genèvekonventioner.
Faktum är att detta område i dag har blivit ett laglöst område där allt tycks vara tillåtet och där en befolkning hålls som gisslan.
För det tredje måste rättvisa skipas för alla dessa brott, oavsett vad de består i och var de begås.
Det kommer aldrig att skapas trygghet utan fred eller fred utan rättvisa.
Övergångsrättvisa finns, den är till för detta och om den inte tillämpas kommer hatet att fortsätta att spridas.
Under de senaste dagarna har vi skapat en kapacitet för hat som kommer att visa sig vara ännu farligare än bomberna.
Europa måste tvinga fram en tillämpning av villkoren i sina partnerskapsavtal, däribland stycke 2 i associeringsavtalet om respekten för mänskliga rättigheter.
Detta är en skyldighet i dessa avtal som det inte kan göras några undantag från.
Sist men inte minst är Israel inte något specialfall utan har sitt ansvar som stat och kan inte vara likställt med Hamas.
När det handlar om internationell rätt finns det inte något ”Du slipper ut ur fängelset”-kort.
På söndagen lämnade vi bakom oss en befolkning i Gaza som var fångad i en fälla, fängslad i ett getto under bomberna, och hundratusentals barn vars framtid i dag ligger i våra händer, och den enda anledningen till att vi kunde ta oss ut ur Gaza var att vi är européer.
De enda palestinierna som lämnar Rafah är de som gör det i ambulans eftersom de är döda eller skadade.
Europa kommer inte längre att vara Europa och ingen medborgare kommer att erkänna sig som europé om vi glömmer dessa grundläggande fakta.
(Applåder)
- (FR) Herr talman, fru kommissionsledamot! Jag vill börja med att upprepa Daniel Cohn-Bendits ord.
I dag grips vi av förtvivlan, detta krig är en tragedi.
Bilderna av lidande och död som oavbrutet har flimrat förbi på våra tv-skärmar i tre veckor är outhärdliga, och det vill jag genast tillägga att alla bilder av krig och alla konflikter är, även dem som det talas allt mindre om, om det överhuvudtaget talas om dem. Några exempel på detta är Kongo, Darfur, Zimbabwe och dessförinnan Tjetjenien, vars fasor ägde rum under en öronbedövande tystnad från medier och, det vill jag framhålla, politiker.
Jag har redan vid ett flertal tillfällen här i parlamentet poängterat det faktum att indignationen hos vissa av mina parlamentskolleger varierar beroende på omständigheterna.
Som Luisa Morgantini ofta har påpekat går det emellertid inte att föra räkenskaper när det handlar om människor som dör, det finns ingen hierarki när det gäller lidande. Varje person som dödas eller skadas, oavsett om det handlar om en man, en kvinna eller ett barn, och oavsett vilken sida offret kommer ifrån, är ett offer för mycket.
Så vad bör vi nu göra för att se till att vår debatt i dag inte blir som den ofta blir - en på något sätt lam och meningslös konfrontation?
Att fortsätta att kasta glåpord efter varandra om de olika parternas historiska ansvar förefaller tycker jag är ett perfekt exempel på sådan meningslöshet.
Jag talar sent i denna debatt, så argumenten har redan nämnts.
Det går att ifrågasätta omfattningen av den israeliska krisen och det israeliska motanfallet, men inte under några omständigheter Israels rätt till säkerhet.
Vilken av våra regeringar i väst skulle finna sig i att se tusentals missiler avfyras mot dess medborgare utan att reagera?
Svaret är självklart.
Utöver uppmaningen om ett nödvändigt framförhandlat eldupphör, och naturligtvis om en garanti om utdelning av humanitärt bistånd och ett slut på leveranserna av vapen via tunnlarna, handlar den faktiska frågan i dag om framtiden.
Fredsfundamentalisterna är välkända. De har redan identifierats vid Taba, Camp David och Annapolis.
Benita Ferrero-Waldner har klargjort detta.
De flesta, men naturligtvis inte alla kort ligger på bordet och detta innebär uppoffringar från båda sidor.
Och när jag talar om uppoffringar är jag överens med Martin Schulz som för närvarande inte befinner sig i kammaren.
Det handlar inte om huruvida en dialog kommer att inledas med Hamas, utan om hur den ska genomföras och på vilka villkor.
De flesta av mina parlamentskolleger har överskridit sin talartid med 50 sekunder, så låt mig avsluta detta, herr talman.
Svaret är det svar som Yasser Arafat gav i maj 1989 när han förklarade sina frihetsförstörande och dödliga stadgar ogiltiga och betydelselösa.
Dessa ord har dessutom blivit en del av det palestinska ordförrådet.
Inter-palestinsk försoning uppnås framför allt till priset av detta, och Europeiska unionens roll är att få förgrundsgestalterna i Palestina och Israel, men även deras arabiska grannar Egypten och Jordanien, att bli samarbetspartner för ett varaktigt fredsavtal.
(Applåder)
(DE) Herr talman! Söndagen den 11 januari besökte vi gränsstaden Rafah på Gazaremsan, som är helt avspärrad.
Detta innebär att civilbefolkningen inte har någon chans att fly från den israeliska arméns dagliga bombarderingar.
Om man inte har sett det med egna ögon går det inte att föreställa sig hur mycket människorna i Gaza lider och hur brådskande det är att nå en fredlig och definitiv lösning på konflikten.
Vi påverkades alla djupt personligt av det oerhörda lidandet hos det palestinska folket och även av förödelsen.
Därför vill jag i starka ordalag upprepa att de israeliska bombningarna måste upphöra omedelbart, precis som Hamas raketeld mot Israel.
Dessutom måste smugglandet av vapen till Gazaremsan från Egypten stoppas. Vidare måste gränserna omedelbart öppnas så att biståndsleveranserna till civilbefolkningen släpps in i området.
Vi träffade även läkare vid gränserna som var redo att resa in i området för att erbjuda hjälp, men som inte kunde det eftersom gränserna var stängda.
Därför vill jag återigen vädja om att gränserna öppnas så att biståndet kan överlämnas.
- (CS) Herr talman! Vem skulle inte lida svåra kval av att se barn dödas av en missil?
Det är en fruktansvärd känsla, men den rättfärdigar inte hyckleri.
Vilka europeiska länder skulle visa lika mycket återhållsamhet som Israel och under flera år finna sig i attacker med fler än 7 000 missiler som hela tiden hotar livet på över en miljon civila?
Invånarna i Gaza är emellertid inte bara oskyldiga offer.
De valde entusiastiskt, medvetet, fritt och demokratiskt Hamas och dess stadgar.
När de talade om befrielse menade de inte befrielsen av Gaza, som redan är fritt, utan om att befria Tel Aviv och Haifa från judar och ödelägga staten Israel.
Det är logiskt att den som väljer brottslingar delar deras öde.
Framför allt när dessa brottslingar gömmer sig bakom kvinnor och barn på samma sätt som de gömmer sig bakom gisslan när de skjuter missiler från skolor och omvandlar moskéer till enorma vapenförråd.
Jag minns bombningen av Dresden 1944 när det brittiska flygvapnet jämnade staden med marken och dödade 92 000 civila, främst kvinnor och barn.
Det förekom inget hyckleri om att man kände anstöt.
Tyskarna valde Hitler av fri vilja och delade hans öde.
Även invånarna i Gaza visste vem de valde och varför.
På samma sätt hamnade en stor andel av de ekonomiska medlen från EU till Gaza i Hamas händer.
Detta kanske var för att invånarna i Gaza, mätta och med stöd av EU, skulle kunna ägna all sin uppmärksamhet åt att gräva tunnlar för att smuggla in allt fler dödliga vapen som används mot den israeliska civilbefolkningen.
Synnerligen proportionerligt!
Herr talman! Det finns två viktiga saker som präglar debatten här idag.
Det ena är att en överväldigande majoritet av detta parlament vill få till stånd ett snabbt eldupphör.
Det andra är att det finns ett överväldigande stöd för att alla parter måste ge staten Israel sin rätt till existens under fredliga gränser.
Detta är en utgångspunkt som är viktig för Europeiska unionen.
Det är viktigt eftersom det är en tragedi som vi ser i Gaza.
Varje liv som går förlorat är en tragedi, oavsett vilken sida om gränsen.
Låt oss inte tro att denna tragedi skulle bli mindre för att de som uppsåtligen vill döda civila skulle lyckas genom raketbeskjutningar ännu längre in bland civila.
Det är en tragedi också för att det skapar hinder för förverkligandet av en palestinsk stat och därmed en fredlig lösning.
Det är en tragedi som också faller på det internationella samfundet, eftersom det som nu händer inte har hänt plötsligt utan har byggts upp genom upprustning, genom smuggling av vapen och genom raketbeskjutning under lång tid.
Det som för oss är viktigt att se är att detta inte är en tragedi som bygger på en konflikt mellan judar och palestinier.
Jag vänder mig mycket starkt mot när man försöker demonisera ett folk.
När jag hörde Chris Davies försöka skuldbelägga ett folk, hör jag toner som jag inte tycker ska höras i detta parlament.
Det är inte en konflikt mellan palestinier och judar, inte en konflikt mellan Israel och den palestinska myndigheten, utan det är en konflikt mellan extremister och moderata krafter i regionen.
Låt oss ge vårt stöd till de moderata krafterna genom att klargöra för var och en som driver hatet och vill eliminera staten Israel att de inte kommer att komma någonvart.
Om Europa ger detta besked stärker vi också de moderata krafterna och lägger en bättre grund för fred.
(PL) Herr talman! Jag vill vända mig till dem som har låtit en laddning i form av bedrägeri och demagogi detonera i parlamentet.
Detta är ett i en rad krig med likheter, men även skillnader.
Den konflikt vi diskuterar i dag är en asymmetrisk konflikt.
Under tre år bombarderades Israel med hemgjorda missiler och inte minsta lilla kritik yttrades i detta parlament mot dem som avfyrade dem. I dag fördömer vi Israel.
Det är lätt att fördöma Israel eftersom landet är medlem i FN.
Det har något att fördöma, det har myndigheter.
Det finns en regering som kan fördömas och kritiseras.
På den andra sidan finns en terroristorganisation vars sanna identitet inte är känd.
En organisation som leker med oskyldiga människors liv genom att agera bakom ryggen på dem.
Ett annat asymmetriskt element är att vi räknar de palestinier som dramatiskt har dödats då de användes som mänskliga sköldar, utan att beakta de israeler som har dödats och de tusentals som lever under hot eftersom blodspillan inte kan kompenseras med ännu mer blodspillan.
Men det allra värsta här i parlamentet är skillnaden mellan ord och handlingar.
Det är lätt för oss att prata, men mycket svårt att vidta effektiva åtgärder.
Utan en internationell närvaro kommer denna konflikt aldrig att lösas.
Slutligen vill jag vända mig till dem som protesterar mot Israels oproportionerliga svarsåtgärd.
Mina damer och herrar! Skulle ni vilja att en terroristorganisation avfyrar 7 000 missiler från Israel till Gaza?
Skulle detta vara proportionerligt?
Eftersom detta är en oproportionerlig konflikt där lagen är ineffektiv måste vi helt enkelt vänja oss. Annars kommer vi bara att gå runt i cirklar och använda ord som inte överensstämmer med verkligheten.
Åsikter som yttras framför tv:n och en varm brasa har inte med sanningen om denna konflikt att göra.
Mina damer och herrar! Jag måste verkligen insistera på att ni håller er till er talartid.
Jag har aldrig avbrutit talare, inte ens när deras talartid har förflutit, men rådets ordförande Karel Schwarzenberg har redan ägnat oss mer tid än vad vi förväntat oss.
Jag har blivit informerad om att han som längst kan stanna till kl. 17.20.
Jag uppmanar er att hålla er till den tid ni har begärt.
I egenskap av general kommer Philippe Morillon att föregå med gott exempel.
- (FR) Herr talman! Det kommer endast att gå att uppnå ett varaktigt lugn i Gaza om en multinationell insatsstyrka sätts in under FN:s kontroll.
För första gången tycks Israel ha funnit sig i denna lösning som palestinierna gång på gång krävt.
Jag vet inte när denna styrka kommer att kunna ingripa. Ett ingripande kommer inte att vara möjligt förrän en överenskommelse har nåtts mellan parterna i konflikten, men vi hoppas alla att detta kan ske så snart som möjligt.
Jag vet emellertid att detta uppdrag kommer att kräva att de som utför det är fullständigt opartiska.
Jag anser därför att Europeiska unionen kommer att ha det bästa utgångsläget för att vidta åtgärder och - varför inte, herr Pöttering? - att göra det inom ramen för Medelhavsunionen.
EU kommer att ha bästa möjliga utgångsläge för att vidta åtgärder eftersom amerikanerna, med rätt eller orätt, anses ha tagit israelernas parti och araberna palestiniernas.
Anser ni inte, herr rådsordförande, att vi bör förbereda oss på detta?
(EN) Herr talman! En långvarig konflikt och ockupation skapar ilska, vrede och besvikelse över myndigheternas ineffektivitet och ger upphov till något vi kallar ”Hamas-effekten”, en viktig faktor.
Arabernas, islamisternas och Hamas förnekande av Israel är oacceptabelt, liksom att använda barn som mänskliga sköldar.
Det ständiga hot som israeliska barn lever under är inte heller acceptabelt.
Frågan är om de nuvarande israeliska ledarna, i denna onda cirkel av våld, kan lära sig av den sex år långa historien i området och applicera den skalpelliknande strategin för två stater.
Jag vet att de fruktar hotet från en aggressiv och oförutsägbar granne som bombar dem med raketer, men i det här avseendet kan det internationella samfundet, inklusive EU, hjälpa till.
Är denna riskfyllda lösning acceptabel, i dag, för Israel?
Men finns det någon annan lösning?
Om den finns, berätta hur den ser ut.
Att förvänta sig att Hamas ska självdö eller försvinna genom att man bombar dem verkar vara en naiv förhoppning och Israel måste därför ha mer mod.
Västvärlden skapade inte två stater 1948, men det bör man göra nu.
Det grundläggande ansvaret försvinner inte.
Låt oss vara modigare i den här strategin.
(SL) Den israeliska staten har beordrat den israeliska armén att krossa Hamas i Gaza.
Den israeliska armén utplånar emellertid Hamas genom att döda palestinier i Gaza.
En tredjedel av alla som dödats är barn och hälften av alla som dödats är kvinnor och barn - men de tillhör inte Hamas.
Det militära våldets omfattning är enorm och oproportionerlig.
Och hur kan eldupphör uppnås när ingen av parterna erkänner den andra partens legitimitet?
Fienden får inte uppfattas som något som ska utsättas för anfall och ödeläggelse, utan som en samarbetspartner som eldupphör kan uppnås med och som ansvarar för att bevara freden i framtiden.
Israel måste erkänna Hamas och inleda en dialog med dem, och vice versa - Hamas måste erkänna Israel.
Det finns inget annat sätt.
Vilken slags fred som helst är bättre än en blodig konflikt.
Det militära våldet måste omedelbart lämna plats för en prioriterad politisk lösning.
Den israeliska premiärministern Ehud Olmert försöker emellertid fortfarande att förbättra sitt dåliga rykte genom att inte tillåta ett eldupphör.
- (CS) Herr talman, fru kommissionsledamot! Låt mig gratulera er till resultatet av era gemensamma förhandlingar, trojkaförhandlingarna i Israel.
Till skillnad från pressen vet vi att det var er delegation som åstadkom att den israeliska sidan övervägde att öppna humanitära korridorer och inleda ett dagligt eldupphör.
Jag tror att detta är första gången som israelerna har accepterat Europa som en betydelsefull samarbetspartner och det tjeckiska ordförandeskapet som en viktig företrädare.
Trots enorma påtryckningar från vänstern enades Europaparlamentet i går om en exceptionell resolution.
Trots de extrema omständigheterna är detta en balanserad resolution, en resolution som kan stödas av högern, en resolution som inte bara är en pamflett eller politisk vinst för vänstern.
Vi har undvikit att infoga ett likhetstecken, oavsett hur abstrakt detta är, mellan en befintlig stat och en terroriströrelse.
Att erkänna staten Israels existens, avstå från våld och inkludera Hamas i avtalen med PLO förblir de viktigaste målen, precis som kravet på att så snart som möjligt uppnå ett permanent eldupphör.
Vi har emellertid inte tillfört något mervärde.
De tre ledande israeliska företrädarna, Barak, Livni och Olmert, är för närvarande oense om under vilka villkor och med vilka garantier de är villiga att genomföra ett eldupphör.
Lösningen är uppenbarligen Egypten och består i en garanti för tunnelkontroller och smugglingskontroller som vore godtagbara för den egyptiska sidan.
Vad gör rådet vid denna tidpunkt?
Hur går det vidare i förhandlingarna med den egyptiska sidan om det tekniska uppdraget, den internationella övervakningen, den tekniska övervakningen och öppnandet av EU BAM Rafah?
Vad kan de parlamentsledamöter som i kväll träffar den egyptiska ambassadören kräva av den egyptiska sidan, eller vice versa, hur kan vi bidra till förhandlingarna med Egypten?
- (CS) Mina damer och herrar! Jag vill uppmana rådet och kommissionen att öka påtryckningarna på båda sidor för att sätta stopp för det pågående våldet.
Vi har säkerhetsrådets resolution 1860 och vi måste följa dess bestämmelser.
Det är nödvändigt att införa garantier för ett långvarigt eldupphör och att låta en humanitär korridor öppnas.
Det har upprepade gånger påpekats att det inte finns någon militär lösning på konflikten mellan Israel och Palestina.
Den enda vägen till varaktig fred går via politiska förhandlingar.
Här är det nödvändigt att Europeiska unionen, i samarbete med USA:s nya regering och Arabförbundet, får en mer framträdande politisk roll än vad som hittills varit fallet.
Den sedan länge pågående konflikten måste stoppas via en politisk överenskommelse som bygger på en tvåstatslösning där israeler och palestinier kan leva tillsammans under fredliga förhållanden med säkra, internationellt erkända gränser och sträva efter att skapa ett fredligt system för regional säkerhet över hela Mellanöstern.
(EN) Herr talman! Vi debatterar ännu en humanitär tragedi i vår närhet - i närheten av mitt eget land - med två av våra partner i Medelhavsregionen.
Tyvärr har palestinierna ännu inte insett att självmordsbomber eller Kassam-raketer aldrig kommer att leda till att ockupationen av deras land upphör.
Israel inser inte att ett så kraftfullt militärt svar ger näring till nya potentiella självmordsbombare och bjuder in nya Kassam-raketer vid första möjliga tillfälle.
Vad händer med de oskyldiga civila, de icke-stridande, kvinnor och barn?
Ingen bryr sig om dem.
Ingen bryr sig om de hundratals barn som dödats, stympats, bränts och skadats - israeliska och palestinska barn.
Vi som sitter bekvämt tillbakalutade framför vår tv mår illa när vi ser det.
Hur ska de som befinner sig på plats må?
Vad kan vi göra?
Att bara försöka skuldbelägga andra hjälper inte de civila.
Att komma med uppmaningar och resolutioner hjälper inte de civila.
Hur kan vi gå från ord till handling?
Det är dags att förhandla med de berörda parterna om att bilda en internationell styrka - vilket andra kolleger föreslagit - som kan gå in i Gaza med en stor polisstyrka som utgörs av arabländer. Där ska den utbilda och hjälpa en polisstyrka från den palestinska myndigheten att i ett brett FN-mandat upprätthålla lag och ordning.
Dessutom behövs en militär europeisk styrka för att säkerställa att raketbeskjutningen och vapensmugglingen upphör och att gränsövergångarna öppnas helt. Vi kan inte längre lägga civilbefolkningens öde i de stridande parternas händer.
(IT) Herr talman, mina damer och herrar! En framstående italiensk antifascist, Piero Gobetti, har sagt att när det bara finns en sanning så är det missvisande att anta en salomonisk ståndpunkt.
Så är fallet med Gaza för närvarande. Jag hoppas att parlamentet kommer att kunna säga de rätta orden för att stoppa Israel.
Om inte kommer det att betraktas som skamligt av historien, palestinierna samt den allmänna opinionen i såväl Europa som arabländerna.
Israel bombar och decimerar ett getto.
Sönerna till dem som tillintetgjorts har blivit de som tillintetgör.
Det finns inga ursäkter för detta, och argumentet att Israel har rätt till sin egen säkerhet är inte godtagbart.
Vem som helst kan om han så önskar se att ingen i dag kan hota Israels säkerhet eller existens.
Detta är uppenbart genom obalansen mellan markstyrkorna, det är uppenbart genom antalet dödade och skadade, det är uppenbart genom det stöd som västländerna fortsätter att överösa Israel med.
Det enda syftet med denna massaker är att förhindra skapandet av en palestinsk stat.
På så sätt förstörs freden och därför måste vi stoppa Israel.
Jag vill tacka rådets ordförande och den tjeckiska utrikesministern för att de fortfarande är hos oss. Vi är inte vana vid en så stark närvaro som det tjeckiska ordförandeskapet i dag visat prov på i denna kammare.
Jag anser att Cristiana Muscardini har rätt. Jag råder dem som inte känner till hur saker och ting förhåller sig i detta område och som måste kunna uttrycka tydliga åsikter att resa dit och se hur saker och ting förhåller sig på plats, genom att antingen resa som turist eller i annat syfte.
Några av oss har varit i Palestina under olika omständigheter, som observatörer vid valet av Abu Mazen eller andra val, och jag anser att man endast kan få en korrekt uppfattning om hur saker och ting förhåller sig genom att personligen vara på plats.
Jag anser att de enda förlorarna under dessa händelser, som härrör från flera decennier tillbaka och inte är något nytt fenomen, är vi i västvärlden eftersom vi aldrig på ett seriöst sätt har tagit itu med problemet och aldrig har försökt lösa det. Vi fortsätter att se det som ett problem mellan två motsatta parter.
Jag har varit i Palestina flera gånger och jag har varit i Israel flera gånger, så jag känner till situationen, om än inte perfekt, så tillräckligt väl, och jag anser att det i realiteten inte är två parter som är inblandade här utan tre.
I detta specifika fall finns det ett problem mellan terroristerna och staten Israel, och det palestinska folket är offren som hamnar i kläm.
Hamas representerar inte det palestinska folket, kanske representerar organisationen en del av dem, men verkligen inte hela det palestinska folket.
Jag kan se en film utspela sig, en film som jag tror att många parlamentsledamöter har sett. Filmen visar alla de israeliska offren, däribland barn och människor i alla åldrar, offer för alla de raketer som har avfyrats och som fortfarande avfyras av Hamas.
Det är ingen slump att det är en stor skillnad mellan Gazaremsan och Västbanken.
Jag riktar denna kommentar till rådets ordförande och till vår utmärkta kommissionsledamot som representerar Europa.
Jag anser att vi måste hantera situationen på rätt sätt.
Jag anser att det viktigaste av allt är att Abu Mazens ställning i dag stärks. Han är den svagaste personen av alla i denna situation, tillsammans med palestinierna, som inte tillmäts något värde i denna fråga.
Jag anser att det är vi alla som är de riktiga förlorarna.
(EL) Herr talman! Den allmänna opinionen i Europa kräver en sak från unionen: att den sätter stopp för slakten på det palestinska folket.
Vi måste fördöma det besinningslösa våldet oavsett varifrån det kommer, men vi måste vara konsekventa och erkänna att Israel svarar med statlig terrorism i en massiv omfattning.
Den asymmetriska vedergällningen, det uppenbara nonchalerandet av alla principer i internationell och humanitär rätt från Israels sida kan inte accepteras.
Det är oacceptabelt att vita fosforbomber och experimentella vapen används mot civila och det är omänskligt att oskyldiga kvinnor och barn blir måltavla.
Om detta skedde i Afrika eller någon annan del av världen skulle vår reaktion vara omedelbar och resolutionen från FN:s säkerhetsråd skulle vara bindande.
När det handlar om Israel inskränker vi oss emellertid till uttalanden och fruktlösa diskussioner.
Jag anser att vi bör använda oss av varje politiskt verktyg, däribland associeringsavtalet, för att övertala Israel att upphöra med det olagliga våldet mot det palestinska folket och att inte längre hindra det humanitära biståndet från att nå fram till de behövande.
Vi kan inte vara passiva åskådare eftersom det gör oss till medbrottslingar i slakten.
Den enda lösningen är ett omedelbart eldupphör, att humanitära korridorer till Gaza öppnas och en dialog med alla parter inleds.
(EN) Herr talman! De fruktansvärda händelserna i Gaza under de senaste två veckorna har lett till ett internationellt fördömande av Israel.
Vi har sett kolleger under dagens debatt stå i kö för att se vem som kan uttrycka starkast vrede över den judiska staten.
För ett land i Mellanöstern är detta dock exakt den händelseutveckling de ville ha: Iran har levererat missiler, krigsmateriel och andra sofistikerade vapen till Hamas i många år.
Landet har försett Hamas stridande med pengar och utbildning.
Målet är att provocera Israel till ett markkrig, och det blodiga resultatet, med fruktansvärda foton av döda barn på tv-skärmar och i tidningar runt om i världen, är bästa möjliga rekryteringsgrund för fundamentalistisk islam och de iranska mullornas vision av en global islamistisk rörelse som står enad mot västvärlden.
Fascistregimen i Teheran är den främsta sponsorn av krig och terror i Mellanöstern och det tragiska resultatet är precis vad Teheran ville ha.
Det avleder uppmärksamheten från den ekonomiska krisen i Iran, som beror på det sjunkande oljepriset, och det avleder den internationella uppmärksamheten från mullornas arbete med att snabbt ta fram ett kärnvapen.
Målet för Irans utrikespolitik är att bli den dominerande regionala makten i Mellanöstern.
Landet vill förena den islamiska världen så att den följer regimens bistra och obehagliga vision av ett totalitärt islamiskt broderskap, där mänskliga rättigheter, kvinnors rättigheter och yttrandefriheten pulvriseras. Skamligt nog har västvärlden inte gjort något för att bemöta eller avslöja den iranska aggressionen.
Västvärlden har ställts inför allt fler bevis på att mullorna sponsrar terror, men har gjort allt för att blidka Teheran och har till och med gått så långt som att gå med på landets krav att avväpna den främsta iranska oppositionsrörelsen, Folkets mujahedin, genom att placera rörelsen på EU:s terrorlista.
Detta måste upphöra.
(EN) Herr talman! Låt oss först och främst vara tydliga med att parlamentet i dag stödjer FN:s säkerhetsråds resolution 1860.
Den måste implementeras utan dröjsmål.
Som en av de parlamentsledamöter som besökt Gaza under blockaden anser jag att ett eldupphör och en reträtt inte räcker.
Självfallet vill vi att raketbeskjutningarna ska upphöra och att terroristerna ska upphöra med sina handlingar, men vi måste få ett eldupphör och ett slut på blockaden så att människorna i Gaza kan börja leva sina liv.
Detta är en fråga om respekt för internationell humanitär rätt.
Human Rights Watch och Islamic Relief har berättat att den dagliga pausen på tre timmar är alldeles för otillräcklig för att kunna gå in och distribuera bistånd.
Det är en fråga om proportionalitet.
Rädda barnen säger att de 139 barn som dödats sedan konflikten började och de 1 271 som skadats inte kan rättfärdigas med att det handlar om självförsvar.
Jag välkomnar uttalandet från EU:s sändebud i Israel, Ramiro Cibrian-Uzal, som i dag sa att EU och Israel nu har fryst förhandlingarna om att uppgradera relationerna av dessa skäl.
Det är inte mer än rätt.
(DE) Herr talman! Först av allt krävs det ett omedelbart och permanent eldupphör på båda sidor - det råder en bred samsyn om detta i parlamentet.
Därefter får vi - EU och det internationella samfundet - emellertid inte låta enbart Hamas och Israel avgöra ödet för människorna på Gazaremsan.
Hamas agerar inte i Gazainvånarnas intresse, eftersom organisationen mycket väl känner till att Israel besvarar ständiga raketattacker - och inte bara under valkampanjer.
Under det senaste året har undersökningar i Gaza visat att det politiska stödet för Hamas har sjunkit till förmån för Fatah.
Det förefaller som om Hamas cyniskt räknar med att det politiska stödet för Hamas kommer att öka igen i och med det stora antalet palestinska offer, på grund av solidaritet med offren.
Israel agerar å andra sidan nästan uteslutande i de egna medborgarnas intresse och därför riktas den internationella kritiken främst mot omfattningen av Israels militära operation och landets acceptans av det stora antalet civila offer.
Därför bör vi européer inte nöja oss med att förhandla fram ett ytterligare eldupphör och finansiera reparationer av infrastrukturen.
Jag kan redan nu se kommissionsledamotens ändringsskrivelse framför mig. Jag är säker på att förslaget redan är slutfört och färdigt att överlämnas till budgetutskottet.
Det räcker inte heller med att bevaka huruvida Egypten stänger tunnelsystemet vid gränsen mot Gazaremsan för vapensmuggling.
Jag uppmanar hela Mellanösternkvartetten att med en stark arabisk närvaro göra ett gemensamt åtagande om att sända trupper med ett starkt fredsbevarandemandat på Gazaremsan och det omgivande området - för att hjälpa människorna i Gaza, Israel och Egypten.
Parallellt med detta måste själva fredsprocessen skyndsamt gå vidare.
Annars befarar jag att vi kommer att få se de slags incidenter som vi har sett i Gaza ännu oftare, och vare sig palestinierna eller israelerna förtjänar detta.
(ES) Herr talman! De spanska ledamöterna i socialdemokratiska gruppen i Europaparlamentet betraktar situationen i Gaza med fasa, smärta och skam, men är även angelägna om att försvara freden, skydda dem som lider mest och upprätthålla värdighet och hopp.
Vår fasa gäller de upprepade scenerna med mördade barn och förtvivlade kvinnor i deras oändliga lidande efter bombningarna av det getto som Gaza har blivit.
Picasso skildrade samma typ av fasa i sin målning Guernica som visar hur vårt Guernica jämnas med marken av junkrarna i Condorlegionen för sju decennier sedan.
Vår smärta gäller det enorma lidandet hos de många offren.
Vår skam gäller oförmågan - hos våra länder, Europeiska unionen och det internationella samfundet - att för det första motverka och för det andra sätta stopp för de brottsliga angrepp som vi fördömer.
Vår skam och ilska gäller de många lögnerna, dubbeltydigheten och det tomma pratet.
Vår skam handlar om att vi vet exakt vad som händer, men ändå inte agerar med den styrka och sammanhållning som krävs.
Historien kommer därför att kräva en förklaring från många av medbrottslingarna, åtminstone när det gäller deras misstag.
Eftersom det alltid är ”bättre sent än aldrig” att agera och det är nödvändigt att hålla dörren till hoppet öppen måste Europeiska unionen stödja den senkomna resolutionen från säkerhetsrådet.
Den måste emellertid se till att denna resolution strikt följs precis som vårt associeringsavtal med Israel också strikt måste följas, vilket innebär att det kan upphävas vid den typ av agerande som nu förekommer.
Är förresten Hamas också ansvarigt för den mörkläggning i medierna som jag ännu inte har hört någon fördöma?
(EN) Herr talman! Jag vill börja med att uttrycka min djupaste sympati för alla oskyldiga människor, både i Israel och i Gaza, som har drabbats under de senaste veckorna och månaderna när konflikten rasat.
Men vi måste se till att vår naturliga mänsklighet, vår högst rimliga oro, inte förvränger vår uppfattning om hur situationen egentligen ser ut.
I Gaza har Hamas skapat ett terrorismens kungadöme: det finns ingen tolerans för opposition mot dess ståndpunkter, man har mördat de palestinier som har opponerat sig, man har splittrat den palestinska myndigheten, man vägrade att upphöra med terrorattackerna mot israeliska civila, man vägrade att erkänna Israels rätt att existera, man vägrade att erkänna de fredsavtal som tidigare framförhandlats.
Jag kommer ihåg vad Hanan Ashrawi sa för tre år sedan, när jag bevakade det palestinska valet.
Hon förutsåg att de mörka krafterna skulle ta över - och hon hade helt rätt!
Vi ska inte vara förvånade över att en Hamas-företrädare är stolt över att säga att döden är en ”industri” för det palestinska folket.
Han syftade på att man använder självmordsbombare och medvetet utnyttjar civila mänskliga sköldar för att skydda potentiella militära mål.
Det är förstås en direkt kränkning av internationell humanitär rätt att använda civila på det här sättet.
Ställd inför en så omedgörlig, förhärdad och hatisk fiende, vad förväntar vi oss att Israel ska göra när landets medborgare hela tiden utsätts för terrorattacker?
Det internationella samfundet uppmärksammade inte detta.
När Israel vidtog fredliga åtgärder, som att införa blockader eller stänga av elektriciteten, fick man kritik.
När nu Israel har vidtagit militära åtgärder som en reaktion på Hamas provokationer drabbas landet av ett kraftfullt internationellt ogillande.
Den sorgliga verkligheten är att det palestinska folket har behandlats illa under många år av dem som har kontroll över den palestinska myndighetens områden, av det internationella samfundet, som har tolererat extremism och korruption, och av arabvärlden som inte har gjort något konkret på flera årtionden för att förbättra deras tillvaro och framtidsutsikter.
Vi behöver en Marshall-plan för Mellanöstern.
Palestinierna behöver inte bara fredsbevarare, utan också en fungerande civil administration, fri från korruption.
Den civila administrationen måste placeras under internationell kontroll, men först måste terroristernas samtliga livlinor - vapen, pengar och politisk släpphänthet - kapas.
(EN) Herr talman! Jag skulle kunna instämma i vad Geoffrey Van Orden säger om Hamas, men faktum är att inget av vad han säger rättfärdigar att Israel bombar civila.
Det är huvudpoängen: vi måste få ett stopp på bombandet, oavsett om det kommer från Hamas eller från Israel.
Jag hoppas att den resolution som följer på den här debatten får starkt stöd i parlamentet i morgon och jag hoppas att det kommer att stärka kommissionen och rådet så att de kan sätta press på både Israel och Hamas att upphöra med dödandet.
Sedan Israel drog sig tillbaka från Gaza har man förvandlat området till det största fängelset i världen och under de senaste tre veckorna har man förvandlat det till ett slakthus. Man använder olagligen terror för att bekämpa terror, dödar civila män, kvinnor och barn och dödar samtidigt möjligheten till en hållbar tvåstatslösning.
Europas relationer med Israel kan inte uppgraderas så länge landet inte kan delta i konstruktiva och väsentliga förhandlingar med sina grannar och alla valda palestinska representanter, inklusive Hamas.
Europa måste göra tydligt att en eskalering av kriget mot Gaza kommer att följas av en eskalering av vår reaktion på kriget.
(HU) Herr talman, kommissionsledamöter, medlemmar av rådet, kära kolleger! Jag uppfattar parternas beteende i Gazakonflikten som cyniskt.
Jag betraktar det som cyniskt och oacceptabelt att Hamas använder civilbefolkningen - till och med barn - som en mänsklig sköld.
Jag uppfattar Israels inställning som cynisk och omänsklig. Landet använder självförsvar som svepskäl för att med oproportionerliga medel skjuta mängder av Gazainvånare, vilket på ett mycket allvarligt sätt drabbar civilbefolkningen, inklusive barn.
Jag betraktar det som cyniskt och lögnaktigt att utländsk diplomati med anmärkningsvärda undantag strävar efter att hålla skenet uppe och till och med efter så många dagar är oförmögen att garantera att civilbefolkningen och biståndsorganen skyddas och dessvärre inte heller kan skydda barnen.
Jag talar för barnens räkning, eftersom det inte finns något ändamål i världen som rättfärdigar att oskyldiga dödas.
Varje barns liv måste vara lika mycket värt, oavsett vilken sida av gränsen barnet befinner sig på.
Detta är det grundläggande axiom som varje part i konflikten måste betrakta som lika viktigt om sann fred någonsin ska kunna uppnås i detta område.
Accepterandet av de värden som handlar om respekt för mänskligt liv, skydd av civila och främjande av humanitärt bistånd kan utgöra grunden till ett varaktigt eldupphör så att fred inom Palestina och mellan Palestina och Israel kan uppnås.
(EN) Herr talman! Hamas bedrev terror mot Israels invånare och har provocerat fram en vedergällning.
På avstånd kan det verka som att en del av dem uppskattar att de får nya civila martyrer - också barn - liksom den publicitet det ger deras sak, oavsett hur obehagligt det är för rättänkande personer att ta in detta.
Jag har aldrig stött terrorism och jag är inte heller någon Israelkritiker. Det är ett land som har rätt till en fredlig samexistens i regionen, men vi skulle vara tokiga om vi inte kände oss känslomässigt berörda och moraliskt skamsna över det som händer i Gaza i dag.
Israels svar är helt oproportionerligt och särskilt dödandet av små barn är en skamfläck.
Jag har hittills inte motsatt mig det nya avtalet mellan EU och Israel.
Jag tror på det råd Dalai Lama gav här i parlamentet förra månaden: det bästa sättet att påverka Kina i Tibet-frågan är att ha goda relationer med dem.
Jag tror att det också gäller relationerna mellan EU och Israel, men hur kan vi få dem att förstå vilken avsmak vi känner inför omfattningen av det som händer?
Jag kan tillägga att i går distribuerades en not om de humanitära behoven i regionen till de av oss som deltog i det gemensamma mötet för utskottet för utrikesfrågor och utskottet för utveckling.
Jag uppmanar kommissionen och rådet att se till att ett fullständigt humanitärt biståndspaket finns redo så att vi kan gå in där och hjälpa de nödlidande vid första möjliga tillfälle.
rådets ordförande. - (EN) Herr talman! Något som nämndes i början var om vi ska kontakta Hamas eller inte.
Jag tror inte att det är dags att göra det ännu.
Under de senaste månaderna har Hamas definitivt fortfarande agerat som en terroristorganisation.
Så länge man agerar så kan organisationen inte kontaktas officiellt av företrädare för EU.
Jag medger att jag är en gammal man och att jag har sett många terroristorganisationer växa fram från början, bli mer eller mindre accepterade och accepteras av det internationella samfundet.
Jag har sett det i Afrika.
Jag har sett det i Irland.
Jag har sett det på många platser.
Det händer.
Men först måste de sluta agera som en terroristorganisation.
Då kommer jag att vara redo att tala med Hamas eller med någon annan, men inte innan de har slutat agera som en terroristorganisation.
Jag tror att det är viktigt att säga detta, eftersom EU inte kan ge upp sina principer.
Det finns olika metoder för att höra vilka idéer de har, det finns indirekta kontakter med politiker i regionen som står i kontakt med dem, vilket är viktigt och bra, men än är det inte dags för EU att ha direktkontakter med Hamas.
Jag menar att vi ska vara orubbliga i detta.
I andra avseenden måste vi hylla Egypten för den viktiga roll landet spelat under de senaste veckorna och dagarna med sina insatser och sitt hårda arbete för att få till stånd ett eldupphör och kanske också en vapenvila som, i processens slut, leder till fred i regionen.
Jag vet hur svår den här frågan är.
Vi står i ständig kontakt med egyptierna.
Vi vet vilket viktigt arbete de gör och jag vill gratulera dem.
Det kom en fråga om hur vi kan bistå i regionen.
För det första, de som befinner sig på plats kan berätta exakt vad de behöver.
Vi ska inte bestämma vad vi ska ge dem.
De måste fråga oss och EU.
Många medlemsstater inom EU har sagt sig vara villiga att hjälpa till på alla möjliga sätt - tekniskt, skicka rådgivare, förbereda det som kan behövas - men detta måste först och främst ske med samtycke från alla berörda stater här.
Det är den första uppgiften som ska genomföras.
Jag hörde ett viktigt förslag som handlade om att ta fram en Marshall-plan för Mellanöstern.
Jag tycker att det är en mycket bra idé och att vi ska följa upp den.
Den här regionen behöver verkligen att man bygger upp nya idéer, på det sätt som hjälpte Europa i så hög grad efter kriget.
Benita Ferrero-Waldner och andra talade om vad man åstadkom under resan.
Jag anser att vi åstadkom mycket och jag vill än en gång berömma Benita Ferrero-Waldner, som gjorde huvudarbetet i vår delegation inom den humanitära sfären, där det vi åstadkom fortfarande fungerar i dag.
Men låt oss vara tydliga med att också dessa mycket svåra förhandlingar i Mellanöstern bygger på den form som redan fanns vid vår delegations besök i Mellanöstern.
Detta handlar i grunden om hur freden ska organiseras och vad som är nödvändigt.
Vår plan bygger på vad vi fick veta då och diskuterade med våra partner.
Det fördes också en diskussion om att uppgradera våra relationer med Israel.
Som ni känner till fattades ett beslut av EU:s ministerråd i juni 2008.
Det kan ändras enbart om ministrarna inom EU bestämmer sig för att ändra beslutet.
Det kan inte ändras, inte ens genom vad en mycket respekterad företrädare för EU säger i Jerusalem.
Jag medger att i den rådande situationen skulle det vara för tidigt att diskutera hur vi ska uppgradera vår relation med Israel och om ett toppmöte ska genomföras under överskådlig tid.
För närvarande har vi betydligt mer brådskande och viktigare frågor att lösa.
Jag vill än en gång betona att beslutet fattats av ministerrådet och att det är det som gäller.
Vad kan göras för att stoppa Israel?
Om vi ska vara ärliga - mycket lite.
Israel agerar som det gör och som en livslång vän av Israel, vilket jag säger helt ärligt i dag, är jag inte så nöjd med det man gör för närvarande.
Jag tror att landets politik också skadar Israel.
Det är en sak, men EU har mycket få möjligheter, annat än att tala mycket tydligt och mycket uppriktigt och be våra partner att sätta stopp.
Våra partner i Mellanöstern måste hitta lösningen: Israel, Egypten och övriga berörda parter.
EU kan hjälpa till här.
EU kan hjälpa till genom att erbjuda all typ av hjälp om man kommer överens om eldupphör för att uppnå de angivna målen: stänga smuggelvägarna, stänga tunnlarna, bevaka havet etc. EU kan hjälpa till i Gaza på flera sätt, t.ex. med återuppbyggnad eller hjälp med humanitärt bistånd.
EU kan göra allt detta, men om man ska vara helt ärlig har vi inte makten och medlen för att säga ”stopp”.
Anser parlamentet att vi kan skicka en jättelik beväpnad styrka till Mellanöstern för att stoppa de stridande parterna?
Nej.
Vi har inte de möjligheterna och både Israel och Hamas är beroende av andra krafter än EU.
Israel har mäktiga allierade också utanför Europa.
Vår möjlighet att uppnå något är begränsad.
Vi kan hjälpa till, vi kan bistå, vi kan erbjuda våra bästa tjänster och vi kan vara djupt engagerade.
I det avseendet har vi åstadkommit en hel del.
Men överdriv inte våra möjligheter.
(EN) Herr talman! Israel säger att man utövar sin rätt till självförsvar.
I så fall måste grundsatserna för ett rättfärdigt krig, inklusive proportionalitet, följas.
Att Israel struntar i detta är uppenbart och att vi struntar i att så är fallet är fel.
Man kan inte använda fosfor mot civila och hävda att detta är ett civiliserat agerande.
Det är uppenbart att EU inte kan lösa detta på egen hand.
Men det finns en vit elefant i rummet.
Vi behöver amerikansk beslutsamhet.
USA:s gensvar har varit en besvikelse eftersom det är obalanserat och orättvist.
Tidpunkten för när de här handlingarna genomförs är strategiskt beräknad från Israels sida, men, herr Obama, det är snart den 20 januari.
Världen väntar och EU är redo att agera partner!
Vill ni återställa de värden som vi delar med er eller kommer ni att tillåta att denna orättvisa får fortgå - än en gång?
Kommer ni att arbeta med oss för att ge alla berörda skydd?
Palestinierna frågar er - hur kan det vara rätt att ert land ber om humanitärt bistånd på plats, men håller tyst när det bara handlar om bomber från luften?
Till de kolleger som vill bryta ner Hamas enbart med militära medel: besök Gaza och Västbanken.
Väck er medmänsklighet till liv så förstår ni varför Hamas bara blir starkare.
Det här är inte rätt sätt att hjälpa Israel eller palestinierna.
Ett omedelbart eldupphör är bara en nödvändig början.
(EN) Herr talman! Det är mycket tydligt att parterna i den här konflikten inte lyckas respektera internationell humanitär rätt och att civilbefolkningen i Gaza därmed betalar ett mycket högt pris.
Ansvar måste utkrävas enligt internationell rätt när krigföringsprinciper som proportionalitet och icke-diskriminering inte respekteras.
En av grundsatserna för ett rättfärdigt krig handlar om att agerandet ska styras av principen om proportionalitet.
Styrkan måste användas i proportion till den kränkning man utsatts för.
Tyvärr har vi sett stor vårdslöshet från israelernas sida.
Även om Hamas började med raketattackerna mot Israel har den israeliska reaktionen, enligt min uppfattning, varit oproportionerlig.
Siffrorna talar för sig själva: drygt 900 palestinier har dödats, men bara ett mindre antal israeler.
Israel måste inse att de har ett ansvar att dimensionera den kraft de använder i enlighet med internationell rätt.
Å andra sidan kan man inte blunda för att Hamas fortfarande är listat som en terroristorganisation av EU och fortsätter att vägra ge upp sin väpnade kamp.
Och inte bara det - Hamas har hela tiden vägrat att erkänna Israels rätt att existera.
Hamas och andra beväpnade palestinska grupper måste inse att människorna i södra Israel har rätt att leva utan att bombarderas.
(EN) Herr talman! För alla som följer konflikten mellan israeler och palestinier kan detta vara en tidpunkt då vi frestas att lyfta händerna i luften och skrika ut vår förtvivlan.
Det tycker jag dock inte att vi ska göra eftersom jag anser att det största provet på vår medmänsklighet i dag är att verkligen förstå de frågor som vi står inför.
Den första frågan handlar om att det inte finns någon hållbar lösning på den här konflikten om inte bombningen av Israel upphör.
Den andra frågan handlar om att det inte finns någon hållbar lösning på den här konflikten om inte Gaza öppnas för humanitärt bistånd.
President Peres har helt rätt när han säger att Gaza ska vara öppet för bistånd och inte avstängt för raketer.
Jag tycker att detta är centralt och alla håller med om detta.
Det går inte att återgå till situationen som den var innan och jag tror att det finns flera saker vi kan göra här. För det första kan parlamentet få båda sidor att mötas för samtal.
För det andra kan vi ställa oss bakom kommissionen och rådet och stödja deras insatser. Och till sist ska vi stödja det egyptiska förhandlingsspåret, eftersom det är det enda spår som kan leda till en lösning och till det eldupphör vi nu alla hoppas på.
(EN) Herr talman! Det är inte bara parlamentsledamöterna som upprörs av utvecklingen i Gaza.
Allmänheten i Europa har också alltför länge upprörts av hur folket i Gazas lider och av den israeliska blockaden.
Till detta kommer de ständiga attackerna och de fruktansvärda israeliska militära angreppen på oskyldiga civila, framför allt kvinnor och barn.
Världssamfundets uppmaningar om ett omedelbart eldupphör hörsammas inte.
Palestinierna behöver omedelbart tillgång till mat, medicinsk hjälp och säkerhet.
Israel måste åtminstone respektera principerna i den internationella rätten.
Om man inte gör det måste Israel förlora det stöd landet fortfarande har från det internationella samfundet.
Det är olyckligt att FN:s resolution har åsidosatts.
Det är beklagligt att EU fortfarande måste hitta sin roll.
Kanske kan man göra det om EU vidtar starkare åtgärder än man hittills har gjort.
Det räcker inte att bara lägga uppgraderingen av relationen på is.
Vi kan påverka.
Vi är en viktig handelspartner.
Vi är en viktig bidragsgivare i regionen.
Vi kan alltså utöva denna roll.
(EN) Herr talman! Är det etiskt acceptabelt och ursäktligt enligt internationell rätt att staten Israel i sina ansträngningar att neutralisera Hamasterrorister kan inleda en större militär terrorkampanj, med allvarliga brott mot FN:s konventioner och de mänskliga rättigheterna mot 1,5 miljoner oskyldiga civila som saknar möjlighet till flykt?
Är sådana handlingar förenliga med EU:s värderingar om rättvisa och demokrati?
Är den israeliska lobbyn så stark att den kan få USA och EU att praktiskt taget stå overksamma och se obeskrivliga grymheter begås i kampen mot terrorismen?
Om svaret på dessa frågor är ja, då bör vi alla prisa den israeliska regeringens agerande i Gaza som modigt. Om svaret är nej bör vi å det starkaste klart och tydligt fördöma Israel, samt snabbt och effektivt vidta åtgärder, till exempel handelssanktioner, för att stoppa blodbadet i Gaza i dag och för all framtid.
Jag håller verkligen inte med ministern som gick i väg, som ansåg att det inte finns mycket vi kan göra.
Vi kan göra åtskilligt, och det är vår skyldighet.
(EN) Herr talman!
Jag valdes till parlamentsledamot för 25 år sedan, men denna är nog den viktigaste debatt som jag deltagit i.
Fru kommissionsledamot! Jag hoppas att ni lyssnade noga till utskottet för utrikesfrågor i går kväll och att ni har lyssnat till parlamentet i dag.
Jag hoppas att ni, till skillnad från rådets ordförande Karel Schwarzenberg, svarar att EU har ett moraliskt inflytande som vi kan utöva på angriparen i det här fallet.
Israels folk är ett rättvist och hedersamt folk som har lidit oerhört under århundraden på vår kontinent.
De kommer att förstå er rekommendation till ministerrådet att EU bör avstå från all kontakt med de israeliska myndigheterna tills de har upphört med bombningarna.
(ES) Herr talman! Vi måste med absolut övertygelse uppmana Israel att upphöra med dödandet och låta de skadade få vård och offren mat.
Vi måste klargöra att Israels inställning till internationell rätt kommer att få konsekvenser för landets förbindelser med Europa.
Jag vill gratulera det fåtal unga europeiska frivilligarbetare som lider tillsammans med folket i Gaza, framför allt Alberto Arce.
De representerar det bästa när det gäller de värden i form av solidaritet och frihet som vårt Europa står för, ett Europa som måste agera därefter i denna fruktansvärda konflikt.
(DA) Herr talman! Jag vill bara säga två saker.
För det första vill jag påminna alla om att det i vårt beslut tydligt anges och upprepas att vi har lagt vårt stöd för uppgradering på is, och jag hoppas verkligen att vi inte kommer att fortsätta som om ingenting har hänt bara för att ordförandeskapet säger att vi ska göra det.
Det andra jag vill påpeka är att Israel inte vid någon tidpunkt har hållit vad man lovade i samband med förhandlingarna.
Det blev inget eldupphör eftersom Israel inte hävde blockaden under denna period, och jag känner att jag även måste nämna Annapolis där Israel lovade att frysa bosättningsverksamheten.
Vad hände i själva verket?
Landet ökade helt enkelt bosättningstakten.
Bosättningstakten har aldrig varit så hög som den varit sedan Annapolis, och jag anser att så länge inga framsteg nås på plats kommer vi aldrig att få Hamas att agera i enlighet med de regler som vi vill att de ska följa. Av denna anledning måste vi se till att Israel uppfyller sin del av avtalet.
(EN) Herr talman! I går genomförde vi ett gemensamt möte med delegationerna för förbindelserna med Israel och med det palestinska lagstiftande rådet, och jag är övertygad om att ni kan föreställa er de häftiga diskussionerna, känslorna och anklagelserna - och föreslagna lösningar - efter 18 dagars krig i Gaza och omkring 1 000 döda.
Faktum är att Israel, efter att ha väntat i åtta år och absorberat ca 8 000 missiler som terroriserat en miljon medborgare längs Gazas gränser, slutligen förlorade tålamodet.
De började värna sina medborgares säkerhet, vilket är deras fulla rätt och ansvar.
Hamas är en terroristorganisation, en otvetydig brottsling och en börda för palestinierna i Gaza.
Lösningen är därför en stärkt kvartett och, framför allt, ett samordnat arbete mellan USA:s nya administration och ett starkare och mer integrerat EU.
Jag välkomnar det tjeckiska ordförandeskapet, dess prioriteringar och dess omedelbara, aktiva engagemang i regionen.
(RO) Denna konflikt, som pågått mycket länge, bygger på problem som handlar om territorium och kulturella skillnader som ibland behandlas på ett överdrivet sätt.
Den långsiktiga lösningen är en skyddad, säker israelisk stat sida vid sida med en godtagbar palestinsk stat.
Denna lösning kan emellertid inte uppnås genom terroristattacker eller väpnade åtgärder.
För att kunna få ett normalt liv måste det palestinska folket bilda en stat som baseras på demokratiska institutioner och rättssäkerhet och som utgör en garanti för ekonomisk utveckling.
De måste avstå från terroristhandlingar och skapa ett normalt politiskt klimat genom att främja valet av politiker som verkligen vill lösa denna konflikt genom förhandlingar.
(GA) Herr talman! Jag vill uttrycka mitt stöd för dem som fördömer attackerna och visa min solidaritet med folket i Gaza.
Minister Schwarzenburg säger att Europeiska unionen inte kan göra så mycket.
Europeiska unionen bör upphöra med uppgraderingen av förbindelserna med Israel, och de avtal som för närvarande tillämpas bör upphävas tills Israel uppfyller sina plikter enligt internationell rätt.
Även innan de omoraliska attackerna, som nyligen genomfördes, upplevde vi år av kollektiv bestraffning av det palestinska folket.
Omfattningen och typen av attacker, som genomfördes i Gaza av en modern armé mot ett belägrat folk, som redan är svagt till följd av isolering och belägring, är helt fruktansvärda.
Det var fel att lägga skulden på dessa människor - vi måste vara tydliga med att säga att de största offren här är människorna, de oskyldiga människorna i Gaza.
(PL) Det är med stor smärta som vi iakttar vad som sker på Gazaremsan.
Vi stöder inte Hamas metoder som handlar om att slåss och provocera, men Israel har valt ett oproportionerligt sätt att lösa sin tvist med det palestinska folket.
Det har förekommit en definitiv kränkning av principerna inom internationell rätt.
Ingen av parterna i konflikten är intresserad av att den motsatta parten ska uppleva fred.
Båda parterna ser endast till sina egna intressen - det är ett exempel på nationell själviskhet.
Den internationella opinionen är emot ett fortsatt krig.
Europeiska unionen och FN, som stöds av många länder, bör ingripa med fasthet.
Det är dags att sätta stopp för detta beklagliga krig.
De israeliska trupperna bör återvända till sina baracker.
Hamas måste upphöra med att avfyra raketer mot Israel.
Vi måste garantera att humanitärt bistånd brådskande ges till civilbefolkningen och att offren, som sägs uppgå till omkring 3 000 människor, erbjuds vård.
Vi måste bygga upp landet och hjälpa det att återgå till ett normalt liv.
Detta är det scenario jag efterlyser hos Europeiska unionens aktuella ledarskap och Europeiska kommissionen.
(EN) Herr talman! Jag undrar bara om vi fortfarande kommer att debattera gasen i dag eller om det strukits från föredragningslistan?
Vi väntar på den debatten.
På föredragningslistan står inte bara en debatt om Mellanöstern, utan även en om gas.
Har den strukits från föredragningslistan?
Det är nästa punkt på föredragningslistan.
(SL) Jag var besviken på det senaste tillkännagivandet från Tjeckiens utrikesminister, som för närvarande leder rådet.
Vi kan naturligtvis sätta allt vårt hopp till vår kommissionsledamot.
Men dödssiffran stiger.
Om vi fortsätter att tala på detta sätt kommer förmodligen 1 500 människor att vara döda om en vecka.
Det är svårt att tala med Hamas.
Organisationen finns på listan över terroristorganisationer och det är svårt att vidta åtgärder mot den.
Israel, å andra sidan, är vår vän, vår samarbetspartner och en viktig medlem av det internationella samfundet.
Israel måste hålla sig till internationella beslut, Förenta nationernas resolutioner och även till rekommendationerna från dess vänner och samarbetspartner.
Om landet inte lyckas med detta måste dess vänner och samarbetspartner kunna fördöma dess handlingar och hota med att vidta sanktioner.
ledamot av kommissionen. - (EN) Herr talman!
Jag kommer att fatta mig kort, eftersom debatten har varit lång.
Låt mig först säga att efter att ha varit medlem av Mellanösternkvartetten i fyra år nu spelar EU en roll. Naturligtvis är vår roll inte den viktigaste.
Det är ibland frustrerande för oss alla, speciellt i den här svåra situationen när man helst vill uppnå en hållbar och varaktig vapenvila som den vi har föreslagit, men detta inte går så snabbt.
Jag skulle vilja ge er den provisoriska information som jag nu har, vilken rapporterats i nyheterna. Källor i Egypten som följer förhandlingarna säger att Hamas reagerar positivt på de senaste förslagen från Egypten.
I varje fall rör saker och ting på sig.
Jag är ännu inte säker på om detta verkligen bekräftats, men Hamas kommer att hålla en presskonferens klockan 20.00 i kväll.
Förhoppningsvis gör vi framsteg.
Det är åtminstone det alla hoppas på.
För det andra har vi, trots all frustration, inget annat alternativ än att fortsätta arbeta för fred, vilket är vad vi kommer att göra.
Det är något jag förbinder mig att göra så länge jag är medlem av Mellanösternkvartetten.
Vi kan bara åstadkomma det tillsammans, och vi måste stödja och förbättra palestinska ansträngningar till försoning eftersom det är enda sättet att stoppa hemskheterna i Gaza.
För det tredje kommer vi, så fort en vapenvila kommer till stånd, att göra allt vi kan för att återställa de grundläggande tjänster till befolkningen som drabbats så svårt.
Framför allt anser jag att det viktigaste nu är att få ett slut på förstörelsen och börja återuppbyggnaden och att försöka åstadkomma fred.
Vi har redan diskuterat detta ämne länge, så jag vill inte dra ut på det mer, men detta är min inställning, och jag hoppas att vi får ett bra tillfälle.
Jag har jag mottagit ett resolutionsförslag, som ingivits i enlighet med artikel 103.2 i arbetsordningen.
Debatten är härmed avslutad.
Skriftliga förklaringar (artikel 142)
Med tanke på den grymhet som det palestinska folket på Gazaremsan har utsatts för, och som skarpt kritiseras och fördöms i den nya resolutionen från FN:s råd för mänskliga rättigheter, krävs följande:
En skarp kritik av kränkningarna av de mänskliga rättigheterna och av de brott som den israeliska armén begår, Israels statliga terrorism!
Ett tydligt fördömande av Israels grymma anfall mot det palestinska folket som ingenting kan rättfärdiga!
Ett slut på anfallet och den omänskliga blockad som befolkningen på Gazaremsan har drabbats av!
Brådskande humanitärt bistånd till den palestinska befolkningen!
De israeliska truppernas tillbakadragande från allt ockuperat palestinskt territorium!
Respekt för internationell rätt och FN:s resolutioner från Israels sida, ett slut på ockupationen, bosättningarna, separationsmuren, avrättningarna, arresteringarna, exploateringen och det oräkneliga antalet förödmjukelser som det palestinska folket utsätts för!
En rättvis fred, som endast är möjlig genom att det palestinska folkets omistliga rätt till en självständig och suverän stat, med gränserna från 1967 och dess huvudstad i östra Jerusalem, respekteras!
I Palestina finns det en kolonisatör och en koloniserad part, en angripare och ett offer, en förtryckare och en förtryckt part, en exploatör och en exploaterad part.
Vi kan inte låta Israel fortsätta på samma sätt ostraffat!
skriftlig. - (EN) Reaktionen på konflikten i Gaza måste bli mer nyanserad än den är i nuläget.
Vi kan inte ursäkta överdrivet våld, men vi måste se mer till konfliktens ursprung.
Att förhandla med Hamas är inte tänkbart.
En terroristgrupp som kallblodigt använder sitt eget folk som skydd mot attacker är inte intresserad av att förhandla fram en verklig fred.
Dessutom måste vi också komma ihåg att Hamas har tagit på sig en viktig roll i den kedja av terroriströrelser som leder till Hizbollah och terroristregimen i Teheran.
Därför måste Hamas ses som en del i bredare ansträngningar för att störa den ömtåliga stabiliteten i Mellanöstern och ersätta den med fundamentalistiska extremistregimer, som i princip inte erkänner Israels existensberättigande.
Vi måste också inse att frågan om Israels säkerhet är kopplad till EU:s säkerhet.
EU måste utöva sitt inflytande för att först och främst åtgärda konfliktens grundorsaker.
För att undvika att fler araber och israeler dödas måste de arabiska parterna ovillkorligen erkänna Israels existensberättigande och bidra till att stoppa infiltrationen från extremiströrelser och införandet av ännu fler dödliga vapen till regionen.
skriftlig. - (FI) Herr talman! Det är ett obestridligt faktum att civilbefolkningen i Gaza och södra Israel har fråntagits rätten till en människovärdig tillvaro.
En nyhetsbyrå återgav historien om två barn som skulle gå över en gata i Gaza.
Barnen tittade varken åt höger eller vänster för att se om något skulle komma - de titta upp eftersom de var rädda för vad som skulle kunna komma från himlen.
Det finns två uppenbart skyldiga parter när det gäller den massiva humanitära krisen i Gaza.
Hamas oansvariga agerande på de palestinska territorierna, deras fega sätt att gömma sig bland civilbefolkningen, och provokationen med raketattackerna visar sammantaget hur instabil den palestinska regeringen är.
Israels oproportionerliga attacker på den redan svaga och desperata palestinska enklaven är ett annat bevis på att landet ställer sig likgiltigt inför internationella humanitära skyldigheter.
Vi måste uppmana parterna att få ett slut på denna vansinniga situation genom ett omedelbart och permanent eldupphör.
Som en första åtgärd bör Israel tillåta humanitär hjälp att komma in i Gaza, där förbättrade levnadsförhållande också skulle bidra till en långsiktig fred.
Mellanösternkvartetten måste vidta åtgärder i rätt riktning, med den nya amerikanska administrationen som vägvisare.
Egypten har ett särskilt ansvar på grund av gränsfrågorna, och landets roll som medlare tillsammans med unionen har ingett oss hopp.
Historien visar att arbete för fred lönar sig i längden.
Vi kan inte ge upp, anpassa oss eller vänja oss vid tanken på en olöst konflikt, eftersom det inte finns någon sådan.
Enligt vinnaren av Nobels fredspris, Martti Ahtisaari, är fred en fråga om vilja.
Det internationella samfundet kan försöka att uppmuntra och främja denna vilja, men bara de berörda parterna kan mobilisera den och skapa en bestående fred.
Fru kommissionsledamot! Skulle ni kunna framföra följande meddelande från EU: ”Folk av det heliga landet, visa att ni vill ha fred.”
skriftlig. - (EN) Det är oroande när en värld förefaller ur stånd att rädda oskyldiga barn från att sprängas i bitar i krig.
Trots allt som sagts har det inte kommit något uppehåll i bombräderna mot Gaza, vilka hittills har lett till att 139 barn omkommit och 1 271 skadats.
Tyvärr kommer dessa upprörande tal att fortsätta stiga.
Hamas raketattacker mot Israel har provocerat det gensvar man avsåg: motattacker och förlusten av civila liv samt ytterligare framflyttning av positionerna.
Jag beklagar djupt att oskyldiga civila används som mänskliga sköldar.
Det måste upphöra.
Jag tänker inte döma i skuldfrågan - båda sidor begår fel, men jag vill betona behovet av att åstadkomma en omedelbar och effektiv vapenvila.
Det är absolut nödvändigt att få till stånd obehindrat tillträde för humanitär hjälp och bistånd till Gaza, utan fördröjning.
Om bara mänskligheten kunde inse hur meningslösa den här typen av krig är!
Varje bild av döda i Gaza upprör människor i hela arabvärlden och jag oroar mig för att den väsentliga grundsatsen i fredsprocessen för Mellanöstern sakta försvinner utom räckhåll: den såkallade tvåstatslösningen, ett självständigt Palestina som existerar sida vid sida i fred med Israel.
Det åligger det internationella samfundet att fördubbla sina ansträngningar för att hitta en lösning.
skriftlig. - (FI) Vi är alla vittnen till de israeliska soldaternas masslakt av civila i Gaza.
Vi, eller närmare bestämt många parlamentsledamöter till höger, blundar för det som sker.
Det skulle inte kunna ske om inte den politiska högereliten i USA och EU blundade för det som sker.
De som blundar är också de som beväpnar dem som dödar civila.
Det är dags att vi tar upp frågan om att bryta de diplomatiska förbindelserna med förövarna av folkmord och etnisk rensning.
skriftlig. - (HU) Situationen i Mellanöstern fyller mig med oro.
Vad kommer det att krävas för att uppnå fred?
Hur många civila döda och sårade kommer det att krävas innan ett verkligt eldupphör kan genomföras? I Bosnien-Hercegovina krävdes det minst 10 000 för att fredsförhandlingar skulle inledas, för att fredsbevarande styrkor skulle komma till platsen och nedrustning påbörjas.
För några dagar sedan hedrade vi minnet av ödeläggelsen av Nagyenyed (Aiud).
För 160 år sedan slaktades flera tusen oskyldiga civila, däribland kvinnor och barn, i denna transsylvanska stad och dess omgivningar.
Sedan dess har det inte varit möjligt att hedra minnet av dessa offer tillsammans med majoriteten av befolkningen.
Det kan komma en tid då israelerna och palestinierna inte bara hedrar minnet av varandras offer tillsammans, utan till och med går samman för att skapa en varaktig fred och framtid.
Fram till dess är det Europeiska unionens uppgift att föregå med gott exempel.
Det återstår mycket att göra för oss också när det gäller att skapa fred inom Europa.
Vi behöver samarbete mellan majoriteter och minoriteter som är likställda med varandra.
Det minsta vi kan göra är att enas och tillsammans hedra minnet av offren.
Det återstår mycket att göra inom EU på området respekt för individers och minoriteters rättigheter.
skriftlig. - (PL) Under plenarsammanträdet i januari antog Europaparlamentet en resolution om konflikten på Gazaremsan.
Båda sidor i konflikten uppmanades att genomföra ett omedelbart och varaktigt eldupphör och att upphöra med den militära verksamheten (Israels militära åtgärder och Hamas raketer), som under en tid hindrat bistånd och humanitär hjälp från att nå fram till medborgarna i det område där konflikten utspelats.
Den har redan kostat tusentals offer i form av civila, däribland kvinnor och barn, som har lidit i nästan tre veckor.
Det råder brist på grundläggande förnödenheter som dricksvatten och livsmedel.
FN:s anläggningar har anfallits.
I resolutionen krävs det att internationell rätt ska följas så att den befintliga konflikten kan lösas.
Israel är vår vän och har rätt att försvara sig självt som stat, men det måste tydligt fastslås och understrykas att de medel som används i detta fall är mycket oproportionerliga.
Israel måste tala och förhandla med Hamas eftersom de tidigare metoderna inte har fungerat.
Europeiska unionen står också inför en svår uppgift. Den måste hitta mekanismer som leder till dialog och förståelse mellan parterna så att konflikten så snart som möjligt kan upphöra permanent.
Bortfallna skriftliga förklaringar: se protokollet
Återupptagande av sessionen
Jag förklarar Europaparlamentets session återupptagen efter avbrottet torsdagen den 5 februari 2009.
Tillämpad forskning inom den gemensamma fiskeripolitiken (kortfattad redogörelse)
Nästa punkt är en kort presentation av ett betänkande av Rosa Miguélez Ramos för fiskeriutskottet, om tillämpad forskning inom den gemensamma fiskeripolitiken.
Herr talman, herr kommissionsledamot, mina damer och herrar! Att förena ett korrekt bevarande av ekosystemen med ett hållbart utnyttjande av marina resurser, förebyggande och kontroll av effekterna av mänsklig aktivitet på miljön, förbättring av kunskaper och teknisk utveckling och förnyelse är uppgifter som vi inte kan lösa om vi inte får stöd av den europeiska forskningsgemenskapen.
Forskning om fiske är också avgörande när vi ska utarbeta rekommendationer och ge lagstiftarna vetenskapliga råd.
Ökade investeringar i forskning och utveckling, och när det gäller insamling och behandling av pålitliga data skulle resultera i en stabilare och hållbarare gemensam fiskeripolitik.
Men även om det jag fick höra av en forskare - ”Det är inte pengarna, utan de mänskliga resurserna som är problemet” - ger en bra bild av situationen, så tänker jag inte säga att forskning om fiskerifrågor har gott om finansiella resurser.
Tvärtom vill jag säga att vi har ett dubbelt problem.
För det första, herr kommissionsledamot, så verkar de belopp som avsatts i sjunde ramprogrammet för marin forskning, som borde vara en sektorövergripande fråga, vara otillräckliga för den integrerade strategi som för närvarande krävs i frågan.
Dessutom, herr kommissionsledamot, har forskarna problem när de skickar in projekt till sjunde ramprogrammet - och jag kan försäkra er att jag talade med många av dem när jag utarbetade mitt betänkande, både före och under processen.
Dessa problem kan delvis tillskrivas det annorlunda fokus som å ena sidan krävs för vattenbruk, som till sin natur i grunden är en industriell verksamhet, och å den andra sidan forskning om fiske och marin vetenskap, som till sin natur är mångdisciplinär och mer långsiktig.
Fram till det sjunde ramprogrammet täcktes båda dessa områden med samma medel, och de rapporterade till generaldirektoratet för fiskerifrågor, vilket gjorde att de kunde komplettera varandra.
För närvarande är det GD Forskning som har ansvaret, och resultatet är att det blir svårare för forskarsamhället att kommunicera sektorns problem och behov till de personer som utarbetar riktlinjerna för förslagsinfordringar.
Den allmänna uppfattningen inom forskarsamfundet är dessutom att generaldirektoratet verkar ha valt att prioritera grundforskning utan att lämna utrymme för forskning som är inriktad på allmänna policyfrågor.
Låt mig lämna ett exempel: att från vetenskaplig synpunkt berika gemenskapens maritima strategi, eller undersöka kopplingarna mellan fiske och klimatförändringar.
Sammanfattningsvis kräver målet för Europeiska unionens marina politik, nämligen att uppnå ett produktivt fiske i en ren marin miljö, att forskarna på detta område har tillgång till horisontella finansieringsmekanismer i sjunde ramprogrammet.
Avslutningsvis vill jag nämna det andra problemet: den oroande bristen på unga forskare inom fiskeriforskningen, vilket verkar vara resultatet av yrkesutbildningar som inte är särskilt attraktiva jämfört med andra basvetenskaper.
Det är viktigt att vi skapar intressanta och givande universitetskurser som erbjuder goda yrkesmöjligheter.
Det verkar också som om vi måste standardisera de olika forskningsmodeller som tillämpas i de olika medlemsstaterna för att vi bättre ska kunna jämföra resultat, ställa samman data och öka samarbetet mellan olika nationella forskningsinstitutioner.
Jag tycker naturligtvis också att det är mycket viktigt att fiskarnas erfarenheter och expertkunnande tas till vara bättre i processen när vi utarbetar vetenskapliga yttranden som är avsedda att utgöra grund för de politiska besluten inom ramen för den gemensamma fiskeripolitiken.
ledamot av kommissionen. - (EN) Herr talman! Jag uppskattar att kunna prata om mitt ansvarsområde.
Kommissionen välkomnar parlamentets betänkande om tillämpad forskning inom den gemensamma fiskeripolitiken och tackar föredraganden Rosa Miguélez Ramos och fiskeriutskottet för ett utmärkt arbete.
Betänkandet kommer lägligt nu när de gemensamma ansökningsomgångarna för havs- och sjöfartsforskning förbereds.
Det sammanfaller också med arbetsprogrammet 2010 för sjunde ramprogrammet och lanseringen av grönboken om en reformering av den gemensamma fiskeripolitiken, som innehåller ett kapitel om forskning.
Kommissionen instämmer i princip med de centrala delarna av betänkandet.
Vi välkomnar att man stöder den europeiska strategin för havs- och sjöfartsforskning, och prioriterar ökad kapacitetsuppbyggnad, ny infrastruktur, nya färdigheter och utbildningsinitiativ, att utveckla samspelet mellan etablerade discipliner för havs- och sjöfartsforskning, samt att främja samverkan mellan medlemsstater och kommissionen och ny forskningsledning.
Kommissionen är medveten om hur viktigt det är att en tillräcklig budget avsätts till forskning inom fiske och vattenbruk i sjunde ramprogrammet, samtidigt som man bör bibehålla en bra balans i förhållande till andra forskningsområden, särskilt inom jordbruk, skogsbruk och bioteknik: tema 2 - KBBE, och tema 6 - miljö.
Årsbudgeten för sjunde ramprogrammet kommer att öka progressivt under programmets tre sista år och både fiske- och vattenbrukssektorn kommer att dra nytta av ökningen.
Kommissionen kommer att forsätta arbetet med att stödja forskningen i linje med betänkandet genom att synliggöra forskningen inom fiske och vattenbruk i sjunde ramprogrammet och skapa en god balans mellan forskning som stödjer politiken och grundforskning, införa mer samhällsvetenskap i arbetsprogrammen, främja spridning av resultat och främja ökad samordning av nationella forskningsprogram.
Slutligen kommer kommissionen att underlätta införlivandet av forskning inom fiske och vattenbruk i sin strategiska forskningsdagordning, det europeiska området för forskningsverksamhet och den nya europeiska strategin för havs- och sjöfartsforskning.
Tack vare de initiativ som jag just har nämnt, känner jag att det finns en fast grund för att förbättra fiske- och vattenbrukssektorn genom innovativ forskning inom ramprogrammet.
Dessa sektorer kommer i sin tur att dra nytta av att den nationella forskningen samarbetar och samordnas på ett bättre sätt, genom de olika initiativen inom det europeiska området för forskningsverksamhet och i samma riktning som den gemensamma fiskeripolitiken.
Om jag får tillägga något mer personligt, kan jag garantera att det inte är mer komplicerat nu än tidigare, helt enkelt beroende på att samma personer arbetar med detta och att vårt samarbete med min kollega Joe Borg går fantastiskt bra.
Det är så forskningen bör bedrivas i framtiden.
Vi samarbetar mellan olika sektorer och det ger bättre resultat, vilket knappast hade varit fallet om det hade gjorts sektorsvis.
Ett stort tack för detta utmärkta arbete.
Punkten är härmed avslutad.
Omröstningen kommer att äga rum på torsdag den 19 februari 2009.
Föredragningslista för nästa sammanträde: se protokollet
18.
Rapport om konkurrenspolitiken 2006 och 2007 (
Inkomna dokument: se protokollet
9. års framstegsrapport om Kroatien (omröstning)
- Före omröstningen om ändringsförslag 13:
för PSE-gruppen. - (DE) Tack, herr talman!
Det har varit många diskussioner mellan grupperna de senaste dagarna, faktiskt ända in i det sista.
Följande ändringsförslag verkar vara det som de flesta i kammaren är överens om och enligt direktinformation som jag har fått har både Kroatien och Slovenien samtyckt till det.
Ändringsförslaget lyder som följer:
för PSE-gruppen.- (EN) ”Europaparlamentet påminner om det informella avtal som Kroatiens och Sloveniens premiärministrar slöt den 26 augusti 2007 om att gränstvisten mellan de båda länderna skulle hänvisas till ett internationellt organ. Parlamentet välkomnar Kroatiens och Sloveniens beredskap att acceptera kommissionens erbjudande om medling och anser att denna medling måste bygga på folkrätten.
Konststudier i Europeiska unionen (kortfattad redogörelse)
Nästa punkt är ett betänkande av Maria Badia i Cutchet, för utskottet för kultur och utbildning, om konststudier inom Europeiska unionen.
Herr talman! Konstutbildning är numera ett obligatoriskt ämne i nästan alla medlemsstater, men det förekommer stora skillnader i hur undervisningen bedrivs.
Tidigare kopplades konststudier till undervisningen av barn och ungdomar, men nu har inriktningen på livslångt lärande och utvecklingen av den nya informations- och kommunikationstekniken (IKT) lett till att konstens och kulturens traditionella utrymme har utvidgats, vilket har gett upphov till nya former av tillgång till och uttryck inom sektorn.
Den kontinuerliga IKT-utvecklingen har även bidragit till att främja en kunskapsekonomi, vilket har lett till att intellektuell och kreativ förmåga har blivit ett viktigt inslag i denna nya ekonomi.
Det förslag till resolution som vi ska rösta om i morgon bygger på tanken att konstutbildning utgör grunden för yrkesutbildningen inom detta område och främjar kreativiteten och den fysiska och intellektuella utvecklingen. Den är också en viktig komponent i barn- och ungdomsutbildningen och konstundervisning i skolan lägger grunden till en verklig demokratisering av tillgången till kultur.
Utbildningen också mycket viktig för framgången för de yrkesverksamma inom den konstnärliga och kreativa sektorn, eftersom konststudier som inriktas på karriär- och yrkesutveckling kräver, förutom talang, att eleverna har en gedigen kulturell grund att bygga på som endast är möjlig att förvärva genom en tvärvetenskaplig och systematisk utbildning.
Detta ökar möjligheten att ta sig in på arbetsmarknaden inom denna sektor eftersom eleverna förvärvar allmänna kulturella kunskaper, forskningsmetoder, företagarkunskaper och affärskunskaper samt kompetenser inom olika verksamhetsområden.
Dessutom ges ett mycket speciellt erkännande av den ekonomiska potentialen hos de företag och industrier som är verksamma inom det kreativa, kulturella och konstnärliga området i EU, som ger ett större bidrag än andra starkt uppmärksammade industrier som kemi- och livsmedelsindustrierna.
Vi får inte heller glömma att konstskolor och konstutbildnings- och formgivningscentrum bidrar till att utveckla nya konstnärliga stilarter och rörelser, samt öppna olika kulturvärldar, vilket förstärker EU:s framtoning i världen.
I förslaget till betänkande betonas att konstämnen bör vara obligatoriska i läroplanerna på alla utbildningsnivåer och medlemsstaterna uppmuntras att samordna sin konstpolitik på EU-nivå och främja både studenters och lärares rörlighet på detta område, samt att i högre grad uppmärksamma frågan om erkännande av kvalifikationer mellan medlemsstater.
Vi uppmanar även rådet, kommissionen och medlemsstaterna att fastställa konstutbildningens roll som ett mycket viktigt pedagogiskt verktyg för att öka kulturens värde, utforma gemensamma strategier för att främja politik för konstutbildning, utbilda ämneslärarna och att erkänna den viktiga roll som konstnärer spelar i samhället, vilket framgick av Europeiska året för kreativitet och innovation.
Slutligen understryks vikten av att utnyttja de resurser som den nya informations- och kommunikationstekniken och Internet erbjuder som kanaler för en modern och nutidsanpassad undervisning när det gäller att införa den konstnärliga dimensionen i läroplanerna. En europeisk portal för konst- och kulturutbildning bör tas fram gemensamt för att garantera utvecklingen och främjandet av den europeiska kulturella modellen.
Av alla dessa skäl uppmanar jag majoriteten att stödja betänkandet som kommer att ge ett tydligt budskap om stöd till yrkesverksamma, studenter och företag inom den kreativa och kulturella sektorn.
Herr talman, mina damer och herrar! Först av allt vill jag tacka Maria Badia i Cutchet för hennes initiativbetänkande om konststudier inom Europeiska unionen.
Konststudier får ett allt viktigare utrymme på EU-nivå.
Vi är alla överens om att kultur och konst är en mycket viktig del av utbildningen.
De bidrar till att utveckla känslighet och självförtroende, nödvändiga egenskaper inte bara för vår roll som medborgare utan också för den ekonomiska aktör som vi alla har inom oss.
Detta råder det ingen tvekan om.
Konstutbildning är en källa till välmående, kreativitet och social integration.
Det är mycket viktigt att denna utbildning främjas i EU:s utbildningssystem från så unga år som möjligt.
Vi delar denna vision och vi gläder oss över att det i ert betänkande hänvisas till flera viktiga initiativ på EU-nivå, t.ex. Europeiska året för kreativitet och innovation.
Konstens och konstutbildningens betydelse för att bygga ett bättre samhälle går hand i hand med dess inverkan på det ekonomiska livet.
Enligt färska beräkningar uppskattas de kulturella och kreativa industriernas bidrag till det ekonomiska välståndet till 2,6 procent av EU:s BNP.
Dessutom kan all ekonomisk verksamhet dra fördel av utbildningen i konst och kultur.
Innovation uppmuntrar till att skapa synergieffekter mellan traditionella verksamhetsområden och mer innovativa sådana.
I dag måste vi kombinera teknik och design samtidigt som vi integrerar principerna om hållbarhet och ekonomisk lönsamhet.
Denna kombination kräver en ny definition av hur kunskap ska överföras och förvärvas.
Dessa olika frågor behandlas i dokumentet om den europeiska referensramen där nyckelkompetenser för livslångt lärande definierades 2006.
Inom denna ram konstateras det att konstnärliga och kulturella uttryck är nödvändiga för att utveckla kreativ kompetens, som är så användbar i arbetslivet.
I den europeiska agendan för kultur presenteras nya metoder, särskilt en strukturerad dialog med det civila samhället och nyligen även nya öppna metoder för kulturell samordning.
Dessa metoder har kunnat tillämpas tack vare en första treårig arbetsplan som rådet antog den 21 maj 2008 och där det anges fem prioriterade insatsområden.
Inom denna ram inrättades en arbetsgrupp av sakkunniga från medlemsstaterna som skulle arbeta på temat synergieffekter mellan kultur och utbildning.
Denna grupp kommer att utforma rekommendationer för att identifiera goda metoder på nationell nivå och även utfärda ett antal rekommendationer till medlemsstaterna och EU-institutionerna.
Dessutom kommer den att ta fram metoder för att bedöma framstegen inom de politikområden som omfattas av dess mandat.
Slutligen bör gruppen kunna ge ett värdefullt bidrag till Europeiskt kulturforum som ska hållas den 29-20 september 2009 i Bryssel.
Jag har precis läst ett svar från min kollega i kommissionen, Ján Figel'.
Punkten är avslutad.
Omröstningen kommer att äga rum tisdagen den 24 mars 2009.
Skriftliga förklaringar (artikel 142)
Europaparlamentets betänkande om konststudier inom EU ingår i de kontinuerliga insatserna för att utveckla den interkulturella dialogen och är mycket viktiga i samband med Europeiska året för kreativitet och innovation.
Konstutbildningen måste utan tvivel ägnas större och mer specifik uppmärksamhet.
Det är viktigt att den är en obligatorisk del av läroplanen så tidigt som möjligt, eftersom den stimulerar den känslomässiga och kulturella utvecklingen hos den unga generationen.
Genom att ge dessa studier ett större praktiskt syfte och införa interaktiv undervisning skulle vi kunna få en djupare förståelse av nationella och europeiska kulturella värderingar.
Genom att ge elever, lärare och yrkesverksamma inom sektorn ökad rörlighet kan vi direkt skapa medvetenhet om den europeiska identiteten och skapa kulturell och religiös tolerans.
Medlemsstaterna måste investera för att skapa bättre möjligheter till informella och oberoende konststudier och förhindra att antalet program på detta område minskar.
Deras stöd till konstnärers yrkesliv skulle öka det allmänna intresset för olika former av konststudier.
Offentlig-privata partnerskap på detta område skulle bidra till att modernisera utbildningsprogrammen och uppmuntra till en mer aktiv integration av ny teknik i undervisningsprocessen.
Större delen av resurserna för en samordnad EU-politik för konststudier utgörs av investeringar för att förstärka EU:s kulturella inflytande globalt, förstärka kreativiteten och, indirekt, EU:s ekonomi.
5.
EU:s prioriteringar för den 64:e sessionen i FN:s generalförsamling (
21.
Ett europeiskt initiativ för mikrokrediter för att främja tillväxt och sysselsättning (
3.
Det europeiska flygsystemets kvalitet och hållbarhet (
- Före omröstningen:
föredragande. - (RO) Parlamentet har enats med rådet. Uppgörelsen stöds av fem partigrupper.
Jag avser här de två följande betänkandena.
Tack vare de ändringsförslag som lagts fram av två ledamöter här - innehållet i ändringsförslagen har förresten redan införts i den kompromiss som vi enats om med rådet - måste vi i dag rösta om flera artiklar.
På grund av regler som jag anser är felaktiga innehåller omröstningsordningen i vissa av artiklarna först texten från utskottet för transport och turism, och sedan kompromisstexten.
Jag vill helst att vi röstar om kompromisstexten i dag, eftersom den har stöd av samtliga fem partigrupper, så att de två förordningarna kan träda i kraft i slutet av denna mandatperiod.
- Tack för era synpunkter.
Vi kommer faktiskt att komma dit ni önskar genom att följa omröstningsordningen och rösta om ändringsförslagen.
20.
Bilindustrins framtid (omröstning)
- Före den slutliga omröstningen:
- (DE) Fru talman! Jag hänvisar till artikel 146 i arbetsordningen och tackar er för ordet.
Jag ber särskilt mina tyska ledamotskollegor om överseende för att jag bett om ordet nu.
När omröstningen började tog Jean-Marie Le Pen till orda.
När han fått ordet upprepade han att gaskamrarna i Auschwitz var en historisk detalj.
Med hänvisning till artikel 146 i arbetsordningen, som fastställer hur ledamöterna ska uppträda i kammaren, uppmanar jag parlamentets presidium att undersöka om ett sådant yttrande är tillåtet i ett parlament där ledamöterna har utfäst sig att uppträda i en anda av försoning, förståelse och aktning för offren, i synnerhet för Hitlers fascism.
Jag skulle uppskatta om parlamentets presidium underrättar oss om vilka åtgärder som bör vidtas.
(Applåder)
- (FR) Jag ber er att visa lite aktning för de offer som dog i Auschwitz och på andra ställen.
Vi har fortfarande två minuter kvar.
Visa lite aktning.
Det enda jag vill säga är att jag helt håller med Martin Schulz, och att vi har fått höra helt omotiverade yttranden här i kammaren i dag.
(Applåder)
- (FR) Fru Wallis, jag tycker att det är väldigt tråkigt att ni gav ordet till Joseph Daul och Martin Schulz, men inte till mig.
Men å andra sidan har ni ju själv i ett betänkande medgett att ni är expert på att tolka arbetsordningens särbehandlande artiklar.
Låt mig därför komplettera Martin Schulz inlägg genom att föreslå att vi döper om Winston Churchill-byggnaden, eftersom Churchill i sina tolv memoarvolymer om andra världskriget inte skriver en rad om gaskamrarnas historia.
Vitbok om skadeståndstalan vid brott mot EG:s antitrustregler (debatt)
- Nästa punkt är betänkandet av Klaus-Heiner Lehne för utskottet för ekonomi och valutafrågor om vitboken om skadeståndstalan vid brott mot EG:s antitrustregler -.
föredragande. - (DE) Herr talman, mina damer och herrar! Låt mig först tacka skuggföredragandena, särskilt Antolín Sánchez Presedo för socialdemokraterna och Sharon Bowles för liberalerna, med vilka jag har haft ett mycket lyckat samarbete om den kompromisstext som läggs fram idag i form av ett betänkande om kommissionens vitbok.
Den här gången har vi lyckats få till stånd en mycket stor majoritet tvärsöver grupperna och en verkligt genomförbar kompromiss som även kan vägleda Europeiska kommissionens, och senare under lagstiftningsprocessen, Europaparlamentets framtida arbete.
Vi har i detta betänkande gjort klart - och detta med rätta - att när det gäller överträdelser av konkurrensreglerna så står parlamentet fast vid sin ståndpunkt att detta enligt europeisk tradition i första hand är en sak för myndigheterna - såväl nationella konkurrensmyndigheter som den europeiska konkurrensmyndigheten - och att det inte handlar om att skapa en andra arm som så att säga står på jämlik fot med myndighetsåtgärder i kampen mot karteller.
I Europa har vi medvetet valt en annan väg än i USA, som man ofta gör jämförelser med.
Det finns en politisk enighet i parlamentet om att vi behöver ett tvistlösningsförfarande för s.k. masskadeståndsanspråk.
Om enskilda personers olagliga beteende skadar ett mycket stort antal människor som har lidit jämförelsevis små förluster behövs en separat lösning för sådana processer eftersom den normala processrätten helt enkelt inte är tillräckligt effektiv.
Inrättandet av ett sådant instrument är också ett led i att göra det möjligt att väcka talan och vidareutveckla den inre marknaden.
Om detta är vi överens.
Det rådde också enighet om att vi inte vill att det ska växa fram en stämningsindustri i Europa liknande den i USA som omsätter 240 miljarder dollar och i slutändan inte gynnar konsumenterna, utan - som var och en vet som har läst de relevanta böckerna - i första hand gynnar de amerikanska advokatbyråerna.
Inget av detta har särskilt mycket att göra med rättssäkerhet och det vill vi inte heller.
Vi enades om att det amerikanska systemets processrättsliga tortyrinstrument inte bör införas i Europa.
Detta gäller i synnerhet bevisupptagning och kostnader.
Det är en mycket viktig punkt.
Vi enades också om att vi i huvudsak anser att lagstiftningen på EU-nivå rent principiellt bara kan vara en lösning baserad på en möjlighet att delta i ett senare skede (opt-in) och att en lösning baserad på en möjlighet att avstå (opt-out) bara kan tillåtas om medlemsstaterna redan har en liknande lösning och detta är tillåtet enligt den nationella konstitutionen.
En möjlighet att delta i ett senare skede är inte tillåten enligt alla länders nationella konstitution och strider också mot principen om den vuxne konsumenten.
Som vi enträget klagar över har Europeiska kommissionen helt glömt bort att behandla frågan om tvistlösning utanför domstolarna i sin vitbok.
Generaldirektoratet för konkurrens och kommissionen går rakt på processandet.
Som vi sedan flera år tillbaka vet till följd av debatterna i detta parlament om politiken i rättsliga frågor är detta emellertid inte alltid det bästa sättet utan tvistlösningsmekanismer utanför domstolarna är ofta mycket lämpligare för att lösa problem.
Det arbete som generaldirektoratet för konsumentskydd har genomfört parallellt om samma fråga har dessutom kommit mycket längre.
Detta generaldirektorat använde en bred marginal för dessa alternativa tvistlösningsinstrument i sin grönbok, som befinner sig i samrådsstadiet före det här.
Vi menar att Europeiska kommissionen omgående måste se över denna fråga.
En sista poäng, som också är avgörande: vi vill inte ha någon fragmentering av lagstiftningen.
Nu rusar konkurrenslagstiftningen iväg och skapar ett sådant instrument.
Konsumentskyddet rullar på beträffande samma fråga.
Vi vet att något liknande förr eller senare kommer att övervägas när det gäller kapitalmarknadslagstiftningen, miljölagstiftningen och sociallagstiftningen.
Vi anser att det är absolut nödvändigt att man även överväger en horisontell strategi och att vi åtminstone stöder de förfarandemässiga instrument som är mer eller mindre identiska inom alla områden med ett horisontellt instrument.
Även detta är av avgörande betydelse.
ledamot av kommissionen. - (EN) Herr talman! Jag välkomnar på kommissionens vägnar det betänkande av Klaus-Heiner Lehne som har antagits av utskottet för ekonomi och valutafrågor (ECON) - antagits som en symbol för en stark enighet mellan de politiska grupperna.
Det gläder oss också att vitboken får starkt stöd i detta betänkande.
Kommissionen noterar att man i betänkandet instämmer med vitbokens slutsatser om att offer för överträdelser av EG:s konkurrenslagstiftning i dagsläget har stora svårigheter att få skadestånd för de förluster som de har lidit.
Vi instämmer i att åtgärder måste vidtas så att dessa offer kan få full ersättning.
Vi delar också uppfattningen att kollektiva prövningsmöjligheter är avgörande för att konsumenter och småföretag ska ha en realistisk och effektiv möjlighet att få ersättning i fall av spridda skador.
Kommissionen instämmer också till fullo med ECON-utskottets betänkande om att ett överutnyttjande eller missbruk av möjligheten till domstolsprövning måste undvikas.
Det måste därför finnas lämpliga garantier i mekanismerna för kollektiv prövning.
Vi instämmer slutligen till fullo med att man måste vara konsekvent när det gäller kollektiva prövningsmöjligheter och att man därför måste se till att initiativ inriktade på olika områden, t.ex. konkurrenslagstiftningen och eller lagar om konsumentskydd, är förenliga med varandra.
Kommissionen välkomnar samtidigt erkännandet att en enhetlig strategi när det gäller kollektiv prövning inte nödvändigtvis innebär att alla områden måste hanteras genom ett enda horisontellt instrument.
Kravet på enhetlighet får inte leda till att utformningen av de åtgärder som bedöms vara nödvändiga för att EG:s konkurrenslagstiftning ska kunna genomföras fullt ut i onödan skjuts upp.
föredragande av yttrandet från utskottet för den inre marknaden och konsumentskydd. - (RO) Utskottet för den inre marknaden och konsumentskydd har formulerat sin ståndpunkt utifrån en viss omständighet: nämligen att de negativa effekterna av överträdelser av antitrustlagstiftningen mycket ofta blir ekonomiskt kännbara i slutet av den kommersiella kedjan genom att drabba slutkonsumenter och småföretag.
I det här fallet är det viktigt men samtidigt svårt att få skadestånd för förluster eftersom det finns många drabbade och det rör sig om små summor.
Vi har därför krävt ett paket bestående av lagstiftning och andra åtgärder som kan bli det verktyg som alla EU-medborgare som hamnar i en sådan situation kan använda för att hävda sin rätt till fullständig och lämplig ersättning.
Vi ställer oss bakom alla åtgärder för att undanröja svårigheterna att nå detta mål: enklare tillgång till handlingar, lägre rättegångskostnader och omvänd bevisbörda.
Vi välkomnar kommissionens förslag att kombinera grupptalan som väcks av behöriga parter och kollektiv talan med uttryckligt medgivande.
Vi anser dock att kollektiv prövning med möjlighet att avstå måste diskuteras ytterligare med tanke på de fördelar som detta medför: en ”en gång för alla”-lösning och mindre osäkerhet.
Trots att det finns ett tydligt förbud mot karteller och andra brott mot konkurrenslagstiftningen i EU-fördraget är det fortfarande svårt för drabbade konsumenter i Europeiska gemenskapen att hävda sin rätt till ersättning.
I Rumänien fick exempelvis en kartell som bildats inom cementindustrin nyligen böta flera miljoner euro.
Men enligt den nuvarande lagstiftningen har de myndigheter som har till uppgift att övervaka konkurrensen ingen skyldighet att hantera frågan om ersättning till drabbade.
Jag vill understryka att dessa myndigheter måste ta hänsyn till den ersättning som betalas eller borde betalas när de bestämmer böter för företag som befinns vara skyldiga till oegentligheter, så att det inte råder en bristande överensstämmelse mellan den skada som åsamkas och det straff som utdöms, och att framför allt se till att skadestånd betalas ut till dem som drabbas av ett sådant agerande.
Jag välkomnar därför kommissionens plan att förbättra metoderna att garantera rättigheterna för konsumenter som drabbas av överträdelser av lagstiftningen över hela Europa.
Parlamentet slog mycket tydligt fast att Europa inte ska ha något system med möjlighet att avstå.
Offren måste därför identifieras så snabbt som möjligt i samband med att det inkommer ett klagomål.
Genom systemet med möjlighet till deltagande i ett senare skede ser man till att de som drabbas av överträdelser av konkurrenslagstiftningen verkligen får ersättning.
Parlamentet vill inte att någon annan, exempelvis advokater, branschorganisationer eller konsumentverket, ska gynnas av en enskild talan.
Jag anser också att parlamentet tillför ett nytt och viktigt inslag som inte fanns med i kommissionens förslag.
Alternativa tvistlösningsmekanismer är i många fall mycket effektivare än rättegångar för offer som har rätt till ersättning.
Jag menar att när ersättning krävs måste man i första hand försöka nå en uppgörelse utanför domstol.
Detta medför betydligt lägre kostnader än en enskild talan eftersom konsumenterna får snabbare ersättning för sina förluster.
för PSE-gruppen. - (EN) Herr talman, herr kommissionsledamot, mina damer och herrar! Detta betänkande har godkänts enhälligt i utskottet för ekonomi och valutafrågor.
Det är inte bara ett fantastiskt resultat utan också, med tanke på hur svåra, komplicerade och kontroversiella dessa frågor är, ett exceptionellt resultat, som bör driva på och fast förankra den nya pelaren för enskild talan, som är absolut nödvändig för att göra principen om gemenskapens behörighet effektiv.
Detta är ett nytt steg i riktning mot en mer avancerad och effektiv ansvarspolitik som i högre grad respekterar offrens rättigheter och på ett effektivare sätt ställer den som gör sig skyldig till överträdelser till svars.
Jag vill därför börja med att gratulera föredraganden Klaus-Heiner Lehne, som har haft det övergripande ansvaret för att ro detta arbete i hamn.
Hans idéers kvalitet, hans öppna sinne och vilja att föra en dialog och hans intelligens när det gäller att finna de bästa kompromisserna har spelat en avgörande roll för detta.
Jag vill gratulera föredragandena av yttrandena, skuggföredragandena och de som har lagt fram ändringsförslag, vars positiva bidrag har förbättrat betänkandet ytterligare.
Kommissionens vitbok om ”skadeståndstalan vid brott mot EG:s antitrustregler” är ett svar på Europaparlamentets begäran i resolutionen om grönboken, vars innehåll parlamentet i stora drag godkände.
Så var t.ex. fallet när man uttalade sig gillande om komplementariteten mellan offentlig och enskild talan och var positiv till kollektiv prövning, men ville undvika de överdrifter som gruppstämningar har lett till i USA, och därmed göra det lättare att få skadestånd, och när man föreslog tillgång till relevant information under domstolarnas kontroll, men inte eftersökningar utan skälig misstanke, och när man erkände och krävde en möjlighet att väcka självständig talan, uppföljande talan eller ett frivilligt ersättningssystem.
Man tar i betänkandet ställning för Europaparlamentets medbeslutande i fastställandet av ett regelverk för skadeståndstalan vid brott mot EG:s antitrustregler.
Detta ska inte tolkas som att man förnekar policyn om gemenskapens behörighet som rättslig grund för lagstiftning, utan som en uppgradering av kraven i det vanliga förfarandet på detta område för att nå upp till de högre värden som erkänns i fördraget.
När en förordning får en betydande inverkan på en grundläggande rättighet, t.ex. medborgarnas rätt till ett effektivt rättsskydd - som ingår i EU:s och medlemsstaternas system - kräver den demokratiska principen och respekten för nationella rättsliga traditioner - enligt vilka dessa frågor bara får regleras genom bestämmelser på rättslig nivå eller, med andra ord, genom att direkta företrädare för allmänheten väcker talan - att Europaparlamentet deltar i lagstiftningsprocessen.
Det fastställs också ett horisontellt och integrerat tillvägagångssätt att hantera gemensamma problem som möjligheten att väcka enskild talan med stöd av konkurrenslagstiftningen kan ge upphov till på andra områden, varigenom man undviker ett splittrat och inkonsekvent angreppssätt.
En privat talan får väckas av ett offentligt organ samt genom en enskild talan eller grupptalan.
Den sistnämnda kan väckas direkt av de drabbade eller indirekt genom behöriga parter utsedda i förväg eller ad hoc, t.ex. konsument- eller branschorganisationer.
Om en talan väcks av en behörig part ska gruppen av offer beskrivas i stämningsansökan, men deras identitet kan anges senare, även om det ska ske så snabbt som möjligt för att undvika onödiga dröjsmål och uppfylla kraven i den befintliga lagstiftningen.
Denna lösning är mycket viktig för fall som rör mindre och spridda skador.
I betänkandet tas frågan om tillgång till information som är nödvändig för att väcka en uppföljande talan upp på ett balanserat sätt.
Skyddet av affärshemligheter måste säkerställas, liksom effektiviteten i programmet för förmånlig behandling, för vilket man vill ha riktlinjer.
Villkor fastställs för att beslut som fattas av en myndighet som ingår i gemenskapens nätverk av konkurrensmyndigheter ska kunna bli bindande i andra medlemsstater och för att man med full respekt för principen om skadeståndsansvar ska kunna tillämpa omvänd bevisbörda, dvs. att man antar att det föreligger en förseelse eller skuld om ett brott har påvisats.
Det är också värt att ta upp godkännandet av försvarsargument om ”övervältrade kostnader” för indirekta offer och ett system som förenklar och minskar rättegångskostnaderna.
Jag vill också betona det positiva samspelet mellan offentlig och privat talan för att både skapa incitament för ersättning till drabbade och när det gäller fastställandet av en femårsperiod för väckande av talan.
Låt mig till sist tacka kommissionen för den dialog som har förts under hela detta förfarande och be kommissionsledamoten att utan dröjsmål lägga fram de initiativ som krävs för att den ska kunna fortsätta.
för ALDE-gruppen. - (EN) Herr talman! Jag vill börja med att tacka Klaus-Heiner Lehne för hans betänkande och bekräfta att min grupp kommer att ge det sitt stöd.
Jag vill också säga att jag tycker att det är lite märkligt att vi har den här debatten sent på kvällen när vi kommer att behandla en fråga om samma ämne i morgon bitti.
Det hade varit en mycket god idé att behandla båda på samma gång.
Låt mig i mitt beröm av betänkandet säga att utgångspunkten för min grupp har varit att ”skipa rättvisa” - att skipa rättvisa för små och medelstora företag och konsumenter över hela EU som ställs inför ett oegentligt och konkurrensbegränsande agerande.
För ett par veckor sedan organiserade min grupp ett seminarium på parlamentet i Bryssel och några av våra besökare som fått känna av de negativa effekterna av ett sådant konkurrensbegränsande beteende, ironiskt nog inom cementindustrin, gjorde ett mycket starkt intryck på mig.
Vad sa de?
Snälla, snälla, se till att driva igenom det här: vi behöver något så att vi kan vidta åtgärder mot dessa oegentliga aktörer på den europeiska marknaden.
Vi vill ha en europeisk lösning och vi vill ha den snabbt, för om vi inte får den är min prognos och varning följande: några av våra medlemsstater kommer att utveckla system som leder till ”forum shopping” till följd av den fria rörligheten för domstolsbeslut.
Så, snälla - ett europeiskt system så snart som möjligt.
- Jag ska se till att er synpunkt beträffande föredragningslistan vidarebefordras till talmanskonferensen som fastställer föredragningslistan - ibland gör de misstag.
för IND/DEM-gruppen. - Herr talman! Den inre marknaden är EU:s absolut förnämsta bidrag till frihet och välstånd i Europa.
Den förutsätter bland annat en effektiv antitrustlagstiftning.
Det vi nu begrundar är frågan om skadeståndstalan vid brott mot antitrustlagstiftningen.
Det finns goda principiella skäl för att medborgare och företag ska kunna kräva skadestånd.
Klaus-Heiner Lehnes betänkande visar, delvis oavsiktligt, på problemen och riskerna.
Vitboken talar om en europeisk rättskultur, men någon sådan finns inte.
Vi ska inte skapa regelverk byggda på önsketänkande.
Föredraganden menar att vi undviker en amerikanisering av skadeståndskulturen.
Det är också ett önsketänkande.
Riskerna för en sådan är tvärtom stora.
Ansvarsfördelningen mellan EU:s institutioner och medlemsländernas förbigås.
Det finns ingen objektiv och förutsättningsanalys av vad subsidiaritetsprincipen säger.
Principen tas helt enkelt inte på allvar.
Det finns också många andra oklarheter och risker för godtycke.
Punkterna 7 och 11 inger tillsammans farhågor.
En självklar utgångspunkt måste vara en skadeståndstalan på grund av brott mot antitrustlagstiftning.
Den kräver att brottet har fastställts i domstol. Därefter måste rimligen res judicata gälla även inom ramen för enskild talan så att domen inte kan omprövas om det gäller samma fall.
Punkterna 15 och 18 tillsammans öppnar för käranden att välja den rättsordning som är mest förmånlig.
Det skapar rättsosäkerhet och det leder till sådan här "form shopping" som blir ett rejält hot.
Informationsassymetrin ska minskas genom att företagen tvingas lämna ut information till käranden.
Det medför en subjektiv hantering av viktig affärsinformation som kan missbrukas.
Det finns alldeles för många oklarheter och risker på detta stadium.
Kammaren bör därför säga nej till detta betänkande och begära en grundligare genomlysning av frågan innan vi går till beslut.
- (DE) Herr talman, mina damer och herrar!
Först ett mycket stort tack till föredraganden Klaus-Heiner Lehne, som har gjort en storartad insats och tillsammans med ledamöterna från de andra grupperna har hittat bra lösningar på en mycket svår fråga.
Det framgår av debatten att vi alla är överens om att vi behöver en horisontell strategi för alla kollektiva skadeståndsanspråk och jag ber därför kommissionen att inte lägga fram separata förslag från olika generaldirektorat för varje enskilt område, utan i stället ge oss en verkligt kollektiv prövningsmekanism som omfattar alla områden för den europeiska inre marknaden och för EU:s medborgare och naturligtvis - som Diana Wallis påpekade - för europeiska små och medelstora företag.
Vi är överens om att man effektivt måste försvara rättigheterna för dem som skadas av karteller och att vi måste införa kartellkontroll i den europeiska ekonomin i enlighet med den sociala marknadsekonomins princip. Vi vill inte heller att olika nationella bestämmelser missbrukas genom ”forum shopping”.
Kvällens debatt har emellertid inte gett mig särskilt mycket information om hur detta bäst kan uppnås, för jag anser att potentialen hos kollektiva prövningsmöjligheter ofta överskattas.
Det är därför viktigt att än en gång slå fast vissa riktmärken mot vilka vi kan mäta alla kollektiva skadeståndsanspråk.
Vi måste besvara frågan om det behövs ett ökat rättsskydd för konsumenter eller offer i massanspråk, gränsöverskridande rättsprocesser och rättsprocesser som berör mer än en medlemsstat.
Vi måste ta hänsyn till medlemsstaternas processrättsliga begränsningar - möjligheten att avstå, frivillig anslutning och flera andra punkter - i det europeiska förfarandet.
Om detta helt enkelt inte går, som kommissionen själv redan delvis har medgett, så måste vi få med oss medlemsstaternas rättsakter och få till stånd ett gemensamt förfarande med medlemsstaternas parlament för att värna de europeiska konsumenternas intressen.
Vi vill absolut undvika kollektiva skadeståndsanspråk i Europa av amerikansk modell.
Vi vill se till att ersättning betalas ut, men bara till dem som verkligen har drabbats av förluster.
Vi vill å det starkaste avråda från ogrundade anspråk och vi vill främja alternativa tvistlösningsförfaranden.
Herr talman! Jag vill också rikta ett tack till Klaus-Heiner Lehne för ett bra och genomarbetat betänkande som tar upp viktiga frågor inom konkurrensrätten och ger stärkt konsumentskydd.
EG-domstolen ger personer och företag rätt till skadestånd vid brott mot konkurrensreglerna, men trots detta har det i praktiken varit så att de personer som lidit skada beroende på brott mot EG:s antitrustregler sällan fått ersättning.
Vi måste därför få till mekanismer som ökar förtroendet och underlättar för personer att kunna hävda sin rätt över gränserna.
Vi vet att konsumenter och småföretag skräms av att inleda processer på grund av oro för långdragna processer och framför allt höga kostnader.
Förändringar i denna riktning kommer att främja handel över gränserna.
Ska vi få en fungerande inre marknad inom hela EU, där personer kan lita på att få sin sak prövad på ett rättssäkert sätt och få full ersättning för den uppkomna skadan, förlusten, då måste vi också hitta nya mekanismer som underlättar grupptalan.
När vi talar om grupptalan kommer alltid USA upp och de amerikanska erfarenheterna och överdrifterna.
Vi måste givetvis dra lärdom av detta, men inte låta oss skrämmas.
Europa ska ha ett europeiskt system, inte ett amerikanskt.
Om vi inte gör någonting kommer situationen bara att bli sämre.
ledamot av kommissionen. - (EN) Herr talman! Tack allihop för mycket intressanta inlägg, i synnerhet Klaus-Heiner Lehnes inledande redogörelse.
Detta var mycket intressant och jag förstår nu varför ni är så eniga och samarbetar om dessa frågor, inte bara i utskottet utan även i parlamentet.
Det finns inte mycket som jag kan tillägga, förutom måhända när det gäller de rättsliga grunderna.
Det beror naturligtvis på målen och innehållet i den föreslagna åtgärden, och jag vill som kommissionsledamot försäkra er - kanske rör det ett annat politikområde, men jag talar på kommissionens vägnar - om att vi principiellt strävar efter ett mycket nära samarbete med parlamentet.
Hur detta ska ske i en praktisk konkret fråga återstår att se, men vi kommer att sträva efter ett nära samarbete eller ett så nära samarbete som möjligt med parlamentet enligt den tillämpliga rättsliga grunden.
När det gäller vad ni sa om fragmentering och en horisontell strategi anser jag att kommissionens svar - och det framgår mycket tydligt i vitboken - är en enhetlig, samstämmig strategi, och jag menar att den europeiska rättstraditionen och vår rättskulturs rötter skiljer sig från det flitigt omnämnda amerikanska systemet.
Jag tror dock att vi kan lära av andra och förbättra vårt system.
När det gäller offentliga myndigheters upprätthållande av lag och rättvisa anser jag naturligtvis att det är mycket viktigt att vi inte går mot en försämring av detta upprätthållande och artiklarna 81 och 82 är förstås mycket viktiga pelare för EU:s inre marknad och inremarknadspolitik.
De handlar om rättsliga frågor och skadeståndstalan är ett komplement till detta upprätthållande.
Sist - men kanske inte minst - det som sas om tvistlösning utanför domstol.
Kommissionen är för detta, men en förutsättning för en sådan strategi, som skulle vara välkommen, är att det finns ett fungerande och effektivt processrättsligt system för skadeståndsanspråk i medlemsstaterna.
Jag tror därför att vi inte bara måste uppmuntra utan även hjälpa våra medlemsstater så att sådana frågor och system finns i EU-27.
Då tror jag att vi även kan ta itu med dessa punkter.
Men låt mig principiellt tacka er så mycket för vad som även för mig har varit en mycket intressant debatt och lycka till!
föredragande. - (DE) Herr talman, herr kommissionsledamot! Låt mig först tacka mina ärade kolleger för deras mycket bra inlägg.
Jag tycker att vi med gemensamma krafter uppnådde ett bra resultat.
Jag vill emellertid också tydligt poängtera för kommissionen, så att det inte råder några missförstånd: ur parlamentets synvinkel är det inte tal om att ni ska anta ett lagförslag som förmodligen redan är helt odugligt.
Absolut inte.
Vi förväntar oss att kommissionen tar hänsyn till det som vi har beslutat idag och integrerar det i det faktiska lagförslaget.
Den horisontella strategin är inte bara en viktig aspekt av de skäl som jag tidigare beskrev närmare. Kommissionsledamoten tog dessutom själv upp frågan om rättslig grund.
Med ett sådant viktigt projekt måste man välja en strategi som i slutändan ser till att parlamentet deltar som lagstiftare på jämlik fot.
Väljer man en strategi som enbart baseras på konkurrensrätten så blir detta inte fallet enligt det nu gällande Nicefördraget.
Detta är också ett mycket grundläggande politiskt argument för varför vi anser att en horisontell strategi är den rätta.
Jag tycker att kommissionen mycket allvarligt ska överväga detta.
En annan avgörande punkt enligt min uppfattning är att vi fortfarande behöver något när det gäller frågan om tvistlösning utanför domstol.
Ni talade tidigare om konvergens med det arbete som har utförts av generaldirektoratet för konkurrens.
Men om man jämför grönboken om konsumentskydd med vitboken om konkurrens får man inte direkt intrycket att det finns någon sådan konvergens.
Det mest påfallande exemplet är skillnaden i behandling - eller närmare bestämt bristen på behandling - av mekanismer för tvistlösning utanför domstol i vitboken.
Det finns fortfarande en rad andra problem som vi förväntar oss ska lösas.
Låt mig bara helt kort ta upp frågan om tillgång till Europeiska kommissionens handlingar.
Det är i alla rättegångsförfaranden som gäller skadeståndsanspråk möjligt att granska den offentliga åklagarmyndighetens ärenden.
Varför gäller inte detta Europeiska kommissionen?
Det övergår mitt förstånd.
Detsamma gäller frågan om fastställande av böter: även detta måste beaktas utifrån synvinkeln att det måste vara möjligt att kräva ersättning i framtiden.
Även här måste kommissionen omgående skriva om texten och lägga fram mer konkreta texter och förslag än de som nu ingår i vitboken.
Låt mig för att undvika missförstånd göra klart att ur parlamentets synvinkel förväntar vi oss mer än vad som ingår i vitboken och vi förväntar oss också att generaldirektoratet för konkurrens som helhet följer våra förslag. Annars kommer det att finnas ett motstånd här i parlamentet.
- Jag tackar för era inlägg i denna viktiga fråga och riktar också ett tack till kommissionsledamoten, personalen och tolkarna.
Debatten är härmed avslutad.
Omröstningen kommer att äga rum torsdagen den 26 mars 2009.
Skriftliga förklaringar (artikel 142)
skriftlig. - (ET) I parlamentets betänkande betonas att sprogram för förmånlig behandling kan vara användbara för att upptäcka karteller och det gläder mig att kunna meddela att det estniska parlamentet just nu diskuterar ett förslag till program för förmånlig program.
Detta bör bli ett viktigt inslag i kampen mot karteller, som är viktig både för att den gemensamma marknaden ska fungera bättre och för att skydda konsumenternas rättigheter, eftersom konsumentpriserna kan stiga med så mycket som 25 procent till följd av karteller.
Jag tror dock att företrädartalan också kan spela en viktig roll för ett effektivt genomförande av konkurrenslagstiftningen och ett bättre konsumentskydd och därför måste vi även uppmärksamma detta, både i Estland och inom EU.
Forskning har visat att företrädartalan skulle öka konsumenternas vilja att hävda sina rättigheter avsevärt och i länder där konsumenterna inte är aktiva på grund av att detta är komplicerat och medför höga kostnader är åtgärder som företrädartalan av avgörande betydelse.
Grupptalan (debatt
Nästa punkt på föredragningslistan är kommissionens uttalande om grupptalan.
ledamot av kommissionen. - (EN) Herr talman! Ända sedan jag tillträdde har jag som ni vet prioriterat möjligheterna till rättslig prövning högt.
Jag anser att de materiella rättigheterna inte visar sin styrka förrän de backas upp av exekutiva åtgärder och faktiska möjligheter för konsumenterna att föra talan.
Allt oftare får stora konsumentgrupper sitta emellan utan att få sin sak prövad till följd av att en handlare tillämpar samma eller liknande olagliga förfaranden.
Kommissionen har granskat de problem som konsumenterna stöter på när de försöker föra grupptalan.
Vi har beställt studier, diskuterat frågan med intressenterna, genomfört undersökningar och haft ett samråd på Internet. Nyligen publicerade vi också en grönbok som vi har fått över 170 reaktioner på.
Trots att samrådet officiellt tog slut den 1 mars 2009 kommer det fortfarande in synpunkter, och jag kan redan berätta att ju mer bevis vi samlar in, desto mer övertygade blir vi om att det finns ett problem.
Därför måste vi hitta en lösning, för att skipa rättvisa och skapa en sund europeisk ekonomi.
I Grönboken om kollektiva prövningsmöjligheter för konsumenter togs olika sätt att komma till rätta med problemet upp.
En preliminär analys av mottagna svar tyder på att intressenterna är medvetna om att situationen i fråga om grupptalan i medlemsstaterna är otillfredsställande.
Det finns en samsyn om behovet av ytterligare åtgärder för att skapa verkningsfulla prövningsmöjligheter för konsumenterna och därmed återställa deras förtroende för marknaden.
Konsumentorganisationerna vill ha bindande åtgärder för nationella system för kollektiv rättslig prövning i alla medlemsstaterna i kombination med andra alternativ, såsom utvidgning av befintliga alternativa tvistlösningsmetoder till att omfatta gruppanspråk.
Företagen förespråkar alternativa tvistlösningsmetoder.
Om några veckor, när vi har analyserat alla svaren ordentligt, kommer vi att offentliggöra dem tillsammans med ett uttalande om den återkoppling vi har fått, och före sommaren kommer vi att skissera olika sätt att ta itu med frågan om gruppanspråk.
Detta blir inte bara en upprepning av de fyra alternativen i grönboken.
Vårt resonemang vidareutvecklas mot bakgrund av svaren på samrådet om grönboken.
Kommissionen kommer att på basis av resultaten av alla samråden göra en noggrann granskning av de ekonomiska och sociala konsekvenserna för intressenterna, däribland kostnader och nytta med olika alternativ.
Den 29 maj kommer vi att ha en utfrågning där vi informerar intressenterna om våra preliminära slutsatser.
Låt mig understryka att vi, oavsett vilken väg vi väljer, inte kommer att följa USA i spåren.
I stället kommer vi att vara våra europeiska rättskulturer trogna och ta hänsyn till gjorda erfarenheter i medlemsstaterna.
När väl alternativen klarnar kommer Europaparlamentet, medlemsstaterna och intressenterna att vara lika övertygade som jag om att vi har ett problem och att en ändamålsenlig lösning måste, och kan, skapas på EU-nivå.
Varför ska hederliga företag lida på grund av ojusta konkurrenter som tjänar pengar när konsumenterna inte gottgörs?
Och jag betonar ”gottgörs”.
Det är just möjligheter till gottgörelse vi eftersträvar.
Varför ska konsumenterna ge upp sina legitima förväntningar på gottgörelse, och varför ska samhället acceptera brister i välfärden och rättvisan?
Jag är säker på att vi kommer att finna en lösning som skapar den rätta balansen mellan att förbättra konsumenternas möjligheter till rättelse och att undvika ogrundade klagomål.
Effektiva prövningsmöjligheter kommer att öka konsumenternas förtroende för den inre marknaden och för vad EU kan göra för dem.
Detta är särskilt viktigt i den bistra verklighet som dagens ekonomiska och finansiella kris har skapat.
Som ni vet kommer det att genomföras många institutionella förändringar under de kommande månaderna, och de kan påverka tidplanen för och presentationen av vårt arbete med grupptalan.
När det gäller kommissionens initiativ om skadeståndstalan vid brott mot EG:s antitrustregler kan jag försäkra er om att kommissionen delar parlamentets inställning att dessa två initiativ som har med grupptalan att göra bör hänga samman.
Konsekvens betyder dock inte att man i olika politiska initiativ måste använda samma verktyg för att nå samma mål.
Jag kan också försäkra er om att jag personligen är engagerad i den här frågan och kommer att fortsätta arbeta med den tills mitt mandat går ut, med samma energi och kraft som hittills, och naturligtvis med välvilligt bistånd och stöd från parlamentet.
för PPE-DE-gruppen. - (EN) Herr talman! Det gläder mig att få välkomna kommissionsledamot Kuneva till kammaren igen.
Jag kan bara upprepa det ni själv sa om hur energiskt och kraftfullt ni försöker tillgodose konsumenternas intressen. Vi på vår sida av kammaren och alla ledamöterna i utskottet, tror jag, beundrar er för det och vill verkligen att ni ska fortsätta så.
När det gäller förslaget om grupptalan tycker jag att ni hanterar det på helt rätt sätt.
Vi har konsekvent sagt att det här är en oerhört komplicerad fråga.
Det handlar inte bara om åtgärder på EU-nivå, utan också om mycket svåra frågor om anknytningen till nationell och regional rätt, och framför allt måste som ni sa konsumenterna stå i centrum.
Ni har verkligen konsekvent hävdat att konsumenternas förtroende för den inre marknaden och gränsöverskridande handel är en av de grundläggande frågor som vi måste ta upp, för annars kan inte konsumenterna utnyttja sin rätt till tillgång och utöva valfrihet över gränserna.
Jag tycker att det är kärnpunkten i det ni sa i dag.
Först och främst anser jag att timingen och lösningarnas komplexitetsgrad är viktiga, för ni har nämnt en lång rad lösningar här, men det står helt klart att lösningar som innebär att nya rättsmekanismer på EU-nivå kan behöva skapas tar mycket längre tid och potentiellt är mer kontroversiella än om man tar till någon av de alternativa tvistlösningsåtgärderna eller använder de befintliga åtgärder för konsumentsamarbete som har införts.
Jag tror att vi alla i utskottet minns att det utökade konsumentsamarbetet var en fråga som utskottet behandlade under parlamentets förra mandatperiod, och vi vill att det blir mer ändamålsenligt.
Jag tror att det kan användas för att ge konsumenterna de prövningsmöjligheter vi efterlyser, inte bara när det gäller grupptalan utan också för att hantera gränsöverskridande anspråk på ett mer verkningsfullt sätt.
Om vi kan göra dessa prioriteringar där och med timing och skyndsamhet snabbt kommer fram till de bästa lösningarna så tycker jag att det är så ni ska gå vidare.
Herr talman, fru kommissionsledamot! Tack för att ni tog fasta på socialdemokratiska gruppens i Europaparlamentet initiativ och tog upp den här frågan, den är viktig för medborgarna.
Jag har min mobiltelefon här.
Jag har hört av många ungdomar att de har en mängd problem till följd av att en summa pengar dras av varje månad i fem, sex, sju eller åtta månader på grund av att de helt ovetande har ingått ett eller annat avtal, till exempel om ringsignaler.
Ingen vänder sig till en domstol för 5 euro, men om en miljon medborgare upplever samma sak och ett företag orättmätigt inkasserar 5 miljoner euro så handlar det om orättvis konkurrens i förhållande till de konkurrenter i Europeiska unionen som uppför sig korrekt.
Därför är det mycket viktigt att vi tar itu med detta.
Det är dock också viktigt att människorna, ungdomarna, föräldrarna som råkar ut för detta får rättsliga instrument som gör att de verkligen får bättre på fötterna.
Vid en tidpunkt då EU växer ihop, när människor handlar på Internet, är det viktigt att vi upprättar dessa som gränsöverskridande instrument så att de faktiskt kan användas ordentligt.
Därför anser min grupp att det just är den grupptalan som sådana instrument möjliggör som måste utredas, så att vi kan se om den kan användas i Europeiska unionen.
Som ni också har sagt, fru kommissionsledamot, måste dock dessa instrument utformas så att vi förhindrar att de ytterligheter som förekommer i till exempel USA smyger sig in, och i stället anpassa instrumenten till vårt eget rättssystem.
Vi måste arbeta på detta, och vi vill driva den här frågan under de närmaste månaderna.
Fru kommissionsledamot! Ni vet att vi står på er sida i den här frågan.
När det gäller att förstärka medborgarnas rättigheter har vi socialdemokrater alltid ett finger med i spelet!
(DE) Herr talman, fru kommissionsledamot! Tack så mycket för att jag fick möjlighet att delta i den här debatten.
Fru Kuneva! Det gläder mig att ni på begäran av gruppen för Europeiska folkpartiet (kristdemokrater) och Europademokrater har bidragit till att utveckla förslaget om grupptalan från GD Konkurrens, som inledningsvis planerade att reglera detta på samma sätt som i USA, till en övergripande metod och faktiskt behandla alla lika i Europeiska unionen - små och medelstora företag, konsumenter, anställda och företagare.
Detta är ett viktigt steg framåt, som vi vill stödja i en mycket konstruktiv och positiv anda.
Vi är medvetna om att gemenskapen i många enskilda fall naturligtvis är bättre på att tillvarata kollektiva rättigheter än individen.
Vi är emellertid övertygade om att grupptalan inte är bästa sättet att skumma av bagatellartade anspråk så att konsumenterna skyddas, utan snarare en offentligrättslig prövning av sådana anspråk, till exempel genom en vinstskumningstalan som i den tyska lagen mot orättvis konkurrens. Enskilda konsumenter skulle då överväga mycket omsorgsfullt om de ska inleda en grupptalan med en advokat om 4,99 euro eller om det faktiskt skulle vara bättre om dessa anspråk till exempel kontinuerligt bevakas av en offentlig ombudsman och genomdrivs med lämpliga medel.
När det gäller hur dessa båda beståndsdelar ska kopplas samman anser jag således att vi noggrant måste överväga hur vi bäst kan hjälpa konsumenterna, för de har ofta inte tid att vända sig till en advokat, utan vill ha hjälp snabbt och lätt.
Det finns en annan sak som jag tycker är viktig - och också här har ert generaldirektorat gjort ett mycket gott arbete. Det mest intressanta inslaget var en diskussion vid den bayerska representationen i Bryssel.
Där svarade en företrädare för ert generaldirektorat på frågan om vi genom att använda EU:s rättsmedel faktiskt kan utesluta den typ av grupptalan som förekommer i USA med att klart säga ”nej, det kan vi inte”.
Det anser vi betyder att vi inte kan bortse helt från denna modell. Vi måste fortsätta att diskutera den, men göra det med stor omsorg och ta med medlemsstaterna och deras lagliga möjligheter i diskussionen så att vi i slutändan uppnår det vi alla vill, det vill säga en verkligt europeisk modell som är särskilt tilltalande för konsumenterna och som också skyddar små och medelstora företag.
(EN) Herr talman! Jag vet att kommissionsledamoten känner till att 4 000 konsumenter kommer att hänvända sig till högsta domstolen i Förenade kungariket i morgon för att söka gottgörelse för allvarliga allergiska reaktioner, sjukhusvistelser och dödsfall till följd av användningen av kemikalier som nu har förbjudits i EU i soffor och hushållsprodukter.
Liknande fall och skador har rapporterats från Frankrike, Sverige och Polen.
I hela EU finns det potentiellt många tusen konsumenter som har lidit allvarliga skador på grund av denna giftiga kemikalie.
Jag tror att medborgarna vill att EU ska ingripa när vi kan ge konsumenterna verklig hjälp med att komma till rätta med verkliga problem.
Verklig hjälp i sådana fall betyder rätt att vidta kollektiva åtgärder, oavsett var man köper varor och tjänster.
Därför lanserade vårt utskott ett samråd på Internet om kommissionens förslag om konsumenträttigheter.
Vi fick många svar och i många av dem framhöll företag och konsumenter att det behövs effektiv tillgång till gränsöverskridande rättsmedel och prövningsmöjligheter.
Jag anser att det finns tillräckligt många fall som liknar fallet med den giftiga soffan och tillräckligt med övertygande bevis för att det behövs möjligheter till grupptalan, inte bara för att förbättra tillgången till rättvisan utan också för att motverka olagliga och orättvisa affärsmetoder.
I vårt utskott vill vi naturligtvis att konsumenterna ska ha tillgång till billiga, överkomliga metoder, såsom alternativa tvistlösningsmetoder, men jag anser att dagens debatt först och främst handlar om att hitta praktiska sätt att ge våra konsumenter och medborgare verklig hjälp, att se till att de får rättvisa lösningar, verkliga prövningsmöjligheter och verkliga rättsmedel.
(DE) Herr talman, mina damer och herrar! Jag vill börja med att säga att också vi i princip välkomnar Europeiska kommissionens förslag och denna grönbok.
Som andra talare har sagt råder det inga tvivel om att det finns ett ”massfenomen” där ett stort antal människor drabbas av relativt små förluster.
De enskilda förlusterna är små, men det sammantagna beloppet är stort.
Vi behöver ett instrument som löser detta problem.
Jag anser att det är rätt att överväga någonting i den här stilen.
För att fortsätta på den positiva sidan välkomnar jag också verkligen att Generaldirektoratet för hälsa och konsumentskydd i sin grönbok betonar frågan om alternativa tvistlösningsmetoder så kraftigt.
Det är en stor skillnad jämfört med vitboken från Generaldirektoratet för konkurrens, som också debatterades i kammaren i går, och i vilken man hittills inte alls tar upp möjligheten till tvistlösning utanför domstol.
Jag anser att Generaldirektoratet för hälsa och konsumentskydd har kommit längre i sin grönbok än kollegerna i Generaldirektoratet för konkurrens.
Jag vill dock slå fast två saker som jag definitivt anser ska betraktas som kritiska kommentarer.
Klockan 12, om några få minuter, kommer parlamentet att anta mitt betänkande om vitboken från Generaldirektoratet för konkurrens.
Med överväldigande majoritet kommer kammaren att kräva att Europeiska kommissionen hanterar den här frågan med en övergripande strategi.
Det får inte bli så att vi får sektorsvisa instrument - ett för konsumentskydd, ett för antitrustlagstiftning, ett annat för kapitalmarknaden, kanske ytterligare ett för miljön, kanske ytterligare ett för sociala frågor - som alla är motstridiga, som alla inkräktar på medlemsstaternas rättssystem och i slutändan leder till en förvirring om rättsläget som ingen jurist längre kan reda ut.
Vi har ofta sett sådana exempel tidigare.
Jag tänker bara på debatten om direktivet om yrkeskvalifikationer, som vi senare också lade ihop till ett enda instrument eftersom denna fragmentarisering inte längre var hanterbar.
Kommissionen bör inte göra samma misstag igen i det här fallet.
Den bör förespråka en övergripande strategi redan från början.
Det är parlamentets tydliga ståndpunkt, vilket kommer att visa sig om några minuter.
En sak till: Jag välkomnar verkligen att vi har kommit överens om att vi inte vill ha en klagomålsindustri efter amerikansk modell med en omsättning på 240 miljarder US-dollar om året, som egentligen bara advokaterna tjänar på medan konsumenterna inte får någonting alls.
Vi vill ha äkta rättssäkerhet i EU och vi vill behålla vårt traditionella system och vårt sätt att betrakta lagen.
(ES) Herr talman! På en marknad utan gränser som EU är det viktigt att vi både garanterar en sund konkurrens och lika nitiskt värnar om konsumenterna.
Under det gångna halvseklet har handelshinder raserats för produkter, men de finns i stor utsträckning kvar för konsumenterna.
Otillåtna affärsmetoder anmäls ofta inte av konsumenterna eller beivras av konsumentorganisationerna på grund av en allmän medvetenhet om att det är svårt att få gottgörelse.
Grupptalan är ett förfarande som underlättar när många människor har drabbats och gör att chanserna att komma fram till en överenskommelse om kompensation ökar betydligt.
Eftersom en stor del av de ekonomiska transaktionerna i Europeiska unionen är gränsöverskridande kan inte denna rätt till kollektiva åtgärder sluta vid landsgränserna.
Vi behöver ett verkligt initiativ som omfattar hela EU och det måste skapa en viss harmonisering eller anpassning av befintliga nationella system för att bli ändamålsenligt.
Den modell vi väljer måste syfta till att ge konsumenterna tillgång till systemet utan svårigheter och att motverka höga kostnader och omfattande byråkrati.
Därför anser jag att vi måste prioritera alternativa konfliktlösningsförfaranden, eftersom de skapar större flexibilitet, samt förenklade och billigare rättsprocesser.
(DE) Herr talman! Det finns en stor samsyn i kammaren om att vi måste erbjuda konsumenterna ett bättre skydd, i synnerhet när små förluster för många enskilda personer sammantagna utgör ett problem, eftersom man inte ser några möjligheter att föra individuell talan på ett meningsfullt sätt.
Frågan är hur konsumentskyddet och förbättringen av detta ska organiseras.
Där anser jag att det är mycket viktigt att vi helt medvetet säger att vi vill utreda alla alternativ och alla aspekter av denna komplicerade fråga och inte fatta beslut om lösningar förrän efter moget övervägande - och det är jag mycket tacksam mot kommissionen för att vi gör.
Jag vill i det här sammanhanget ta upp en sak som ännu inte har nämnts.
Vi har redan konstaterat att möjligheterna att föra grupptalan håller på att bli ett sätt för många icke-statliga organisationer och konsumentskyddsorganisationer att marknadsföra sig, och så kan det bli än mer i framtiden.
Denna risk bör vi mycket medvetet ta med i våra beräkningar så att det inte slutar med att vi hjälper dem som inte behöver någon hjälp medan de som faktiskt behöver hjälp blir utan.
kommissionsledamot. - Herr talman! Jag skulle vilja tacka er för alla era värdefulla synpunkter.
På ett sätt känner jag väl till de flesta av dem eftersom vi har diskuterat igenom de viktigaste aspekterna av era betänkligheter och förhoppningar vad gäller att införa grupptalan i Europa, punkt för punkt.
Jag skulle återigen vilja understryka att jag håller helt med er om att det inte ska införas någon USA-liknande grupptalan i den europeiska kulturen.
Jag vet att detta är något av det som oroar er mest.
Som Arlene McCarthy också påpekade handlar det här om skadestånd.
Detta förekommer redan i Storbritannien, men det har ingenting att göra med vad vi diskuterar här och vad jag föreslår som våra framtida åtgärder i den här riktningen.
I det hänseendet skulle jag vilja understryka följande: Kontrollerar vi om det finns ett verkligt behov av grupptalan?
Ja, det gör vi och vi kommer också att fortsätta att göra detta efter grönboken.
Respekterar vi de konstitutionella begränsningarna? Ja.
Undviker vi en USA-liknande grupptalan? Ja.
Ser vi till att det utgår ersättning för skadestånden som omfattar konsumentens samtliga kostnader, men samtidigt utesluter något inslag av straffskadestånd? Ja, det tänker vi göra.
Motverkar vi oberättigade anspråk, som Reinhard Rack tog upp? Ja.
Främjar vi alternativa tvistlösningsmetoder? Självklart, eftersom detta kostar mindre tid och pengar och är lättare att hantera för både konsumenter och företag och även följer subsidiaritetsprincipen.
Med dessa få ord skulle jag vilja säga att vi är fullt medvetna om utmaningarna och att vi är redo att ta oss an dem och steg för steg lägga fram ett bra förslag genom att uppnå samförstånd med er.
Vad jag verkligen uppskattar här i dag är att vi alla inser att vi har ett problem och att vi är redo att ta itu med det problemet.
Det är verkligen en mycket bra utgångspunkt för nästa diskussionsfas.
Eftersom det är en utmaning som vi står inför skulle jag framför allt vilja understryka det som Klaus-Heiner Lehne tog upp - den gemensamma strategin, den övergripande strategin med kommissionsledamot Kroes.
Kommissionsledamot Kroes och jag och våra båda enheter samarbetar mycket nära för att våra initiativ ska vara enhetliga och ge synergieffekter.
Principen om enhetlighet utesluter inte nödvändigtvis att särskilda situationer kräver särskilda lösningar.
Vart och ett av de båda initiativen har en specifik inriktning.
I grönboken för konsumenter behandlas talan som rör överträdelser av konsumentskyddslagstiftningen, medan vitboken om konkurrens uteslutande handlar om överträdelser av konkurrenslagstiftningen.
En annan betydande skillnad mellan de båda initiativen är att grönboken för konsumenter endast avser konsumenters möjlighet till prövning, medan den prövningsmekanism som föreslås i vitboken om konkurrens är tänkt att gynna både konsumenter och företag.
Så min utmaning är att uppnå en effektiv prövningsmöjlighet för våra konsumenter och därigenom ge dem förnyat förtroende för marknaden.
Från tidigare diskussioner vet jag att Europaparlamentet stöder oss i våra försök att uppnå detta mål.
Låt mig återigen understryka att parlamentet tillsammans med medlemsstaterna och aktörerna kommer att bli övertygade inte bara om att vi har ett problem, utan också om att det är nödvändigt och möjligt att nå fram till en effektiv och välavvägd lösning på EU-nivå.
Jag skulle vilja tacka er för denna givande diskussion och era värdefulla synpunkter och jag ser fram emot att samarbeta med er kring det här ärendet under de kommande månaderna.
Debatten är avslutad.
Skriftliga förklaringar (artikel 142)
Jag skulle vilja framföra mina lyckönskningar när det gäller Europeiska kommissionens insatser för att förbättra konsumenternas möjligheter att tillvarata sina rättigheter i hela EU.
De alternativ som presenteras i grönboken måste diskuteras ingående.
Men en sak som redan är säker är att alternativ nr 4 - som innebär att det skulle införas en kategori av opt out-åtgärder som ger konsumentorganisationerna en andel av gottgörelsebetalningarna - inte är möjligt (genomförbart).
Om vi vill öka konsumenternas förtroende för den inre marknaden måste vi överväga en kombination av alternativ 2 och 3.
Vi måste med andra ord skapa ett europeiskt nätverk av nationella verkställande offentliga myndigheter som får utökade befogenheter att vidta effektiva åtgärder i samband med internationella anspråk (utomlands).
Vidare måste vi se över alternativa mekanismer för att lösa befintliga tvister samt vid behov införa en ny mekanism som gör att konsumenternas rättigheter kan tillämpas (utövas) mer efffektivt även utanför domstolarna.
Jag skulle vilja avsluta genom att understryka att vi måste se till att tillämpa ett övergripande synsätt när det gäller mekanismen för grupptalan, så att vi undviker en fragmentering av den nationella lagstiftningen och upprättar ett enda, gemensamt instrument för samtliga medlemsstater.
(Sammanträdet avbröts kl. 11.35 och återupptogs kl. 12.05.)
Justering av protokollet från föregående sammanträde: se protokollet
15.
Förslag till ändringsbudget 2/2009 (
Valprövning: se protokollet
8.
Skyddstiden för upphovsrätt och vissa närstående rättigheter (
- Före omröstningen:
(EN) Herr talman! Jag beklagar att jag måste besvära kollegerna under ett långt omröstningspass, men det har ånyo angetts i omröstningslistan att ändringsförslag 80 till ett skäl faller om ändringsförslag 37 går igenom.
Den första hälften av ändringsförslaget är exakt densamma, men den nya biten - den andra delen - är följdriktig.
Det har inte angetts att ändringsförslag 81, som är motsvarande ändringsförslag för artikeln, faller om motsvarande ändring av artikel 55 antas.
Därför yrkar jag på att vi röstar om ändringsförslag 80 som ett tillägg till ändringsförslag 37 om ledamöterna tillstyrker det - vilket är en annan sak - eftersom det tydligen är vad vi kommer att göra med ändringsförslag 81.
Tack, fru Bowles.
Nu vore det bra att få höra vad föredragande Crowley anser.
föredragande. - (EN) Herr talman! Jag tycker inte att det kan tas som ett tillägg.
Det bör behandlas separat.
Rättelser/avsiktsförklaringar till avgivna röster: se protokollet
Frågestund (frågor till rådet)
Nästa punkt på föredragningslistan är frågestunden med frågor till rådet (B6-0227/09).
Vi ska nu behandla en rad frågor till rådet.
Angående: Antilissabonretoriken
Den globala finanskrisen har visat hur viktigt det är med ett starkt EU.
Vi i Irland har snabbt lärt oss att myter och vilseledande information om Lissabonfördraget är en klen tröst i en krympande ekonomi och ökande arbetslöshet.
När nu Tjeckien är ordförandeland, och landets egen president anslutit sig till antilissabonretoriken, hur tänker då rådet hantera dessa signaler när det står helt klart att behovet av samarbete inom EU är större, inte mindre?
rådets tjänstgörande ordförande. - (CS) Fru talman, mina damer och herrar! Rådet har alltid klargjort sitt fasta beslut att stärka samarbetet inom EU, i synnerhet i krissituationer.
Under det tjeckiska ordförandeskapet, som bygger vidare på föregångarnas arbete, arbetar vi hårt på att lösa de problem som orsakas av den rådande finansiella och ekonomiska krisen och har i detta sammanhang beslutat om åtgärder på olika nivåer. En gemensam ram för medlemsstaterna har etablerats, såsom kan ses exempelvis från bankräddningsplanen, den ekonomiska återhämtningsplanen för Europa och reglering och tillsyn av finansmarknaderna.
Europaparlamentet har också bidragit till åtgärderna genom att stötta investeringar i infrastrukturen, inte minst genom sina internationella insatser. Vid mötet den 19 och 20 mars var rådet helt inriktat på att övervinna finanskrisen och problemen med realekonomin och klargjorde mycket tydligt att EU kan bemästra problemen och stoppa den rådande krisen endast genom en enad och samordnad handling inom ramen för den inre marknaden och EMU.
Vid mötet den 19 mars beslutade rådet att en nära samordnad EU-respons inom ramen för den ekonomiska återhämtningsplanen för Europa ska innehålla mobilisering av alla tillgängliga instrument, inklusive gemenskapsmedel och att fullständigt integrerade strategier för tillväxt, sysselsättning, social integration och socialförsäkring ska ingå.
Beträffande Lissabonfördraget uppnådde rådet en överenskommelse om ytterligare framsteg, i december 2008.
På Irlands begäran har medlemsstaterna gått med på att åstadkomma specifika lagliga garantier gällande de problem som var en källa till oro under förra årets folkomröstning i Irland.
Rådet har också gått med på att om Lissabonfördraget träder i kraft, kommer man att efter grundläggande rättslig prövning anta ett beslut om de respektive medlemsstaternas fortsatta nationella representation i kommissionen.
Med undantaget att specificerad, relaterad verksamhet i frågan ska slutföras under mitten av 2009 och förutsatt att genomförandet blir tillfredsställande är den irländska regeringen samtidigt fast besluten att arbeta för en ratificering av Lissabonfördraget mot slutet av kommissionens innevarande mandatperiod.
Under mötet den 19 och 20 mars informerades Europeiska rådet om den rådande situationen i frågan och man beslöt att ta upp frågan på nytt under mötet i juni 2009.
(EN) Fru talman! Jag vill tacka ministern för hans svar.
Jag tycker att vi är alltför defensiva här i kammaren - och i institutionerna i allmänhet - när det gäller Lissabon och EU i allmänhet.
Det är dags att vi sätter dem som attackerar Europa på defensiven.
Var skulle vi vara utan Europeiska centralbanken?
Var skulle vi vara - de av oss som tillhör euroområdet - utan euroområdet?
Det enda vi saknar är en igenkännbar ledare för Europeiska rådet som kan tala om frågor som rör den ekonomiska återhämtningen, och jag tycker att det är uppenbart att den bestämmelse i Lissabonfördraget som möjliggör att en sådan person utses verkligen är avgörande.
Om vi hade haft en sådan person nu hade vi sluppit sicksackandet mellan de sex månader långa ordförandeskapen.
Kanske ministern i sitt svar skulle kunna uttala sig om sin syn på utsikterna för en ratificering av fördraget i Tjeckien.
rådets tjänstgörande ordförande. - (CS) Jag kommer att besvara alla frågor senare, i en följd.
Enligt vår normala arbetsordning ska ni först svara frågeställaren och dennes följdfråga och sedan, vanligtvis, kommer jag - och så har jag valt att göra - att samla ihop de andra följdfrågorna och ställa de till er.
Får jag be er att svara först.
rådets tjänstgörande ordförande. - (CS) Tack, fru talman!
Mina damer och herrar! Jag ska nu besvara frågan.
Vad beträffar ratificeringen av Lissabonfördraget vill jag framhålla att Republiken Tjeckiens tvåkammarparlament, som utgörs av representanthuset och senaten, arbetar mycket hårt på fördraget och att det godkändes av representanthuset den 18 februari i år.
Här måste jag betona att det enligt tjeckiska grundlagar krävs en konstitutionell majoritet för att fördraget ska gå igenom.
Det tjeckiska parlamentets senat kommer förmodligen att rösta om fördraget den 6 maj, men senaten har som villkor för godkännandet krävt ett utkast till en lämplig lag enligt vilken överföring av behörighet kräver omröstning med kvalificerad majoritet och godkännande från parlamentets båda kamrar.
Detta innebär ett så kallat villkorat mandat.
Den tillämpliga lagen har redan utarbetats och godkänts och vi förväntar oss att senaten kommer att rösta om lagen den 6 maj och att Lissabonfördraget kommer att ratificeras av parlamentet så snart som lagen har antagits.
(EN) Håller inte det tjeckiska ordförandeskapet med om att problemet när det gäller Lissabonfördraget i första hand inte handlar om bristen på information om det, eftersom det finns gott om information tillgänglig, utan om den betydande mängd felaktig information som avsiktligt sprids av fördragets motståndare?
Håller det inte också med om att de nationella regeringarna måste göra mycket mer för att motverka de myter och den felaktiga information som Gay Mitchell talade om och få ordning på denna mycket viktiga debatt om Europas framtid, med tanke på att fördraget inte skrivs under av de europeiska institutionerna utan förhandlades fram av medlemsstaterna?
(EN) Herr minister! Jag är säker på att i ert land, liksom i Irland, uppfattar väljarna för närvarande och oroar sig för ett orwellskt EU.
De är inte dumma, och de vet att kommissionen manipulerade sitt lagstiftningsprogram så att inga dåliga nyheter nådde de irländska medierna.
Det är synd att Gay Mitchell, Richard Corbett och de andra är så förblindade av lockelsen i att bli framgångsrika eurokrater att de inte förstår vad frågan handlar om: att det irländska folket har meddelat sitt beslut.
Kanske ni kan få rådet att ge kommissionen i uppdrag att stoppa den stora ökningen av sina avdelningar för kommunikation och information - det vill säga propaganda - och låta det resultat som det fantastiska irländska folket har meddelat visa att demokratin lever i EU.
rådets tjänstgörande ordförande. - (CS) Jag vill betona att vi alla bör ha kurage nog att medge för oss själva att EU-medborgarna har mycket dålig kännedom om hur EU fungerar.
EU påverkar oftast medborgarna på ett abstrakt sätt och EU:s institutioner är mycket svåra att förstå.
Enligt min mening skulle felaktig information och lögner inte kunna få fäste om vi tog itu med bristen på demokrati och det faktum att medborgarna inte alltid identifierar sig med EU och dess institutioner.
Jag är av den bestämda uppfattningen att regeringarna i EU:s medlemsstater har en grundläggande skyldighet att motarbeta felaktig information och osanningar.
Det är min absoluta mening att vi endast då kan uppnå verkliga demokratiska framsteg.
Angående: Dubbelbeskattning
I ljuset av den senaste rättspraxisen från EG-domstolen vad avser dubbelbeskattning, vilka åtgärder avser rådet vidta för att harmonisera EU:s skatterätt så att europeiska skattebetalare inte behöver betala skatt två gånger för samma sak?
rådets tjänstgörande ordförande. - (CS) Fru talman, mina damer och herrar! Vad beträffar det rådande tillståndet inom gemenskapen har man på gemenskapsnivå ännu inte godkänt några åtgärder för att ta bort dubbelbeskattningen inom området direktbeskattning, med undantag av rådets direktiv 90/435/EEG av den 23 juli 1990 om gemensamma beskattningssystem för moderbolag och dotterbolag hemmahörande i olika medlemsstater, konventionen från den 23 juli 1990 om undanröjande av dubbelbeskattning vid justering av inkomst mellan företag i intressegemenskap och rådets direktiv 2003/48/EG av den 3 juni 2003 om beskattning av inkomster från sparande i form av räntebetalningar.
Det beror på att området i fråga är medlemsstaternas ansvar, förutsatt att de tillämpar gemenskapslagstiftningen.
Överenskommelser om att undanröja dubbelbeskattning som enligt de tidigare nämnda autonoma befogenheterna och i enlighet med provöverenskommelsen med OECD, ingås bilateralt mellan medlemsstaterna, tycks inte räcka till för att undanröja all juridisk dubbelbeskattning inom EU.
Kommissionen, som har den exklusiva rätten att initiera lagar inom gemenskapen i samband med direktbeskattning, föredrar för närvarande helt klart en pragmatisk strategi i den här frågan, med tanke på subsidiaritetsprincipen, som tillämpas på gemenskapslagstiftningen inom området direktbeskattning och med tanke på kravet på enhällighet.
Denna pragmatiska strategi borde uppmuntra medlemsstaterna att samarbeta för att se till att de inhemska beskattningssystemen, inklusive de bilaterala beskattningsavtalen, fungerar smidigt.
Detta omnämns, bland mycket annat, i kommissionens meddelande om samordning av medlemsstaternas direktbeskattningssystem inom den inre marknaden, särskilt i den slutliga versionen av dokumentet.
Rådet har bekräftat kommissionens samarbetsbaserade strategi i slutsatserna från den 27 mars 2007.
Det betonades att den inre marknadens funktion inom beskattningsområdet kan förbättras genom samarbete på medlemsstatsnivå och, där så är tillämpligt, på EU-nivå med beaktande av medlemsstaternas behörighet.
Rådet förklarade att godtagbara lösningar kan ha olika utformningar, i enlighet med subsidiaritetsprincipen.
(ES) Herr talman! Den information som ni ger oss är korrekt men vi som parlamentsledamöter, och definitivt EU-medborgarna, har ett intryck av att det finns en mycket farlig lucka i gemenskapsrätten.
Eftersom skattekraven hela tiden ökas i samtliga medlemsstater är rörlighet för närvarande i det närmaste omöjligt.
När vi ber kommissionen förklara den pragmatiska strategin verkar det som om kommissionen inte har något stöd i rådet.
Vi tycks ha hamnat i en ond cirkel där kommissionen hänvisar oss till rådet och rådet hänvisar oss tillbaka till kommissionen, samtidigt som verkligheten är den att medborgarna i det EU som vi försöker bygga upp inte kan välja att bosätta sig eller ha kontakter i olika länder, på grund av den tunga skattebörda som orsakas av skattesystemets brist på harmonisering.
Kan rådet göra något för att få slut på den här onda cirkeln?
rådets tjänstgörande ordförande. - (CS) Först och främst vill jag betona att det långsiktiga målet är en lösning i form av ett direktiv eller multilateralt fördrag.
Bara på det sättet kan vi utveckla systemet effektivt med utgångspunkt från rättsprinciper.
Kommissionen ska föreslå en lösning på de mest överhängande problem som uppkommer i samband med den inre marknaden, genom ökad samordning av medlemsstaternas skattelagstiftning och bättre beslutsprocesser.
Kommissionen föreslår i sitt meddelande om samordning av medlemsstaternas direktbeskattningssystem inom den inre marknaden att inrätta en mekanism för en effektiv lösning av tvister i samband med problem med internationell dubbelbeskattning inom EU, men på grund av otillräckligt stöd från medlemsstaterna, som Paul Rübig nämnde, har kommissionen övergett frågan till förmån för andra initiativ.
Kommissionen är fullt medveten om hur dubbelbeskattningsavtal påverkar den inre marknaden och kommer att förbereda offentliga samråd under 2009. Med utgångspunkt från samråden ska kommissionen utarbeta ett meddelande om vad man kommit fram till samt ett förslag på en godtagbar lösning på de existerande problemen.
Rådet har gång på gång brottats med det här problemet inom ramen för olika initiativ.
Första gången gällde det expansion av ramarna för direktiv 90/435/EEG om ett gemensamt beskattningssystem för moderbolag och dotterbolag, genom rådets direktiv 2003/123/EG, som undanröjer den ekonomiska och juridiska dubbelbeskattningen av gränsöverskridande flöden av utdelningar inom ramen för gemenskapen.
1990 antogs ett skiljedomsfördrag med syftet att undanröja den dubbelbeskattning som uppkommer genom att man fastställt internpriser mellan närstående företag.
Det visade sig emellertid att direktivet inte var så effektivt, delvis eftersom det har karaktären av internationellt avtal som ingåtts mellan medlemsstater och inte karaktären av en gemenskapsrättsakt.
År 2003 antogs direktiv 2003/49/EG, vilket undanröjde dubbelbeskattning av räntor och royalties som betalas mellan närstående bolag i olika medlemsstater och som innebär att endast det land där förmånstagaren för utbetalningen är bosatt, har rätt att beskatta betalningen.
Frågan om att expandera ramarna för detta direktiv bör bli föremål för fortsatta förhandlingar i rådet.
I samband med kommissionens båda meddelanden om samordning av medlemsstaternas direktbeskattningssystem och sociala avgifter inom den inre marknaden, har Ekofin antagit rådets resolution från december 2008 om sociala avgifter. Resolutionen syftar till att undanröja dubbelbeskattning och samordna statliga förfaranden inom området för sociala avgifter på så sätt att, vid överföring av ekonomisk verksamhet från en stat till en annan, när fysiska eller juridiska personers tillgångar överförs från en stat som tillämpar beskattning vid utflyttning, ska den mottagande staten tillämpa den utväxlade tillgångens marknadsvärde vid tidpunkten för överföringen från utflyttningsstaten som en kostnad när tillgången säljs.
(EN) Vi förstår alla att dessa skattefrågor kan vara mycket tekniska, men kan ministern ändå rent allmänt hålla med om att alla som förstår dessa frågor säkerligen inser att en skatteharmonisering inte är avgörande för att dubbelbeskattning ska kunna undvikas?
Allt som krävs - jag vet att det är rätt tekniskt - är en vilja till bättre samarbete mellan medlemsstaterna.
Med tanke på de stora belopp som regeringarna i nuläget tar från hårt pressade skattebetalare är det väl säkerligen dags att uppmuntra mer skattekonkurrens för att minska bördan för arbetande familjer i hela EU.
(DE) Herr ordförande! Jag anser att det tjeckiska ordförandeskapet har en mycket positiv och proaktiv inställning i denna fråga.
Det gratulerar jag er till, för det är naturligtvis viktigt att skydda medborgare och små och medelstora företag så att också de kan få in sina inkomster när de tillhandahåller tjänster.
Det finns överhuvudtaget inget som gör dubbelbeskattning socialt berättigat.
Därav min fråga: anser ni att EG-domstolen kan fastställa krav på detta område?
rådets tjänstgörande ordförande. - (CS) Fru talman, mina damer och herrar! EG-domstolen har slagit fast att det faktum att gemenskapens lagstiftning, den fria rörligheten och principerna om icke-diskriminering är direkt tillämpliga inte innebär att medlemsstaterna måste avskaffa laglig dubbelbeskattning som beror på en ömsesidig påverkan mellan olika skattesystem i gränsöverskridande situationer i gemenskapen.
Denna ståndpunkt grundar sig på EG-domstolens dom i mål C-513/04, Kerckhaert Morres.
Domstolen har redan avgjort denna fråga och här tror jag faktiskt att möjligheterna är mycket begränsade.
Enligt EG-domstolens rättspraxis måste fördrag om avskaffande av dubbelbeskattning uppfylla den inre marknadens krav och de får i synnerhet inte leda till diskriminering eller skillnader när det gäller de grundläggande rättigheter som slås fast i fördraget om upprättandet av Europeiska gemenskaperna.
Å andra sidan anser jag att risken för dubbelbeskattning gör att skattesystemen blir enormt komplicerade och inte minst gör saker och ting komplicerade för små och medelstora företag, som ibland har mycket svårt att förstå de komplicerade system som lyder under enskilda länders lagstiftning.
Denna risk är störst just för små och medelstora företag, som får högre kostnader på grund av att de inte har råd att anlita dyra konsult- och advokatbyråer på samma sätt som stora företag - inte minst multinationella företag. De komplicerade skattesystemen är därför en större börda för små och medelstora företag.
Jag är personligen övertygad om att det mest rättvisa vore att alla medlemsstater hade enklast tänkbara och mest insynsvänliga system för direktbeskattning och, enligt min personliga uppfattning, så låga skatter som möjligt.
Angående: Fjäderfäkött
Kommissionen har lagt fram ett förslag till rådets förordning om ändring av förordning (EG) nr 1234/2007 om upprättande av en gemensam organisation av jordbruksmarknaderna, vad gäller handelsnormerna för fjäderfäkött.
Håller det tjeckiska ordförandeskapet, mot bakgrund av detta förslag och med hänsyn till konsumenternas hälsa, livsmedelssäkerheten, spårbarheten och produktkvaliteten, med om att märkningen ”färskt” i fråga om fjäderfäkött måste vara en garanti för att köttet just är färskt?
Instämmer ordförandeskapet i att fjäderfäkött som slaktas och fryses in i ett tredjeland och som sedan transporteras och tinas upp, och ibland även bearbetas, i en av EU:s medlemsstater och som sedan marknadsförs och säljs som ”färskt” kött producerat i EU utgör ett allvarligt problem?
Håller ordförandeskapet med om att detta inte är acceptabelt, att det missleder konsumenterna och att det är orättvist mot producenter inom gemenskapen som tillämpar EU:s stränga riktlinjer?
Vilka åtgärder vidtar det tjeckiska ordförandeskapet i dagsläget för att se till att förordningen införs på ett smidigt sätt?
rådets tjänstgörande ordförande. - (CS) Fru talman, mina damer och herrar! Ordförandeskapet kan försäkra ledamoten om att vi fäster stor vikt vid att det ska finnas en stark livsmedelssäkerhet och ett starkt konsumentskydd i gemenskapen, oavsett om livsmedlen produceras lokalt eller importeras från tredjeländer.
I detta sammanhang kan ordförandeskapet hänvisa till slutsatserna från rådets möte den 18-19 december 2008 om säkerheten hos jordbruksprodukter och livsmedelsprodukter som importerats till gemenskapen.
I sina slutsatser uppmanade rådet i enlighet med gemenskapens regler kommissionen att före utgången av 2010 lägga fram en rapport till rådet och Europaparlamentet om effektiviteten hos och tillämpningen av sanitära och fytosanitära kontroller av importerade livsmedel.
Till följd av sin skyldighet att säkra ett starkt skydd för människors hälsa i genomförandet av gemenskapens politik förkastade rådet i december 2008 kommissionens förslag till rådets förordning om genomförande av rådets förordning (EG) nr 853/2004 vad gäller användning av antimikrobiella ämnen för att avlägsna ytkontaminering från slaktkroppar av fjäderfä.
Rådet ansåg att det skulle vara möjligt att dölja dålig sanitär praxis genom att använda sådana ämnen.
Europaparlamentet motsatte sig förslaget i en resolution av den 19 juni 2008 och bad rådet att förkasta det.
När det gäller kommissionens förslag om handelsnormer för fjäderfäkött kan ordförandeskapet bekräfta att förslaget för närvarande är föremål för förhandlingar inom rådet och att målet är att säkra ett starkt konsumentskydd och förhindra att fjäderfäkött som har varit djupfryst säljs som färskt.
Ordförandeskapet kan försäkra ledamoten om att man gör allt för att denna förordning snabbt ska kunna antas så snart Europaparlamentet har avgett sitt yttrande.
(EN) Jag vill tacka ordförandeskapet för detta svar eftersom det tjeckiska ordförandeskapet, om jag har förstått saken rätt, kommer att vidta åtgärder i denna fråga.
Det gläder mig att höra att rådet diskuterar att vidta åtgärder för att förhindra att fjäderfäkött fryses och därefter säljs som om det vore färskt, eftersom detta naturligtvis innebär att många EU-producenter inte bedriver sin verksamhet på lika villkor - i själva verket gör ingen det.
Därför är min fråga till ordförandeskapet: När kan vi förvänta oss något svar från rådet om detta, och kan ni säga någonting om vilka särskilda åtgärder ni skulle kunna vidta i denna fråga?
rådets tjänstgörande ordförande. - (CS) Fru talman, mina damer och herrar! Detta problem har nu lösts av rådets arbetsgrupper i samband med förhandlingarna om förslaget till rådets förordning om ändring av förordning (EG) nr 1234/2007 om upprättande av en gemensam organisation av jordbruksmarknaderna, vad gäller handelsnormerna för fjäderfäkött.
Det tjeckiska ordförandeskapet har föreslagit en kompromisstext som har fått stöd av en majoritet i rådets jordbrukskommitté.
Texten kommer att läggas fram för bedömning av WTO i samband med samråden med handelspartner.
Om resultatet blir positivt och Europaparlamentet godkänner sitt betänkande vid plenarsammanträdet, vilket verkar bli fallet, kommer det tjeckiska ordförandeskapet att överlämna kompromisstexten till rådet.
Rådet har en formell skyldighet att invänta Europaparlamentets yttrande, även om man inte behöver hänvisa till det i sitt beslut.
I kompromisstexten sägs att när det gäller produkter som framställs av färskt fjäderfäkött i enlighet med denna förordning får medlemsstaterna föreskriva vissa variationer i temperaturkraven, vilka får tillämpas under en minimal tidsperiod och bara i den mån det är nödvändigt för att möjliggöra hantering och styckning i bearbetningsanläggningar i samband med produktionen av produkter av färskt fjäderfäkött.
Vi förväntar oss att rådet kommer att ta upp detta förslag i maj och tror mot bakgrund av de förhandlingar som hittills har förts att resultatet kommer att bli positivt.
(EN) Efter BSE-krisen i nötköttssektorn för några år sedan införde vi fullständig identifiering och spårbarhet för nötköttsprodukter i Europa.
Håller inte rådet med om att vi måste agera snabbt, inte bara när det gäller fjäderfäkött utan även fårkött och griskött, för att ge konsumenterna samma information och tillhandahålla samma spårbarhet om något skulle gå fel?
Renate Sommers betänkande om information till konsumenterna behandlas i parlamentet för närvarande, och kanske kan rådet hålla med om att man skulle kunna uppnå detta med hjälp av utökad märkning - vilket skulle öka spårbarheten.
rådets tjänstgörande ordförande. - (CS) Fru talman, mina damer och herrar! I december förra året enades Europeiska rådet om en europeisk plan för ekonomisk återhämtning.
Planen omfattar konkreta åtgärder för att stödja små och medelstora företag, varav de viktigaste är åtgärderna för att förbättra tillgången till finansiering och minska den administrativa bördan för företag.
Europeiska rådet uttryckte samtidigt sitt stöd för ökade insatser av Europeiska investeringsbanken under perioden 2008-2011, i synnerhet i form av lån till små och medelstora företag, som skulle öka med 10 miljarder euro jämfört med den nuvarande utlåningen till denna sektor.
Europeiska rådet har vidare gett sitt stöd till att tröskelvärdena för statligt stöd tillfälligt får överskridas under minst två år när det gäller belopp på högst 500 000 euro, och till att regelverket för statligt stöd anpassas för att stimulera stöd till företag och framför allt till små och medelstora företag.
Europeiska rådet krävde också att de påskyndade förfaranden som är tillåtna enligt gemenskapsrätten skulle tillämpas i samband med offentlig upphandling och att de administrativa bördorna för företag ska minska.
Europeiska rådet stöder också ett fullständigt genomförande av kommissionens handlingsplan för småföretagsakten, som antogs av rådet den 1 december 2008.
Handlingsplanen för småföretagsakten bör hjälpa små och medelstora företag under den ekonomiska turbulensen genom att förbättra deras möjligheter att få lån, minska de administrativa bördorna, hjälpa dem att dra nytta av den inre marknadens fördelar och öka deras konkurrensförmåga på utländska marknader.
Den 5 mars slog rådet fast att handlingsplanen bör genomföras fullt ut så snart som möjligt på EU-nivå och i medlemsstaterna i enlighet med subsidiaritetsprincipen.
Rådet tog dessutom än en gång upp vikten av att förbättra möjligheterna att skaffa finansiering ännu mer - jag tänker här på lån, garantier, mezzaninfinansiering etc. - eller riskkapital för nyetablerade innovativa företag och små och medelstora företag, om det är nödvändigt på grund av effekterna av den nuvarande finanskrisen.
Vi måste förbättra små och medelstora företags marknadstillträde genom framför allt ökad övervakning av marknaden och av enskilda branscher så att hinder på den inre marknaden kan upptäckas och åtgärdas.
Redovisningskraven bör i hög grad förenklas och det bör gå snabbare att starta nya företag.
Vid sitt möte den 19-20 mars enades Europeiska rådet om följande åtgärder: att undanröja befintliga hinder och förhindra att nya uppstår, att uppnå en fullt fungerande inre marknad, att minska de administrativa bördorna ytterligare, att förbättra ramvillkoren för näringslivet i syfte att upprätthålla en stark industriell bas för företagen med särskild inriktning på små och medelstora företag och innovation, att uppmuntra till partnerskap mellan olika affärsområden, forskning och utbildning, samt att öka kvaliteten på investeringar i forskning, kunskap och utbildning.
Mina damer och herrar! Jag vill även påpeka att rådet den 10 mars 2009 uppnådde en politisk överenskommelse om att det genom en ändring av direktiv 2006/112/EG ska bli möjligt för alla medlemsstater att permanent införa lägre moms på ett antal arbetsintensiva tjänster, och det handlar förstås i hög grad om tjänster som tillhandahålls av små företag.
Bland övriga lagförslag som har uppstått till följd av initiativ i samband med småföretagsakten bör rådet anta en förordning om stadgan för det europeiska privata aktiebolaget, som skulle göra det lättare för små och medelstora företag att bedriva verksamhet över gränserna.
Rådet kommer även att överväga en revidering av direktivet om sena betalningar så att små och medelstora företag får betalt i tid för sina affärstransaktioner.
När det gäller agendan för bättre lagstiftning lade kommissionen förra året fram elva nya påskyndade åtgärder för att minska de administrativa bördorna för företag och har satt som mål att de nuvarande bördorna till följd av EU:s lagstiftning ska minskas med 25 procent fram till 2012.
Beräkningar visar att detta kan leda till besparingar på omkring 30 miljarder euro och fördelarna skulle vara störst för små och medelstora företag.
Den 10 mars i år uppmanade rådet kommissionen att lägga fram förslag till nya särskilda åtgärder för att minska bördorna inom vart och ett av de 13 viktiga prioriteringsområdena i handlingsplanen.
Exempel på faktiska åtgärder i detta sammanhang är antagandet av förslag för att förenkla det tredje och det sjätte direktivet om fusioner och upplösning av handelsföretag i samband med den första behandlingen i Europaparlamentet, samt godkännandet av revideringen av det fjärde och det sjunde direktivet.
Detta viktiga arbete bör emellertid fortsätta så att de administrativa bördorna kan minskas med 25 procent och kommissionen bör snarast möjligt slutföra sin översyn av alla befintliga lagbestämmelser.
(EL) Fru talman! Jag tackar ministern för hans svar, i vilket han räknade upp alla åtgärder som planeras.
Nu gäller det förstås att tillämpningen av dessa åtgärder också leder till konkreta resultat för alla i EU som i dag har små och medelstora företag som har drabbats av krisens följder och för alla som vill starta nya små och medelstora företag.
Det är just på denna punkt som jag skulle vilja att ministern anger om det finns statistik över nya företag som startas, samt statistik över företag som försvinner.
Jag tycker att det vore intressant att få dessa jämförande siffror, om inte i dag så i ett svar framöver.
rådets tjänstgörande ordförande. - (CS) Fru talman, mina damer och herrar! I slutsatserna från mötet den 19-20 mars 2009 slog rådet fast att det kommer att krävas betydande interna och externa finansieringskällor, såväl offentliga som privata, för att finansiera åtgärder för begränsning och anpassning, särskilt i de mest utsatta utvecklingsländerna, och att EU kommer att bidra med en rimlig del av finansieringen av sådana åtgärder i utvecklingsländerna.
Kommissionens beräkningar baserade på de senaste studierna visar att de tillkommande offentliga och privata investeringarna måste öka till nästan 175 miljarder euro fram till 2020 om utsläppen ska minskas till en nivå som är förenlig med EU:s mål.
Färska undersökningar visar också att mer än hälften av dessa investeringar måste göras i utvecklingsländerna.
Sekretariatet för FN:s ramkonvention om klimatförändring beräknar vidare att anpassningskostnaderna i utvecklingsländerna år 2030 kommer att ligga på mellan 23 och 54 miljarder euro om året.
När det gäller finansieringen av begränsningsåtgärder i utvecklingsländerna har rådet intagit en tydlig ståndpunkt.
Utvecklingsländerna bör med de utvecklade ländernas hjälp upprätta strategier och planer för att etablera en ekonomi med låga koldioxidutsläpp.
I dessa strategier och planer bör man skilja mellan åtgärder som kan vidtas för sig, eftersom de inte medför några eller mycket låga kostnader eller till och med en nettovinst på medellång sikt, och åtgärder som kommer att leda till ytterligare kostnader som inte enkelt kan finansieras av de enskilda länderna själva.
För att genomföra Köpenhamnsöverenskommelsen krävs ett stöd som är tillräckligt, förutsägbart och ges i rätt tid.
Den internationella finansiella struktur som förmedlar detta stöd måste baseras på principer om effektivitet, lämplighet, jämlikhet, öppenhet, ansvar, sammanhållning, förutsägbarhet och god ekonomisk förvaltning.
När det gäller finansieringskällorna godkände rådet alternativ som man kan titta närmare på i internationella förhandlingar, däribland en strategi som bygger på medverkan i enlighet med en överenskommen skala, marknadsbaserade metoder som bygger på auktionsarrangemang, eller en kombination av dessa och andra alternativ.
Under övergången till en global marknad för handel med koldioxidutsläpp kommer dessutom flexibla mekanismer, mekanismen för ren utveckling och gemensamt genomförande att fortsätta att spela en viktig roll för att finansiera utsläppsminskningar i utvecklingsländer och övergångsekonomier.
Det kommer i detta sammanhang att vara viktigt att stärka integriteten i ett miljöperspektiv, bidraget till hållbar utveckling och en rättvis geografisk fördelning.
Marknaden för handel med koldioxidutsläpp måste dessutom utvidgas för att skicka en tydlig signal om vad koldioxidutsläppen kostar.
Det är ett av de mest kostnadseffektiva sätten att minska utsläppen samtidigt som det tydligt uppmuntrar en övergång till en ekonomi med låga koldioxidutsläpp.
Rådet har i samband med EU:s överenskommelse om klimat- och energipaketet även betonat hur detta paket bidrar till EU:s försök att finansiera åtgärder inriktade på att begränsa klimatförändringarna och anpassa sig till dem.
Det står klart att vi måste göra mycket mer på finansieringsområdet.
Rådet har beslutat att ta upp denna fråga igen under mötet i juni för att förtydliga sin ståndpunkt ytterligare i de pågående internationella förhandlingarna.
(EN) Jag vill tacka det tjeckiska ordförandeskapet för ett utförligt svar.
Jag fick det faktiskt skriftligt tidigare i dag eftersom de inte trodde att vi skulle hinna med fråga 10.
Kan jag utgå ifrån att detta verkligen är den tjeckiska regeringens åsikt, som ni just har framhållit, jag skulle verkligen känna mig uppmuntrad om jag trodde det?
Jag vill tacka er, för det innebär att den tjeckiska regeringen har kommit långt i frågor som rör klimatförändringar sedan ordförandeskapet inleddes.
Om man bortser från rådsmötet i juni, kan ni säga något om resten av tidsplanen när det gäller att nå en överenskommelse om EU:s ”rättmätiga del” när det gäller att finansiera tredjeländernas mildrande av och anpassning till klimatförändringen?
För övrigt instämmer jag helt med vad ni säger om koldioxidmarknaden och dess bidrag.
Tack, fru Doyle.
Det förvånar mig att ni hade fått svaret i förväg.
Jag har väldigt länge velat uppmuntra detta både från rådets och kommissionens sida, därför vill jag gratulera er båda för att ni har lyckats med det.
(Utrop från Avril Doyle: ”Det var för att de inte trodde att vi skulle hinna fram till fråga 10!”)
rådets tjänstgörande ordförande. - (CS) Mina damer och herrar! Ju mindre tid som återstår av det tjeckiska ordförandeskapet, desto snabbare tycks den gå och det är kanske därför vi försöker snabba på och hinna med allt det administrativa i tid.
Jag vill som svar på ledamotens fråga säga att rådet kommer att diskutera denna fråga på nytt i juni i år.
Enligt rådets uppfattning är det viktigt att inrikta sig mer på de finansiella mekanismerna i kampen mot klimatförändringarna.
Inför Köpenhamnsmötet kommer rådet att offentliggöra hur man ställer sig till olika sätt att finansiera begränsnings- och anpassningsåtgärder, stödja ny teknik och skapa de rätta förutsättningarna för ett genomförande av dessa planer.
Rådet kommer även att visa hur EU ska bidra konkret till dessa planer och förklara hur kostnaderna ska fördelas mellan medlemsstaterna, samt insatserna för att uppnå dessa mål.
Allt kommer att baseras på faktiska förslag från kommissionen.
När det gäller vissa andra problem som rör finansieringen av det globala avtalet om bekämpning av klimatförändringarna har EU gjort klart att man här vill ta på sig en proportionerlig del av ansvaret.
EU har dessutom fastställt grundläggande principer när det gäller finansieringen och har gjort klart att man tänker diskutera dessa alternativ med sina globala partner.
Men det är förstås för tidigt att lägga korten på bordet genom att offentliggöra vissa siffror.
Det vore inte klokt och förnuftigt. Det vore inte taktiskt.
Vi har en uppfattning om hur mycket pengar som kommer att krävas för att genomföra den globala planen.
Men vi behöver åtminstone på ett ungefär veta vilket slags begränsningsåtgärder som tredjeländerna planerar att genomföra.
Jag vill i detta sammanhang påpeka att EU år 2007 gjorde ett frivilligt åtagande om att minska utsläppen med 20 procent - eller, om man lyckas uppnå ett globalt avtal, med 30 procent - och detta var långt innan något annat land i världen hade offentliggjort några förslag om begränsningar överhuvudtaget.
Nu när tillfälle gavs vill jag framhärda eftersom jag tycker att om svaren på de frågor vi inte tror att vi ska hinna med kan ges på förhand så finns det ingen anledning till att svaren på de frågor som vi kommer att hinna med inte ska kunna ges på förhand, så att vi - precis som vi fick nu - kan få ett bättre och mer givande utbyte.
Jag vill tacka er båda för att ni har visat detta, och därmed belyst något som många av oss länge har velat föra fram.
Frågor som inte har besvarats på grund av tidsbrist, kommer att få skriftliga svar (se bilagan).
Frågestunden är avslutad.
(Sammanträdet avbröts kl. 20.10 och återupptogs kl. 21.00.)
Arbetstidens förläggning för personer som utför mobilt arbete avseende vägtransporter (debatt)
Nästa fråga är betänkandet av Marie Panayotopoulos-Cassiotou, för utskottet för sysselsättning och sociala frågor, om arbetstidens förläggning för personer som utför mobilt arbete avseende vägtransporter - C6-0354/2008 -
föredragande. - (EL) Fru talman! Direktivet 2002/15/ΕG behövde verkligen revideras, och efter ett betänkande som Europeiska kommissionen var skyldig att presentera lade man fram lämpliga ändringsförslag för att hjälpa denna industri, för att skydda dess arbetstagares hälsa och säkerhet och samtidigt främja en sund konkurrens.
Utskottet för sysselsättning och sociala frågor godkände yttrandet från utskottet för transport och turism och avvisade, trots min rekommendation, kommissionens förslag. Med andra ord gick utskottet inte med på att förare som är egenföretagare ska undantas från direktivets tillämpningsområde.
Jag måste påpeka att direktivet från 2002 innebar att förare som är egenföretagare ska omfattas från och med den 23 mars 2009.
Utvecklingen är inte alltid som den ter sig i kölvattnet av de intryck och den upphetsning som orsakades av debatten om ett direktiv om vägtransport.
När det gäller körtider och viloperioder har det skett en stor utveckling sedan 2002, eftersom förordning (EG) nr 561/2006, som trädde i kraft 2007, gäller alla lastbilsförare och innebär en garanti för att de har lämpliga körtider och viloperioder.
Om förare som är egenföretagare skulle omfattas av ett direktiv om arbetstid vore det därför ett bevis på att man missuppfattat begreppet egenföretagande eftersom en egenföretagare bestämmer över sin egen arbetstid. Detta vore därför en allvarlig och skadlig åtgärd mot små och medelstora företag.
Det skulle begränsa den frihet som är förknippad med att vara företagare och bidra till att skapa ytterligare administrativa bördor Och det skulle skapa ett prejudikat för att inleda en debatt om att integrera egenföretagare inom andra sektorer och därigenom begränsa deras möjlighet att arbeta så länge de vill.
Detta medför ett allvarligt problem: vem är egenföretagare och vem är ”falsk” egenföretagare?
Det är uppenbart att vissa förare utger sig för att vara egenföretagare, men inte är det.
Europeiska kommissionen föreslog att vi skulle fastställa kriterier så att vi kan skilja mellan ”falska” egenföretagare och riktiga egenföretagare.
Detta är emellertid inte möjligt eftersom kontrollerna fortfarande utförs nationellt.
Om det därför skulle fastställas vem som är ”falsk” egenföretagare och vem som inte är det i EU-lagstiftningen skulle detta inte upptäckas vid nationella kontroller.
Därmed har vi alltså möjlighet att genom våra nya förslag på medlemsstatsnivå fastställa vem som ska och vem som inte ska omfattas av direktivet om personer som utför mobilt arbete avseende vägtransporter.
I våra förslag uppmanar vi även Europeiska kommissionen att på nytt fastställa resultatet av tillämpningen av direktivet.
Jag uppmanar mina parlamentskolleger att avvisa ändringsförslaget, vars syfte är att återförvisa förslaget till utskottet, och stödja min grupps förslag, som även stöds av gruppen Alliansen liberaler och demokrater för Europa och gruppen Självständighet/Demokrati.
Fru talman, ärade parlamentsledamöter! Ni vet att vägsäkerhet är en av de prioriterade frågorna i mitt arbete som kommissionsledamot för transport.
Det är även viktigt att från början betona att även om vägsäkerhet naturligtvis är en grundläggande aspekt vid diskussioner om frågor såsom förares arbetstid handlar inte dagens debatt om vägsäkerhet utan om social lagstiftning, inte om körtid utan om arbetstid.
Den fråga vi måste besvara i dag är denna: bör entreprenörer som är egenföretagare omfattas av restriktioner i fråga om arbetstid enligt samma villkor som anställda?
Detta är något vi måste undersöka mycket noggrant, eftersom det inte någonstans i EU-lagstiftningen fastställs hur länge en egenföretagare får arbeta på ett kontor eller i ett laboratorium.
År 1998, när rådet och parlamentet för första gången debatterade direktivet om arbetstid för mobila arbetstagare, såg situationen inom vägtransport helt annorlunda ut än vad den gör i dag. Som föredraganden Marie Panayotopoulos-Cassiotou sa var det vid den tidpunkten praxis att smita från de regler som gällde körtid, vilket innebar att yrkesförare tillbringade alldeles för lång tid vid ratten.
Utifrån den föregående förordningen om körtid, som infördes 1985, var det nästan omöjligt att kontrollera körtid på ett effektivt sätt.
När det gäller detta diskuterade lagstiftarna mellan 1988 och 2002 ett kommissionsförslag vars syfte var att reglera arbetstiden, inte bara för anställda förare utan även för förare som var egenföretagare.
Som ett resultat av denna diskussion antogs sektorsdirektivet om arbetstid för mobila arbetstagare.
Förhoppningen var att minska de negativa konsekvenser som otillräckliga bestämmelser om körtid medförde för vägsäkerheten genom att utöka tillämpningsområdet för lagarna om arbetstid så att även förare som var egenföretagare omfattades.
Problemet löstes emellertid inte och efter ett förlikningsförfarande mellan parlamentet och rådet uppmanades kommissionen att väga fördelarna mot nackdelarna med att utöka bestämmelserna om arbetstid till att omfatta egenföretagare och lägga fram ett förslag 2008.
Kommissionen tillmötesgick denna begäran och offentliggjorde en detaljerad undersökning 2007 med följande slutsatser:
För det första får arbetstid inte förväxlas med körtid.
När det gäller detta har situationen förändrats radikalt.
Som ni känner till har parlamentet tillsammans med rådet antagit nya bestämmelser om körtid.
Dessa bestämmelser innebär bland annat att en digital färdskrivare, en ytterst tillförlitlig övervakningsanordning, ska användas och att ett särskilt genomförandedirektiv ska upprättas.
De nya bestämmelserna som trädde i kraft 2007 gäller alla lastbilsförare, däribland förare som är egenföretagare.
Med den nya digitala färdskrivaren, som registrerar alla lastbilens rörelser minut för minut, kan en förare inte köra mer än nio timmar om dagen och i genomsnitt 45 timmar i veckan.
Kontentan är att det nu är möjligt att övervaka tillämpningen av dessa bestämmelser mer noggrant än vad det var 1985.
För det andra finns det ingenting i gemenskapens sociala lagstiftning som styr egenföretagares arbete.
En arbetstagare som är egenföretagare kan i själva verket inte tvingas arbeta övertid såtillvida att han per definition är fri att organisera sitt arbete såsom han önskar.
Vidare är det så gott som omöjligt att i praktiken styra arbetstiden för denna grupp av människor.
För det tredje är den övergripande balansen mellan för- respektive nackdelarna med att utöka reglerna om arbetstid till att omfatta egenföretagare mycket osäker, och det är inte möjligt att visa att en tillämpning som omfattar förare som är egenföretagare kommer att ge tydliga fördelar.
Dessutom är det mycket viktigt att påpeka att tillämpningen av bestämmelser om arbetstid på förare som är egenföretagare är ineffektiv och mycket svår att genomföra, eftersom dessa förare inte måste registrera arbetstiden av löneskäl, för att inte nämna det faktum att de administrativa kostnaderna med att tillämpa sådana bestämmelser skulle kunna bli mycket höga.
För det fjärde finns det emellertid en aspekt där ingripande krävs, nämligen när det gäller förare som är ”falska” egenföretagare, dvs. förare som formellt sett är egenföretagare, men som i själva verket inte är fria att organisera sin egen verksamhet eftersom de helt och hållet är beroende av ett enda företag som de får inkomst och beställningar ifrån.
När det gäller sociala villkor är de sårbara.
Nu omfattas de i teorin av direktivet, men genom att det inte tillämpas är det inte så i praktiken.
Kommissionens förslag är därför att intensifiera genomförandet av direktivet och erbjuda förare som är ”falska” egenföretagare det sociala skydd de behöver.
Att under en ekonomisk kris införa ytterligare en administrativ och ekonomiska börda för små och sårbara företag, som drabbas av recessionens konsekvenser, vore oklokt.
Av detta skäl välkomnar kommissionen de ändringsförslag som gruppen Europeiska folkpartiet (kristdemokrater) och Europademokrater, gruppen Alliansen liberaler och demokrater för Europa och gruppen Självständighet/Demokrati har lagt fram och som överensstämmer med den gemensamma ståndpunkt som antogs vid det senaste mötet med rådet (transport), och sänder genom dessa ändringsförslag ett tydligt budskap till industrin: fenomenet med förare som är ”falska” egenföretagare kommer inte att tolereras, och lagstiftarna kommer att se till att bestämmelserna tillämpas över hela Europa.
föredragande för yttrandet från utskottet för transport och turism. - (NL) Fru talman! Sanningens ögonblick närmar sig.
I morgon eftermiddag röstar vi om Marie Panayotopoulos-Cassiotous betänkande.
Föredraganden och jag som föredragande för yttrandet från utskottet för transport och turism har samma perspektiv när det gäller fri företagsamhet. Därför har vi tillsammans undertecknat ungefär tio ändringsförslag som rådet också kan acceptera.
Jag är tacksam över att kommissionsledamot Tajani kan stödja dem.
I morgon måste vi först av allt hantera det ändringsförslag som lades fram av utskottet för sysselsättning och sociala frågor med innebörden att man vill avvisa förslaget.
Jag är fortfarande mycket upprörd över detta ändringsförslag.
Förra veckan förvandlades emellertid denna upprördhet till fasa när jag såg de europeiska fackliga organisationernas positionsdokument.
Av rädsla för vilsna rumänska eller bulgariska förare som är egenföretagare dammas osanning efter osanning av för att övertala parlamentsledamöterna att rösta mot kommissionens förslag.
I dokumentet antyds att förare som är egenföretagare arbetar 86-timmarsveckor.
Förare, både anställda och egenföretagare, får köra i genomsnitt 45 timmar per vecka under en tvåveckorsperiod, vilket kommissionsledamot Tajani också har påpekat.
Ska vi alltså utgå från att de ägnar 41 timmar i veckan åt att arbeta med sina företag?
Inte heller dokumentets argument om vägsäkerhet är hållbart.
Det finns inga belägg för att det finns något samband mellan vägsäkerhet och ett undantag för förare som är egenföretagare från bestämmelserna om arbetstid, tvärtom.
I förbigående kan påpekas att positionsdokumentet tydligt visar att de fackliga organisationerna är fullt medvetna om att deras position är mycket svag.
Miljön och den inre marknaden dras in i detta under protest, förmodligen för att visa att vi bör rösta för förslaget om avvisande när kommissionens mycket omfattande konsekvensanalys visar att förslaget kommer att gynna den inre marknadens funktion, transportsektorn och miljön.
Därför måste vi i morgon rösta mot det ändringsförslag som lagts fram av utskottet för sysselsättning och sociala frågor, där man vill avvisa förslaget, och i stället rösta för föredragandens ändringsförslag.
Jag litar på att det sunda förnuftet kommer att segra vid omröstningen.
Avslutningsvis vill jag tillägga att jag anser att det e-postmeddelande som Stephen Hughes skickade i lördags är djupt olämpligt.
Att göra politik av dödsoffren i...
(Talmannen avbröt talaren.)
för PPE-DE-gruppen. - (FI) Fru talman, mina damer och herrar! Begränsningar av arbetstiden bör inte omfatta entreprenörer och förare som är egenföretagare och lyckligtvis har både kommissionen och rådet kommit fram till denna slutsats.
I mitt hemland Finland skulle en begränsning av arbetstiden få mycket negativa följder för förare som är egenföretagare.
Förare i Finland är ofta entreprenörer som verkar i liten skala.
Mer än hälften av dem äger det fordon de kör.
De sköter därför allting själva: de underhåller sina fordon och sköter sin egen redovisning.
Förare som är egenföretagare omfattas redan nu av samma begränsningar när det gäller körtid och obligatoriska viloperioder som förare som är anställda.
Detta är viktigt inför framtiden.
Körtiderna bör inte i sig utökas, men om detta ändringsförslag från gruppen De gröna/Europeiska fria alliansen och Socialdemokratiska gruppen i Europaparlamentet skulle träda i kraft skulle förarna exempelvis inte kunna underhålla sina fordon eller sköta sin redovisning under sin lediga tid.
Hur skulle efterlevnaden av en sådan förordning förresten övervakas?
Under en ekonomisk kris är det ytterst viktigt att stödja sysselsättningen och entreprenörskapet.
Jag hoppas att alla kommer att enas med kommissionen och transportministrarna om att förare som är egenföretagare inte ska omfattas av tillämpningsområdet för reglerad arbetstid enligt detta direktiv.
för PSE-gruppen. - (NL) Fru talman, mina damer och herrar! Socialdemokratiska gruppen i Europaparlamentet anser att förslaget till revidering av bestämmelserna om arbetstid inom vägtransport inte är tillräckligt genomtänkt och att det dessutom är inkonsekvent.
Bristfälligt införlivande och bristfällig efterlevnad av lagstiftningen får inte vara en anledning till att mjuka upp bestämmelserna.
Som kommissionen säger kan lagstiftningen endast bli effektiv om den omfattar alla berörda parter.
I mina frågor till kommissionen har jag strävat efter att få klarhet i vilka åtgärder kommissionen planerar att vidta mot användningen av förare som är ”falska” egenföretagare.
När det gäller detta har rådet nu uttryckt avsikten att inte bara undanta förare som är egenföretagare från tillämpningsområdet utan att även undvika att vidta tillräckliga åtgärder mot ”falska” egenföretagare, vilket inte vunnit gehör hos PSE-gruppen.
Verksamheten för både förare som är anställda och förare som är egenföretagare är lika viktig för deras egen som för andra människors säkerhet.
Att göra skillnad mellan dem är uteslutet för vår grupp.
Jag måste stödja kommissionsledamoten: det är inte första gången som även egenföretagare har omfattats av samordningen av säkerheten, det har även skett på byggarbetsplatser för att garantera deras egen och andras säkerhet.
Under denna mandatperiods sista sammanträde måste parlamentet anta direktivet om arbetstid för mobila arbetstagare.
Som föredragande för gruppen Alliansen liberaler och demokrater för Europa anser jag att det vore oansvarigt för oss att stödja avvisandet av kommissionens text i sin helhet, vilket har föreslagits.
Vi liberaler stöder och står bakom de tiotusentals mobila arbetstagare som är egenföretagare och som vill behålla sina konkurrensfördelar eftersom de är en del av syftet med att vara egenföretagare.
Den aktuella situationen är oroväckande.
Genom det nuvarande direktivet försvinner en grundläggande princip för den fria marknaden, nämligen entreprenörskap och stöd till detta.
Det är oacceptabelt för oss att behandla dem som arbetar enligt ett anställningsavtal likadant som dem som är egenföretagare.
Till skillnad från avlönade arbetstagare arbetar egenföretagare inte ett fastställt antal timmar, utan arbetstiden avgörs av vilka varor de hanterar samt antal och typ av partier.
Att låta dem omfattas av det nya direktivet skulle i praktiken förstöra deras entreprenörskraft.
En lag som reglerar arbetstiden för egenföretagare skulle utgöra ett farligt och omotiverat prejudikat.
Det finns ingen liknande lagstiftning i någon annan sektor.
Att anta ett sådant beslut skulle ha en negativ effekt på den europeiska ekonomin.
Definitionen av nattarbete är också av stor praktisk betydelse.
För närvarande kan medlemsstaterna definiera nattarbete själva.
På så sätt blir det möjligt för dem att maximera antalet arbetstimmar för transport av passagerare och varor enligt det skiftande dagsljuset.
Som ni känner till är natt i Finland inte samma sak som natt i Italien.
Genom att tillämpa flexibilitet kan trafikstockningar vid rusningstid, liksom en majoritet av de skadliga utsläppen från trafiken, minskas.
Avslutningsvis vill jag tillägga att liberalerna som stöds av gruppen Europeiska folkpartiet (kristdemokrater) och Europademokrater och många andra ledamöter vill fortsätta debatten om direktivets grundläggande element.
Med andra ord stöder vi den flexibla, pragmatiska ståndpunkt som godkändes i rådet och föreslogs av Europeiska kommissionen när det gäller att undanta egenföretagare från direktivet.
Jag uppmanar er verkligen att rösta för detta.
Fru talman! Den oro som råder världen över och alla de åtgärder som för närvarande vidtas för att bekämpa svininfluensan saknar, i likhet med de åtgärder som vidtogs för några år sedan mot fågelinfluensan och galna kosjukan, helt proportioner med tanke på de bristfälliga ansträngningarna när det gäller det mycket högre antalet dödsfall på vägarna.
Fyrtiotusen människor dör varje år på vägarna i Europeiska unionen.
Många människor skadas eller handikappas för livet.
Detta accepteras helt enkelt som ett exempel på force majeure.
Alla vet att antalet lastbilar som är inblandade i allvarliga vägolyckor är oproportionerligt.
De vanligaste orsakerna är för hög hastighet, att föraren är uttröttad och alkohol.
Detta direktiv är ett steg mot att förhindra att förare blir uttröttade.
Inte bara körtider, som övervakas med hjälp av färdskrivaren, utan även lastnings- och avlastningstider bör nu betraktas som arbetstid för alla.
Detta är den rätta lösningen.
Om en förare redan har arbetat i flera timmar när han sätter sig bakom ratten på en 40-tonslastbil kommer han att vara trött och ha svårt att koncentrera sig.
För mig är det fullkomligt obegripligt att denna förordning endast ska gälla förare som är anställda av andra och inte egenföretagare.
Den enda ursäkten är att det är svårare att övervaka arbetstiden för egenföretagare.
Detta må vara sant, men utgör en förare som är egenföretagare en mindre risk bakom ratten när han är uttröttad än en anställd företagare?
(EN) Fru talman! Vi måste förkasta detta förslag från kommissionen av tre uppenbara anledningar.
För det första hävdar de att förordning (EG) nr 561/2006 om körtid och viloperioder omfattar alla och att det därför inte finns något problem med att egenföretagare utesluts.
Det är felaktigt.
Körtiden utgör i genomsnitt bara halva arbetstiden för en förare.
De som inte omfattas skulle i realiteten kunna få arbeta 86 timmar per vecka, alla veckor under året.
För det andra omfattas inte de hundratusentals förare som kör fordon på under 3,5 ton av bestämmelserna.
Om de undantas från detta direktiv kommer det inte att finnas någon gräns alls för deras arbetstid, vilket är än värre.
För det tredje skiljer kommissionen mellan egenföretagare och ”falska” egenföretagare, och säger att den gör detta eftersom man inte kan inspektera eller kontrollera egenföretagares arbetstid.
Om så är fallet, hur kommer de att kontrollera arbetstiden för de ”falska” egenföretagarna?
Detta är att undgå sitt ansvar och det är en öppen inbjudan för skrupulösa arbetsgivare att ständigt leta efter nya former av ”falskt” egenföretagande för att undvika lagen.
Vi måste förkasta detta förslag från kommissionen.
(FI) Fru talman! Jag vill börja med att tacka kommissionsledamot Tajani för ett utmärkt arbete och för att han i sitt tal alldeles nyss mycket lovvärt påpekade att detta i mindre grad handlar om säkerhet och antalet timmar som ägnas åt körning än om antalet timmar som ägnas åt arbete.
Vi måste respektera det faktum att det i Europa finns små och medelstora företag som sköter sitt arbete och skapar arbetstillfällen och att detta vore ett slag i ansiktet på entreprenörer som verkar i liten skala, framför allt under den rådande ekonomiska situationen.
För ungefär två veckor sedan hade vi en häftig debatt här om att det är de små och medelstora företagen som håller igång hela den europeiska ekonomin.
Nu ställs vi inför det praktiska problemet att bestämma om vi ska stödja dem eller inte.
Kommissionsledamot Tajani klargjorde vad vi bör övervaka och vad vi behöver göra för att se till att dessa förare som är egenföretagare kan fortsätta att arbeta efter de timmar de ägnat åt att köra.
Fru talman, mina damer och herrar! Jag vill lugna de ledamöter som har uttryckt oro angående den text vi debatterar.
Vägsäkerheten står definitivt inte på spel. Jag upprepar att det är en av mina prioriteringar att arbeta för att minska antalet vägolyckor.
Jag anser att vi inte bör blanda ihop arbetstid med körtid.
Jag kan mycket väl förstå det ni sa om att en egenföretagare kan arbeta först och sedan vara trött när han sätter sig bakom ratten, men jag tror inte att en egenföretagare kan styras oavsett vilket arbete han har. Naturligtvis är egenföretagaren också medveten om vad han gör.
Han kan till exempel lasta en lastbil och sedan vila i två, tre eller fyra timmar och därefter sätta sig bakom ratten igen och vara i utmärkt skick att köra ur säkerhetssynpunkt.
Faktum är att det är mycket svårt att styra någon typ av egenföretagare, hantverkare eller entreprenör i liten skala.
Dessutom är det dessa män och kvinnor som utgör ryggraden i EU:s ekonomi.
Samtidigt vill jag påpeka att vi alla är angelägna om att garantera hälsa och säkerhet för de anställda och för de arbetstagare som utger sig för att vara egenföretagare, men som i allt väsentligt är anställda.
Därför vill kommissionen - och jag tror att föredraganden delar vår ståndpunkt när det gäller detta - att den verksamhet som ”falska” egenföretagare utför också ska vara föremål för lagstadgad kontroll.
Så jag anser att detta är en viktig signal. Denna lagstiftning uppfyller verkliga krav och jag anser att det är rätt att återigen betona hur viktigt det är att ytterligare framsteg görs på detta område.
Därför vill jag be Socialdemokratiska gruppen i Europaparlamentet och gruppen De gröna/Europeiska fria alliansen att fundera över de kommentarer som har fällts och att inse att vad kommissionen anbelangar så är och förblir vägsäkerheten en prioritering. Lagstiftningen omfattar emellertid inte denna sektor, utan syftar snarare till att på ett bättre sätt reglera i synnerhet arbetstiden för alla som arbetar inom vägtransportsektorn och införliva de ”falska” egenföretagarna med de anställda eftersom de i realiteten inte är egenföretagare utan de facto anställda.
Så låt mig återigen lugna dem som uttryckt oro, eftersom jag anser att den text som kan antas är en bra text och ett steg i rätt riktning när det gäller att värna EU-medborgarnas intressen.
föredragande. - (EL) Fru talman! Jag tackar kommissionsledamoten för att han i sitt tal uttryckte sig så tydligt och för de förtydliganden han gjorde i efterhand, dvs. hans försäkran om att det viktigaste målet är vägsäkerheten och att samtidigt skydda den europeiska ekonomins konkurrenskraft samt att stödja små och medelstora företag.
Jag tackar alla mina parlamentskolleger för deras synpunkter och jag vill påpeka att det är just denna dialog vi vill lämna öppen genom att röst mot ändringsförslag 54 där kommissionens förslag avvisas.
Jag uppmanar därför alla mina parlamentskolleger att avvisa ändringsförslag 54, så att dialogen förblir öppen och så att vi kan hjälpa de arbetstagare som utnyttjas och som utger sig för att vara egenföretagare fast de i själva verket är ”falska” egenföretagare.
Vi vill bidra till att förbättra sysselsättningen inom vägtransportsektorn genom att skydda vägsäkerheten enligt den förordning som omfattar alla och värna om arbetstiderna i det direktiv som vi har framför oss.
Jag vill påminna ledamöterna om att jag skickat dem en artikel från en tysk dagstidning där exemplen tydligt visar att risken vid bilkörning inte är att föraren har arbetat för mycket utan att varje person utnyttjar den tid han eller hon har till sitt förfogande på ett dåligt sätt, oavsett om han eller hon är anställd eller egenföretagare, vilket i själva verket är irrelevant.
Det som är viktigast är att varje person tar ansvar för sina åtgärder och kör på ett omdömesgillt sätt samt uppfyller sina skyldigheter som samhällsmedborgare.
Vi kommer inte att uppnå detta genom att skapa hinder mot arbete.
När Jan Cremers nämnde byggindustrin avslöjade han avsikten hos alla dem som stöder dessa åsikter i upptakten till valet.
Debatten är härmed avslutad.
Omröstningen äger rum på tisdag den 5 maj 2009.
8.
Program för att bidra till ekonomisk återhämtning genom finansiellt stöd från gemenskapen till projekt på energiområdet (
för PPE-DE-gruppen. - (DE) Fru talman! Efter ett kort samråd med föredraganden enades vi om att punkterna 2, 3 och 5 i lagstiftningsresolutionen skulle ändras.
Jag föreslår följande engelska text till punkt 2:
(EN) ”Europaparlamentet anser att det referensbelopp som anges i lagförslaget är förenligt med den reviderade fleråriga budgetramen.”
I punkt 3 bör den första meningen strykas och resten kvarstå oförändrat: ”Europaparlamentet påminner om att man måste undvika alla omfördelningar som kan få negativa konsekvenser för andra politikområden inom EU genom att leda till en minskning av de tilldelade anslagen”
Punkt 5: ”Europaparlamentet noterar att lagstiftningsförfarandet kan slutföras så snart som finansieringen av programmet godkänts”
Kommissionens åtgärder till följd av parlamentets åtgärder och resolutioner: se protokollet
Presentation av det svenska ordförandeskapets program (debatt)
Nästa punkt är ett uttalande från rådets ordförandeskap om offentliggörandet av det svenska ordförandeskapets arbetsprogram.
rådets ordförande. - Herr talman, ärade ledamöter! Låt mig först gratulera er till valet av ny talman.
Jag ser fram emot att samarbeta med Jerzy Buzek under det svenska ordförandeskapet - och naturligtvis också tiden därefter.
Det är en ära för mig att tala inför Europaparlamentet som ordförande för Europeiska rådet.
Jag vet att uppemot hälften av er är invalda till denna församling för första gången.
Tillsammans ger ni alla röst åt 500 miljoner européer.
Det finns stora förväntningar på er.
Jag talar till er i utmaningarnas tid.
Sällan har EU-samarbetet stått inför svårare prövningar och av så olika slag.
På kort sikt har vi ambitionen att säkerställa en smidig övergång till ett nytt fördrag - Lissabonfördraget.
Nu och på lite längre sikt måste vi fortsatt hantera den ekonomiska och finansiella krisen.
Under ytan hotar en växande klimatkris som på lång sikt är den största av våra utmaningar.
En sak är klar.
För att lyckas med de många utmaningar som väntar det svenska ordförandeskapet måste vi arbeta sida vid sida med er - ni som verkar i kärnan av den europeiska demokratin.
Vi hoppas på ert stöd och samarbete, och att ni är redo att anta utmaningarna tillsammans med oss.
När vi talar om EU:s historia brukar vi framhålla att samarbetet skapat grund för fred i ett Europa som så ofta har kännetecknats av det motsatta.
Jag vill berätta för er att min farfar var svensk beredskapssoldat vid norska gränsen under andra världskriget, ett krig som Sverige stod utanför.
Det närmaste min farfar kom kriget var att då och då få en skymt av det - på betryggande avstånd.
Sådan var länge Sveriges relation till Europa: på avstånd betraktande.
När Europa stod i ruiner efter andra världskriget var Sverige orört.
Vi var ekonomiskt rikare - men fattiga på europeisk gemenskap.
För 20 år sedan kapades taggtråden mellan Österrike och Ungern.
Berlinmuren revs, och Europa ändrades nästan över en natt.
Då påbörjade flera länder den resa som ledde till att det i dag sitter representanter från 27 länder i denna sal.
Sverige var ett av dessa länder.
Den som startar sent behöver tid för att hinna ikapp.
Under det sena 80-talet börjar vårt politiska engagemang i Sverige för Europa att mogna fram.
Långsamt växer insikten om Sveriges närhet och beroende av Europa.
I arbetet med att föra Sverige in i det europeiska samarbetet, dvs. att bejaka öppenhet, globalisering och frihandel, spelade utrikesminister Carl Bildt en avgörande roll, driven av en fast övertygelse om att Sverige hörde hemma i Europa.
För 18 år sedan lämnade vi in vår ansökan om medlemskap i Europeiska unionen.
Till slut hade vi mognat i övertygelsen om att människors vardag och vår framtid bäst formas i samarbete och i gemenskap med andra, att vi hade något att bidra med - och att vi hade mycket att lära.
Nu var vi inte längre rädda för samarbete.
Vi vågade vara en del av Europa.
Dessa för Sverige omvälvande år, från mitten av 1980-talet och framåt, löpte parallellt med att mitt eget politiska engagemang fördjupades.
Längtan efter Europa var stark hos mig och hos många i min generation av svenska politiker.
Jag minns hur jag som ung och ny riksdagsledamot välkomnades att besöka Europaparlamentet.
Det var ett tecken på parlamentets öppenhet och tillgänglighet - trots att Sverige då stod utanför unionen.
Några år senare, 1997, efter det att Sverige blivit medlem, var jag med om att bygga upp PPE-gruppens ungdomsorganisation, Youth of EPP, och jag blev själv dess förste ordförande.
På det sättet fick jag se hur det europeiska samarbetet fungerade i praktiken.
Gemensamt sökte vi europeiska lösningar på europeiska problem.
Vi lärde inte bara känna varandra utan också varandras historia och kultur.
Det fick mig att lära känna Europas huvudstäder - och det antal kyrkor jag genom det besökt i Europa är inte lätta att räkna.
På 20 år har Sverige gått från att på avstånd betrakta till att vara en aktiv del i Europasamarbetet.
Det har i sin tur påverkat svenska folket.
För tio år sedan tyckte var tredje svensk att medlemskapet i EU var bra för vårt land, men lika många tyckte tvärtom.
I dag har det vänt.
Nästan två av tre svenskar menar att EU-medlemskapet är bra för Sverige.
I valet till Europaparlamentet i juni gick över 45 procent av svenskarna iväg för att rösta.
Det är åtta procentenheter fler än 2004, och det är mer än genomsnittet i Europa.
I dag är Sverige ett land som uppskattar och bejakar EU-medlemskapet.
Vi vaknade sent, men vi har flitigt arbetat oss ikapp.
Det är en seger för alla oss som tror på Europasamarbetet.
(Applåder)
Herr talman, ärade ledamöter! Vi står inför vår generations ödesfråga, ett samhällsproblem som olikt många andra växer långsamt - och bara i fel riktning.
Vår värld har feber.
Febern stiger - och det ligger på oss att reagera.
Grönlandsisen minskar med mer än 100 kubikkilometer varje år.
Istäcket i Västantarktis smälter allt snabbare.
Vi vet att enbart den minskande Grönlandsisen kan leda till en höjning av havsnivån på upp till två meter.
Effekterna blir dramatiska.
Om havsnivån skulle stiga bara en meter världen över, skulle ett hundratal miljoner människor behöva flytta bara i Asien.
Värst utsatta är människorna i Bangladesh, i östra Kina och i Vietnam.
Vi står emellertid också inför andra allvarliga konsekvenser.
Vädret kommer att förändras, och många växt- och djurarter riskerar att utrotas.
Detta även om vi håller oss inom det tvågradersmål som FN har satt upp, och som i förra veckan såväl G8 som Major Economies Forum i L'Aquila ställde sig bakom.
Vårt klimat hotas av vårt användande och vårt beroende av fossila bränslen.
Det är de dåliga nyheterna.
Så vilka är då de goda?
Även om tiden är knapp är den fortfarande på vår sida.
Vi måste dock agera nu.
Redan i dag har vi förutsättningarna för utbyggnad av förnybar energi och tekniken för energieffektivisering.
Enligt internationella energiorganet, IEA, kan mer än hälften av de åtgärder som krävs för att inte överstiga tvågradersmålet vidtas med den teknik vi redan har.
Dessutom följs åtgärder mot klimatförändringarna av mycket värdefulla sidoeffekter, effekter som i sig motiverar åtgärderna.
När vi förbrukar mindre energi, sparar vi pengar.
Vi förbättrar de offentliga finanserna samtidigt som hushållen får mer resurser.
När vi investerar i förnybar energi och energieffektiviserar, förbättrar vi vår energisäkerhet.
Vi blir mindre beroende av import från länder som ibland är både politiskt och ekonomiskt instabila.
Investeringarna i den gröna ekonomin kommer att skapa nya arbetstillfällen och driva på tillväxten under de kommande årtiondena.
Låt mig ge ett konkret exempel.
Många EU-länder drabbades i januari av gaskrisen i Ukraina.
I förra veckan pratade jag med president Jusjtjenko om hur vi ska försöka undvika en liknande händelse.
Samtidigt är det viktigt att kunna vrida på perspektiven.
Om Ukraina investerade i energieffektivitet så att landet nådde samma nivå som Tjeckien eller Slovenien, skulle det översatt i sparad mängd energi motsvara hela landets gasimport för eget bruk från Ryssland.
Ukraina skulle kunna bli helt oberoende av gasimport från Ryssland och dessutom spara mycket pengar - bara genom att öka sin egen energieffektivitet.
Det är så vi måste söka klimatsvaren.
(Applåder)
För tolv år sedan byggdes i Kyoto en koalition av frivilliga.
Bara frivillighet räcker emellertid inte.
Om vi ska lyckas få en global klimatöverenskommelse på plats, då måste resan från Kyoto till Köpenhamn gå från de frivilligas koalition till att bli allas ansvar.
Hur når vi då dit?
Europa måste agera gemensamt och samlat.
Vi måste visa ledarskap och stå vid våra löften.
Europa är avgörande för att få med andra i en global överenskommelse.
Världen över måste vi sätta ett pris på utsläppen.
Vi måste börja använda nationella koldioxidskatter och utsläppshandel.
Då växer de miljövänliga alternativen fram.
Sätts priset på användande av fossila bränslen utan hänsyn till klimatpåverkan, kommer den globala uppvärmningen att fortsätta.
Alternativen växer inte fram.
Åtgärder för att öka energieffektiviteten kommer inte att bli ekonomiskt lönsamma.
Det räcker emellertid inte.
Vi måste ha ett bredare svar på frågan ”hur?”.
Det räcker inte med att begränsa utsläppen i en krets av länder som frivilligt tar på sig reduktioner, men som tillsammans bara står för 30 procent av utsläppen.
Inte heller räcker det med lösningar som bara bygger på begränsningar i de mest utvecklade länderna.
För även om de så kallade Annex I-länderna skulle minska sina utsläpp till noll skulle utvecklingsländernas snabbt växande utsläpp ändå leda oss över tvågradersmålet.
Därför måste vi diskutera finansieringen av investeringar i utvecklingsländerna.
Vi behöver säkra en snabb tekniköverföring, och vi behöver se till att också utvecklingsländerna gör åtaganden för att bryta den utveckling de nu har framför sig.
Vi kommer dessutom att kräva tydliga åtaganden på medellång sikt även för länder utanför Europa.
Ansvar av några måste nu bli allas ansvar.
Jag vet att Europaparlamentet kommer att ta sitt ansvar.
Det svenska ordförandeskapet ser er som våra allierade.
Nu vill vi skriva historien om hur klimathotet avvärjdes, och vi vill skriva den tillsammans med er.
Herr talman, ärade ledamöter! Den ekonomiska och finansiella krisen spreds som en löpeld över världen inom loppet av några veckor.
Några hade varnat, men för de allra flesta kom den som en överraskning, framför allt dess omfattning och djup.
I en global värld sprider sig även problem snabbt till andra.
Kraften i nedgången är av det slaget att ingen har någon mirakelkur för att snabbt ta sig ur den.
Ett samordnat agerande från EU:s sida är det bästa verktyg vi har för att möta krisens utmaningar.
Mycket kan dessutom fortfarande gå snett.
Givet omständigheterna lyckades EU visa ledarskap genom prövningarna.
Vi enades om garantier och trafikregler för att stödja bankerna.
Vi enades om en gemensam återhämtningsplan för att stimulera ekonomin.
President Sarkozy och det franska ordförandeskapet spelade en viktig roll i arbetet, men jag vill också framhålla att Europaparlamentet var pådrivande.
Nu behöver vi ägna hösten åt att diskutera fortsatta åtgärder för att ta oss genom krisen.
Det ekonomiska läget är fortfarande kärvt, och de offentliga finanserna är nu ansträngda i alla medlemsländer.
Enligt kommissionens prognoser kommer underskotten inom EU att överstiga 80 procent av BNP nästa år.
Det går inte att blunda och låtsas att det inte är ett problem.
Mitt i allt detta får vi inte heller glömma att det bakom dessa siffror finns människor som känner oro för sina jobb, och som undrar hur de ska klara av att betala sitt boende och att upprätthålla sin levnadsstandard.
Det är vår uppgift att svara.
När miljontals européer förlorar sina jobb och hamnar i utanförskap hotas hela vår välfärd. Detta i ett läge där trycket på vår välfärd redan är stort.
Vi lever längre, samtidigt som vi arbetar kortare och föder färre barn.
Om 50 år kommer det att finnas dubbelt så många äldre människor som barn i Europa om denna trend håller i sig.
Så vad kan vi då göra?
Vi måste återupprätta förtroendet för finansmarknaderna.
Vi måste snabbt få en fungerande tillsyn på plats för att förhindra att liknande kriser uppstår i framtiden.
Det svenska ordförandeskapet arbetar för att rådet ska kunna enas om detta innan årets slut.
Vi hoppas på er hjälp att föra det snabbt och slutgiltigt i hamn.
Våra medborgare kommer inte att acceptera att skattemedel används fler gånger för att rädda finansinstitut som har agerat oansvarigt.
Vi måste snabbt ta oss ur de växande offentliga underskotten genom en samordnad exit strategy och en stegvis återgång till stabilitetspaktens regler.
Annars följs kortvariga obalanser av kroniska underskott.
Då väntar stora nedskärningar, som ju redan är en realitet i delar av EU, och som vi har tidigare erfarenhet av i Sverige.
Då väntar massarbetslöshet, social oro och stigande skattetryck.
Vi måste säkerställa en social dimension i Europapolitiken som bygger på sunda offentliga finanser och på att få in fler på arbetsmarknaden.
Det är det absolut bästa sättet att värna våra välfärdssystem.
Jag vet att inte minst här i Europaparlamentet är detta en mycket viktig fråga.
Det är ohållbart att tre av tio européer i arbetsför ålder står utanför arbetsmarknaden.
Målet måste vara en aktiv arbetsmarknadspolitik som tillsammans med väl fungerande trygghetssystem effektivt kan hantera omställningar.
Vi måste stärka den enskildes anställningsbarhet och möjlighet att göra sig gällande på arbetsmarknaden.
Vidare måste vi aktivera och återaktivera arbetslösa.
Med fler i arbete kommer det att finnas mer till stöd för dem som står utanför.
Vi måste också satsa på reformer, modernisering och anpassning till en ny verklighet.
Världen utanför EU står inte stilla.
Den rör sig framåt i en fantastisk fart.
Det är något vi bör bejaka och anamma.
En översyn av EU:s Lissabonstrategi kan bidra till en nödvändig reformagenda.
Den diskussionen kommer vi att inleda under hösten.
I den ekonomiska krisens spår kan vi se idéer om ökad protektionism.
WTO bekräftar att antalet handelsbegränsande åtgärder ökat avsevärt under de senaste tre månaderna.
Därför välkomnar jag L'Aquila-överenskommelsen om en nystart av Doharundan - för att se till att världens länder återigen slår in på den frihandelsvänliga väg som vi vet gynnar oss alla i längden.
Målsättningen måste vara ett EU som kommer stärkt ur krisen.
Herr talman, ärade ledamöter! När jag reser omkring i Sverige och pratar om EU-samarbetet får jag få frågor om EU:s institutioner.
Det handlar snarare om krokiga gurkor, snus och andra vardagsnära frågor.
Icke desto mindre: det institutionella ramverket är viktigt, eftersom det definierar vad vi kan göra och på vilka områden.
Därför är ratificeringen av Lissabonfördraget så central.
Fördraget kommer att göra EU mer demokratiskt, mer transparent, mer effektivt och mer inflytelserikt på den internationella arenan.
Allra viktigast dock att med Lissabonfördraget på plats sätts punkten för en inåtvänd fas i EU-samarbetet.
Det är nu dags för EU att blicka utåt och framåt.
Det svenska ordförandeskapet är redo att genomföra allt förberedande arbete för att säkerställa en smidig övergång till ett nytt fördrag, men det förutsätter förstås att fördraget har ratificerats av alla medlemsländer.
Låt oss hoppas att det ska bli verklighet inom de kommande månaderna.
Den internationella brottsligheten växer sig allt starkare.
Kriminella nätverk ser inte längre några gränser för sin verksamhet.
Vi ser hur handel med narkotika och med människor breder ut sig.
Det hotar våra demokratiska värden, och det hotar våra medborgare.
Samtidigt är friheten att röra sig fritt över våra gränser grundläggande för vår gemenskap - att studera, arbeta och leva i ett annat EU-land.
En ny tid kräver emellertid nya svar.
Därför kommer vi att utarbeta ett nytt program på området under hösten, nämligen det som vi kallar Stockholmsprogrammet.
Stockholmsprogrammet vässar de instrument som skapar säkerhet i EU, och som bekämpar organiserad brottslighet och terrorism.
Samtidigt skapar vi en bättre balans mellan dessa instrument och de åtgärder som säkerställer rättssäkerhet och som skyddar individens rättigheter.
Det ser också till att den som söker asyl i EU möts med ett gemensamt och rättssäkert system - mer lika mottagning och asylprövning, mer lika återvändandepolitik.
Drömmen om en framtid i Europa är stark hos många.
Samtidigt blir Europas befolkning äldre och äldre.
Genom ett flexibelt system för arbetskraftsinvandring kan dessa två realiteter mötas.
Herr talman, ärade ledamöter! För drygt 50 år sedan lade sex länder grunden för det europeiska samarbetet.
I dag är vi 27.
Vi har vuxit i styrka och inflytande, och vi har vuxit i välfärd och i mångfald.
Europa har berikats.
Därmed står vi också bättre rustade för att tillvarata såväl globaliseringens möjligheter, som för att möta dess utmaningar.
Ensam är inte stark.
Det heter ”förhandlingar” om medlemskap.
Ytterst handlar medlemskapet emellertid om att dela en gemensam värdegrund och följa gemensamma regler.
Det här begrundas nu av dem som står utanför - från Reykjavik, till Ankara, över västra Balkan.
De båda ledarna på Cypern står inför en historisk möjlighet att enas om en lösning för att återförena den ö som under alltför lång tid varit delad.
För dem som är innanför kan det locka till att låta medlemskapsprocessen bli tillfället att lösa långdragna tvistefrågor.
I sådana fall måste vi hitta lösningar som kan gynna bägge sidor och öppna vägar framåt.
Annars äventyras framsteg i målen om fortsatt europeisk integration.
Det svenska ordförandeskapet kommer att verka för att föra utvidgningsprocessen framåt enligt de åtaganden som EU gjort, och på strikt basis av de kriterier som gäller.
Vi ska agera ”honest broker”.
Herr talman, ärade ledamöter! Med styrka och inflytande följer ett globalt ansvar, som vi fortfarande strävar efter att axla.
På det följer en skyldighet att använda det ansvaret för allas bästa.
EU ska arbeta för fred, frihet, demokrati och mänskliga rättigheter.
Vi har ett ansvar att stödja de fattigaste och mest utsatta länderna i världen, ett ansvar att leva upp till FN:s millenniemål.
Vi har ett ansvar att stödja FN-arbetet också i andra delar, att arbeta tillsammans med våra strategiska partners, att engagera oss i världens krishärdar - oavsett om det gäller fredsprocessen i Mellanöstern, Iran, Afghanistan, Pakistan, Nordkorea eller de stora utmaningarna på den afrikanska kontinenten.
Vi har emellertid också ett ansvar för regionala initiativ som Medelhavsunionen och det östliga partnerskapet som skapar stabilitet och samverkan mellan grannländer med olika förutsättningar.
Jag är särskilt tacksam för Europaparlamentets drivande roll vad gäller Östersjösamarbetet.
Redan 2005 presenterade parlamentet ett förslag till en strategi för regionen.
Nu hoppas vi att detta initiativ kan krönas med antagandet av en Östersjöstrategi vid Europeiska rådets möte i oktober.
Konflikterna på Balkan på 90-talet blev en början på EU:s engagemang som krishanterare, ett engagemang som nu stadigt växer.
I dag deltar EU i ett tiotal krisinsatser världen över.
I vår tid knackar världens problem på EU:s dörr.
Över hela vår värld - och inte minst i vårt närområde - knyts många människors förhoppning om sin egen utveckling till samarbetet.
Låt oss tillsammans motsvara de förväntningarna.
(Applåder)
Herr talman, ärade ledamöter! Det europeiska samarbetet har gjort att vår kontinent i dag lever i fred och i välstånd, under frihet och stabilitet.
Vi har öppna gränser och en social modell som kombinerar marknadsekonomi med omtanke om varandra.
Detta är vårt gemensamma Europa.
Våra medborgare vill emellertid också känna att Europa bärs av idéer för framtiden och att samarbetet inte bara har ett historiskt syfte utan är framåtblickande.
Därför har vi som folkvalda ett ansvar för att tala om vad vi vill med Europa.
Låt mig berätta hur jag ser på framtidens Europa.
Jag vill se ett Europa som med kraft agerar för demokrati, fred, frihet och mänskliga rättigheter på den globala arenan, och som vågar ta plats på den utrikespolitiska scenen.
Bland oss har vi nämligen erfarenheter av hur det är att leva utan demokrati och frihet. Därmed har vi också trovärdigheten att agera.
Jag vill se ett Europa som tar ledningen i kampen mot klimathotet, och som ser bortom lockelsen att konkurrera med en industri som inte betalar för de utsläpp som förstör vårt klimat, och som ställer om incitamenten så att grön teknik lönar sig, för att våra barn och deras barn ska få uppleva naturen som vi känner den.
Jag vill se ett Europa som tar ansvar för ekonomin. Lending for spending kan inte vara den enda devisen.
Inte heller kan det vara så att ”vinster är privata och förluster statliga”.
Låt oss bygga upp de offentliga finanserna igen.
Reglera sunda finansmarknader. Säkra de ekonomiska reformer som vi behöver för tillväxt och en industri som är konkurrenskraftig även i framtiden.
Jag vill se ett Europa som vidareutvecklar sin sociala modell, ett Europa som kombinerar ett väl fungerande välfärdssystem med tillväxt - med social sammanhållning, ett Europa som genom arbete, företagande och sunda offentliga finanser skapar utrymme för att upprätthålla och utveckla våra välfärdsmodeller, med alla våra medborgares bästa för ögonen.
Jag vill se ett Europa som inte låter sig lockas av protektionismens kortsiktiga korståg, ett Europa som slår vakt om den inre marknad som lagt grunden för vårt EU-samarbete, och som låter varor och tjänster strömma fritt över våra gränser, till förmån för oss själva och för resten av världen.
Jag vill se ett Europa som är ödmjukt inför olikheter, öppet för andras argument och som har en stark vilja att finna kompromisser, med det gemensamma bästa för sinnet.
Ett sådant Europa står sig starkt i alla tider.
(Applåder)
Herr talman, ärade ledamöter! Det är en ära för mig att stå här tillsammans med er och representera den europeiska demokratin.
Många har sagt mig att detta blir det svåraste ordförandeskapet på många år.
Prövningarna är många, och vi måste förbereda oss på det oväntade.
Många frågar sig om ett land av Sveriges storlek kan axla detta ansvar.
Inte ensamma, men tillsammans kan vi anta utmaningarna.
Låt oss göra det med visioner och handlingskraft, med insatser och mod.
Europa behöver det.
Människorna i Europa behöver det.
Europaprojektet handlar om drömmen om att gemensamt lösa människors problem.
Den drömmen gör Europa starkt.
Detta år, 2009, är ett ödesår för Europasamarbetet.
Nu har vi chansen att ta nästa steg.
Det svenska ordförandeskapet är redo att anta utmaningen.
Låt oss anta den tillsammans!
(Kraftiga applåder)
kommissionens ordförande. - (EN) Herr talman! Dessa tider är inte vanliga tider och detta kommer inte att vara något vanligt ordförandeskap.
Förutom det vanliga lagstiftningsarbetet kommer det svenska ordförandeskapet att ha andra typer av högst politiska utmaningar, och ingen är bättre lämpad att hantera dessa utmaningar än statsminister Fredrik Reinfeldt och det svenska ordförandeskapet.
I dag vill jag belysa två av de största politiska utmaningar som EU står inför under de kommande sex månaderna, nämligen att hantera den ekonomiska krisen och att förhandla fram en ambitiös internationell överenskommelse om klimatförändringarna i Köpenhamn.
Den värsta finansiella och ekonomiska krisen i mannaminne fortsätter att ha förödande effekter för våra samhällen och familjer. Särskilt arbetslösheten fortsätter att växa.
Att få ekonomin tillbaka på rätt spår är den främsta prioriteringen.
EU:s gemensamma åtgärder har lett till en exempellös finansiell insats som ger konkreta resultat.
Vi har också visat solidaritet mellan medlemsstaterna, till exempel genom att fördubbla taket för betalningsbalansstöd till medlemsstater som inte ingår i euroområdet, till 50 miljarder euro.
Vi behöver nu till fullo genomföra återhämtningspaketet i alla dess aspekter och se till att det tar sig uttryck i skapande av arbetstillfällen och främjande av grundläggande ekonomisk verksamhet.
Jag ser det som nödvändigt att prioritera åtgärder som begränsar arbetslösheten och som ser till att folk kommer tillbaka till arbetsmarknaden.
Här kan vi bygga vidare på resultaten från sysselsättningstoppmötet i maj, som var en del av kommissionens initiativ tillsammans med det tjeckiska, svenska och spanska ordförandeskapet.
Vi behöver omsätta det gemensamma åtagandet för ungdomar och sysselsättning i praktiken.
Naturligtvis ligger ansvaret för arbetsmarknadspolitiken hos medlemsstaterna, men vi kan och bör använda befintliga EU-instrument för att hjälpa medlemsstaterna upprätthålla sysselsättningen och utbilda medborgarna för framtidens jobb.
Därför kommer kommissionen att lägga fram ett förslag för att förenkla förfarandena för strukturfonderna och undanröja behovet av nationell medfinansiering i fråga om Europeiska socialfonden för 2009 och 2010.
Vi kommer också att omplacera resurser för att finansiera ett nytt mikrokreditsystem för sysselsättning och socialt deltagande.
Jag hoppas att Europaparlamentet kommer att stödja dessa förslag.
Kommissionens förslag utifrån ”de Larosière-rapporten”, som jag beställde i oktober förra året, kommer att utgöra grunden för en stärkt tillsyn och reglering av finansmarknaden.
Med de förslag som redan lagts fram - många av dem är redan godkända av parlamentet och av rådet, vissa är fortfarande under behandling i vår beslutsprocess - tar vi verkligen ledningen globalt i reformen av det internationella finansiella systemet.
Jag är säker på att vi kommer att fortsätta så vid G20-mötet i Pittsburgh i september.
Att göra framsteg med alla dessa frågor under de kommande sex månaderna är avgörande för att kunna bygga upp en ny ekonomi, eftersom ekonomin efter krisen definitivt inte kan och inte kommer att vara densamma som ekonomin före krisen.
Vi behöver omforma vår ekonomiska modell och åter sätta värderingarna i centrum för vår sociala marknadsekonomi, där de hör hemma.
Vi måste bygga upp en ekonomi och ett samhälle som grundas på möjligheter, ansvar och solidaritet, en ekonomi som kommer att behöva hitta nya vägar till tillväxt eftersom vi inte alltid kan förlita oss på monetära och finansiella stimulansåtgärder.
Vi måste bygga upp ett EU med öppna och väl fungerande marknader, ett EU med smart, miljövänlig tillväxt, ett EU med effektivare reglering och tillsyn av finansmarknaderna, ett EU som fördjupar sin inre marknad och till fullo utnyttjar dess potential, ett EU som motstår tendensen till splittring och protektionism.
När det gäller klimatförändringarna är EU redan den första regionen i världen som genomför långtgående, rättsligt bindande klimat- och energimål.
Jag är stolt över hur kommissionen arbetade med det förra parlamentet och rådet för att införa denna lagstiftning och jag vill ha ett nära samarbete med er och med ordförandeskapet under tiden före toppmötet i Köpenhamn.
Vår ledarroll uppskattades i hög utsträckning vid förra veckans möten i L'Aquila med G8 och i Major Economies Forum.
Ni har hört om de framsteg som gjordes vid dessa möten.
För första gången åtog sig alla deltagare att sätta ett tak på 2°C för temperaturökningen för att respektera klimatforskningen.
Detta är utan tvivel ett välkommet framsteg men vi får inte lura oss själva. Vår ambition och vårt åtagande matchas ännu inte av de andra.
EU ligger långt före genomsnittet i resten av världen och, uppriktigt sagt, då det är 145 dagar kvar till Köpenhamnstoppmötet oroar det mig.
Under de kommande veckorna kommer vi att trappa upp vårt arbete med internationella partner för att se till att tydliga åtaganden görs i Köpenhamn.
Vi behöver också göra framsteg i fråga om nödvändiga medel för att stödja utvecklingsländer och främja tekniköverföringar.
I september kommer kommissionen att lägga fram sina finansieringsförslag så att vi kan nå ett europeiskt samförstånd och förhandla med andra.
Dagordningen för klimatförändringarna är naturligtvis nära knuten till en annan prioritering: trygg energiförsörjning.
I dag kommer kommissionen att anta förslag för att stärka våra regler angående säkra gasleveranser och stärka solidariteten mellan medlemsstaterna, och jag litar på att det svenska ordförandeskapet kommer att arbeta vidare med dessa med ert stöd.
Dessa är de viktigaste prioriteringarna - vilket är helt i sin ordning.
Men det finns många andra saker som behöver göras under de kommande sex månaderna.
Låt mig bara flagga för Stockholmsprogrammet, där kommissionen nyligen har lagt fram en ambitiös vision som sätter medborgaren i centrum för vår politik om rättvisa, frihet och säkerhet, och där man balanserar säkerheten mot skyddet av de medborgerliga friheterna och de grundläggande rättigheterna.
Under större delen av detta årtionde har EU ägnat sig åt inre institutionella debatter.
Förändringar i vårt viktigaste fördrag är helt nödvändiga för att ge det utvidgade EU förutsättningar att kunna arbeta demokratiskt och effektivt.
Jag hoppas att ratificeringen av Lissabonfördraget kommer att ske under de närmaste månaderna så att vi kan omsätta dess bestämmelser i praktiken och gå vidare med den politiska dagordning som jag just har skisserat.
Det är viktigt att diskutera förfaranden men jag anser att det är ännu viktigare att diskutera innehållet.
Det svenska ordförandeskapet och det kommande spanska ordförandeskapet kommer förhoppningsvis att behöva övervaka en komplex övergång till det nya fördraget där kommissionen och parlamentet kommer att behöva spela en viktig roll.
EU har konstant förnyat sig, från den ursprungliga uppgiften att läka en krigshärjad världsdel till byggandet av den inre marknaden och senare vidare till Europas återförening.
Under de senaste 50 åren har EU konsekvent överträffat förväntningarna och fått farhågorna att komma på skam.
Jag är säker på att vi också kommer att klara den nya utmaning som vi står inför, dvs. att lägga grunden för en smart och miljövänlig ekonomi för framtiden.
Vi kommer att lyckas om vi beaktar den viktigaste lärdomen från ett halvt århundrade av europeisk integration: EU går framåt när alla dess delar samarbetar i en anda av öppenhet, tillit och partnerskap.
I det svenska ordförandeskapets program erkänns detta. Kommissionen är redo att spela sin roll och jag är säker på att även Europaparlamentet är det.
(Applåder)
för PPE-gruppen. - (FR) Herr talman! Jag vänder mig normalt inte till er men i dag ska jag för första gången ägna er en minut.
För det första, herr Buzek, hyllar jag er som motståndsman och som en av grundarna av Solidarnoœæ, som den man från Schlesien som aldrig glömde sina rötter, sin historia eller sina värderingar.
Inom Europeiska folkpartiets grupp (kristdemokrater) är vi också stolta över att ha övertygat det stora flertalet ledamöter i Europaparlamentet från alla politiska bakgrunder - även Martin Schulz - att göra er till talesman för 500 miljoner medborgare.
Valet av er som talman är en symbol för detta öppna Europa, för detta toleranta Europa, för detta politiska Europa som förespråkas av PPE-gruppen och av de flesta ledamöter här i parlamentet.
Herr rådsordförande, herr kommissionsordförande! Vad vi förväntar oss av er att ni kommer att göra handling till det ledande temat för det svenska ordförandeskapet under de kommande sex månaderna - med andra ord, inför den dubbla utmaningen med ekonomin och klimatförändringarna menar vi att vi måste göra mer, och snabbare, för att ta oss ur krisen, genom att fullständigt tillämpa vår sociala marknadsekonomi.
Jag tror definitivt att det är ekonomins livskraft och endast detta som kommer att möjliggöra för oss att föra den verkligt sociala politik som vi behöver.
Om vi vill ha en återhämtning och om vi vill att den kommer från EU och inte från Asien, vilket kan väntas, måste vi utan tvekan skynda på saker i dag.
När krisen är över kommer vinnarna att vara de som satsade på innovation, på utbildning - kort sagt, på handling.
I detta avseende föreslår PPE-gruppen bland annat att man ska öka stödet till små och medelstora företag, som är centrala för att bevara och skapa arbetstillfällen.
Jag vill också framhålla att den ekonomiska krisen inte fordrar ett nationellt svar utan ett europeiskt svar. Våra medborgare är övertygade om detta.
Man behöver bara se på opinionsundersökningarna i de olika länderna. Över 66 procent av tyskarna och över 70 procent av EU-medborgarna är övertygade.
Mer handling och snabbare handling, herr Reinfeldt, herr Barroso, det är också vad PPE-gruppen förväntar sig av er i kampen mot den globala uppvärmningen.
Det är EU:s ansvar att under er ledning leda världen i denna process, och alla här medger att det är en brådskande och högt prioriterad process.
Vilket tillfälle är bättre för att agera och skynda på saker än den konferens om klimatförändringarna som ska hållas i december i Köpenhamn, det vill säga på vårt eget territorium!
När det gäller klimatförändringarna har vi i EU visat bortom alla tvivel att vi kan vidta åtgärder bara vi vill.
Uppgiften är nu att utnyttja detta för att få de andra världsmakterna att ansluta sig.
Jag tänker naturligtvis på Förenta staterna, som måste omsätta ord i handling, men jag tänker också på tillväxtländerna, vare sig det är Kina, Indien eller Brasilien, som inte längre kan bortse från att de i stor utsträckning bär ansvaret för den globala uppvärmningen.
Vi ska därför bedöma det svenska ordförandeskapet efter hur det klarar krisen och mot bakgrund av dess resultat i miljöfrågorna.
Avslutningsvis måste EU, för att agera kraftfullt på dessa båda fronter, vara utrustat med lämpliga institutioner.
Det senaste året har tydliggjort att det med samma fördrag och med samma föråldrade enhällighetsprincip var möjligt att göra framsteg med EU men att det också var möjligt att hamna i ett dödläge.
Det handlar om politisk vilja, herr Reinfeldt och herr Barroso. Snabba på.
Det är var PPE-gruppen ber er göra under de kommande sex månaderna, och vi har förtroende för det svenska ordförandeskapet.
Snabba på.
Det är vad EU-medborgarna önskade när de valde detta parlament och det är det vi måste ge dem om vi vill se fler av dem dyka upp vid valet om fem år.
(Applåder)
Herr talman, premiärminister Reinfeldt, mina damer och herrar! Det svenska ordförandeskapet inträffar under en period när institutionerna får en nystart.
Det är inte bara Europaparlamentet som börjar på nytt.
EU är inne i en övergångsperiod mellan Nicefördraget och Lissabonfördraget. Som vi alla vet är det en tid av osäkerhet, men inte desto mindre behöver vi klarhet i fråga om politiska beslut om ekonomiska och finansiella frågor, arbetsmarknadsfrågor och klimatfrågor i EU och dess medlemsstater.
Ni har talat om detta och jag håller med i mycket av det ni sade.
Klimatförändringarna är naturligtvis den viktigaste frågan och ni har gett den rätt prioritering.
Jobbkrisen kräver naturligtvis också en omedelbar och ändamålsenlig lösning.
Därför ber vi er att under ert ordförandeskap uppmana medlemsstaterna att ta investeringsplanerna och de ekonomiska återhämtningsplanerna på större allvar än de hittills gjort.
Vad vi främst behöver är att bevara arbetstillfällena - nu, inte nästa år, eftersom hotet mot jobben finns här och nu.
Anställningstryggheten är avgörande för samhällets inre stabilitet.
Därför förväntar vi oss att ni ger högsta prioritet åt arbetstillfällen och anställningstrygghet på något sätt, till exempel genom att kombinera miljöskydd och industripolitik, vilket är en mycket intelligent lösning.
När det gäller anställningstrygghet vill jag säga er detta, herr Reinfeldt: vad som på allvar äventyrar EU:s arbetstillfällen och i ännu högre grad äventyrar den sociala sammanhållningen är EG-domstolens rättspraxis.
Som ni just har sagt reser ni mycket i Sverige och i Europa.
Det gör vi också och vad vi hör från våra medborgare är att de inte vill ha ett EU där företag flyttar från land till land och sänker lönenivån.
Därför behöver vi initiativ från EU.
(Applåder)
Vi behöver dessa initiativ till följd av EG-domstolens domar i målen Laval, Viking, Rüffert och Luxemburg.
Dessa är åtgärder som ni behöver hantera under ert ordförandeskap, och ni i synnerhet, eftersom Sverige drabbas av denna missriktade politik och denna missriktade rättspraxis.
Ni behöver också hantera en annan institutionell fråga, nämligen frågan om hur nästa kommission ska utses.
Här måste jag säga att jag på sätt och vis får det allmänna intrycket att inte bara ni utan också alla era kolleger i rådet har påverkats av den nya starten för institutionerna och ovissheten om vilket fördrag vi faktiskt bör ha som grund för våra åtgärder, och att ingen riktigt vet var vi står.
Det är lite som Astrid Lindgrens Pippi Långstrump i hennes Villa Villekulla - jag ska göra världen som jag vill att den ska vara.
Underbart!
Om vi utser kommissionens ordförande på grundval av Nicefördraget kommer vi att ha 20 kommissionsledamöter.
I detta fall skulle jag vilja veta vilket land som inte kommer att ha någon kommissionsledamot.
Här kommer rådet naturligtvis att säga ”nej, vi vill definitivt inte starta ett blodbad bakom lyckta dörrar.
Så vi har en perfekt lösning - inledningsvis utser vi kommissionsledamoten på grundval av Nicefördraget.
Det kommer att ta ett par månader för kommissionen att installeras och vid det laget kommer irländarna att ha röstat och vi kommer att ha Lissabonfördraget.
Då kan vi rösta om allt annat på grundval av Lissabonfördraget.
Toppen!”
Vi är en rättsligt grundad gemenskap - det är åtminstone vad jag trott hittills - där grundvalen är den gällande rätten.
Den gällande rätten är Nicefördraget.
För övrigt finns det någon som, i egenskap av fördragens väktare, först av allt måste förtydliga vilken rättslig grund som ska tillämpas.
Det är kommissionens ordförande, men jag har inte hört ett ord från honom i denna fråga.
Därför vill jag säga mycket tydligt vad vi förväntar oss.
Mitt förslag, herr statsminister, var att ni inte skulle ta beslutet om formalisering omedelbart, utan först skicka er kandidat till parlamentet så att han kan berätta för oss vad han vill göra för att återställa ekonomin, bevara arbetstillfällena, bekämpa klimatförändringarna, införa en sysselsättningspakt, ta initiativ till ett direktiv om offentliga tjänster och till att förbättra direktivet om utstationering av arbetstagare samt inrätta en garanti mellan kommissionen och parlamentet i fråga om utvärderingen av de sociala följderna av kommissionens initiativ.
Vi kunde redan ha diskuterat allt med kandidaten för flera veckor sedan för att se om han skulle få en majoritetsröst i parlamentet på grundval av sina förslag.
Sedan skulle ni ha kunnat fatta ett beslut om formalisering.
Ni valde i stället en annan väg.
Ni sade ”nej, vi kommer först att fatta beslut om formalisering och sedan skicka kandidaten”.
Jag är rädd för att detta var ytterligare ett misstag och jag är också rädd för att denna kandidat, om han inte gör en avsevärd ansträngning, inte kommer att få någon majoritetsröst här i parlamentet.
(Applåder)
Jag vill verkligen tydliggöra detta så att vad som troligen kommer att bli den största tvistefrågan under ert ordförandeskap är helt klart mellan oss redan från början.
Vi förväntar oss institutionell tydlighet, vi förväntar oss ett socialpolitiskt åtagande och jag räknar med att vi kommer att hålla med er när det gäller klimatpolitiken.
Herr talman! Bara för er skull har jag hållit min talartid exakt.
Ni kommer att se att mina sex minuter tar slut om några sekunder.
Ni kommer inte att behöva tillrättavisa mig - jag visste att det var det ni tänkte göra och jag ville inte ge er det nöjet.
(Applåder)
Herr talman! För det första vill jag säga till Fredrik Reinfeldt att gruppen Allianser liberaler och demokrater för Europa till fullo ställer sig bakom det svenska ordförandeskapets prioriteringar, det vill säga ratificeringen av Lissabonfördraget, som vi naturligtvis förväntar oss ska genomföras snabbt och fullständigt, förberedelserna inför toppmötet om klimatförändringar i Köpenhamn som redan har nämnts och som är en prioritering som vi helt delar, och slutligen också Stockholmsprogrammet.
Dessutom, och detta är temat för mitt anförande, herr Reinfeldt, vill jag hänvisa till en fråga som tas upp i varje inlägg här i parlamentet - kampen mot den ekonomiska och finansiella krisen - för att säga till er att ni kommer att leda Europeiska rådet vid en mycket bestämd tidpunkt.
Det är bra att det är Sverige som är ordförande för rådet eftersom ni har särskild erfarenhet på detta område.
Under 1990-talet upplevde Sverige exakt samma ekonomiska kris som vi nu upplever i hela Europa och i hela världen.
Ni har upplevt en kris inom fastighetssektorn.
Under 1990-talet hade ni också en finanskris och ni löste alla dessa problem genom att direkt ta itu med problemen inom finanssektorn.
Mitt budskap till er är att ni måste agera på precis samma sätt i dag på EU-nivå, eftersom det är vad vi saknar.
Vi försöker bekämpa den ekonomiska och finansiella krisen genom 27 olika strategier i de olika länderna. Det kommer aldrig att lyckas.
Vi förväntar oss att ni använder er erfarenhet från Sverige, eftersom det Sverige gjorde var en framgång, till skillnad från Japan, som har varit ekonomiskt stillastående under lång tid.
Sverige tog sig ur krisen eftersom ni omedelbart hanterade problemen inom finanssektorn, något som för närvarande inte görs i EU.
Tanken är att Storbritannien kan nationalisera sina banker medan andra - särskilt Frankrike - kan rekapitalisera dem.
I Tyskland pågår arbetet med att skapa avvecklingsenheter, ”bad banks”, medan man i Beneluxländerna gör lite av varje på samma gång.
Resultatet är att det inte finns någon enhetlig strategi.
Förenta staterna stabiliserar sina banker och undanröjer de dåliga verksamheterna samtidigt som vi fortsätter att ha problem.
Min uppmaning till er är därför att ni använder er erfarenhet för att presentera en enhetlig räddningsplan för EU:s finanssektor som ska utgöra grunden för den ekonomiska återhämtningen.
Utan en sådan plan kommer det aldrig att ske någon ekonomisk återhämtning, bankerna kommer inte att börja låna ut pengar igen, och så vidare.
Detta måste vara er främsta prioritering.
(EN) Den andra punkten är att vi hoppas att ni, tillsammans med kommissionen, också kan lägga fram en ny återhämtningsplan, eftersom 27 olika återhämtningsplaner inte kommer att leda till de resultat som behövs under de kommande åren.
Det är helt nödvändigt att rådet och kommissionen tillsammans tar ledningen i detta.
Jag vet att det nu finns 27 återhämtningsplaner på nationell nivå men vi ser ett antal protektionistiska åtgärder inom dessa nationella planer.
Det är ert ansvar, herr Reinfeldt, att säga till era kolleger att ett bättre sätt att hantera detta är att tillsammans med kommissionen utarbeta en enhetlig återhämtningsplan och att investera i hållbar energi och i den nya ekonomin.
Med er erfarenhet från Sverige under 1990-talet är ni rätt man på rätt plats för att göra det som vi hittills inte har gjort, det vill säga att utarbeta en enhetlig EU-strategi för att bekämpa denna ekonomiska och finansiella kris.
(Applåder)
för Verts/ALE-gruppen. - (DE) Herr talman, herr Reinfeldt, herr Barroso! Min kollega Martin Schulz sade allt som finns att säga om de institutionella betänkligheter som min grupp länge har haft när det gäller det kommande valet av kommissionens ordförande.
Vi instämmer i vad han sade.
Vi vill att hela kommissionen och all personal på hög nivå inom EU ska väljas enligt villkoren i Lissabonfördraget och vi kommer inte att vika en tum på denna punkt.
Emellertid, herr Barroso, vill jag passa på att förklara de politiska skälen bakom min grupps tvivel och dess åsikt att ni ur politisk synvinkel inte är kapabel att göra vad som krävs i den aktuella situationen i EU.
Ta till exempel det ofta nämnda behovet av en ny reglering av finansmarknaderna.
Vi har haft G8-toppmöten, G20-toppmöten, förlängda G8-toppmöten, EU-toppmöten.
Hur långt har vi kommit?
Vi kan se på var vi står i dag och jämföra med monopolspelet, som vi alla känner till. Bankerna har återupprättats, de har passerat ”gå” och kom inte i fängelse, de har tagit hundratals miljoner med offentligt godkännande och började sedan helt enkelt spela från början.
Jag tror inte att folk är domedagsprofeter när de menar att nästa krasch blir oundviklig som en följd av detta.
Herr Barroso! Vad hände med er kraftfulla insats?
Var är era konkreta resultat?
Vi har inte sett något prov på dem.
(Applåder)
När det gäller klimatpolitiken, vet ni att vi inom gruppen De gröna/Europeiska fria alliansen under hela vår EU-kampanj har förespråkat en ”Green New Deal”.
Vi är fullständigt övertygade om att det är helt fel att göra som ni upprepade gånger har gjort under de gångna fem åren, nämligen att spela ut ekonomiska strategier mot miljö- och klimatstrategier.
Vi anser att detta verkligen hör hemma i det förgångna och att det måste upphöra.
Vi måste tänka på ekonomisk utveckling på ett hållbart sätt och vi måste se till att klimatskyddsmålen är anpassade till miljömålen.
Detta kommer att gynna ekonomin och det kommer att skapa tusentals eller till och med miljontals arbetstillfällen.
Andris Piebalgs har än en gång, i sin undersökning under de senaste månaderna, visat att detta gäller för energisektorn.
Enligt vår erfarenhet har ni inte förutsättningar att kunna utveckla denna ”Green New Deal”.
Sammanfattningsvis kan jag bara säga att européerna under de senaste månaderna har haft en framträdande plats på den internationella arenan, i frågan om klimatskyddet. En anledning är att de har börjat tveka - hur långt vill vi egentligen gå med minskningsmålen?
En annan anledning är också deras nya snålhet och detta gäller tyvärr också Sverige.
Inrättandet av den internationella klimatskyddsfonden för de fattigare länderna har gått extremt dåligt. Det är fortfarande en hemlighet att Sverige vill ta pengar från utvecklingsmedlen, bland annat, för att använda för detta klimatskydd.
Det är ett nollsummespel och ur de fattigare ländernas synvinkel är det totalt oacceptabelt. Vi måste snabbt komma till rätta med denna nya snålhet och tvekan inom EU.
(Applåder)
Slutligen, herr Reinfeldt, kan jag säga något positivt.
Vi är beredda att kämpa tillsammans med er om den nya definitionen av Lissabonstrategin och att samarbeta med er om detta.
Ni har sagt att ni kommer att göra detta innan året är slut.
Vi ska hjälpa er med detta.
Vi kommer också att stödja er om ni vill göra mer när det gäller Östeuropa och Ryssland, men inriktningen för en verklig klimatpolitik får inte bara vara en fråga om rubriker, det måste också korrigeras i den finstilta delen av Sveriges program.
(Applåder)
Herr talman! Först vill jag uppriktigt gratulera till gårdagens val, valet av en utmärkt talman - parlamentets nye ledare.
Ni vet mycket väl att jag gör det som polsk politiker men också som privatperson.
Som ni vet var det tack vare er som jag träffade min fru och det är ändå det viktigaste som hänt mig i mitt liv.
Jag gratulerar och önskar er stor framgång i ert arbete.
Gruppen Europeiska konservativa och reformister lyssnade noga till ert tal, herr statsminister, och jag är glad över att kunna säga att vi delar era synpunkter i väldigt många frågor.
Särskilt viktigt är ert tillkännagivande av aktiva åtgärder för att hantera krisen.
Den ekonomiska krisen, som är den värsta kris som vår civilisation har upplevt sedan 1930-talet, skapar obefogad ängslan i hela Europa - i fattigare länder och i rikare, i länder i norr och i söder.
Jag är glad över att ni har tillkännagett en aktiv kamp mot krisen och jag är glad över att ni kan se prioriteringar som vi också delar - större frihet för marknaden, mindre reglering, större ekonomisk frihet, större öppenhet för frihandel.
Det handlar här om recept på ekonomisk tillväxt för vår världsdel, för vårt EU.
Vi delar också er övertygelse om att hanteringen av klimatförändringarna är en viktig fråga.
Jag vet att ni har djärva åsikter i denna fråga och jag vill uppmuntra er att vara djärv på detta område.
Klimatförändringsfrågan visar mycket tydligt att vi i dag inte bara lever i ett enhetligt EU utan också i en enhetlig värld där hoten är gemensamma för alla och måste hanteras effektivt.
Jag är mycket glad över att ni tog upp kampen mot brottsligheten som ett allvarligt problem i EU.
Då Sverige redan är en betydande kraft när det gäller deckarromaner, är jag övertygad om att vi under er ledning också kommer att kunna bekämpa brottsligheten med framgång.
Det är ytterst viktigt och jag är glad över att både ni och er utrikesminister nyligen har nämnt att ni vill vända blicken mot våra grannländer och ha vad jag hoppas kommer att bli en välvillig syn på EU:s utvidgning.
Vi får inte glömma att det på andra sidan av EU:s östra gränser finns länder som har rätt till att vara en del av det område av demokrati och välstånd som vi i dag är en del av.
Jag måste tyvärr säga att det finns en punkt där min grupp inte är överens med er.
Detta rör frågan om ratificeringen av Lissabonfördraget.
Ni talade om demokrati i samband med Lissabonfördraget och det gjorde ni rätt i.
Man bör komma ihåg att det var i en demokratisk folkomröstning som irländarna förkastade Lissabonfördraget.
Eftersom vi har respekt för demokratin bör vi respektera irländarnas röst.
Herr statsminister! Jag hoppas att era prioriteringar, som i mycket stor utsträckning delas av ECR-gruppen, kommer att göra det möjligt för er att effektivt leda EU och att effektivt hantera den kris som i dag är vårt största problem.
(Applåder)
för GUE/NGL-gruppen. - (DE) Herr talman, statsminister Reinfeldt, mina damer och herrar! Det svenska ordförandeskapet har lagt fram ett ambitiöst arbetsprogram som inkluderar ett förslag om större öppenhet.
Öppenhet krävs särskilt när man bekämpar den kris som vi för närvarande genomgår.
Många tror att krisen har orsakats långt borta i USA, av några bankdirektörer som sägs vara giriga.
EU-medlemsstaternas regeringschefer verkar inte ha haft något att göra med krisen.
De är oskyldiga i sammanhanget.
De som gottar sig åt att vara oskyldiga gör inget för att bekämpa krisen.
Jag anser att öppenheten också bör handla om att man talar om de politiska misslyckanden som bidrog till krisen och även om bankdirektörer, givetvis.
Öppenhet är modernt i kasinokapitalismen.
Vi är ivriga att se vad som sker med Östersjöstrategin och jag ställer mig bakom rådsordföranden om han väljer att fokusera på dialog med Ryssland.
Vi vill också att EU stöder president Barack Obamas och president Dmitrij Medvedevs utfästelser om kärnvapennedrustning.
EU bör dra nytta av denna nya möjlighet till nedrustning.
Det svenska ordförandeskapet vill ytterligare harmonisera asylrätten och göra EU mer attraktivt för migrerande arbetstagare.
Asylpolitiken ska vara nära kopplad till utvecklingspolitiken.
Detta är bra enligt vårt synsätt, men vid EU:s rigoröst vaktade yttre gränser, särskilt vid Medelhavet, dör tusentals människor varje år när de söker en fristad från förföljelse, fattigdom, naturkatastrofer och krig.
Trots kostsamma gränskontroller och övervaknings- och datainsamlingssystem för att förhindra olaglig invandring, efterlyser gruppen Europeiska enade vänstern/Nordisk grön vänster en mänsklig behandling av flyktingar och invandrare och en förändring i ekonomi- och handelspolitiken för att effektivt bekämpa de faktorer som får folk att bli flyktingar över huvud taget.
Det svenska ordförandeskapet fokuserar på mer inkluderande arbetsmarknader för att skapa full sysselsättning och vill därför inleda reformer av arbetsmarknaden och vidta åtgärder för jämställdhet mellan könen.
Också vi är positiva till en strategi för goda arbetsrutiner, där man kommer att stödja löneökningar och införa en lagstadgad minimilön för alla i de 27 medlemsstaterna.
Vi vill se att EU enas om mål för minimilönen som uppgår till minst 60 procent av den nationella genomsnittslönen, för att förhindra att folk hamnar i fattigdom trots att de har ett inkomstbringande arbete.
Jag välkomnar särskilt vad ni sade om Cypern och jag önskar er all framgång i genomförandet av era ambitiösa klimatmål.
Herr talman, mina damer och herrar! Jag uppskattade att det svenska ordförandeskapet betonade frågor som berör medborgarna, våra väljare, nämligen miljön och klimatförändringarna, finanskrisen, bevarandet av arbetstillfällen och kampen mot brottslighet.
För att göra ett bra arbete måste vi vara i harmoni med dem som röstade för oss. Vi är vare sig bättre eller sämre än våra väljare men jag menar att det är viktigt att agera i enlighet med deras önskemål och dessa punkter verkar vara i linje med vad jag nämnde.
När vi går vidare måste vi naturligtvis omsätta förslagen i konkreta åtgärder och här kommer vi att konfrontera varandra framför allt i medbeslutandeförfarandet, eftersom vi i parlamentet och ni i rådet ska fastställa de regler som kommer att styra våra väljares liv, angelägenheter och intressen. Jag anser att det är vår grundläggande uppgift som lagstiftare.
Vi måste övervinna den förtroendekris som utan tvekan finns.
Den dåliga uppslutningen vid valet till Europaparlamentet är en följd av denna kris, och för att lösa detta problem måste vi agera helt enligt våra väljares vilja. Vi kanske också måste undvika att göra jämförelser.
Jag bor nära Schweiz. De ligger utanför EU men de mår bra ändå.
De har samma problem, men de har det inte sämre än vi. Här är det viktigt att inse och visa att EU är något värdefullt.
Jag ser detta som en stor utmaning, men jag tror samtidigt att vi med allas hjälp kan visa att EU inte är något som ska uthärdas utan att det bör vara en möjlighet för befolkningen och medborgarna.
(NL) Det nederländska frihetspartiet har kommit in i Europaparlamentet för att kämpa för nederländska medborgare och för att ta tillbaka det alltför höga belopp som Nederländerna har betalat till detta pengafrossande och byråkratiska EU.
Frihetspartiet valdes in i Europaparlamentet av nederländska väljare för att tydliggöra de nederländska medborgarnas åsikt att EU:s utvidgning redan har gått för långt.
Herr talman! Europaparlamentet ägnar sin tid åt att reglera frågor som bör avgöras i medlemsstaterna.
Vårt parti anser att EU bara bör ägna sig åt frågor som gäller ekonomiskt och monetärt samarbete.
Det är med nederländska intressen i tankarna som vi kommer att hålla ögonen på det svenska ordförandeskapet, eftersom det inte gör något för de nederländska medborgarna.
Ni vill bara gå vidare med EU-konstitutionen, som nederländska väljare förkastade och som är till 99 procent identisk med Lissabonfördraget.
Ni gör heller inget åt den oerhört dyra förflyttningen varje månad från Bryssel till Strasbourg.
Ni har inte ens satt upp frågan på dagordningen.
Varför inte?
Det kostar tusentals miljoner euro och de enda som uppskattar detta är kanske de på IKEA, som får en chans att sälja flyttlådor och extra skåp.
Vi vill också att förhandlingarna med Turkiet omedelbart upphör.
Turkiet är ett muslimskt land och den muslimska ideologin står helt i strid med vår västerländska kultur.
Dessutom är Turkiet inte alls ett europeiskt land utan ett asiatiskt land, och Turkiets medlemskap skulle än en gång kosta de nederländska medborgarna en massa pengar.
Turkiet kan vara en bra granne men det hör inte hemma inom den europeiska familjen.
Frihetspartiet står för ett EU med självständiga stater, men det som sker under det svenska ordförandeskapet är ytterligare steg mot en federal superstat där medlemsstaterna får bestämma mindre och mindre över sina egna frågor.
Därför hoppas vi att irländarna kommer att ha mod nog att åter rösta nej till Lissabonfördraget.
Irlands befolkning har nu möjlighet att agera som en röst för EU:s befolkning.
rådets ordförande. - Herr talman! Låt mig först gratulera er alla kollektivt till att ha blivit valda till gruppledare.
Jag vet att flera av er har blivit valda med mycket starkt stöd.
Jag vet t.ex. att Martin Schulz blev omvald med mycket starkt stöd i den socialdemokratiska gruppen.
Det är viktigt att starkt kunna representera sina respektive grupper.
Jag har väldigt mycket välkomnat den dialog som vi har haft och de konsultationer som jag fick i uppgift av Europeiska rådet under junimötet att inleda.
Det har gjorts av EU-minister Cecilia Malmström.
Det har också gjorts av mig själv både i telefonkontakter och också vid det möte som vi hade på en skärgårdsbåt när vi rörde oss genom vatten i Stockholm och då satt och diskuterade den uppkomna situationen.
Jag hade fått i uppdrag att undersöka möjligheten att välja José Manuel Barroso, utpekad av Europeiska rådet, till kommissionens ordförande för en andra mandatperiod.
Flera av de frågor som ni berörde är de huvudfrågor som vi vill arbeta med under det svenska ordförandeskapet.
Låt mig säga att vi sätter jobben främst.
Vi vill se ett Europa där fler får arbete.
Diskussionen måste utgå från hur man åstadkommer det.
Jag tror precis som Joseph Daul påpekade att det handlar om innovation och utbildning, dvs. det som i grunden driver företagandet och möjliggör anställningsbarhet.
Jag tror att Martin Schulz har rätt i att vi ska akta oss för att få ett Europa där vi konkurrerar med dåliga villkor.
Den diskussionen har vi i Sverige, och den har vi runtom i Europa.
Det är ingen bra utgångspunkt att försöka möta konkurrens med att ha låg eller ingen lön, utan det är med bra villkor som vi vill möta framtida konkurrens.
Låt mig nämna några andra saker som jag ser som mycket viktiga för att styra Europa genom krisen.
Jag har sett hur kommissionen - och tycker själv att det är viktigt - har fått försvara den inre marknadens princip i en tid då många försöker rucka på den och få in protektionism.
Det är så lätt att lyssna till dem som säger ”Varför räddade ni inte jobben i just det här landet?”, utan att se konsekvenser av om alla skulle agera likadant.
Då skulle vi i grunden släcka ner frihandeln och möjligheten att ha gränsöverskridande handel.
Det som i grunden har skapat rikedom och välstånd skulle mycket snabbt gå förlorat om vi inte på detta sätt har stått emot ropen på protektionism.
Att slå vakt om den inre marknaden och den fria rörligheten tror jag är en viktig utgångspunkt för att säkerställa jobben.
Jag tror också mycket på det som har nämnts av flera av er, t.ex. att investera i människors kunskaper och säkerställa att det finns rörlighet i arbetsmarknaden.
Jag tror exempelvis att just den fria rörligheten, också över gränser, är ett sätt att hantera det.
Jag tror precis som Martin Schultz, Rebecca Harms och Joseph Daul nämnde att det här också är tillfället att möta detta med en grön utveckling, att få fram de lågutsläppsekonomier som vi talar om världen över som ett sätt att också komma ur krisen.
Det är viktigt hur vi styr finansiering och hur vi investerar.
Jag vill också säga - jag håller med Guy Verhofstadt på den punkten - att våra svenska erfarenheter av vår krishantering under 90-talet var att inte tro att detta på ett bra sätt blandar sig med att tappa greppet om de offentliga finanserna.
Jag har lärt mig att när underskotten blir stora och när det ska saneras är det människor med små marginaler och de som är mest beroende av välfärdsinstitutioner som får stå tillbaka.
Därför är en politik som är aktsam om de offentliga finanserna en bra politik för människor som är fattiga eller som lever med små marginaler.
När det gäller klimatfrågan, som kommer vara vår huvudfråga att arbeta med inför Köpenhamnstoppmötet, vill jag säga att det stämmer att det finns mycket kvar att göra.
Tiden är knapp.
Jag vill säga till Rebecca Harms att det är ovanligt att vi i Sverige får kritik för våra biståndsåtaganden.
I Europa går i genomsnitt 0,4 procent av bruttonationalinkomsten till sådana åtaganden.
Sverige är ganska unikt på så sätt att en procent av vår bruttonationalinkomst går till utvecklingsstöd.
För mig hänger dessa frågor ihop.
Vi har haft en egen genomgång under ledning av vår biståndsminister inom ramen för FN:s insatser.
Vi har då analyserat just hur vi måste tänka klimatomställning i vårt utvecklingsarbete.
Det går inte att bedriva utvecklingsinsatser om man inte samtidigt ser klimatomställningen och hur den redan påverkar fattiga delar av vår jord.
Därför kan vi inte separera och säga att här är utvecklingspolitiken och där borta är klimatpolitiken, utan de hänger ihop och måste samverka.
När det gäller fördraget och till Martin Schulz vill jag säga att min roll är att se till att det finns ett fungerande europeiskt ledarskap i en svår tid.
Vi måste kunna leverera svar till de medborgare som vill se oss agera mot finanskris och i klimatfrågor.
Vi är alla politiskt verksamma och vet att i den politiska miljön, där vi blir inåtblickande och diskuterar namn och ledarskap, så uppfattar våra medborgare det som om vi har vänt ryggen mot dem.
Vi tittar inåt.
Därför gör jag vad jag kan i min roll.
Jag har i uppdrag från Europeiska rådet att säkerställa att vårt samarbete och vår respekt för den integritet som finns hos Europaparlamentet förenas av att vi är tydliga - det gäller både i form av Nice- och Lissabonfördrag - och nominerar en kandidat till posten som kommissionens ordförande.
När det gäller José Manuel Barroso är det viktigt att konstatera att han hade ett enhälligt stöd i Europeiska rådet, att han var välkänd som kandidat och presenterad för väljarna redan före valet.
Det gjorde det naturligtvis enklare för mig att agera - naturligtvis med respekt för att Europaparlamentet kommer att få tillfälle, när ni anser er vara redo att fatta beslut, att säga ja eller nej till den nominerade kandidaten från Europeiska rådet.
Under tiden finns det tid för diskussioner, vilket jag vet att även José Manuel Barroso har förklarat, och för att föra den typ av samtal om hur den europeiska politiken ska utvecklas under de kommande åren.
Jag hoppas att detta nu ska kunna gå att förena enligt den överenskommelse som har slutits.
Det är vad Europas väljare nu förväntar sig, och därmed kan vi agera starkt tillsammans.
kommissionens ordförande. - (FR) Herr talman! Några viktiga frågor har ställts.
För det första Martin Schulz' viktiga fråga angående fördragen.
Han berörde särskilt kommissionens roll som fördragens väktare.
Vi i kommissionen anser att de gällande fördragen bör respekteras.
Det gällande fördraget är Nicefördraget.
Alla ni som sitter här valdes enligt Nicefördraget.
Om kommissionens ordförande väljs nu kommer han naturligtvis att väljas liksom er, enligt Nicefördraget.
Med detta sagt hoppas jag att vi kommer att få Lissabonfördraget.
De nödvändiga anpassningarna kommer att behöva göras när det gäller parlamentets sammansättning, som inte längre kommer att vara densamma med Lissabonfördraget, eftersom det kommer att bli vissa förändringar, och samma sak kommer att behöva göras med kommissionen.
Inte desto mindre följde Europeiska rådet alla aspekter av ert betänkande - Jean-Luc Dehaenes betänkande - som antogs med en överväldigande majoritet.
Innan Europeiska rådet formaliserade sitt beslut genomförde det samråd, där man också - för första gången - beaktade resultatet i valet till Europaparlamentet, för att inte nämna att det hade varit en kandidat som stöddes av en politisk kraft.
Uppgiften är nu att få Europaparlamentets godkännande.
Jag vill i dag upprepa vad jag redan har uppgett i en skrivelse till Europaparlamentets talman. Jag är redo att diskutera innehållet i riktlinjerna för nästa kommission med alla politiska grupper som vill diskutera dem.
I vilket fall som helst är detta är min hållning i de institutionella frågorna.
På ett politiskt plan vill jag betona en mycket viktig punkt.
Jag ser det som viktigt att koppla valet av kommissionens ordförande till det demokratiska val som har ägt rum, ert val.
Ni har valts genom Nicefördraget och det är min åsikt att kommissionens ordförande också bör ha denna legitimitet, vilket på sätt och vis bör vara en följd av detta demokratiska val.
Mot bakgrund av den ekonomiska och finansiella krisen - och jag tror absolut att de som är för ett starkt EU och en stark kommission kommer att instämma - bör frågan om kommissionens ordförande inte lämnas olöst i väntan på den slutliga ratificeringen av Lissabonfördraget, som vi alla vill ha - åtminstone en majoritet av oss - eftersom vi inte vet när detta fördrag kommer att träda i kraft.
Att lämna Europeiska kommissionen och dess ordförandeskap i ett tillstånd av ovisshet under en ekonomisk kris, en finansiell kris och en social kris, då vi har mycket viktiga förhandlingar framför oss i Köpenhamn, förefaller inte vara särskilt klokt.
Hur som helst är det upp till Europaparlamentet att fatta beslut och jag är redo att delta i en demokratisk debatt såsom jag faktiskt gjorde för fem år sedan.
(EN) På den andra frågan om finans och ekonomi och med tanke på vad Guy Verhofstadt sade kan vi alla ha högre ambitioner. I denna fråga delar jag er ambition.
Men vi kan inte säga att vi inte antog någon europeisk ekonomisk återhämtningsplan, och det var vad medlemsstaterna maximalt accepterade.
Kommissionen föreslog mer, men detta var vad våra medlemsstater accepterade.
Jag vill uppmärksamma er på att vissa medlemsstater - som inte var mindre inflytelserika i den begynnande krisen - föreslog att vi inte skulle ha någon samordningsplan alls.
Andra medlemsstater föreslog en finanspolitisk stimulans på 1 procent, kommissionen kom omedelbart med förslaget på 1,5 procent och de automatiska stabilisatorerna var i realiteten på omkring 5 procent.
Frånsett detta fattade vi dessa viktiga beslut om betalningsbalansstöd till vissa medlemsstater som inte ingår i euroområdet och även om vissa initiativ på global nivå.
Så ni kan räkna med att kommissionen gör allt den kan för att främja EU-nivån och en gemensam strategi. Det får inte råda några tvivel om detta.
Men låt oss samtidigt vara ärliga mot oss själva. Vi är inte Förenta staterna - vi är inte en integrerad nationalstat - så naturligtvis har vi olika situationer.
Man kan inte begära att Tyskland och Lettland ska göra samma sak.
Vi har länder i EU som mottar betalningsbalansstöd, så naturligtvis kan vi inte ha en strategi som passar för alla.
Vi måste ha en gemensam strategi men med specifika nationella svar eftersom det är den verklighet som vi står inför i EU och som vi kommer att stå inför i framtiden.
Vi har i huvudsak nationella budgetar.
Så jag delar ert synsätt om att ha en mer samordnad europeisk plan för att komma ur denna kris och skapa den typ av smarta miljövänliga tillväxt som vi vill ha. Men samtidigt måste vi acceptera att vi har 27 olika nationella budgetar, vi har 27 finansministrar, vi har 27 nationella banker utöver vår Europeiska centralbank och det är mycket viktigt att stärka euron och att föra en hållbar ekonomisk och finansiell politik.
Om inte kommer vi att utsätta euron, en av den euroepiska integrationens största framgångar, för risker.
Slutligen, i fråga om klimatförändringarna kan vi än en gång alltid ha högre ambitioner.
Men för mig var det mycket viktigt att statsminister Fredrik Reinfeldt var med mig nyligen i L'Aquila, när vi hörde FN:s generalsekreterare säga: ”Ni är ett lokomotiv för världen”.
Vi kan alltid ha högre ambitioner, men EU leder kampen mot klimatförändringarna i världen.
Ingen är mer ambitiös än vi, så visst skulle jag åtminstone förvänta mig ett ord av erkännande för det arbete som kommissionen har gjort, tillsammans med våra medlemsstater, för att lägga fram ambitiösa förslag.
Låt oss nu försöka övertyga andra, eftersom vi behöver andra, eftersom problemet med klimatförändringarna inte bara är ett europeiskt problem, utan ett problem för hela vår jord.
Med ert stöd tror jag att vi kan uppnå goda resultat vid Köpenhamnskonferensen.
(Applåder)
Herr talman! Som svensk är det med stolthet som jag lyssnar på det svenska ordförandeskapets prioriteringar och dessutom kan hälsa Sveriges statsminister välkommen tillbaka hit än en gång.
De utmaningar vi har är rätt betydande.
Vi har 20 år av fantastisk mirakulös omvandling av Europa bakom oss, som har lett till att vi idag har en av de tidiga företrädarna för frihetsrörelsen Solidaritet som talman för Europaparlamentet.
Det är ideal som demokrati, frihet, rättsstat, marknadsekonomi som har gett oss 20 år av fantastisk utveckling.
Nu lever vi i en ny omvandlingens tid med ett nytt fördrag, klimatfrågan som ställer krav på en konsekvent politik som kan ha global genomslagskraft och den ekonomiska krisen.
Då är det viktigt att vi har ett ordförandeskap, men också ett parlament, som är förmöget att se till att vi får stabilitet när det gäller offentliga finanser, stabilitet när det gäller den inre marknaden och stabilitet när det gäller öppenhet för handel och rörelse över gränserna som kan bidra till att få oss ut ur krisen.
Jag skulle vilja sätta perspektivet ytterligare ett steg framåt.
De beslut som vi nu lägger grunden för genom det svenska ordförandeskapet och i detta parlament kommer också att avgöra hur Europa och Europeiska unionen kommer att se ut efter krisen - vilken dynamik vi kommer att ha på de finansiella marknaderna och vilket förtroende och trovärdighet de kommer att ha och vilket utrymme vi kommer att ha för innovation och företagande, för investeringar och nya jobb.
Om det var en sak som valet till Europaparlamentet visade så är det att Europas medborgare vill ha mindre byråkrati och regleringar och mer öppenhet - över gränserna och ut gentemot världen.
Det är den öppenheten som kommer att vara avgörande för Europas förmåga att vara en ledande kraft för de värden som för 20 år sedan började omvandla Europa och som vi kan bidra till i världen med.
(Applåder)
Herr talman! Jag vill först tacka den svenske statsministern för presentationen av vad han och hans regering vill göra under det närmaste halvåret.
Vi vet att utgångsläget är tufft, krisen är djup.
Det handlar om jobben, det handlar om dramatiskt växande klyftor, det handlar om en ungdomsgeneration som går rakt ut i arbetslöshet och det handlar förstås om miljö- och klimatkrisen.
Det här har också beskrivits av statsminister Fredrik Reinfeldt, men det som överraskar är slutsatserna.
Det som lyfts fram som den centrala frågan för det svenska ordförandeskapet är inte jobb eller investeringar, utan medlemsländernas förmåga att upprätthålla budgetdisciplin.
På väg mot 27 miljoner öppet arbetslösa i EU så är det alltså det tydligaste beskedet från det svenska ordförandeskapet: budgetdisciplin.
Det är illa, och också oroande.
Här har Reinfeldts parti - i motsats till vad som tidigare sagts här - ett historiskt inrikespolitiskt tungt bagage att bära på.
Den förra konservativa svenska regeringen ledde Sverige in i ett ekonomiskt sönderfall, och det var en socialdemokratisk regering som fick ägna tio år till att sanera de offentliga finanserna.
Men gamla inrikespolitiska tillkortakommanden kan ju inte få bestämma dagordningen för hela EU i ett läge när vi befinner oss i allvarlig kris.
Det som krävs är stora investeringar i jobb, utbildning och grön omställning, inte att man med budgetdisciplin sätter anorektiska ekonomier på svältkur.
Europafackets generalsekreterare John Monks har också uttryckt oro över att den sociala dimensionen i det svenska ordförandeskapet är så lågt prioriterad.
Mest vackra ord, säger Monks, väldigt lite av reella planer.
Vi känner samma oro i min partigrupp och det omfattar också löntagarnas fackliga rättigheter, som Martin Schulz redogjorde för i sitt inlägg.
Efter Lavaldomen och efter Viking-, Rüffert- och Luxemburgdomarna så har löntagarnas villkor försämrats.
Deras rättigheter har försvagats.
Vad jag och min grupp vill ha från det svenska ordförandeskapet är ett konkret åtagande om att EU:s löntagare ska få sina fulla fackliga rättigheter tillbaka.
De fackliga rättigheterna måste gå före den fria rörligheten.
Det måste vara väldigt tydligt.
Vi vill inte leva i ett Europa där krisen möts med budgetdisciplin och med konfrontation.
Står denna fråga på dagordningen över huvud taget, vill jag fråga den nye ordföranden, statsminister Fredrik Reinfeldt.
(FR) Herr talman! Vi står inför två frågor.
Den första frågan är krisen.
Som alla vet behöver vi ett konsekvent och gemensamt svar på den ekonomiska och sociala krisen, det vill säga en europeisk återhämtningsplan för att öka investeringarna och främja sysselsättningen.
I dag måste EU verkligen visa att det är mer uppmärksamt och närmare våra medborgare när det gäller deras problem.
EU måste göra mer för att hjälpa dem som drabbas av krisen.
I detta perspektiv är situationen brådskande.
Den andra frågan handlar om den nya utvecklingsmodell som måste komma efter krisen.
Det måste vara en enklare, mer rättvis och mer hållbar modell, där vi ser till att finansen tjänar realekonomin, utvecklar nya former av solidaritet mellan européerna, tar hänsyn till de sociala och miljömässiga utmaningarna i den internationella handeln och radikalt reformerar våra förbindelser med världens fattigaste länder, och här tänker jag särskilt på Afrika.
Utöver dessa båda viktiga frågor finns det ett demokratiskt krav som gäller den process där ni, det svenska ordförandeskapet, har ansvaret.
Cecilia Malmström - som jag är glad över att välkomna i dag - vet bättre än någon annan att det finns vissa betydande skillnader mellan Nicefördraget och Lissabonfördraget i fråga om utnämningsförfarandet: enkel majoritet å ena sidan och kvalificerad majoritet å andra sidan, en utnämning å ena sidan och en nominering å andra sidan, samt ett annat antal kommissionsledamöter beroende på fördrag.
För min del ber jag er verkligen att se till att fördragens anda och ordalydelse respekteras.
Detta faller inom ert behörighetsområde och det är mycket viktigt för våra institutioners trovärdighet.
Tack på förhand.
Herr talman! Gratulationer till er utnämning!
Jag vill först berömma regeringen för att ni har ett ärligt engagemang för Östersjön och där hoppas jag att vi kommer vidare.
Ni har också en förvånansvärt bra klimatretorik.
Vad jag nu efterlyser är givetvis klimatpraktik också.
Ni talar ofta om att Europa och Sverige står för en liten andel av jordens utsläpp, men om vi bara är åtta procent av jordens befolkning i EU-länderna, och släpper ut 30 procent, då är det också vårt ansvar att ta en stor del av klimatarbetet på allvar.
Det är här jag saknar de konkreta frågorna.
Hur går ni vidare med IPPC-direktivet om industriella utsläpp?
Hur går ni vidare med illegal avverkning?
Hur går ni vidare med energieffektivitetsnormer för byggnader och hur går ni vidare med att flyget inte kan fortsätta att släppa ut och slippa betala de 14 miljarder euro i energiskatt som de borde betala?
Sen vill jag också ta upp Stockholmsprogrammet och Acta.
Beträffande Acta måste se till att här blir öppenhet.
Tyska författningsdomstolen har sagt att länderna måste få mer inflytande, att parlamenten måste få mer inflytande.
Vi behöver öppenhet i Acta-förhandlingarna.
Vi kan inte gå ensidigt mot övervakning.
Samma sak gäller min hemstad, och Stockholmsprogrammet.
Låt det bli ett namn som förknippas med EU:s övergång från terrorparanoia till mänskliga fri- och rättigheter och med att asylrätten förstärks och integriteten skyddas.
Då har vi nått framgång med det.
(EN) Herr talman! Jag vill gratulera det svenska ordförandeskapet för att det prioriterar de ekonomiska utmaningarna.
När vi har en ekonomisk osäkerhet är vår förmåga att möta andra utmaningar uppenbart försvagad.
Ni gör rätt i att prioritera behovet av att återupprätta de offentliga finanserna.
De ovanligt höga statsskulderna utgör stora och långsiktiga hot som kan kvarstå under många årtionden om vi inte tar itu med dem nu.
Men att återställa finansinstitutionernas hälsa är också väsentligt för att återupprätta konsumenternas förtroende och återställa den ekonomiska tillväxten, för att inte tala om skattebetalarnas pengar.
I samband med era prioriteringar tar ni upp vikten av tillsynssystem.
Jag skulle vilja tillägga att tydliga regler är avgörande.
Som vi alla vet är dessa industrier globala industrier.
Kapitalet, talangen och de enskilda företagen är mycket flytande.
De behöver fungerande och bestämda lagstiftningsprogram, prioritering av lagstiftningen och tillfredsställande samråd.
Jag välkomnar ert åtagande att arbeta parallellt med G20. Om vi kommer ur takt och går framåt på ett ensidigt sätt inom EU riskerar vi att inte bara att utsätta låntagare och investerare för en konkurrensnackdel utan också att industrier utlokaliserar sin verksamhet utanför ...
(Talmannen avbröt talaren.)
Herr talman! Först vill jag naturligtvis gratulera till talmansuppdraget och samtidigt tacka för de intressanta åsiktsutbyten vi hade under valperioden.
Herr statsminister och kolleger! Jag tackar för redogörelsen för ordförandeskapets program.
Jag är övertygad om att det svenska ordförandeskapet organisatoriskt kommer att bli en stor framgång och att det kommer att skötas alldeles utmärkt av den kompetenta svenska statsförvaltningen.
Politiskt delar jag naturligtvis ordförandeskapets uppfattning om de två stora kriserna - den ekonomiska krisen och klimatkrisen - och det är de prioriterade frågorna, självklart.
Men det jag saknar är en analys.
Den ekonomiska krisen och klimatkrisen är ingen förutbestämd ödesutveckling.
Kriserna har sin grund i politiskt fattade beslut.
Det är positivt för det innebär att vi också kan lösa kriserna genom politiska beslut, men jag saknar en annorlunda, förändrad politik från ordförandeskapet.
Det är samma ekonomiska politik som inte tar social hänsyn eller miljöhänsyn.
Det jag gemensamt med många av medborgarna saknar i programmet är löntagarnas rättigheter, som har fokuserats efter domarna i domstolen, och de sociala frågorna, där vi inte får några svar.
Inte heller den välkända, progressiva jämställdhetspolitiken har vi hört någonting om.
När det gäller Stockholmsprogrammet säger man att det ska skapa trygghet, men i praktiken är det ett kontrollsamhälle som växer fram, som hotar den personliga integriteten.
Vi kan aldrig acceptera inskränkningar i asylrätten eller att våra fri- och medborgerliga rättigheter inskränks i det här programmet.
Vi kräver en human asyl- och invandringspolitik.
(FI) Herr talman, mina damer och herrar! Sverige har alltid respekterat de mänskliga rättigheterna och demokratin.
För ett tag sedan röstade svenskarna mot euron och ni har respekterat det beslutet trots att ni själv var klart positiv till euron.
Därför är det ganska märkligt att Irland nu genast måste rösta igen om exakt samma fördrag.
Det nordiska och det svenska sättet innebär att man respekterar folkets röst.
Jag önskar er lycka och framgång i den utmaning som ni nu står inför.
Jag hoppas att ni kommer att respektera den nordiska demokratins värderingar när den är som bäst: inte genom tvång utan genom samarbete.
Jag är mycket glad över att ni nämnde Östersjön och jag stöder er till fullo i denna fråga.
Östersjön har svårigheter. Den dör och den måste räddas.
Den nordliga dimensionen har dock saknats i allt detta och jag hoppas att ni kommer att göra mycket för att främja den, trots att ni inte nämnde det.
(DE) Herr talman! Vi behöver en demokratisk revolution.
Vi behöver djärva demokrater och i denna nya period behöver vi brådskande ett spännande, demokratiskt och verkligt effektivt EU.
Kreativa konstnärer och i synnerhet frilandsskribenter kommer att spela en roll i fastställandet av värderingarna för detta nya EU.
Deras ocensurerade fantasi kommer att kunna stoppa tillbaka den byråkratiska ande som vill förstöra demokratin i sin flaska.
När allt kommer omkring är det spännande idéer som ligger till grund när sociala förändringar föds.
De som kan erbjuda hoppfulla visioner som låter dessa idéer komma in i folks medvetande - svenskarna har varit särskilt bra på detta tidigare och i detta avseende har jag det största förtroende för min tidigare kollega Cecilia Malmström - kan också väcka deras intresse för socialpolitiska frågor.
På detta sätt formulerade jag det avslutande stycket i min nya bok i början av den senaste valkampanjen, som förde med sig stora förändringar och som är kopplad till stora förhoppningar om att särskilt ni från Sverige med er goda demokratiska tradition och öppenhet nu kommer att uppmärksamma tidens tecken.
Vi står inte bara inför den ekonomiska krisen, och här har svenskarna visat sin skicklighet genom att i stor utsträckning undvika denna. Vi har också behövt hantera en relativt hotfull svängning till höger.
Därför tror jag fullt och fast att vi demokrater tillsammans måste stå upp för verklig öppenhet och särskilt måste vi vara samlade i kampen mot extremhögern.
(NL) Varmt tack för de ambitiösa planer som ni har lagt fram för de kommande sex månaderna.
Vi har höga förväntningar på er eftersom ni ända från början har ansetts försvara den europeiska integrationen och våra europeiska värderingar.
Det är viktigt att de lösningar som vi lägger fram och som ni arbetar med för att ta oss ur denna ekonomiska kris stärker vår sociala marknadsekonomi.
Det är också viktigt att dessa lösningar inte bara främjar våra medborgare i dag och i morgon, utan också sörjer för våra barns framtid.
Det är därför mycket viktigt att fortsätta utvecklingen mot en hållbar ekonomi och mot att förhindra klimatförändringarna.
Det är bra att ni prioriterar detta så pass högt i ert program.
Jag hoppas verkligen att era insatser på detta område bidrar till att få medlemsstaterna att närma sig varandra och att ni inför Köpenhamnskonferensen också lyckas få de största aktörerna på världsarenan att verkligen göra sitt för att hitta en lösning på klimatförändringarna.
Herr talman! Den sociala marknadsekonomin är också viktig när det gäller hållbara statsfinanser eftersom underskott i den offentliga sektorns finanser utgör en börda för kommande generationer.
Därför är det viktigt att respektera stabilitets- och tillväxtpakten och det är bra att ni har sagt detta uttryckligen.
Ironiskt nog har finanskrisen fört Island närmare EU.
Jag hoppas att det svenska ordförandeskapet är välkomnande mot Island men att det samtidigt också noga ser till att Island följer anslutningskraven och att landet uppfyller skyldigheterna i fråga om EU:s lagstiftning och skyldigheterna mot medlemsstaterna.
(DE) Herr talman, herr statsminister! Jag hoppas att ni i detta sammanhang låter mig tala särskilt till Carl Bildt, eftersom jag först av allt vill beröra ämnet utvidgning, särskilt när det gäller Balkan.
Ni nämnde att denna utvidgningsprocess kommer att bli långsammare än vad många på bägge sidor skulle ha önskat.
Det är dock mycket viktigt att ge tydliga signaler.
Jag förväntar mig att det svenska ordförandeskapet särskilt hjälper människorna i sydöstra Europa att övervinna de problem som de står inför där - inklusive mellanstatliga problem - så att de kan känna sig förhoppningsfulla över att vägen mot EU inte kommer att blockeras utan att framstegen kan fortsätta, även om det kanske tar lite längre tid.
Men dessa länder måste naturligtvis göra de förberedelser som krävs.
För det andra vill jag gärna beröra ett annat ämne som ni nämnde, nämligen frågan om ekonomisk omstrukturering och sammankopplingen av den ekonomiska politiken och miljön.
Det har redan sagts att ni har vårt fulla stöd i detta.
Jag anser att detta är en viktig uppgift för EU.
Det är sant att vi i detta avseende i stor utsträckning går i spetsen, men det finns fortfarande mycket kvar att göra.
Samtidigt ökar också arbetslösheten.
Arbetslösheten i EU har ännu inte nått sin högsta nivå.
Läget kommer tyvärr att försämras ytterligare.
Det är därför ytterst viktigt att nämna den andra dimensionen, den sociala dimensionen. Endast om folk känner att deras sociala behov och krav tas på allvar kan vi få ett brett stöd för den miljövänliga ekonomiska omstruktureringen.
Särskilt de nordiska länderna har många bra exempel på en aktiv arbetsmarknadspolitik.
Vi kan inte skapa arbetstillfällen, vare sig som EU eller som enskilda medlemsstater, men vi kan hjälpa folk som har förlorat jobbet att hitta jobb igen så snabbt som möjligt.
Det är vad vi avser med ett socialt Europa - denna aktiva arbetsmarknadspolitik som vi behöver i de enskilda medlemsstaterna, där EU och särskilt rådet måste sända ett tydligt budskap.
Den miljövänliga omstruktureringen av ekonomin kommer i slutändan att leda till lägre, inte högre, arbetslöshet.
Det är vad vi efterlyser.
Herr talman! Herr rådsordförande!
Gott att se er här! Utmaningarna är många i denna stormiga tid: en svår ekonomisk nedgång, osäkerheten kring Lissabonfördraget och förhandlingarna inför klimatmötet i Köpenhamn.
Ni har att göra.
Herr statsminister, några viktiga punkter.
Ni har också att övertyga era kolleger i rådet att protektionism är en styggelse.
EU:s styrka är öppna gränser och fri handel.
Statsstöd för att rädda bilindustrin är inte lösningen.
Finanskrisen pockar på en global nyordning, men regelverket måste vara balanserat utformat utan överreglering.
I höst, som några har sagt här, måste EU komma en bit närmare en anständig asylpolitik.
Energipolitiken, precis som några har sagt, kräver både realism och solidaritet.
Inga nya gaskriser, inget ensidigt beroende.
Internet var en viktig fråga i valrörelsen.
Sverige har här ett stort ansvar för att föra det s.k. Telekompaketet i hamn.
Rättssäkerheten ska gälla också i den virtuella världen.
Jag hade hoppats att parlamentet under denna session skulle godkänna utnämningen av José Manuel Barroso för en ny femårsperiod som ordförande för kommissionen.
Nu blir det inte så, det beklagar jag.
Nu är inte tid för EU att ägna sig åt institutionella maktstrider.
Nu är tid för politiskt ledarskap och handlingskraft.
Euron har visat sin styrka.
När tror statsministern att vi i Sverige är beredda att bli fullvärdiga EU-medlemmar och ha euron också i våra fickor?
Tack, och som vi säger i mitt parti: Lycka till!
(FI) Herr talman, mina damer och herrar! Sverige har nu ett enormt ansvar för mänsklighetens framtid.
Statsminister Reinfeldt! Ni talade med rätta om klimatkrisen.
Vi vet att den teknik som vi behöver under kommande årtionden finns och att den finns tillgänglig till ett rimligt pris, men den mest problematiska frågan är den oerhörda utmaning som klimatskyddet utgör för det mänskliga samarbetet.
Tyvärr liknar de förhandlingar som för närvarande pågår mer en kombination av kurragömma och en tävlig i självbelåtenhet.
EU måste våga lägga fram ett förslag som inte bara gäller EU:s egna utsläppsminskningar utan också principen om delade bördor, där alla industriländer uppnår minskade utsläpp enligt riktlinjerna från Mellanstatliga panelen för klimatförändringar (IPCC).
Det viktigaste är att vi uppnår målen för minskade utsläpp för 2020.
För det andra måste vi inse att utvecklingsländerna inte kommer att kunna anpassa sig till ett system med avpassade utsläppsgränser om vi inte stöder dem finansiellt på en helt ny nivå. EU bör kunna komma med förslag också om detta.
(PL) Herr statsminister! Vi lyssnade på ert tal med stor uppmärksamhet och hoppas att de viktigaste punkterna i programmet kommer att förverkligas på ett bra sätt.
Emellertid vill jag uppmärksamma tre utmaningar.
Den första av dessa är den europeiska solidariteten, som är särskilt viktig under en finanskris.
Vi kan inte tillåta att situationer uppstår där olika EU-länder inte behandlas likvärdigt.
Vi kan inte acceptera en situation där vissa länder tillåts subventionera sin banksektor medan andra fördöms för att de har försökt stärka sin varvsindustri.
Det är inte solidaritet, det är hyckleri.
För det andra är vi glada över att Östersjöstrategin är en av det svenska ordförandeskapets prioriteringar.
Det är ett viktigt område för det makroregionala samarbetet.
Östersjöns ekosystem bör skyddas från risker såsom det mycket riskabla och finansiellt orimliga Nord Stream-projektet.
Behovet av att diversifiera energikällorna bör också nämnas.
För det tredje, låt oss komma ihåg att Moskva inte inskränker sig till att vrida av kranen, vilket Georgien upptäckte.
När Sverige tar rodret för EU under de kommande sex månaderna hoppas jag att det kommer att vara lika beslutsamt som minister Carl Bildt, som fördömde det ryska angreppet mot Georgien.
Jag är säker på att det svenska ordförandeskapet kommer att kunna klara dessa utmaningar.
Det kan räkna med stöd från oss.
(DA) Herr talman! Två saker slog mig när jag läste det svenska ordförandeskapets arbetsprogram.
För det första alla löften om hur EU kommer att användas för att skapa en bättre ekonomi för att lösa klimatproblemen och andra problem, samtidigt som det inte sägs ett enda ord om de problem som EU skapar - de problem som EU har skapat på våra arbetsmarknader, de problem som EU har skapat inom vår fiskesektor, i vår ekonomi, i samband med kampen mot brottslighet ... Jag skulle kunna fortsätta.
Det är den första viktiga observation som vi kan göra när vi läser det svenska ordförandeskapets arbetsprogram - att EU bara företräder lösningar och att EU inte är ett problem.
Det säger mer om det svenska ordförandeskapet än det säger om EU.
För det andra nämns det inte att den 2 oktober kommer att vara en av de viktigaste dagarna i hela EU:s historia, och detta kommer att inträffa under Sveriges ordförandeskap.
Jag syftar naturligtvis på den andra folkomröstningen.
Det sägs inte ett ord om vad det svenska ordförandeskapet ska göra för att se till att de så kallade garantier som har getts till irländarna också kommer att betraktas som sådana.
Vi har tidigare sett hur folk har vilseletts - vilseletts i fråga om folkomröstningar och i fråga om demokratin.
Vad kommer det svenska ordförandeskapet göra för att se till att detta inte sker igen?
(DE) Herr talman, herr rådsordförande, herr kommissionsordförande! Jag välkomnar svenskarna och gratulerar dem till att de - som statsministern sade - slutligen har hittat fram till EU efter en lång process.
Vi är mycket nöjda över att se att svenskarna i dag är bland de bästa EU-medlemmarna.
Ni har presenterat ert program och det är mycket ambitiöst.
Emellertid vill jag be er överväga om Sverige skulle ha modet att ansluta sig till euron, särskilt efter erfarenheten med krisen på finansmarknaden och särskilt eftersom ni sade att stabilitets- och tillväxtpakten måste respekteras.
Ni har ju ingen undantagsklausul som till exempel Storbritannien och Danmark och ni uppfyller nu alla villkor.
Kommer ni att ha modet under ert ordförandeskap att stabilisera EU ytterligare och ansluta er till euroområdet?
Jag stöder er prioritering av klimatpolitiken och Östersjöstrategin, men när det gäller ert program i dess skriftliga form har jag en förfrågan. Var vänlig och lägg större omsorg är vad som har föreslagits på att bekämpa krisen på finansmarknaden.
Inget av de andra projekten kommer att ha en chans om krisen på finansmarknaden och inom ekonomin inte blir löst så snabbt som möjligt.
För detta behöver vi tydliga regler.
Det duger inte att City of London än en gång anger riktningen.
Vi behöver tydliga regler i den sociala marknadsekonomin, eftersom en marknadsekonomi utan regler inte kan fungera och inte kommer att få majoritetens stöd.
Därför bör ni än en gång överväga - fastän vi till fullo stöder ert program - huruvida ni inte bör ge frågan om att lösa krisen på finansmarknaden högre prioritet än vad ni hittills har gjort.
Tack så mycket och lycka till i en svår och omvälvande period.
(Applåder)
(ES) Herr talman, herr rådsordförande! Vi har alla lyssnat på det svenska ordförandeskapets program med stort intresse och stor uppskattning.
Dess tydliga prioriteringar är ekonomin och energin, eftersom EU:s prioritering är att bidra till en nystart för ekonomin, skapa sysselsättning, stävja arbetslösheten och se till att mötet i Köpenhamn i december 2009 blir en framgång.
Emellertid vill jag rikta uppmärksamheten mot ett politiskt, medborgerligt och demokratiskt mål som handlar om att ersätta Haagprogrammet med det program som ska uppkallas efter Sveriges huvudstad, Stockholm.
Programmet kombinerar det som uppnåtts på området frihet, säkerhet och rättvisa under de senaste fem åren, vilket har varit mycket betydande i termer av harmonisering, ömsesidigt erkännande samt principen om tillit i samband med grundläggande rättigheter och rättsligt skydd, men också i samband med aktivt samarbete.
Jag uppmanar er att vara ambitiös på detta område. Såsom inom alla områden som gäller förvaltningen av de yttre gränserna, invandring, asyl, flyktingar och kampen mot olaglig handel, organiserad brottslighet och terrorism, är det - när det gäller politikens innehåll - lätt att närma sig reaktionära synsätt som strider mot det regelverk av grundläggande rättigheter som bör särskilja EU och som Sverige identifierar sig med så mycket, i egenskap av ett land som respekterar öppenhet och demokratiska principer.
Jag uppmuntrar er att också vara ambitiösa när det gäller politikens form, eftersom det svenska ordförandeskapet med största sannolikhet kommer att bana väg för Lissabonfördraget, som för det första innebär att vi inte längre kommer att ha de dubbla procedurreglerna inom den tredje och den första pelaren, vilka ofta är förvirrande.
Viktigast av allt är dock att parlamentet därmed också kommer att ha större kapacitet att övervaka de lagstiftningsinitiativ som det svenska ordförandeskapet genomför som en del av Stockholmsprogrammet.
Detta innebär att vad som hittills ofta har setts som en brist hos Bryssel eller hos rådet också kommer att bli parlamentets ansvar.
Självklart är jag mycket glad och stolt över att se min regering i det svenska ordförandeskapet och jag tycker också att det i programmet finns mycket bra när det gäller lösning av klimatjobb, finanskrisen, Köpenhamnskonferensen, Östersjöstrategin, gemenskapspolitiken, utvidgningen, Island, Kroatien, Turkiet osv. Men jag tänkte att jag ser en annan fråga, en viktig framtidsfråga, dvs. det öppna Europa, integritet och yttrandefrihet.
I dag möts ministrarna i Stockholm för att diskutera Stockholmsprogrammet.
Det som är bra är att detta är strategin för den lagstiftning som nu ska utarbetas.
Det finns delar i förslagen som vi har längtat efter länge.
Det blir äntligen en ratificering, hoppas jag, av den europeiska konventionen om mänskliga rättigheter.
Barns rättigheter och brottsoffers rättigheter. Det går att göra något väldigt bra av detta, men det finns också nackdelar, nämligen det hot mot det öppna samhället som finns i Stockholmsprogrammet.
Hot mot det öppna samhället måste bekämpas med det öppna samhällets metoder.
Delar av det som finns i Stockholmsprogrammet är varken liberalt, humant eller framsynt.
Att registrera vårt resande, att masslagra personliga kännetecken och systematisk kartläggning av ekonomiska transaktioner är varken liberalt, tolerant eller framsynt.
Låt Stockholm stå för öppenhet, frihet och tolerans. Inte registrering, övervakning och intolerans.
För övrigt anser jag att vårt arbete i Strasbourg ska läggas ner.
Innan jag ger ordet till Theodor Stolojan vill jag välkomna en gäst, ett barn som sitter på stol 505.
Jag är särskilt glad över att se barn som visar intresse för EU-frågor och för våra institutioner. Det är viktigt att växa upp som europé från tidig ålder.
(RO) Jag önskar det svenska ordförandeskapet all framgång och jag anser att de prioriteringar som har beskrivits överensstämmer med våra förväntningar.
De kommande sex månaderna är avgörande för EU:s medborgare och för EU.
De är avgörande för om våra länder ska komma ur den ekonomiska krisen nästa år eller om ett stort frågetecken ska fortsätta hänga över ekonomin i ett år till.
Många förslag och nya program läggs fram.
Jag anser dock att det är dags för oss att bedöma vilken inverkan det ekonomiska återhämtningsprogram som lanserades av kommissionen i början av året har, om det har någon inverkan alls, och ta en nära titt på EU:s budget för detta år för att se vilka verksamheter som har upphört och vilka resurser som vi kan fortsätta att använda för att komma med nya åtgärder.
Vi har också planerade investeringsprojekt för energisektorn som redan har godkänts från detta belopp på omkring 3 miljarder euro.
Vi kommer att behöva vidta särskilda åtgärder för att genomföra dessa projekt.
Jag vill tacka ordförande José Manuel Barroso för hans särskilda bidrag för att Nabucco-projektet skulle komma igång.
Slutligen skulle jag vilja att ni kommer ihåg EU:s politiska åtagande för att andra länder också ska kunna ansluta sig till EU.
(EN) Herr talman! Vi kommer inte att ta oss ur den djupa kris som drabbat finansmarknaden, ekonomin och arbetsmarknaden - eller lösa problemet med klimatförändringarna - som självständiga, protektionistiska stater.
Utan EU och euron är kontinenten illa ute, men vi kan inte heller fortsätta som union som om vårt enda problem vore några giriga bankdirektörer. Budgetdisciplin kommer inte att lösa problemet.
Systemet är bristfälligt och måste genomgå en grundlig förändring.
De finansiella institutionerna spjärnar redan emot de regler vi behöver för att förhindra en framtida härdsmälta.
Vi behöver få en bättre integration av vår politik som rör sociala, ekonomiska samt klimat- och energirelaterade frågor för att kunna behålla och skapa arbetstillfällen med goda levnads- och arbetsvillkor.
Vi behöver ett genombrott vid toppmötet om klimatförändringarna i december.
Nu behöver vi mer än någonsin förnya vårt åtagande för millennieutvecklingsmålen och om jag ska vara direkt, herr rådsordförande, tycker jag att det är synd att ni inte krävde ett omedelbart hävande av ockupationen av Gaza eller visade något intresse för att ta nya tag i fredsprocessen tillsammans med president Barack Obama.
Som en av de irländska ledamöterna vill jag påminna parlamentet om att politisk ironi är mycket uppskattat på Irland.
Jonathan Swift, författaren till Gullivers resor, föreslog en gång till den brittiska regeringen att den, för att lösa fattigdomsfrågan på Irland, skulle uppmana irländarna att äta sina barn.
Jag tror inte att irländarna kommer att missa den historiska ironin i förslaget från UK Independence Party om att komma till Irland och propagera för Storbritanniens självständighet i förhållande till EU, utan de kommer att få sig ett gott skratt.
Det kommer att vara en syn för gudar att se Nigel Farage utstyrd i sin Union Jack och sin irländska hatt gå arm i arm med IRA:s forne ledare Gerry Adams och Joe Higgins, min kollega där borta, och uppmana irländarna att rösta nej till Lissabonfördraget, var och en med sina egna ideologiska baktankar, som är helt oförenliga med varandra.
Jag är helt säker på att irländarna kommer att säga till den här cirkusen som de sade till Libertas: Försvinn härifrån!
(Applåder)
(EL) Herr talman! Det svenska ordförandeskapets program omfattar verkligen alla viktiga frågor som är aktuella just nu, både i nuet och i framtiden.
Jag ska börja med recessionen.
Jag antar att det svenska ordförandeskapet kommer att undersöka den här frågan mer ingående.
Den sociala marknadsekonomin behöver investeringar i realekonomin och inte bara i den typ av finansiella produkter som gjorde att vi hamnade i den här situationen från början.
Frågan om klimat och hållbar utveckling, som även inbegriper social utveckling, samt sysselsättningsfrågan är självklart oerhört viktiga.
Men även här behöver vi verkliga investeringar i ekonomin, i kombination med större kontroll.
En marknadsekonomi som försöker närma sig en strategi i stil med laisser faire - laisser passer är inte vad EU behöver.
Frågor som brottslighet och rättsliga och inrikes frågor är något som verkligen berör oss alla.
Den organiserade brottsligheten är inte vad den var tidigare, och den har helt säkert koppling till terrorism och alla andra typer av olaglig verksamhet.
Därför krävs det en annan strategi.
Jag anser att det viktigaste är att vi även undersöker, med tanke på det stora antalet invandrare från tredjeländer, om EU:s utvecklingspolitik verkligen har varit framgångsrik, och i så fall på vilka områden.
Det svenska ordförandeskapets program är verkligen mycket ambitiöst, särskilt när det gäller den transatlantiska dialogen, bland annat.
Men här måste vi fråga oss om det är ändamålsenligt för EU att bara bry sig om utveckling och om det är ändamålsenligt för USA att bara bry sig om säkerhet.
(ET) Mina damer och herrar! Som företrädare för Estland, ett av Sveriges grannländer, med Östersjön som binder oss samman, vill jag tala om en av ordförandeskapets prioriterade frågor, nämligen Östersjöstrategin.
Denna strategi - som infördes med det aktiva stödet från min socialdemokratiska kollega från den tidigare mandatperioden, den nuvarande presidenten Toomas Hendrik Ilves - är mycket viktig för hela EU, och jag vill tacka ordförandeskapet för att det har gjort den till en prioriterad fråga.
Det är även ett gott exempel på hur initiativ som läggs fram från parlamentsledamöter kan få konkreta resultat.
Jag vill uppmana det svenska ordförandeskapet att genomföra Östersjöstrategin och utnyttja detta gyllene tillfälle.
För att kunna göra det måste vi bidra med finansiering till den i nuläget tomma budgetposten i EU:s budget.
Jag hoppas att strategin antas i Europeiska rådet under det svenska ordförandeskapet. Det finns två andra områden som är viktiga för mig.
Som före detta finansminister anser jag att det är mycket viktigt att vi hanterar den ekonomiska krisen och skapar insyn i finanssektorn ... (Talaren avbröts.)
(LV) Herr talman, herr Barroso, herr Reinfeldt! Först och främst vill jag gratulera den svenska regeringen till de mål den har satt upp för sitt ordförandeskap.
Det är ingen lätt tid för EU, det är en tid full av utmaningar.
Bland de många viktiga frågor som Sverige har prioriterat inför sitt ordförandeskap vill jag lyfta fram EU:s strategi för Östersjöområdet, och särskilt den del som rör trygghet på energimarknaden.
Gemensam trygghet för EU:s energimarknad är en omöjlighet så länge problemet är uppdelat och ömsesidigt isolerade marknader förekommer i EU, både när det gäller el och gas.
Av historiska skäl är detta problem särskilt tydligt i Östersjöområdet.
För att lösa problemet och fördela riskerna med elförsörjningen behöver vi en gemensam EU-politik på energifronten.
Grundstenarna i en sådan politik får inte bara vara energieffektivitet och förnybara resurser, utan vi måste även inrätta en gemensam el- och gasmarknad med ett nätverk för verksamheten inom EU.
EU:s Östersjöstrategi är ett steg i rätt riktning.
Den syftar till att gradvis koppla upp områdets energimarknader, få bukt med brister i nätet och skapa gemensamma marknadsmekanismer.
Det arv vi bär på efter Sovjetunionens ockupation av Östersjöområdet är en splittrad och delvis isolerad marknad som ökar riskerna i vår elförsörjning.
Vår utmaning för framtiden ligger i att förändra denna situation, och genom att göra det kommer vi att förbättra vår energitrygghet.
Jag önskar det svenska ordförandeskapet lycka till med att få en kraftfull start på denna viktiga uppgift.
Tack för er uppmärksamhet.
Herr statsminister! För att det ska bli ett bra internationellt klimatavtal måste vi lyssna även på andra länder.
Gör man det inser att man att det krävs för det första att EU och andra länder tar ett större ansvar för att minska våra utsläpp på hemmaplan, och för det andra att EU och andra i-länder konkretiserar hur vi ska bidra ekonomiskt till fattigare länders klimatarbete.
Att den svenska regeringen hittills har motarbetat detta har dessvärre undergrävt möjligheterna till ett bra avtal i Köpenhamn.
Detta måste också ministerrådet inse, och jag vill därför ställa följande två frågor: Är det svenska ordförandeskapet berett att bidra till ett bra internationellt klimatavtal genom att göra en större del av EU:s utsläppsminskningar på hemmaplan?
När tänker man presentera konkreta förslag till finansiering av fattiga länders klimatarbete?
(EN) Herr talman! Jag vill gratulera det svenska ordförandeskapet till detta historiska tillfälle att styra EU mot ett genomförande av Lissabonfördraget.
Jag vill säga tre saker.
För det första är det oerhört viktigt att den nya kommissionen kommer igång med sitt arbete så snart som möjligt.
Institutionell osäkerhet får inte utnyttjas som en ursäkt för att försena bildandet av den nya kommissionen.
Dessa argument låter väldigt hycklande.
För att ta oss igenom den ekonomiska krisen och skapa nya arbetstillfällen behöver vi mer än någonsin en stark, självständig och nytänkande kommission.
För det andra vill jag berömma det svenska ordförandeskapet för att det har tagit initiativet att genomföra Östersjöstrategin, som föreslogs av parlamentet.
Men det finns även en särskild budgetpost för den här strategin som fortfarande är tom. Vi kan inte förvänta oss några positiva miljömässiga förändringar i Östersjön om vi bara förlitar oss på enskilda projekt.
Vi behöver även ett samordnat stöd från EU:s budget.
För det tredje är Stockholmsprogrammet viktigt för Estland.
Det bör även inbegripa ett program för användandet av modern informationsteknik.
Jag undrar om inrättandet av en byrå för verksamhetsstyrningen av storskaliga IT-system inom området med frihet, säkerhet och rättvisa skulle bidra till att genomföra denna strategi.
Herr talman! Gratulationer till utnämningen!
Jag vill också tacka Fredrik Reinfeldt för en utomordentlig genomgång och redogörelse.
Vi förväntar oss nu alla att stordåd ska ske i Köpenhamn, trots att detta också ska betonas vara ett internationellt arrangemang.
Förväntningarna skruvas verkligen upp, men jag vågar säga att om inte alla grupper blir nöjda med resultatet så kommer inte jorden att gå under av den anledningen.
Den ekonomiska krisen har här lyfts fram, självklart.
De stora koncernerna, de stora företagen får alltid uppmärksamhet.
Jag skulle vilja understryka att också de små lojala underleverantörerna inte får glömmas när de finansiella frågorna är på tapeten.
Jag vill också understryka Östersjöstrategins konkreta värden.
Jag tror att Östersjöstrategin kan bli ett legitimitetslyft för hela EU.
Europas största innanhav kan, och måste, räddas.
Östersjöstrategin kan också medverka till att brottsutveckling och trafficking hejdas.
Detta är också en viktig miljöfråga som kanske man kan säga kräver sitt Köpenhamnsmöte.
Det gläder mig att arbetet med en gränslösning mellan Kroatien och Slovenien är aktuellt och att Cypernfrågan också blir löst.
Det är vi alla angelägna om.
Vi får också så småningom, tror jag, se Norden utvidgas här i EU med Island och, gissar jag, också inom en icke avlägsen framtid med Norge.
President Barack Obama höll ett utomordentligt anförande i Afrika om Afrika häromdagen.
Jag har anledning att stryka under att Sverige kan känna sig stolt över sina insatser och jag hoppas att vi kan hålla den solidariska fanan högt fortsättningsvis.
(NL) Jag anser att vi och EU-projektet står vid ett verkligt vägskäl.
Lissabonfördraget, klimatkonferensen i Köpenhamn och en kraftfull strategi för att hantera den finansiella och ekonomiska krisen är tre stora frågor som ni kommer att behöva ta itu med under de kommande sex månaderna, och om vi kan få ett lyckat resultat skulle EU verkligen kunna ta ett stort steg framåt.
Ni är säkert medvetna om att en stor majoritet av ledamöterna är beredda att stödja ert program, och jag vill uppmana er, med glimten i ögat, att låta kritikerna och olyckskorparna föra sitt oväsen vid sidan om.
Låt dem inte avleda er från ert uppdrag, ert syfte.
Jag anser att vi måste koncentrera oss på de viktigaste frågorna.
Låt mig bara påpeka en sak, herr Reinfeldt.
Det är oerhört viktigt att vi koncentrerar oss på en av våra viktigaste prioriteringar, nämligen en ambitiös framtidsplan för bilindustrin i EU.
Enligt min åsikt har vi hittills inte haft en sådan plan - eller så har den varit otillräcklig - jag tror att ni kan hålla med mig om det.
Det är absolut inte för sent.
Räddningsplanen för Opel är redan i full gång, och världen, till och med EU, har fortfarande protektionismen kvar att kämpa emot.
Den ligger och lurar under ytan, och Sverige är precis lika drabbat som Belgien, eller som Frankrike, Tyskland och Slovakien.
Vi sitter alla i samma båt.
Vad vi behöver är att ha en solidarisk inställning till varandra och anta en samordnad strategi i stället för en strategi som går ut på att ”var och en är sig själv närmast”. Det är viktigt att vi inte försöker hålla varandra tillbaka.
Jag anser att ni har fått en unik möjlighet att samarbeta med kommissionens ordförande - detta är även en tydlig signal till kommissionen - för att upprätta en gemensam plan, en gemensam plan, herr Barroso, för våra bilfabrikers framtid. På så sätt kan ni föra dem in i 2000-talet.
Vi anser att det är möjligt att framställa energieffektiva och miljövänliga bilar i de bilfabriker som redan finns i EU, och vi räknar med att ni, herr Barroso och herr Reinfeldt, står på vår sida.
(HU) Enligt vår mening är Sverige synonymt med EU.
Det är ett land med välgång, trygghet och frihet, där frågor som rör de mänskliga rättigheterna och friheterna är lika viktiga som frågor om ekonomi och klimatförändringar.
Sedan har vi det parlament i en av EU:s medlemsstater som antog en ny lag den 30 juni 2009 där det fastslås att om någon, inklusive alla er, inte kallar landets huvudstad vid det namn den har i landets officiella språk, Bratislava, utan använder det tyska namnet Presburg eller det ungerska namnet Pozsony, kan personen i fråga bli tvungen att betala 5 000 euro i böter.
I motiveringen till ändringen av språklagen står det att skyddet av det nationella språket ibland går före yttrandefriheten och rätten till personlig integritet.
Ett EU där sådana lagar antas är inte längre ett frihetens EU.
Jag ber det svenska ordförandeskapet att göra sitt yttersta för att se till att den här lagen upphävs och att den slovakiske statschefen inte undertecknar den.
(HU) Jag vill lyfta fram två av det svenska ordförandeskapets prioriteringar som det gladde mig mycket att se på listan.
Den första av dessa prioriteringar är det otvetydiga ställningstagandet mot diskriminering, rasism, antisemitism, främlingsfientlighet och homofobi.
Jag anser att den här frågan är särskilt viktig med tanke på att vi såg hur tydligt stödet var för högerextremistiska partier i flera EU-länder i valet till Europaparlamentet.
Därför har vi alla ett ansvar, även parlamentet och det nuvarande ordförandeskapet, att se till att de mest utsatta grupperna inte hamnar i svåra situationer.
Vi måste i synnerhet göra allt vi kan för att se till att det inte förekommer något samarbete mellan de partier som gör anspråk på att vara demokratiska och extremistpartierna.
Ett mycket gott exempel på detta är den slovakiska språklagen som redan har nämnts flera gånger i dag, som är gravt diskriminerande, precis som man har beskrivit.
Den andra prioritering som jag vill välkomna är den uppsättning EU-åtgärder som inriktas på att integrera romerna.
(PL) Herr talman! EU:s fortsatta utvidgning och Lissabonfördragets framtid finns med bland det svenska ordförandeskapets mål.
Den tyska författningsdomstolen bedömde nyligen att Lissabonfördraget endast kan godkännas på villkor att Bundestag och Bundesrat får behålla sin företrädesrätt, vilket ifrågasätter EU-federalismen.
Lissabonfördraget har därför visat sig vara ett rättsligt monster, vilket inte bara tyskarna har insett, utan även irländarna i folkomröstningen samt Tjeckiens och Polens presidenter.
Mot bakgrund av detta bör det svenska ordförandeskapet inleda en debatt i hela EU om vilken roll de 27 medlemsländernas parlament ska spela och ta fram en samarbetsmodell mellan suveräna EU-stater.
Därför hoppas jag att det svenska ordförandeskapet, som jag önskar all framgång, kommer att lyssna mer uppmärksamt till medborgarnas röst.
(MT) Jag vill också visa min uppskattning för statsminister Fredrik Reinfeldt för att han stannade hos oss ända till slutet av denna diskussion.
Vi kommer att räkna med att ordförandeskapet driver igenom dessa tre viktiga prioriteringar.
Den första är Stockholmsprogrammet för ett område med frihet, säkerhet och rättvisa.
Vi måste få igenom en överenskommelse om programmet så snart som möjligt.
Den andra prioriteringen är genomförandet av pakten för invandring och asyl.
Vi kommer att förvänta oss av er, herr statsminister, att ni tillämpar den pakt som vi kom överens om förra året.
För det tredje nåddes vid Europeiska rådets möte en överenskommelse om pilotprojektet för ansvarsfördelning i invandringsfrågor.
Ni har mycket arbete som väntar, och vi och vår president kommer att följa er noggrant för att se till att detta arbete utförs.
(PT) Sedan Dag Hammarskjölds tid har Sverige varit en framstående medlem i FN.
Därför vet svenskarna att det, utan organ med allmänt erkänd legitimitet och representativitet, inte kommer att finnas någon politisk kraft för att fullfölja Kyoto2, Doharundan och millennieutvecklingsmålen. Vi kommer inte att kunna reglera den globala ekonomin, och inte heller försvara de mänskliga rättigheterna.
Det är beklagligt att det svenska ordförandeskapet begränsar sig till den informella och omtvistade ramen för G20-mötena.
Det är tragiskt att EU - detta världslokomotiv enligt José Manuel Barroso som citerade FN:s generalsekreterare - varken har någon ledning eller strategisk vision på detta område, samtidigt som president Barack Obama kungör sitt engagemang för det globala styret.
I stället har vi för vår del endast hört påven insistera på det akuta behovet av att omorganisera FN:s säkerhetsråd och Bretton Woods-institutionerna.
Herr rådsordförande, varför vägrar det svenska ordförandeskapet leda EU till att tvinga fram en reform av FN:s säkerhetsråd genom att kräva att EU ska få en plats vid bordet i och med att Lissabonfördraget träder i kraft?
(GA) Herr talman! Den folkomröstning om Lissabonfördraget som kommer att hållas på Irland den 2 oktober i år kommer att vara en av de viktigaste händelserna under det svenska ordförandeskapet.
Irland har fått rättsliga garantier på en rad politiska områden, och detta är till stor hjälp för att minska den oro som folket visade vid folkomröstningen förra året.
Nu måste vi som tror att Lissabonfördraget kommer att gynna Irland arbeta för att driva igenom denna nya överenskommelse i mitt land.
Om Lissabonfördraget ratificeras - och jag hoppas att folkomröstningen kommer att ge ett positivt resultat - kommer de olika länderna att få nominera en medlem till kommissionen.
De som är för fördraget kan inte tillåta sig att vara självbelåtna på något sätt.
Vi måste göra vårt yttersta för att se till att det lyckas.
(Talmannen avbröt talaren.)
(PL) Herr talman! Jag vill mycket gärna tacka statsminister Fredrik Reinfeldt för att han tog med behovet av att utveckla samarbetet med våra grannländer i öst bland sina prioriteringar.
Jag vill även tacka honom för Sveriges engagemang i utvecklingen av det östliga partnerskapet.
Mot bakgrund av detta vill jag påpeka att vi som union och Sverige som ordförandeskap under de kommande sex månaderna kommer att bli tvungna att ta itu med problem som rör åsidosättandet av de mänskliga rättigheterna i Vitryssland.
I sex månader nu har tre entreprenörer, Nikolaj Avtukhowich, Jurij Leonov och Vladimir Osipienko, hållits häktade och inte kunnat få en rättvis dom.
Utav tolv unga aktivister som deltog i en demonstration i januari 2008 har elva fått fängelsestraff och för ett antal dagar sedan dömdes en av dem till ett års fängelse.
Får jag be er, herr statsminister, att under de kommande sex månaderna hålla ett vaksamt öga på brotten mot de mänskliga rättigheterna i Vitryssland.
rådets ordförande. - Herr talman! Jag hoppas kunna återlämna lite av den tid jag lånade tidigare.
(Talmannen avbryter kort.)
Jag vet att ni väntar på en omröstning.
Låt mig tacka er alla för att ni har företrätt era respektive partigrupper på ett mycket bra sätt.
Jag noterar er iver och den förväntan som finns på det svenska ordförandeskapet, er önskan om att vi ska vara mer pådrivande i klimatförhandlingar och agera mot finanskris och ekonomisk nedgång.
Ni har noterat vår Östersjöstrategi, vårt Stockholmsprogram, vår fortsatta strävan att driva på i fråga om utvidgningen, och jag vill tacka er alla för det stöd vi känner för det.
Jag vet också att övergången till Lissabonfördraget kommer att göra att vi träffas igen, och att vi har väldigt mycket att göra tillsammans under denna höst.
Flera av statsråden i min regering finns med mig här i dag.
Vi har noterat och noga följt era frågor och synpunkter.
Jag hoppas på ett nära samarbete och ett återseende under hösten.
Vi räknar även med en ständig diskussion och regelbunden kontakt med ordförandeskapet.
Det är mycket viktigt för Europaparlamentet.
Vi är i början av vår mandatperiod och vi har mycket att göra, och det svenska ordförandeskapet är en mycket bra utgångspunkt.
Tack så mycket, herr statsminister.
Jag vill även tacka kommissionens ordförande.
(Applåder)
Debatten är härmed avslutad.
Skriftliga förklaringar (artikel 149)
Jag välkomnar det svenska ordförandeskapets förslag om att vi bör inrikta oss på politiska frågor i stället för på konstitutionella frågor under Sveriges ordförandeskap.
Men rådet har bestämt sig för att ignorera irländarnas demokratiskt uttryckta vilja, och det har beslutat sig för att tvinga igenom Lissabonfördraget.
Tyvärr är den politiska ram de eftersträvar samma misslyckade agenda för avreglering och liberalisering.
Det är inte det rätta sättet att hantera den ekonomiska krisen.
Tvärtom, det är en fortsättning på den politik som utlöste krisen och det är samma politik som stärks ytterligare i Lissabonfördraget.
Vi får höra att vi behöver Lissabonfördraget eftersom det har tagit många år att utforma det.
Men Lissabonfördraget utarbetades och godkändes före den ekonomiska krisen, och det grundas på en politik som bidrog till att utlösa krisen.
Att tvinga fram denna förlegade politik nu skulle vara en katastrof, eftersom det skulle förvärra krisen ytterligare.
Vi behöver en ny politik för en ny tidsepok.
Vi behöver ett nytt fördrag för en ny tidsepok.
När det gäller klimatförändringarna är det viktigt att det svenska ordförandeskapet gör sitt bästa för att uppnå en stabil överenskommelse i Köpenhamn.
skriftlig. - (EN) Det kommande svenska ordförandeskapet har många utmaningar framför sig, men den största utmaningen är att se till att EU respekterar medlemsstaternas suveränitet och inte trampar på EU-medborgarnas demokratiska rättigheter.
Alltför ofta förbises våra medborgares oro och intressen i den besinningslösa brådskan att driva fram en federalistisk agenda som har sitt exempel i Lissabonfördraget.
När det gäller de förändringar som vi står inför kommer förberedelserna inför reformen av den gemensamma jordbrukspolitiken 2013 att vara en viktig fråga under detta ordförandeskap.
Vi måste lyssna på rösterna från de områden som är starkt beroende av jordbruket, exempelvis Nordirland, i diskussionerna och debatten om reformen av fiskeripolitiken.
Vi har ett stort ansvar för att hjälpa och skydda våra väljare i den rådande finansiella turbulensen.
EU får inte ställa ytterligare hinder i vägen för ekonomisk tillväxt och stabilitet.
skriftlig. - (PT) Det svenska ordförandeskapets antisociala program är ett farligt steg mot utbredandet av den nyliberala politiken.
Det är ett bevis på EU:s kapitalistiska ledares outtröttliga strävan efter denna politik.
Trots att det svenska ordförandeskapet i presentationen av sitt program nämnde medborgarna och problemen med arbetslöshet, nämnde det inte en enda åtgärd för att ändra den befintliga politik som har orsakat dessa problem.
Tvärtom.
Ordförandeskapet framhävde särskilt politiken för fri konkurrens på en lång rad områden, inklusive tjänster och utrikeshandel.
Det har satsat alla sina kort på finansmarknadens återhämtning, ett återupptagande av stabilitetspaktens synsätt och försvaret av nyliberalismen, vilket säkert kommer att leda till nya attacker mot sociala rättigheter och arbetstagarnas rättigheter.
Ordförandeskapet såg också till att insistera på en ny folkomröstning på Irland om förslaget till Lissabonfördraget, som redan har planerats till den 2 oktober. Man fortsätter att bedriva utpressning mot irländarna för att snabbt kunna gå vidare med förstörandet av de offentliga tjänsterna och inskränkningen av de sociala rättigheterna, bland annat inom områden som social trygghet, hälsa, vatten, socialt skydd och arbetstagarnas rättigheter.
Det är lätt att förutse att man kommer att lägga fram förslag till nya direktiv där man försöker driva igenom samma förslag som förkastades under den tidigare valperioden.
Jag välkomnar det kommande ordförandeskapet och jag vill uttrycka min förhoppning om att Sverige, den tredje medlemmen av rådets trojka, kommer att fortsätta det arbete som påbörjades under de tjeckiska och franska ordförandeskapen i fråga om romernas sociala integration.
Flera faktorer hindrade det föregående tjeckiska ordförandeskapets arbete, men på det stora hela ser vi positivt på utvecklingen i romerfrågorna.
Den romska plattformen hade faktiskt sitt första möte i april i Prag, och i juni förstärkte Europeiska rådet sina allmänna mål om att ge romerna jämlika förutsättningar genom att uppmana kommissionen och medlemsstaterna att bekämpa romernas fattigdom och sociala utanförskap.
I samma dokument antog rådet de gemensamma grundprinciper som fastställdes i Prag för att uppnå social integration för romer, med en uppmaning till offentliga beslutsfattare att de ska ta hänsyn till dessa principer och följa dem.
Med tanke på de resultat trojkan hittills har uppnått, hoppas jag att det svenska ordförandeskapet åtminstone ska ägna mer uppmärksamhet än tidigare åt romerfrågorna.
Jag hoppas till exempel att frågan om EU:s största minoritet kommer att prioriteras vid den kommande konferensen om den inkluderande arbetsmarknaden i oktober och toppmötet om jämställdhet i november.
Om man ser till befolkningsmängd är denna minoritet betydligt större än befolkningen i hela Baltikum, som har angetts vara en av ordförandeskapets prioriteringar.
Jag hoppas att det svenska ordförandeskapet kommer att gå längre än de teoretiska strategier som redan har antagits och de organisationsfrågor som redan har retts ut, och börja vidta konkreta åtgärder och på så sätt omsätta denna ram i praktiken.
Stockholmsprogrammet, som är en av det svenska ordförandeskapets prioriteringar, måste ge stöd till främjandet av området med frihet, säkerhet och rättvisa och gynna den ekonomiska verksamheten under den rådande krisen, särskilt med tanke på möjligheten att Lissabonfördraget kommer att träda i kraft.
Om Stockholmsprogrammet lyckas kommer EU att bli mer tillgängligt för sina medborgare.
Denna framgång kommer att märkas i stärkandet av rörelsefriheten för alla EU-medborgare och den omfattande tillämpningen av principen om ömsesidigt erkännande i civilrättsliga frågor och brottmål på EU-nivå.
Det svenska ordförandeskapet måste fortsätta det arbete som påbörjats av de franska och tjeckiska ordförandeskapen, som prioriterade att ge alla arbetstagare i EU full tillgång till gemenskapens arbetsmarknad, en frihet som i allra högsta grad symboliserar EU-medborgarskapet.
För att göra detta måste medlemsstaterna delta aktivt genom konkreta åtgärder i avskaffandet av de virtuella gränser inom EU som begränsar medborgarnas rörelsefrihet eftersom de drabbas av administrativa och rättsliga problem när de lever och arbetar i en annan medlemsstat.
Rörelsefriheten måste vara en verklighet för alla EU-medborgare, särskilt under den rådande ekonomiska krisen som förstärker behovet av att stödja fri rörlighet för arbetskraften.
Denna rörlighet kan vara självreglerande och ge flexibilitet och minska mängden oredovisat arbete och den naturliga arbetslösheten.
EU står inför enorma utmaningar just nu: den ekonomiska och finansiella krisen, den oroväckande ökningen av arbetslösheten och klimatförändringarna.
Arbetslösheten i EU ligger på 8,9 procent just nu, och 19 procent av ungdomarna under 16 år samt 19 procent av de äldre riskerar att hamna i fattigdom.
Människor förlorar sina arbeten, många företag går i konkurs och det finns stora underskott i de statliga budgetarna.
EU:s svenska ordförandeskap har ett enormt ansvar gentemot sina medborgare.
Det måste återupprätta hoppet om ett drägligt liv och lägga grunden för ekonomisk återhämtning genom att få alla att hjälpas åt.
Det svenska ordförandeskapet prioriterar åtgärder som att öka energieffektiviteten, använda energi från förnybara källor och förbättra EU:s energitrygghet.
Jag hoppas att EU:s svenska ordförandeskap kommer att bli början på en period av välstånd som tryggar den ekonomiska tillväxten för de kommande 40-50 åren.
Jag anser att vi nu, mer än någonsin, behöver investera i utbildning, forskning, energieffektivitet och framför allt i människorna.
Sverige är känt för sin sociala politik och sin höga levnadsstandard.
Därför vill jag, tillsammans med mina kolleger i parlamentet och alla EU:s medborgare, önska er all framgång, och vi hoppas att den här perioden kommer att bli en språngbräda in i en ny framtid.
skriftlig. - (EL) Det svenska ordförandeskapets prioriteringar är en upptrappning av EU:s gräsrotsfientliga kampanj vars syfte är att trygga den fortsatta lönsamheten med det EU-omfattande kapitalet genom att lämpa över den kapitalistiska recessionen på arbetarklassen och vanliga medborgare.
Det svenska ordförandeskapet vill skynda på kapitalistiska omstruktureringar inom ramen för Lissabonstrategin.
I centrum för denna attack mot arbetstagarna ligger nedskärningar av löner och pensioner, ett fullständigt raserande av arbetsrelationerna, arbetstagarnas rättigheter, socialt skydd och försäkringssystem samt en allt större privatisering av hälso- och sjukvården och av utbildningsväsendet.
Den ”gröna ekonomin” är utformad så att nya, lönsamma verksamhetssektorer kan öppnas för kapital, under förespeglingen att bekämpa klimatförändringarna.
Med Stockholmsprogrammet försöker man, genom att påstå sig bekämpa terrorism och organiserad brottslighet, ytterligare förstärka det borgerliga politiska systemet så att de kan kväva reaktioner på gräsrotsnivå och trappa upp de diskriminerande åtgärderna mot invandrare.
Östersjöstrategin har banat väg för en mer aggressiv strategi från de EU-omfattande monopolen i EU:s östliga länder som försöker stärka sin position i den imperialistiska dragkampen.
Genom att använda ”garantier” som en dimridå och genom att utöva uppenbart tvång, försöker man roffa åt sig irländarnas röster för att genomföra det gräsrotsfientliga Lissabonfördraget.
Meddelande om förslag från talmanskonferensen: se protokollet
Meddelande från talmannen
(efter Rebecca Harms inlägg, se punkt 4.1).
Ja, fru Harms.
Jag vill informera er om att talman Jerzy Busek har gjort ett offentligt uttalande om den fråga ni just nämnde. Jag kommer att läsa upp det för er.
Det är med mycket stor sorg jag har hört om Natalja Estemirovas tragiska död, som bortfördes tidigare i dag i Grozny.
Jag vill på Europaparlamentets vägnar uttrycka vår medkänsla och sända våra kondoleanser till den avlidnas familj och vänner.
Natalja Estemirova var en människorättsaktivist och en ledande forskare i Tjetjeniens historiska minne.
År 2005 tilldelades hon Robert Schuman-medaljen av PPE-gruppen i Europaparlamentet.
Vi i Europaparlamentet har uppskattat hennes arbete med mänskliga rättigheter, främjande av demokratisk ansvarsskyldighet och upprätthållande av rättsordningen.
Vi uppmanar på det bestämdaste myndigheterna i Ryssland att inleda en ingående utredning av hennes död och göra sitt yttersta för att ställa de ansvariga för denna tragiska död inför rätta.
Europaparlamentet står i främsta linjen för främjandet av demokrati, upprätthållandet av rättsordningen och försvaret av de mänskliga rättigheterna.
Det är därför vår skyldighet att stödja och visa vår solidaritet med alla dem som kämpar överallt i världen för samma värden, vilket Natalja Estemirova gjorde.
(Applåder)
Fru Harms! Ordförandeskapet instämmer i ert förslag om att hålla en tyst minut till Natalja Estemirovas minne.
(Parlamentet höll en tyst minut.)
Begäran om upphävande av parlamentarisk immunitet: se protokollet
Anföranden på en minut om frågor av politisk vikt
Vi ska nu övergå till anförandena som får vara högst en minut långa.
Talarlistan är mycket lång.
Detta visar att det finns ett stort intresse av att delta, vilket hedrar denna kammare.
Jag kommer dock inte att kunna ge ordet till alla de som vill tala, eftersom 100 begäranden skulle ta en och en halv timme medan vi däremot bara har en halvtimme till förfogande.
(GA) Herr talman! Eftersom detta är första gången som jag får tala i parlamentet skulle jag vilja inleda på mitt modersmål.
Som ni vet pågår kampanjen inför folkomröstningen om Lissabonfördraget för fullt i Irland just nu och vi hoppas på ett positivt resultat den 2 oktober.
En av de saker som gör en stor skillnad den här gången är de garantier som Europeiska unionen har gett den irländska regeringen när det gäller skatter, aborter och försvar.
Något som inte nämndes överhuvudtaget förra gången och som också är mycket viktigt är befogenheterna inom idrott som nu har införlivats i Lissabonfördraget.
(EN) Jag har alltid varit idrottsengagerad: Jag har spelat på olika nivåer och varit aktiv i styrelser.
Jag anser därför och av andra mer uppenbara skäl, till exempel de hälsorelaterade, sociala och fysiska fördelarna med idrott, att det är viktigt att man efter Lissabonfördraget ger betydande resurser till...
(Talmannen avbröt talaren)
(RO) Herr talman! Jag anser att det finns vissa olikheter mellan strukturproblemen inom Rumäniens jordbrukssektor och de som finns i andra medlemsstater.
Jag måste understryka att Europeiska unionen borde utnyttja sitt politiska och ekonomiska inflytande för att lägga större vikt vid förvaltningen av det jordbruksstöd som ges till de nya medlemsstaterna.
Min åsikt är att man också kan lösa problemet genom att stödja en hållbar jordbrukssektor med en lämplig budget efter 2013. Detta skulle ge jordbrukarna framtidsutsikter på medellång och lång sikt och tillräckliga resurser så att det rumänska jordbruket kan komma i nivå med europeiska standarder.
(SK) Mina damer och herrar! Ungern och de ungerska minoriteterna tar ständigt upp frågan om nationella minoriteter.
Genom att ta till halvsanningar och ibland även lögner försöker de manipulera den allmänna opinionen inom EU till deras fördel.
Vad är sanningen egentligen?
Under de senaste 80 åren har de nationella minoriteterna i Ungern nästan utplånats samtidigt som EU tigande har sett på.
Den slovakiska minoriteten har även den minskat från 300 000 till 10 000 medlemmar.
Antalet medlemmar i de ungerska minoriteterna i de angränsande länderna, däribland Slovakien, har förblivit oförändrat.
Under de två senaste åren har sex romska medborgare mördats i Ungern och dussintals har blivit allvarligt skadade.
Det finns en rädsla för attacker mot judar samtidigt som andra former av extremism ökar och sprider sig över gränserna.
Ungern hanterar inte denna typ av aggression på rätt sätt och landet måste fördömas.
EU-institutionerna borde inta en mer bestämd hållning mot dessa tecken på extremism.
(PT) Den kupp som ägde rum i Honduras den 28 juni var ett angrepp mot det honduranska folkets politiska yttrandefrihet och de mest grundläggande demokratiska rättigheterna.
Sedan dess har regeringen faktiskt vidtagit repressiva åtgärder mot gräsrotsrörelsen. Denna har demonstrerat på gatorna och infört ett system med medietystnad, begränsade friheter, förföljelse, olaga frihetsberövande, försvinnanden och till och med mord på medlemmar i den organiserade motståndsrörelsen mot kuppen.
Vi kunde bevittna allt detta under det besök som nyligen gjordes av en delegation från Europeiska enade vänstern/Nordisk grön vänster i Honduras och Nicaragua där vi träffade landets lagligt valda president, Manuel Zelaya. EU-institutionernas reaktioner på dessa omständigheter är minst sagt tvetydiga.
Medan några är oacceptabelt tystlåtna vädjar andra till båda parter att göra allt som står i deras makt för att nå en politisk lösning så fort som möjligt.
De drar alla över samma kam och struntar i vem som är skyldig. Det är precis som om det inte fanns någon demokratiskt vald president på ena sidan och en olaglig regering på den andra vilken presidenten frihetsberövades och landsförvisades av när den på olaglig väg övertog makten.
Den mest grundläggande respekten för demokrati kräver att EU-institutionerna tydligt och kraftigt måste fördöma kuppen och genomföra åtgärder på internationell nivå för att isolera och öka trycket på den olagliga regering som är vid makten.
De får inte heller erkänna eller stödja några val som hålls innan den demokratiska legitimiteten har återupprättats i landet.
(EN) Herr talman! Som en ny ledamot av detta parlament anser jag att ett av de största problem som jordbrukare i Wales och resten av Storbritannien står inför är den föreslagna elektroniska identifieringen av får som kommer att införas den 1 januari 2010.
Saken är den att skanningsutrustningen inte är tillförlitlig.
Om jag har förstått det rätt har den bara en tillförlitlighet på 79 procent vilket kommer att leda till stora problem för jordbrukare i hela Storbritannien.
Jag uppmanar kommissionen att ompröva dessa bestämmelser och bara införa detta på frivillig grund för lantbrukarna.
Jag är rädd för att den otillförlitliga utrustningen kommer att skada många jordbrukare och att det samlade gårdsstödet kommer att minskas.
I allra värsta fall kan det minskas med 100 procent.
De eftergifter som redan har gjorts är till stor hjälp men otillräckliga.
Jag tycker att det rent av är förvånande att kommissionen vill införa elektronisk identifiering med en utrustning som har så pass stora brister.
En förnuftig lösning vore att införa elektronisk identifiering endast på frivillig grund från januari nästa år.
Jag ber ledamöterna i detta parlament att stödja mig i denna oerhört viktiga fråga för jordbruksnäringen i hela EU.
(EN) Herr talman! Jag skulle vilja uppmana parlamentet att vidta omedelbara och effektiva åtgärder för att rädda de små jordbruken och familjejordbruken i de nya medlemsstaterna, framför allt i Öst- och Centraleuropa och då särskilt i mitt eget land, Ungern.
Vad har dessa jordbrukare råkat ut för?
Som en följd av att vi anslöt oss till Europeiska unionen var vi tvungna att ”erbjuda”, så att säga, 100 procent av vår marknad och i utbyte fick vi ett stöd på motsvarande 25 procent.
Detta är inte bara orättvist och oberättigat utan även olagligt: Det har gjorts en tydlig överträdelse av Romfördraget.
Eftersom jordbrukarna har försökt konkurrera på dessa orättvisa och olagliga villkor har de tvingats ta enorma lån för att inte konkurreras ut.
Nu har de försatts i konkurs och måste sälja sin mark under omständigheter som påminner om kolonisering. Vi måste nämligen upplåta marken till länder som har 10 gånger högre BNP än vad vi har.
Jag begär att Köpenhamnsavtalet omprövas omedelbart.
(Talmannen avbröt talaren)
(RO) Herr talman! Jag skulle precis som mina medledamöter vilja ta upp ett problem inom jordbrukssektorn.
En artikel som nyligen publicerades i Wall Street Journal har särskilt fångat mitt intresse och därför ser jag det som en hedersplikt att presentera denna för parlamentet och framföra skribenternas önskemål.
Artikeltiteln, som jag tycker förmedlar vad artikeln handlar om, löd ”Barroso, ta bort hindren för småföretagarna”.
Artikeln är helt enkelt en vädjan till den framtida Europeiska kommissionen att koncentrera sina åtgärder på att ge stöd till små och medelstora företag, som är mycket sårbara i kristider, och att inte på något sätt kompromissa om genomförandet av 2008 års Small Business Act.
Europaparlamentet har en skyldighet att se till att dessa åtgärder genomförs på ett vederbörligt och effektivt sätt eftersom de behövs för de över 20 miljoner små och medelstora företagen i Europeiska unionen.
(BG) Herr talman! I början av augusti ägde en oerhört dramatisk händelse rum i f.d. jugoslaviska republiken Makedonien som chockade allmänheten i Bulgarien.
Spaska Mitrova, en 23-årig medborgare i f.d. jugoslaviska republiken Makedonien och mamma till ett litet barn som då fortfarande ammades, fördes med våld till polisstationen och förflyttades sedan till det ökända fängelset Idrizovo samtidigt som hon fråntogs sitt barn.
Polisen tog tag i hennes hår och drog ner henne från översta våningen till bottenvåningen av byggnaden eftersom hon inte ville skiljas från sitt barn.
Hon dömdes till tre månaders fängelse eftersom hon inte kunde ge sin före detta make en sovplats i deras barns sovrum.
Ni kan föreställa er följderna av detta.
Vidare fick Spaska Mitrova bulgariskt medborgarskap tidigare i år.
Detta verkar vara den främsta orsaken till den omänskliga behandling som hon utsattes för, och detta fall är inte det första.
För cirka två år sedan frågade jag den nuvarande utrikesministern i f.d. jugoslaviska republiken Makedonien om varför det finns så mycket hat mot människor från f.d. jugoslaviska republiken Makedonien med bulgariskt medborgarskap.
Han svarade att de är spår från det förflutna.
Eftersom de ansträngningar som har gjorts av den bulgariske presidenten och den bulgariska regeringen inte har lett till något resultat ber jag kommissionsledamot Olli Rehn att personligen sätta sig in i detta fall som kännetecknas av uppenbar orättvisa i ett land som vill inleda anslutningsförhandlingar.
(SL) Italien vill anlägga en gasterminal utmed kusten på gränsen till Slovenien utan samråd.
Europeiska unionen grundades dock på ömsesidigt förtroende och goda grannskapsrelationer.
Miljöskadliga energikällor kräver särskilda miljöskyddsåtgärder men i grund och botten även grundläggande ärlighet.
Italien försöker undanhålla Slovenien information om de skadliga konsekvenserna för den gränsöverskridande miljön. Italien skadar på så sätt alla inblandade, inklusive sig självt men framför allt de människor som bor i närheten av den omtvistade anläggningen.
Allmänheten och regeringen i Slovenien motsätter sig starkt denna terminal.
Att ljuga inför kamerorna kan mycket väl vara Berlusconis taktik för politisk överlevnad i Italien.
Ett sådant beteende får och borde dock inte accepteras som en medveten handling inom Europeiska unionen.
Det är oacceptabelt.
Det hela utgör en uppenbar överträdelse av Europeiska unionens principer och Italien utövar en manipulativ taktik vilket skadar mänskligt liv och miljön.
Det vore internationellt sett vårdslöst att försöka bygga en kustterminal vid Žavlje (Aquilinia) i Triestebukten som redan är extremt trång.
Det förstör miljön, raserar framtidsutsikterna för kommunalt samarbete vid gränsen och utgör ett mycket dåligt exempel för kommande medlemsstater.
(PT) Herr talman! Det som händer med den före detta tyska skotillverkaren, Rhode, i Santa Maria da Feira, som nu heter Sociedade Luso-Alemã de Calçado, är mycket oroande.
Företaget hade en gång i tiden nästan 3 000 anställda men efter problemen i Tyskland har företaget tagit bort flera arbetstillfällen och har nu runt 1 000 anställda.
Merparten av dem är kvinnor som de flesta har fått gå ned i timmar och lön.
Man fruktar nu att företaget kommer att läggas ned när det portugisiska valet är över.
Arbetslösheten i kommunen fortsätter att öka och drabbar nu tusentals anställda, särskilt inom sko- och korktillverkningsindustrin.
Med tanke på detta ber vi om att särskilda nödåtgärder vidtas för att förhindra ännu ett allvarligt slag mot tillverkningen och arbetstillfällena i ett område som har drabbats så pass hårt av arbetslöshet.
(EN) Herr talman! Jag accepterar inte parlamentets eller någon annan EU-institutions behörighet att stifta lagar för Storbritannien.
Mina väljare har sänt mig hit för att tala om för er att de inte vill att 45 miljoner brittiska pund av deras pengar ska användas varje dag på Europeiska unionen.
Vi vill att dessa pengar ska användas inom Storbritannien, på våra skolor, våra sjukhus och vår infrastruktur, och inte kastas bort på era korrumperade räkenskaper under 14 års tid.
Jag har helt enkelt följande budskap från de som har valt mig till kommissionen: Fortsätt ni med er byråkrati och var beredda på Storbritanniens utträde ur den korrupta och dödsdömda röra som Europeiska unionen är.
(EN) Herr talman! Detta parlament stod nyligen enat inför ett globalt terrorhot.
I min valkrets i Nordirland vet vi vad terrorism kan orsaka.
Ja, vi har sett en förändring i Nordirland de senaste åren men det finns fortfarande de som gärna skulle vilja se blod flyta.
Förra veckan utplacerades en bomb på ca 275 kilo av oliktänkande republikaner i South Armagh.
Om den inte hade upptäckts hade många människor mist livet.
I Nordirland har vi inte glömt de som föll offer för vårt förflutna och för terrorism och därför skulle jag vilja be parlamentet om att stödja kravet på ersättning från Libyen.
Libyen tillhandahöll IRA vapen.
Dessa vapen dödade många människor och skadade andra.
Landet måste hållas ansvarigt för detta.
(SK) Så här i början av en ny mandatperiod bör vi tänka på vårt gemensamma ansvar för en fredlig utveckling i Europa, så att våra medborgare kan leva ett fridfullt och angenämt liv.
Vi måste även visa våra medborgare att vi är här för deras skull, för att tillvarata deras intressen.
Vi måste alltid ha detta i åtanke, även när det uppstår problem mellan två parter i vår politiska familj.
Det europeiska sättet att lösa problem är att föra en dialog i sann partnerskapsanda, i syfte att nå förnuftliga lösningar, och inte att ignorera den andra parten eller lägga fram frågor direkt till EU-institutionerna, som det här är ett exempel på.
En ständig, förnuftig och ömsesidig dialog är också den rätta vägen för att motverka extremister på båda sidor, och på så sätt kväva eller strängt begränsa eventuella farliga handlingar som de kan begå i framtiden.
(RO) Kampen mot rasism utkämpas genom kraftfull EU-politik, och ändå har på mindre än en vecka tyska och brittiska politiker varit inblandade i smutskastning av rumänska arbetstagare, antingen på grund av okunnighet eller på grund av en drivkraft att kunna vinna sympatier och röster från befolkningen.
Mycket oroande är makabra uttalanden som att rumäner skulle sticka en kniv i dig så snart de fick syn på dig, vilket yttrades på ett offentligt möte i Storbritannien, och kommentarerna från en tysk politiker om att rumäner inte kommer till arbetet klockan sju på morgonen och inte heller vet vad de ska göra.
Vi utarbetar EU-politik för att motverka rasism.
Det är vårt gemensamma mål.
Men vad gör vi om våra politikerkolleger från stora EU-medlemsstater uttalar sig på det här sättet?
(ES) Herr talman! Förra veckan blev tre baskiska tonfiskfartyg från Bermeo återigen hotade av somaliska pirater.
Vi är oroade över de upprepade angreppen mot fiskefartyg i området och över att offren känner sig otrygga, samtidigt som den spanska regeringen inte gör någonting.
Dessa angrepp kan förvärras när monsunen kommer, precis som yrkesfiskarna säger.
Innan det är för sent vill jag därför här i kammaren säga att vi snarast behöver beväpnat militärt skydd ombord på dessa fartyg.
Några av de europeiska regeringarna har redan föranlett detta, till exempel Frankrikes och Italiens regering, vilket har varit framgångsrikt.
Kommissionen bör därför rekommendera att alla medlemsstaterna omedelbart vidtar liknande kraftfulla åtgärder.
Vi måste snarast utöka de skyddskriterier som har upprättats för handelsfartygens sjövägar till fiskeområdena.
Parlamentet har ett problem, vilket fastställdes i resolutionen om kapningar till sjöss av den 23 oktober förra året.
Avslutningsvis vill jag på nytt upprepa vår övertygelse att Europa behöver en gemensam utrikes- och säkerhetspolitik som gör EU-institutionerna mer effektiva och trovärdiga när det gäller att ta itu med sådana här kriser.
(EL) Herr talman! Den 4 september 2009 utförde de tyska trupper som utgör en del av den ockuperande armén i Afghanistan tillsammans med Förenta staterna, EU och Nato dödliga attacker i regionen Kunduz, som visade sig bli en massaker med över 135 civila dödsoffer och dussintals skadade, däribland många barn, vilket är en krigsförbrytelse mot det afghanska folket.
Det här angreppet var givetvis inte ett angrepp mot talibanerna, utan mot 500 civila medborgare.
Det dagliga blodbadet, det organiserade våldet och de korrupta valen för att sätta marionetter för den afghanska ockupationen på plats liksom den fattigdom och misär som hemsöker det afghanska folket visar att de imperialistiska angrepp som Förenta staterna, EU och Nato har genomfört under förevändningen att de ska motverka terrorism i detta ockuperade land - och även i en rad andra länder - har fått katastrofala följder för människorna.
Både uttalandena från Natos nye generalsekreterare Anders Fogh Rasmussen och från EU:s utrikesministrar syftar till en enda sak: att fortsätta ingripa mot folket.
Människorna i varje land och i varje EU-medlemsstat måste kräva och insistera på att dessa trupper lämnar deras länder och återvänder hem.
(EN) Herr talman! Den 2 oktober kommer Irland att hålla en ny folkomröstning om Lissabonfördraget.
Lissabonfördraget är i stort sett identiskt med den konstitution för Europa som fullständigt förkastades av Frankrike och Nederländerna.
Lissabonfördraget har redan förkastats av Irland en gång, men ”nej” är alltid fel svar när det gäller EU och fortsatt politisk integration.
Därför måste irländarna hålla en ny folkomröstning så att de kan komma fram till det enda svar som är godtagbart i EU - nämligen ett ”ja”.
EU håller på att förstöra demokratin i medlemsstaterna.
EU bygger på felaktiga påståenden, bedrägerier och lögner.
I Storbritannien har vår föraktliga regering och politiska fraktion sagt nej till en folkomröstning, just på grund av att de vet att resultatet skulle bli ett rungande ”nej”.
Men oavsett hur resultatet blir i Irland kommer Storbritannien en dag att lämna EU och återvinna sin nationella självständighet.
Jag är stolt över att kunna använda min tjänsteställning för att förorda Storbritanniens ovillkorliga utträde ur EU.
Tack, herr Batten.
Jag gav er 14 extra sekunder även om ni sade en sak som inte stämmer, nämligen att Lissabonfördraget är samma sak som konstitutionen.
(RO) Herr talman!
Jag vill tala om ett EU-projekt som kallas ”Voices of Youth” och som jag har fått äran att ansvara för.
Unga människor från alla medlemsstaterna kan delta i det här projektet och målet är att de ska hitta och föreslå lösningar på sociala problem som de stöter på.
Jag ber inte bara er, herr talman, utan även Europeiska kommissionens ordförande att se till att vi bättre uppmärksammar de förslag som de kommer med.
Det är vårt ansvar i dessa svåra tider att se till att Europa och framför allt unga europeiska medborgare får tydliga möjligheter.
Min generation har varit tillräckligt lyckligt lottad för att ta del av återuppbyggnaden av ett enat Europa.
Unga människor som utgör dagens Europa och särskilt morgondagens har rätt att skapa det Europa som de vill ha. Tack.
Må Guds hjälp vara med oss.
Tack, och tack även för det kortfattade anförandet.
(HU) Spöket av den vänster- och högerextremistiska ideologi som återspeglar de två diktaturer som dominerade Europa under 1900-taler har återvänt för att hemsöka 2000-talets EU.
Vi har ett fall där en EU-medborgare har förbjudits att resa till ett annat land, vilket innebär att rörelsefriheten för denna person har begränsats.
I ett annat fall ville en EU-medlemsstat arrestera 15 medborgare, anklaga dem för förräderi och förbjuda dem att lämna landet eftersom de skulle diskutera minoritetsfrågor med likasinnade landsmän i ett forum för ungerska parlamentsledamöter från Karpaterna.
I det berörda landet bestraffas människor för att de inte talar landets officiella språk ordentligt på sjukhus, polisstationer, ålderdomshem och mödravårdscentraler.
Inte ens immigranter behandlas på det här sättet i EU, än mindre människor som har levt här under tusen år, där en ny stat bildades för bara 17 år sedan.
Därför är det viktigt att EU inför en gemensam lag som skyddar minoriteter och som är bindande för alla länder.
(EN) Herr talman! Jag vill informera parlamentet om att den brittiske justitieministern i förra veckan bad en av mina väljare om ursäkt, nämligen Michael Shields, som har släppts fri från fängelse efter att ha suttit fyra och ett halvt år för ett brott som han inte har begått.
Michael Shields fick en ursäkt på grund av bevis som tydligt visar att han är moraliskt och tekniskt oskyldig till brottet.
Shields arresterades, anklagades och dömdes 2005 på mindre än åtta veckor för ett brutalt överfall mot Martin Georgiev, en bulgarisk kypare, trots att det saknades rättsliga bevis, att identifieringsförfarandet genomförts bristfälligt och att en annan man, Graham Sankey, undertecknat en bekännelse av brottet.
Jag vill i dag tacka talman Josep Borrell Fontelles och talman Hans-Gert Pöttering samt parlamentets utskott för framställningar för deras stöd till Michael Shields kamp för rättvisa.
Än är det hela dock inte över, och jag ber ordföranden för utskottet för framställningar att fortsätta att stödja Michael Shields kamp för rättvisa och snarast uppmana de bulgariska myndigheterna att granska bevissamlingen.
Detta är mycket viktigt för att var och en av våra medborgare ska kunna ha tillit till och förtroende för det rättsliga och politiska samarbetet i Europa.
(ET) Bankväsendet kräver övervakning.
Det är Europeiska rådets och Europeiska kommissionens ståndpunkt.
Europeiska kommissionens konsumentskyddsundersökning, som offentliggjordes i februari, avslöjade flera allvarliga negativa tendenser inom bankväsendet.
Som vald företrädare från Estland vill jag ge några exempel från Estland för två svenska banker som har verksamhet i Estland.
Problemet är att dessa banker behandlar kunder i Estland annorlunda än kunder i det egna hemlandet.
Både priserna för banktjänster och räntesatserna är betydligt högre för de estniska kunderna.
Räntesatserna skiljer sig exempelvis mellan 0,21 % i Sverige och 12,2 % i Estland - vilket är 600 gångers skillnad.
Att använda finanskrisen för att rättfärdiga olika behandling strider mot EU:s värderingar.
Jag skulle vilja fråga Sverige, som för närvarande är EU:s ordförandeland, vad man har att säga om detta och hur länge det kommer att vara på det här sättet med deras banker i Estland.
(DE) Herr talman! Jag har tidigare sagt att vi behöver en demokratisk revolution, och nu står vi alla som av egen fri vilja inte företräder någon politisk grupp i parlamentet inför en ohållbar situation.
Jag vill be presidiet att finna en vänskaplig lösning på problemet med samordnare.
I det här avseendet är vi diskriminerade eftersom vi inte får delta i samordnarnas sammanträden i de olika utskotten och vara vederbörligen aktiva.
Jag vill gärna medverka till att undvika att rättegångsförfaranden i EG-domstolen resulterar i ett utslag att alla beslut som har fattats hittills av samordnarna ogiltigförklaras, så som tidigare har skett i kölvattnet efter diskrimineringsmålet från 2001.
Det skulle inte bara vara till enorm skada för parlamentet, utan det är även onödigt från politisk synpunkt.
Jag ber därför presidiet att snarast vidta lämpliga åtgärder för att sätta stopp för denna diskriminering av grupplösa ledamöter och återgå till de solida arbetsmetoder som vi haft under de senaste tio åren.
(ES) Herr talman!
Den här sommaren har terroristgruppen ETA mördat tre människor i Spanien som försvarat rättvisa och frihet, nämligen en polisman från den nationella poliskåren och två befäl inom civilförsvaret.
Jag vill uttrycka vårt deltagande, vårt stöd och vår omsorg till deras familjer.
ETA är en kriminell grupp som inte hör hemma i Europa, eftersom det i EU inte finns utrymme för radikalism, totalitarism eller terroristmord.
Europaparlamentet och alla EU-institutionerna bör av denna anledning fortsätta att fördöma ETA-terrorister och arbeta för att undanröja och utrota den cancersvulst som ETA:s terroristattentat utgör och deras medverkan till brott från vår kontinent.
I mitt första anförande vid denna mandatperiods första ordinarie plenarsammanträde i Europaparlamentet vill jag därför påminna om och uppmärksamma alla dem som fallit offer för ETA:s terrorism, och fördöma terroristorganisationen ETA här i kammaren.
(EN) Herr talman! För sex månader sedan chockades världen av den död och ödeläggelse som Israel utsatte Gazaremsan för.
När kamerorna nu har stängts av fortsätter den ekonomiska belägringen.
Mindre än en fjärdedel av de material och förnödenheter som människorna är i behov av kommer igenom gränsövergångarna - bara 18 artiklar allt som allt.
Ingenting för återuppbyggnad, ingenting för affärslivet, ingenting som skapar arbetstillfällen eller inger hopp.
Israel håller praktiskt taget en och en halv miljon människor i ett slags fångläger, omgivet av murar och övervakat av beväpnade vakter.
Jag ber er, herr talman, att uppmana ordföranden att besöka Gaza snarast möjligt för att bedöma läget på egen hand.
Om han anser att en sådan kollektiv bestraffning inte kan godtas bör han uttala sig till förmån för alla oskyldiga.
- (DE) Herr talman! Den ekonomiska krisen har slagit hårt mot jordbruksproduktionen.
Situationen har försämrats drastiskt särskilt för mjölkproducenterna de senaste 20 månaderna.
Med priser under 0,21 euro tvingas jordbrukarna sälja sin mjölk till ett pris som är lägre än deras produktionskostnader.
Överlevnaden för många av de familjedrivna jordbruken i EU är allvarligt hotad, och i dagsläget kan många av dem bara överleva genom privata besparingar, vilket naturligtvis inte är hållbart.
Kommissionens siffror ger en dramatisk bild över prisfallet för mjölk och mjölkprodukter.
Åtgärder till stöd för mjölkproducenterna är av största vikt för att undvika en kollaps inom jordbruket.
Kvalitet har som bekant sitt pris, men den principen tycks inte gälla längre inom jordbrukssektorn.
För närvarande står producenternas pris inte i relation till konsumenternas pris.
Våra familjedrivna jordbruk behöver snarast marknadsstödsåtgärder.
Det handlar om att säkra livsmedelsförsörjningen i Europa.
Framför allt får vi inte glömma bort att hundratusentals arbetstillfällen i Europa är beroende av ett fungerande jordbruk.
(EN) Herr talman! Jag vill ta upp fallet med John Zafiropoulos, som sitter i fängelse i Grekland.
Hans familj, som tillhör min valkrets, är övertygad om att han är oskyldig.
I början av det här året skrev jag till justitieministern i Aten angående fallet.
Jag fick inget svar, så i ett anförande på en minut här i maj tog jag upp det i kammaren.
Omedelbart efter att jag hade talat kom Greklands ständiga representation skyndande till mitt kontor och lovade mig att snarast komma med ett svar från ministern personligen.
Fyra månader senare har ingenting hänt.
Om Greklands ständiga representation lyssnar på oss nu i kammaren vill jag uttrycka min förvåning och bestörtning över att ingenting har hänt.
Jag ber om ett svar från ministern och att John Zafiropoulos fall ska undersökas på nytt.
(EN) Herr talman! Under den turiska ockupationen av Cypern 1974 fotograferade en turkisk journalist 14 cypriotiska soldater som överlämnades till den turkiska armén.
Fotografiet blev en symbol för sökandet efter de saknade personerna.
För ett par veckor sedan identifierades soldaternas kroppar genom DNA, 35 år efter att de dödats och blivit nedslängda i en grav i den ockuperade norra delen av ön.
Detta är ett bevis för en uppenbar överträdelse av Genèvekonventionen av den turkiska armé som var ansvarig för de fångar som överlämnades till dem.
Jag uppmanar parlamentet att uppmana Turkiet att samarbeta med FN:s kommitté för saknade personer genom att ställa sina förteckningar till förfogande och öppna de båda platser som nyligen har pekats ut i Lapithos, vilka betecknas som ”skyddade militära områden”, där man tror att ytterligare 800 fångar ligger begravda.
(EN) Herr talman! I parlamentet kommer vi att ha många viktiga diskussioner och beslut att fatta i budgetfrågor.
För närvarande behandlar vi givetvis budgeten för 2010, och fortfarande är det många problem som måste lösas innan vi kan enas om den.
Parlamentet kommer snart också att börja diskutera den nya budgetplanen för tiden efter 2013.
Samtidigt har vi även halvtidsöversynen av budgeten, och jag tycker att det verkar som om vi nästan har glömt bort det.
Vi får inte glömma den, eftersom den ger oss stora framtida möjligheter.
Vi kommer att kunna granska våra prioriteter på nytt.
Vi kommer exempelvis att kunna tilldela den nya ekonomiska återhämtningsplanen för Europa mer stöd.
Vi kommer kanske också att kunna avsätta mer medel till de åtgärder som Köpenhamnskonferensen leder fram till i slutet av året.
Jag anser att parlamentet måste hålla ett öga på det här.
Parlamentet bör fortsätta att utöva påtryckningar på rådet och kommissionen, så att de återigen granskar halvtidsöversynen och vi får möjlighet att framföra våra prioriteringar.
(HU) Herr talman! Yttrandefrihet och frihet att välja vilket språk man vill tala är grundläggande mänskliga rättigheter.
Ett språk är en symbol av största vikt för alla som talar det och själva grunden för deras självidentitet.
Alla som tänker så om sitt eget språk måste respektera andra folkgruppers olika språk.
Nyligen har emellertid ett av EU:s officiella språk angripits i Slovakien, nämligen ungerskan, på ett sätt som fullständigt strider mot det europeiska tänkesättet.
Slovakiens språklag innebär en uppenbar diskriminering av rättigheterna för den ungerska befolkningsgruppen i landet, dit en halv miljon människor hör, att använda sitt eget språk.
I vissa fall kan personer dömas till böter på 5 000 euro.
EU har förpliktigat sig till att verka för kulturell och språklig mångfald. Till och med en kommissionsledamot för flerspråkighet har utsetts.
Europeiska stadgan för regionala språk och minoritetsspråk, som även Slovakien har ratificerat, utgör en garanti för medborgarnas rättigheter att använda sitt eget modersmål på alla utbildningsnivåer, för administrativa ändamål, på offentliga institutioner och i officiella handlingar.
EU-institutionernas enda stöttepelare kan inte tillåta att en av medlemsstaterna uppenbart strider mot grundläggande EU-normer och går till angrepp mot minoriteters rättigheter, utan att göra sin röst hörd.
(PL) För ett par månader sedan debatterade vi här i kammaren situationen inom den polska fartygsindustrin, och nådde en överenskommelse.
Martin Schulz, ordföranden för vår politiska grupp, intygade på vår grupps vägnar att parlamentet inte samtyckte till att tiotusentals arbetstillfällen på skeppsvarven och deras leverantörsföretag skulle försvinna.
Martin Schulz intygade att parlamentet inte samtyckte till att avskaffa denna industrigren i Polen, eller till att Europas industriella kapacitet stadigt minskar.
Sex månader har förflutit och nu är läget följande: Regeringen har inte kunnat privatisera skeppsvarven, kommissionen har inte tagit någon som helst hänsyn till parlamentets ståndpunkt, skeppsvarven har ingen produktion, framtiden är osäker och människorna har förlorat sina jobb och lämnats i ovisshet.
Nog måste vi alla vara överens om att kommissionen helt saknar uppfattning om en europeisk industripolitik och att den inte har insett att fartygen behövs - de har behövts tidigare, de behövs nu och de kommer att behövas även framöver.
(EN) Herr talman! Den 23 augusti 2009 inföll 70-årsdagen för den illa beryktade pakt mellan nazisterna och Sovjetunionen som en gång delade Europa.
Jag anser att detta är ett chockerande exempel på hur nära till synes motsatta politiska ytterligheter kan komma varandra.
Både Moskva och Berlin enades då om att det första steget vore att störta den demokratiska politiska ordningen i Europa. Både Moskva och Berlin ville få herraväldet över världen.
Följaktligen får vi inte glömma att det krävdes två diktatorer för att starta andra världskriget.
Fyra dagar innan Stalin undertecknade pakten förklarade han själva poängen för sina kamrater. Han sade att det låg i Sovjetunionens intresse att det utbröt krig mellan Tredje riket och det kapitalistiska anglo-franska blocket.
Allt skulle göras för att kriget skulle vara så länge som möjligt, för att de båda sidorna skulle bli utmattade.
Därefter skulle Stalin och hans anhängare ha en stor arena för att utveckla världsrevolutionen.
Jag vill påminna ledamöterna om Europaparlamentets resolution från april om att göra den 23 augusti till en gemensam minnesdag för att hedra offren för alla totalitära regimer.
(SK) Både under parlamentets förra session och under den nuvarande har vi hört anföranden från många ungerska parlamentsledamöter som kritiserar den slovakiska språklagen.
Jag vill samtidigt nämna att ni alla har skickat dokument med åtskilliga argument, som i de flesta fall är feltolkningar, förvrängningar eller rentav rena lögner, för att säga det rent ut.
Den slovakiska språklagen är fullt förenlig med alla mänskliga rättigheter och rättigheter som skyddar minoritetsspråk.
Enligt min mening är det en mycket farlig politik som de ungerska parlamentsledamöterna bedriver, genom att klart och tydligt provocera extremism, både i Ungern och i grannländerna omkring.
Jag tycker att de borde inse att denna politik är mycket farlig och sätta stopp för lögnerna, precis som vi har hört här tidigare i dag.
(SL) Jag har blivit ombedd av flera slovenska och italienska medborgare att uppmärksamma parlamentet på Italiens avsikter att bygga en gasterminal i Triestebukten.
Jag delar oron med de slovenska och italienska miljöorganisationerna över att denna gasterminal kan utgöra en stor börda för området, som redan är mycket miljökänsligt.
Jag tänker på Triestebuktens vatten och dess tätbebyggda inland.
Miljöorganisationerna har också framfört sina tvivel på att de handlingar som använts vid miljökonsekvensbedömningen har varit riktiga.
Jag uppmanar även den italienska och slovenska regeringen att samarbeta i det här projektet i enlighet med det samförståndsavtal som de undertecknade i september förra året.
Med andra ord så uppmanar jag dem att samarbeta vid alla miljökonsekvensbedömningar i norra Adriatiska havet, särskilt i Triestebukten.
Jag förväntar mig att regeringarna till följd av sådan miljökonsekvensbedömning kommer att enas om en bättre lämpad plats för denna gasterminal än Triestebukten.
(FI) Herr talman! Jag håller med min estniska kollega Siiri Oviir om att den ekonomiska krisen är långtifrån över.
En besynnerlig optimism framträder överallt i Europa, fastän arbetslösheten ökar, de nationella ekonomierna har skulder, befolkningen blir äldre och ett slags tredelad giljotin hänger över Europa. Trots allt detta förklaras lågkonjunkturen vara över.
En strategi för att ta sig ur krisen är under planering, vilket gör att vi inte behöver bry oss om att fortsätta med återhämtningsstrategin.
Europa började mycket bra med återhämtningsstrategin och med att ta sig an den ekonomiska krisen på ett exemplariskt sätt, i sådan utsträckning att Förenta staterna drog lärdom av EU och följde dess exempel. Men därefter har EU:s ansträngningar fullständigt stannat av.
Denna falska optimism leder även till felaktiga lösningar.
Än har den ekonomiska krisen inte övervunnits.
(RO) Bildandet av alliansen för europeisk integration, i kölvattnet efter de tidiga valen i juli 2009, bekräftar återigen de moldaviska medborgarnas positiva inställning till europeiskt engagemang.
Ett mycket viktigt steg har tagits, som Moldavien och EU inte har råd att missköta.
Den politiska situationen är fortfarande känslig.
Därför är framgångarna för alliansen, och indirekt för ett demokratiskt Moldavien, starkt beroende av stödet från dess europeiska partner.
Moldavien har åtagit sig att slå in på en EU-vänlig kurs och EU:s ansvar är att underlätta för Moldavien att följa denna kurs.
Även på politisk nivå är det nu tydligt att det moldaviska folket har valt det europeiska alternativet.
Vi måste därför ge vårt ovillkorliga stöd till alliansen för europeisk integration i Moldavien, eftersom den enda chansen att gradvis, men ändå snabbt, integrera landet i den europeiska familjen är genom alliansen.
Jag uppmanar kommissionen att förhandla om undertecknandet av en ny överenskommelse med Moldavien som en brådskande angelägenhet och att använda alla resurser som krävs för att hjälpa denna republik ut ur sin svåra finansiella situation.
(HU) EU:s trovärdighet undergrävs fullständigt om vi enbart uttalar oss om brott mot mänskliga rättigheter utanför EU och inte protesterar vid allvarliga överträdelser av mänskliga rättigheter inom EU, till exempel av de slag som precis har inträffat i Slovakien till följd av den nationella språklagstiftningen, och som har gett upphov till spänningar utan tidigare like mellan de största och minsta grupperna i samhället.
Minoritetsspråket har underordnats huvudspråket, som OSSE:s höge kommissarie för nationella minoriteter Knut Vollebæk har uttryckt det.
Jag vill påpeka för min kollega Boris Zala att vi gärna hade sluppit att ta upp den här frågan i Europaparlamentet.
Jag har gjort det enbart till följd av att en lag har trätt i kraft i Slovakien som innebär att minoritetsspråkens användning strikt begränsas och att den ungerska befolkning som lever där diskrimineras.
Därför hör det till nästa kommissions och ordförande José Manuel Barrosos ansvar att skapa forum där dessa fall kan undersökas, som Leonard Orban också har framfört i sin skrivelse.
Slovakien måste stå fast vid sina internationella åtaganden, ramkonventionen om skydd för nationella minoriteter och den europeiska stadgan om landsdels- eller minoritetsspråk.
(PL) Herr talman! Jag bad om ordet med hänvisning till uppdraget i Afghanistan.
Ett ämne som är svårt för alla inblandade och som påverkar både Nato och EU.
Jag vill särskilt uppmärksamma kravet på humanitärt, socialt och ekonomiskt bistånd till det afghanska folket, som tyvärr har varit utsatta för krig i 30 år.
Anledningen till att jag tar upp det här ämnet är en ökning av attacker mot soldater i samband med presidentvalet.
Som vi alla vet har dessa attacker blivit allt vanligare och våldsammare under valslutspurten.
Ett sådant bistånd är särskilt viktigt för att skapa förtroende och för att återuppbygga landet.
Kapten Daniel Ambroziński i den polska militärstyrkan förlorade nyligen livet i Afghanistan.
Det verkar som att hans död främst orsakades av brister hos den afghanska militären och polisen, vilka givit efter för mutor.
Det är välkänt att den afghanska armén och polisstyrkan befinner sig i en svår ekonomisk situation.
Enligt media tjänar afghanska soldater 20 US-dollar om de har tur.
Det är viktigt att den militära insatsen åtföljs av socialt, humanitärt och ekonomiskt bistånd.
Tjugo sekunder till Seán Kelly för en mycket kort kommentar.
(EN) Herr talman! Jag vill bara mycket kortfattat säga att ett felaktigt och något nedlåtande uttalande gjordes i kväll om Lissabonfördraget i Irland, av en brittisk kollega.
Ingen har tvingat Irland till att rösta om fördraget en andra gång.
Det var ett beslut som fattades av det irländska parlamentet, och kommer att verkställas av det irländska folket.
I själva verket har vi inte blivit tvingade till att göra någonting sedan vi vann vår självständighet från Storbritannien 1922.
Mina damer och herrar! Vi har haft 39 anföranden under 45 minuter.
Det anser jag vara en utmärkt prestation. Det har varit en bra debatt och jag vill framför allt gratulera de som har hållit sitt första anförande.
Jag vill särskilt betona vikten av att kommissionen tar hänsyn till kommentarerna i debatten, annars blir parlamentet bara en plats för att lufta åsikter.
Jag märkte att kommissionen var uppmärksam, och de kommer med all sannolikhet att göra en uppföljning av alla våra ledamöters kommentarer.
1.
Avtal mellan EG och Mongoliet om vissa luftfartsaspekter (
5.
Förslag till ändringsbudget nr 6/2009 (
Skogsbränderna sommaren 2009 (ingivna resolutionsförslag): se protokollet
8.
De institutionella aspekterna av inrättandet av den europeiska avdelningen för yttre åtgärder (
Herr talman! Jag vill lägga fram ett muntligt ändringsförslag till De gröna.
Om de godtar förslaget vill jag rekommendera att man röstar ”ja”.
Om vi inför meningen ”There should be no duplication of external service in the Council or in the European Council” rekommenderar jag att parlamentet röstar ja till detta.
(EN) Herr talman!
Vi skulle kunna rösta i block.
Jag föreslår att vi röstar från 56 till 28.
(Applåder)
Välkomsthälsning
Mina damer och herrar! Jag ber att få säga varmt välkommen till den delegation från senaten i Malaysia som sitter på åhörarläktaren.
Delegationen leds av Hans Excellens Datuk Wong Foon Meng, ordförande i senaten.
Jag vill upplysa om att Europaparlamentet och det malaysiska parlamentet har en regelbunden och givande kontakt.
Malaysias samhälle präglas av aktivitet, ekonomin blomstrar och landet har en viktig roll inom Sydostasiatiska nationers förbund (Asean).
Därför har jag och parlamentet nöjet att ännu en gång få välkomna våra vänner och kolleger från senaten. Vi hoppas att ni får ett mycket givande besök.
Öppnande av sammanträdet
2.
Statistik om bekämpningsmedel (
Jag vill bara förklara att det här är det sista av tre betänkanden om användningen av bekämpningsmedel.
Tidigare i år, under förra mandatperioden, antog vi en förordning om utsläppande av växtskyddsmedel på marknaden.
Vi antog då även ett direktiv om en hållbar användning av bekämpningsmedel. Föreliggande förordning om statistik om bekämpningsmedel är den tredje delen.
Detta förslag fick behandlas i förlikningskommittén eftersom någonting gick fel under förra mandatperioden.
Ett stort antal personer var inte där, och vid andra behandlingen närvarade alltför få personer för att få tillräckligt med röster för att slutföra den andra behandlingen.
Jag vill därför tacka det svenska ordförandeskapet och, framförallt det tjeckiska ordförandeskapet, eftersom de helt kunde ha förstört den andra behandlingen: De kunde ha vägrat att låta förslaget gå till förlikning.
Tack vare deras goda förbindelser med parlamentet, och tack vare ordförandena för de politiska grupperna som tillsammans med mig skrev ett brev till ordförandeskapet direkt efter valet, har det gått att rädda betänkandet och, genom förlikningsförfarandet, se till att vi idag kan rösta om texten i den form som vi kom överens om vid andra behandlingen.
Jag vill tacka alla inblandade.
2.
Avtal om tekniskt och vetenskapligt samarbete EG/Ukraina (
2.
För en politisk lösning beträffande piratverksamhet utanför Somalias kust (omröstning)
EU-instrument för mikrokrediter för sysselsättning och social inkludering (Progress) (debatt)
Nästa punkt är ett betänkande av Kinga Göncz, för utskottet för sysselsättning och sociala frågor, om förslaget till Europaparlamentets och rådets beslut om inrättande av ett EU-instrument för mikrokrediter för sysselsättning och social inkludering (Progress-instrument för mikrokrediter) - C7-0053/2009 -.
(FR) Fru talman! Jag noterade att ni under föregående debatt kallade den debatt som nu ska äga rum för en debatt om Progress-instrumentet.
Men enligt parlamentets beslut som bekräftats av talmanskonferensen kommer vi bara att rösta om instrumentet för mikrokrediter.
Därför tycker jag att det är viktigt att klargöra att den här debatten handlar om mikrokrediter och inte om Progressprogrammet.
Tack så mycket, fru talman! Jag är också tacksam för detta klargörande, eftersom det är oerhört viktigt att vi nu ska tala om mikrokreditinstrumentet.
Jag vill också hälsa kommissionsledamot Vladimír Špidla välkommen till den debatt som följer.
Inledningsvis vill jag säga att när jag blev föredragande för det här programmet trodde jag att jag skulle få en mycket enkel uppgift med tanke på det breda samförstånd och stöd som finns i frågan, något som också bekräftades under debatten.
Stödet har varit brett i många avseenden.
För det första kommer detta krishanteringsinstrument att hjälpa just dem som läget är mest hopplöst för, som har förlorat sitt arbete och som på grund av den ekonomiska krisen heller inte kan få lån eller stöd.
För det andra är det här ett exempel på instrument som inte ger folket fisk utan lär dem att fiska.
Det skapar just den sortens kreativitet som vi bäst behöver för att få ett positivt slut på krisen.
För det tredje ökar EU:s resurser, vilket enligt min uppfattning är en finansministers högsta dröm.
Vissa av resurserna är bidrag från Europeiska investeringsbanken och en del kommer från andra kommersiella banker, eftersom EU står för det primära risktagandet vilket underlättar för övriga aktörer att ta risker.
Som jag nämnt finns det ett brett stöd för innehållet i programmet.
Tack vare dessa tre aspekter tror jag att den fråga som ledde till debatt under diskussionerna med rådet och kommissionen hade att göra med vilka resurser EU ska använda i finansieringen av just detta primära risktagande.
Den andra tvistefrågan var storleken på de resurser som kan användas som stöd till vid inrättandet av instrumentet och som faktiskt kan förväntas dra till sig andra betydelsefulla resurser.
Rådet och kommissionen föreslog först att 100 miljoner euro skulle komma från Progressprogrammet, vilket främst syftar till att utarbeta åtgärder för att motverka socialt utanförskap och stödja lika möjligheter.
Vi i parlamentet har redan från början sagt att Progressprogrammet inte på något sätt får äventyras, eftersom det behövs mer än någonsin i den nuvarande krisen.
Vi godtar inte heller att man mixtrar så mycket med Progressprogrammet att hela programmet faktiskt kan sättas på spel.
Parlamentet har i högsta grad varit redo att kompromissa under debatten.
Vi har också fört tre informella trepartssamtal, varav ett pågick ända in på småtimmarna, där vi föreslår att vi skulle kunna tänka oss att laborera med Progressprogrammet, bara inte dess funktion äventyras.
Vi har föreslagit att vi med hänsyn till det ursprungliga förslaget till och med skulle kunna tänka oss att använda 100 miljoner euro i stället för 150 miljoner euro till att inrätta programmet.
I parlamentets budgetförslag för 2010 finns resurser på 25 miljoner euro, vilket gör det möjligt att sätta igång programmet redan i början av 2010, och dessa resurser är tillgängliga utan att man rör Progressprogrammet 2010.
Vi har också begärt att denna punkt ska avföras från dagens dagordning eftersom vi misslyckats med att komma överens om den.
En annan fråga som vi uppfattat som ett problem är att ordförandeskapet kom till trepartssamtalen utan mandat vid alla tre tillfällena, vilket gjorde det mycket svårt att överväga våra förslag på lämpligt sätt.
Jag tycker att det är viktigt att parlamentet röstar så snart som möjligt i denna fråga, kanske till och med den här veckan, så att projektet kan inrättas i början av 2010 med 100 miljoner euro i finansiering. På så vis förmedlas budskapet att detta är ett krishanteringsinstrument där snabbt agerande fyller en mycket viktig funktion.
Jag hoppas verkligen att kommissionsledamot Vladimír Špidla kan hjälpa oss att få kommissionen att återkalla sitt första förslag om att ta de 100 miljonerna från Progressprogrammet, så att programmet kan sättas igång så snart som möjligt.
ledamot av kommissionen. - (CS) Mina damer och herrar! Jag vill börja med att betona vikten av detta initiativ på området mikrokrediter.
I samband med den nuvarande krisen ökar arbetslösheten väsentligt i alla medlemsstater, vilket tyvärr leder till att de mest utsatta personerna i vårt samhälle drabbas värst.
Mikrokreditinstrumentet syftar särskilt till att hjälpa dessa grupper av medborgare att hitta annan sysselsättning och själva bli mikroentreprenörer.
Jag vill gratulera utskottet för sysselsättning och sociala frågor till det enastående arbete de åstadkommit på området, och i synnerhet välkomnar jag Kinga Gönczs bidrag till initiativet.
Jag är medveten om de insatser som gjorts i förhandlingarna mellan parlamentet och rådet i syfte att nå en överenskommelse vid första behandlingen.
Med hänsyn till att båda organen stöder mikrokreditinstrumentet har man kommit en god bit på väg med de grundläggande formuleringarna i förslaget.
Framgången återspeglas i hög grad av de ändringsförslag som lagts fram i dag.
Naturligtvis handlar den svåraste frågan om budgeten.
Även om båda organen antagligen kommer att godkänna en övergripande budget på 100 miljoner euro till detta instrument består det huvudsakliga hindret fortfarande i att hitta finansieringskällorna.
Som ni vet ingår förslaget till mikrokrediter i ett paket som innebär att 100 miljoner euro överförs från Progressprogrammet.
Ni har bestämt er för att inte rösta om detta andra förslag den här veckan.
Överföringen av medel från Progressprogrammet stöds av rådet och ses i många av medlemsstaterna som en grundläggande del av hela paketet.
Om vi inte enas om hur området ska finansieras kommer vi inte att nå målet om ett snabbt genomförande av instrumentet.
Men i dag diskuterar vi texten till det beslut som ska ligga till grund för instrumentet.
Slutligen vill jag ännu en gång hylla föredraganden för hennes arbete med betänkandet och ändringsförslagen som gör det möjligt för de båda lagstiftningsorganen att koncentrera sig det huvudproblem som återstår att lösa, nämligen finansieringen.
föredragande för yttrandet från utskottet för ekonomi och valutafrågor. - Fru talman! Om arbetslösheten ska kunna sänkas så måste EU tillsammans med medlemsländerna ta ett större ansvar.
Förslaget om mikrokrediter är ett initiativ där parlamentet varit pådrivande.
Det handlar om att ge arbetslösa en ny start och att öppna dörren till företagande för några av de mest utsatta grupperna inom EU, bland annat ungdomar.
Förslaget ska underlätta småskaliga investeringar och ge mikroföretag möjligheter att växa.
Efter en del smärre förändringar och förtydliganden fick förslaget ett brett stöd i utskottet för ekonomi och valutafrågor.
Den fråga som har skapat debatt är finansieringen, vilket också nämnts här.
Kommissionens förslag var att inga extra pengar skulle skjutas till utan att medlen skulle tas från programmet Progress.
Denna uppfattning delades dock inte av det ansvariga utskottet som någon felaktigt hävdat.
Detta är läget i dag.
Jag måste säga att jag tycker att det är konstigt att rådet så envist säger nej till vårt förslag om 150 miljoner under perioden - njuggt och snålt i dessa svåra tider!
för PPE-gruppen. - (HU) Herr kommissionsledamot, mina damer och herrar! Även vid tidigare debatter har vi upplevt att frågorna om den ekonomiska krisen, och hur vi ska ta oss ur den, engagerar oss alla och har fått stor uppmärksamhet.
I egenskap av samordnare från Europeiska folkpartiets grupp (kristdemokrater) i utskottet för sysselsättning och sociala frågor vill jag bara bekräfta vårt stöd till en av de frågor som är viktigast för oss i vart och ett av de dokument som framlagts, nämligen att trygga sysselsättningen och skapa nya arbetstillfällen.
Låt mig påminna er om att Europeiska folkpartiets grupp (kristdemokrater) länge har varit positiv till mikrokrediter.
Det var faktiskt min före detta kollega Zsolt Becsey som i sitt initiativbetänkande 2009 var först med att ta upp ämnet i parlamentet.
Det byggde på Ungerns tidigare och dåvarande erfarenheter av det instrument som kallades Széchenyi-kortet och hade samma syfte som i nuläget, nämligen att ge små kortfristiga lån till mikroföretag.
Låt oss tänka på slaktare, bagare, grönsakshandlare eller kanske till och med apotekare.
De påverkas också av krisen.
Enormt många människor är anställda i dessa företag.
I vissa länder finns så många som 90 procent av de anställda inom denna sektor.
Så är det t.ex. för mer än 90 procent av företagen i Ungern.
De behöver inga stora belopp, och de vill heller inte betala några höga räntor.
I vissa fall behöver de tillfälliga driftskrediter och tillfälligt stöd.
I kommissionens förslag tar man upp just detta problem och som föredraganden sagt finns det verkligen ett brett stöd och samförstånd bakom förslaget.
Därför tycker jag att det är viktigt att vi också enas om finansieringen så snart som möjligt.
Vi stöder även de 35 förslag som Europeiska folkpartiets grupp (kristdemokrater) lagt fram tillsammans med socialdemokraterna, liberalerna och de konservativa, eftersom vi anser att villkoren då är uppfyllda för att vi ska kunna godkänna instrumentet vid första behandlingen och införa det så snart som möjligt.
Fru talman! Jag är ganska förvånad.
Vi ska anta ett instrument som är ett innovativt redskap, ett nödvändigt redskap, för att hjälpa dem som drabbats hårdast av krisen att hantera den och skapa sina egna jobb i framtiden.
Det här instrumentet ska antas genom medbeslutandeförfarandet, men rådet är inte närvarande.
Det måste vara därför som rådet inte har något att säga oss i frågan och inte anser sig vara förbundet till Europaparlamentets ståndpunkt.
Det är i vart fall är det intryck som vi har fått vid flera tillfällen under förhandlingarna.
Europaparlamentet kommer att ta sitt ansvar.
Tack vare samarbetet och den konstruktiva dialogen mellan alla grupperna kan vi anta mikrokreditinstrumentet, vilket är på ett konsekvent sätt hänger samman med åtgärderna under många år, vilket Csaba Őry påmint oss om.
Men jag vill också framhålla de pilotprojekt som vi har tagit initiativ till.
Vi vet att de mest utsatta i detta krisläge, nämligen de som inte kan finansiera sin verksamhet med lån från de stora bankerna, med hjälp av detta redskap kan utveckla sina egna strategier och på sätt och vis sina egna jobb.
Jag ska inte upprepa innehållet i, förloppet för och räckvidden av de förhandlingar som har ägt rum.
Förhandlingarna hölls under lämpliga förhållanden.
Frågan om finansiering är svårare.
I samband med José Manuel Barrosos initiativ hösten 2008 att organisera Europas återhämtning betraktades det som viktigt att använda detta redskap för att förverkliga EU:s strategi.
Men kommissionen har föreslagit att vi enbart ska finansiera ett nytt projekt med pengar från att annat viktigt projekt som redan föreslagits.
Vi hade ett projekt som skulle gynna stödnätverk för de mest utsatta - Progressprojektet - och som det fanns ett starkt stöd för i parlamentet, men kommissionen föreslår nu att vi ska finansiera mikrokrediterna genom att helt enkelt ta av de resurser som avsatts till Progressprogrammet.
Det är denna nonchalans som parlamentet inte godtar, och det är därför som vi inte har slutfört förhandlingarna.
Det är därför som vi intar en ansvarsfull hållning och talar om att vi är redo att behandla vårt förslag under det spanska ordförandeskapet i början av januari: 40 miljoner euro tas från budgetmarginalerna och 60 miljoner euro tas från Progressprogrammet, med en omfördelning av 20 miljoner euro, så att bördan kan fördelas rättvist.
Sedan ska vi ta vårt ansvar i utskottet för sysselsättning och sociala frågor och se över hur ett sådant program kan genomföras i var och en av medlemsstaterna, så att samverkanseffekter skapas mellan de olika experiment som ska utföras i medlemsstaterna - det är vi säkra på - när paketet antas i sin helhet i januari.
för ALDE-gruppen. - (EN) Fru talman! Det är glädjande att få tillfälle att säga några ord om det föreslagna mikrokreditinstrumentet.
Tidigare talade vi om Europeiska fonden för justering för globaliseringseffekter och hur den kan användas till stöd för de anställda som blivit övertaliga i vissa sektorer.
Mikrokreditinstrumentet är en annan del av pusslet, där EU i detta fall försöker erbjuda mikrokrediter till dem som inte kan få sådana lån från det som brukar kallas finansinstitut i vanlig mening.
På så vis skulle entreprenörskap främjas och dessa personer skulle få möjlighet att starta egna företag.
I detta sammanhang är det glädjande att kunna konstatera att fonden kan förvaltas av kreditföreningar, kooperativa banker och andra gemensamma finansinstitut, eftersom de ofta står närmare dem som kan tänkas vilja få tillgång till just detta instrument.
Jag känner verkligen inte till förhållandena i andra länder, men i Irland är det bara kreditföreningsrörelsen som lyckats klara verksamheten utan pengar från skattebetalarna, och detta är ett icke-vinstdrivande institut som drivs av medlemmarna.
När vi talar om social inkludering inom ramen för EU:s socialpolitik måste vi se till att vi genom våra åtgärder integrerar social inkludering i de beslut vi fattar, och social inkludering står skrivet över hela det här programmet.
I samband med detta vill jag framföra hur oerhört besviken jag är över att vi efter tre trepartssamtal fortfarande inte kunnat enas om finansieringskällan till det här instrumentet.
Jag anser att det svenska ordförandeskapet inte verkade ha möjlighet att föra meningsfulla förhandlingar i frågan.
Jag vet inte hur det är med er, men som jag sade är jag mycket besviken över att det inte var mer än 40 miljoner euro fördelat på tre år och 27 medlemsstater som hindrade oss från att komma överens.
Uppenbarligen var det många finansministrar som inte ville ha någon riktig förhandling.
Jag kan inte rå för att jag tror att många av dessa ministrar gav miljarder i stöd till bankerna men inte kunde stödja andra finansinstitut, som skulle ge mikrokrediter till dem som förlorat sina jobb och som skulle få svårt att låna från samma banker som räddats med offentliga medel.
Fru talman, herr kommissionsledamot, mina damer och herrar! Mikrokrediter och småskaliga lån kan vara till hjälp för personer som inte anses kreditvärdiga på den vanliga lånemarknaden.
På så vis kan, vilket redan nämnts, även dessa personer starta företag och använda sina idéer till att skapa ett arbete.
Personer med denna förmåga kan ta sig ur en kris med hjälp av sådana lån.
Mikrokrediter är dessutom ett viktigt sätt att stödja samhällsekonomin.
Olika former av mikrokrediter har sedan 2000 varit ett erkänt sysselsättningspolitiskt instrument på lokal nivå i EU.
Och därför beslutade parlamentet klokt nog 2006 att medel från Europeiska socialfonden även ska kunna betalas ut i form av mikrokrediter eller räntesubventionerade lån, detta i enlighet med artikel 11 i förordningen om Europeiska socialfonden.
Men i Europeiska socialfonden finns 76 miljarder euro att tillgå, och med samfinansiering blir det 118 miljarder euro!
Om man bara skulle ta en tiondel av detta fick man 11 miljarder euro att använda i medlemsstaterna.
Men de används inte till mikrokrediter!
Därför har kommissionen genomfört en testperiod för mikrokrediter med hjälp av instrumentet Jasmine, även detta finansierat med EU:s strukturfonder.
Och eftersom det föll så väl ut ska ytterligare ett instrument inrättas efter detta, dock inte med hjälp av strukturfonderna, där det finns miljarder att tillgå, utan genom det minsta av alla EU:s program, nämligen fattigdomsprogrammet Progress, som bara omfattar 743 miljoner euro under en sjuårsperiod.
Det är avsett för icke-statliga organisationer som bygger upp nätverk i medlemsstaterna i syfte att skapa en lobbygrupp för de fattigaste av de fattiga.
Europeiska informationskontoret för romer finansieras till hälften av Progressprogrammet.
Verksamheten går ut på att bygga upp nationella och regionala informations- och rådgivningskontor och att ge den romska minoriteten en röst, särskilt i de östeuropeiska staterna.
De gröna/Europeiska fria alliansen kommer inte att godkänna instrumentet om parlamentet gör som rådet vill och kallar detta för ett Progress-instrument enligt de kompromisser som föreslås av Europeiska folkpartiets grupp (kristdemokrater), Progressiva alliansen av socialdemokrater och demokrater i Europaparlamentet samt Alliansen liberaler och demokrater för Europa.
Sådana trolleritrick går inte an - att först ta pengar från de fattiga och sedan betala ut ...
(Talmannen avbröt talaren.)
för ECR-gruppen. - (CS) Mina damer och herrar! I det finansiella och ekonomiska krisläge som fortfarande råder behövs det inte bara stöd till banker och storföretag utan även till småföretag och egenföretagare.
Vi är alla medvetna om att det är i dessa småföretag, bland annat familjeägda företag, som det skapas och finns ett stort antal arbetstillfällen.
Vi stöder det nya finansieringsinstrumentet för mikrokrediter för sysselsättning och social inkludering, som i samarbete med Europeiska investeringsbanken ska göra det lättare att få lån för just egenföretagare, nystartade småföretag och familjeföretag.
Vi samtycker till förslaget om att satsa 100 miljoner euro på att trygga dessa småskaliga lån under en begränsad period.
Vi ser programmet som ett effektivt och bra instrument för en aktiv sysselsättningspolitik och som ett bra sätt att använda så kallade EU-pengar, med andra ord våra pengar.
Vi ger vårt fulla stöd till att de resurser som behövs för detta finansieringsinstrument tas från de medel som ursprungligen var avsedda för Progressprogrammet.
Vi håller inte med om att mikrokreditinstrumentet bör finansieras med reserver eller med medel från andra budgetposter.
Medlen i Progressprogrammet uppgår till 700 miljoner euro, om jag inte missminner mig, och används till att bygga upp nätverk för undersökningar och analyser.
Inga av Progressprogrammets resurser har öronmärkts för direkt stöd till personer som söker jobb eller skapar arbetstillfällen.
Jag tvivlar inte på att man behöver bygga upp nätverk och göra analyser och undersökningar.
Men i det svåra läge som råder för entreprenörer och arbetstagare bör man prioritera att använda EU:s budgetmedel till program riktar sig direkt till arbetsgivare och arbetstagare.
för GUE/NGL-gruppen. - (DE) Fru talman, mina damer och herrar! Ett mikrokreditinstrument för arbetslösa, för dem som riskerar att bli arbetslösa och framför allt för dem som inte har tillgång till den vanliga kreditmarknaden visar på goda avsikter och stöds i princip av vår grupp.
Men det som kommissionen och rådet hittills har åstadkommit i frågan är helt enkelt otillräckligt och i vissa avseenden fel, och vår grupp kan inte stödja det.
För det första är vi kritiska till det totala belopp som anslås.
Det totala anslag som föreslås är inte rimligt för ett program för bekämpning av arbetslöshet, och det kan knappast kallas mikrokreditprogram - det är i bästa fall ett nanokreditprogram!
För det andra är vi av principskäl mot denna typ av trolleritrick som inte har den minsta effekt och som finansieras på bekostnad av andra program och därför bara rinner ut i sanden.
För det tredje anser vi att det absolut behövs mentorskap och vägledning för att den här typen av program ska lyckas och vara hållbart.
Många nystartade företag misslyckas, särskilt i samband med mikrokrediter, och detta måste man ta hänsyn till i programmet.
För det fjärde måste man se till att betalningen av sociala avgifter i medlemsstaterna inte upphör för dem som drar nytta av programmet, annars får det ingen effekt.
Arbetslösheten går inte att bekämpa långsiktigt på detta sätt.
Vi säger nej till programmet i dess nuvarande form.
Fru talman, mina damer och herrar! Det förslag till beslut som Europaparlamentet och rådet har lagt fram om att inrätta ett europeiskt instrument för mikrokrediter på området sysselsättning och social inkludering är i grunden ett förslag där det ursprungliga Progressprogrammet anpassas till den ekonomiska verklighet som råder i ett Europa märkt av den finansiella och ekonomiska krisen.
Kommissionen föreslår stöd i form av mikrokrediter till småföretag som stimulansåtgärd för att upprätthålla och öka sysselsättningen i krisdrabbade regioner.
Men för att nå detta mål måste vi se till att de ekonomiska resurser som satsas inte går till sociala förmåner eller konsumtion.
De får endast gå till vettig och hållbar företagsverksamhet genom tillämpning av objektivt mätbara kriterier och förfaranden öppna för insyn.
Därför är det mycket viktigt att kräva att de slutgiltiga långivarna gör en noggrann utvärdering av ansökarnas affärsplaner, riskerna i samband med det affärsprojekt som presenteras och även av avkastningen på investeringarna.
Därför tycker jag att det är ytterst viktigt att stödja och komplettera de ändringsförslag som lagts fram av utskottet för ekonomi och valutafrågor, som ger vettiga ramar åt kommissionens förslag.
(FI) Fru talman, herr kommissionsledamot, mina damer och herrar! Det framstår som märkligt att det skulle finnas motstånd i parlamentet mot det här utmärkta och viktiga programmet med tanke på att läget på arbetsmarknaden blir allt sämre.
Prognosen om att ytterligare tio miljoner människor kommer att vara utan arbete i Europa nästa år och att svårare tider väntar dem som har sämre status på arbetsmarknaden.
Dessa uppgifter stärker skälen att investera i entreprenörskap.
Det är alltid de nystartade företagen som har störst svårigheter att få banklån.
Exempelvis är mer än 93 procent av företagen i Finland mikroföretag med färre än tio anställda, och ändå sysselsätter dessa småföretag 46 procent av den förvärvsarbetande befolkningen.
Därför är det inte mer än rätt av EU att inrätta ett instrument för mikrokrediter som svar på sysselsättningskrisen och på så vis även stödja enskilda medlemsstaters program med samma mål.
Men jag vill betona att det krävs en övergripande strategi för det här programmet.
De system för sociala förmåner, semester och pension som gäller i småföretagen behöver också utvecklas i linje med övriga sektorer.
I Europa råder det särskilt brist på högriskfinansiering och sådana personer, affärsänglar, som är beredda att investera i företag som befinner sig i ett tidigt skede.
Dessutom bör man på alla utbildningsnivåer stödja entreprenörskapsutbildning och kontakter med arbete och sysselsättning, och det bör finnas mer av seminarier och företagskuvöser för unga och mer resurser till sådant.
Mikrokrediter fungerar bara som en komponent i den här typen av övergripande strategi, som skapar verkliga tillfällen till en framgångsrik och vinstbringande verksamhet för nya småskaliga entreprenörer och hela den miljö de verkar i.
(EN) Fru talman! Jag välkomnar verkligen detta initiativ.
Arbetslösheten är det största problemet vi står inför just nu, och allt vi kan göra för att lindra dess effekter är viktigt för välståndet i våra samhällen.
Men jag tycker att det med tanke på den ökande arbetslösheten saknas tillräckliga ambitioner i förslaget om att tillföra 100 miljoner euro under en treårsperiod.
Likaså är jag förvånad över att de pengar som föreslås inte är nya pengar, så att följden blir att vi tar av det ena för att betala det andra, vilket redan har sagts, nu när alla resurser som finns i Progressprogrammet bör användas enligt den befintliga planen.
Vi måste göra allt vi kan för att snabbt komma överens under det spanska ordförandeskapet, så att programmet kan sättas igång snarast möjligt.
Rådet har lika stort ansvar för att enas och ta hänsyn till parlamentets synpunkter.
Det här är inte rätt tillfälle för rådet att köpslå om småsummor.
(Talaren godtog en fråga ställd i enlighet med blåkortsförfarandet i artikel 149.8 i arbetsordningen.)
(EN) Herr De Rossa! Har ni tänkt på att arbetslösheten i Irland har oerhört mycket att göra med Irlands medlemskap i valutasamarbetet, vilket innebär att Irland varken kan devalvera, sänka räntesatserna eller införa några kvantitativa lättnader?
Har ni aldrig tänkt på att det kanske vore bättre om Irland gick ur valutasamarbetet i stället för att sträcka ut en tiggande hand mot de EU-länder som bidrar?
(EN) Fru talman! Jag har inte alls några problem med att svara på det vanliga struntpratet från den yttersta högern i parlamentet.
Utan euron skulle Irlands ekonomi befinna sig i helvetet.
Som jag sade tidigare är det inte rätt tillfälle för rådet att köpslå om småsummor med tanke på jobbkrisens omfattning och den totala budgetens storlek, särskilt med tanke på det stöd som medlemsstaterna och Europeiska centralbanken gett till banksektorn - en banksektor som händelsevis inte vill låna ut till de personer som vi försöker hjälpa.
Jag tror helt och fullt på att vi kan komma överens utifrån föredragandens pragmatiska ansats, om rådet visar vilja till samförstånd.
Jag hoppas verkligen att det sker snabbt.
(PL) Fru talman, herr kommissionsledamot! I ljuset av den här debatten bör vi fästa uppmärksamheten vid att man i kommissionens strategi helt och hållet bortser från sysselsättningen inom sjöfartsekonomin.
Avsaknaden av en samordnad havspolitik har i många år varit orsaken till denna sektors systematiska sönderfall i EU, trots att vi borde tänka på att det är en enorm arbetsmarknad.
Dessutom ger kommissionen inte heller något stöd till den marginaliserade varvsindustrin, som i princip är utslagen i Europa till följd av den dumpningspolitik som förs av länderna i Fjärran östern.
Bara i mitt hemland, Polen, har kommissionens åtgärder lett till att varvsindustrin har kollapsat och att tusentals personer som var sysselsatta i sektorn förlorat sina jobb. Dessutom har det lett till nästan 80 000 indirekt förlorade arbetstillfällen.
Men denna sektor kommer inte att försvinna från världsekonomin.
I enlighet med de senaste årens utveckling kommer den att flytta till länderna i Fjärran östern på bekostnad av arbetstillfällen i Europa.
Det är extremt riskfyllt att inte ha en strategi för hur man ska återföra fartygen till sina nationsfärger.
Den här politiken leder till enorma oåterkalleliga inkomstförluster för Europa, pengar som i stället strömmar till skatteparadisen.
En annan mycket viktig del av kommissionens politik är fisket, som för ovanlighetens skull är den enda sektor som gynnar icke-industrialiserade områden i EU.
Kommissionen koncentrerar sig främst på att minska storleken på fiskeflottorna, men misslyckas samtidigt med att förhindra massimport till EU från Fjärran östern, exempelvis av hajmal som har mycket negativa effekter.
I dessa kristider måste kommissionens politik vara utgångspunkten för ekonomins utveckling och inte någon snabbåtgärd mot följderna av en felaktig strategi.
(PT) Fru talman, herr kommissionsledamot, mina damer och herrar! Jag vill gratulera föredraganden till hennes arbete med det här betänkandet och till det anförande hon gjorde nyss.
Det nya mikrokreditinstrumentet gör det möjligt att bevilja mikrokrediter till småföretag och personer som har förlorat sina jobb och vill starta sin egen verksamhet och skapa sina egna jobb.
Det är mycket viktigt nu när den ekonomiska krisen väntas leda till 3,5 miljoner förlorade arbetstillfällen bara i EU.
I och med den ekonomiska nedgången har bankerna slutat bevilja lån för att starta företag och skapa jobb, och det har blivit svårare att få lån just när det skulle behöva vara lättare.
Men det nya mikrokreditprogrammet kommer att vända den nuvarande trenden med begränsat kreditutbud, så att det blir lättare att skaffa resurser för att starta företag och skapa nya arbetstillfällen.
Kommissionen föreslår att 100 miljoner euro överförs från Progressprogrammets budget till detta finansieringsinstrument.
Vi instämmer inte med det förslaget.
Den finansiella och ekonomiska krisen är också en social kris.
Att ta resurser från Progressprogrammet, som riktar sig till de mest utsatta grupperna, är verkligen inte den lämpligaste lösningen.
Därför förordar vi att man skapar en egen budgetpost för att finansiera instrumentet samt ökar anslaget till 150 miljoner euro.
Vi håller också med om behovet av att göra det tydligare i själva lagstiftningen att målgruppen är alla utsatta grupper som har svårt att komma in på eller komma tillbaka till arbetsmarknaden och som riskerar att drabbas av socialt utanförskap.
Hänvisningen till specifika grupper bör därför strykas.
Slutligen vill jag betona att det är nödvändigt att de som får ekonomiskt stöd även bör få lämplig utbildning.
Den djupa ekonomiska krisen har mycket allvarliga effekter på sysselsättningen, med många arbetstagare som riskerar att förlora sina jobb samtidigt som det finns massor av unga som inte kommer in på arbetsmarknaden. Mot bakgrund av detta är det nödvändigt att EU och medlemsstaterna vidtar åtgärder, med hjälp av både övergripande strategier och riktade instrument.
Mikrokreditinstrumentet är just ett sådant riktat instrument, vilket syftar till åtgärder för alla dem som står utanför bankernas kreditmarknad och har svårigheter att komma in på arbetsmarknaden men som vill starta ett projekt, en ekonomisk verksamhet, vilket kan leda till egen försörjning och därmed bidra till den allmänna tillväxten.
Om vi vill att mikrokreditinstrumentet ska vara effektivt och ge varaktiga resultat är det särskilt viktigt att medlemsstaterna förbereder sig tillräckligt och bland annat skapar förbindelser på lokal administrativ nivå, där man har närmare kontakt med konkreta sociala krisförhållanden, och spelar en aktiv roll i att göra det nya instrumentet lättillgängligt.
Det är viktigt att betona att de långsiktiga effekterna av verksamheter finansierade genom mikrokreditinstrument och möjligheten att nå fullständig social integration i stor utsträckning är beroende av att det samtidigt finns väglednings-, mentors- och utbildningsprogram som måste samordnas med mikrokrediterna.
Mot bakgrund av de mål som ska nås med hjälp av mikrokreditinstrumentet är det nödvändigt att samtidigt betona en avgörande åtgärd, nämligen aktivt främjande av att män och kvinnor får lika tillgång till mikrokreditprogrammen.
Det är faktiskt kvinnor som är särskilt missgynnade när det gäller tillgång till såväl arbetsmarknaden som den konventionella kreditmarknaden.
Generellt sett är det betryggande att se att parlamentet är enat och ställer sig positivt till mikrokrediter och negativt till en sådan socioekonomisk bakgrund som denna.
Det är upp till rådet och medlemsstaterna att visa att de är seriösa och engagerade och staka ut riktningen så att det ekonomiska läget kan vändas rätt.
(ET) Fru talman, herr kommissionsledamot, mina damer och herrar! Kommissionen har lagt fram ett förslag om att skapa ett nytt finansieringssätt - mikrokreditinstrumentet.
Initiativet är viktigt och bra, men man har föreslagit att medlen till detta ska tas från Progressprogrammet, som redan är igång, och detta är inte godtagbart.
Jag vill påminna rådet och kommissionen om att vi inte blev valda till det här parlamentet för att vara en gummistämpel.
I slutet av 2006 när vi antog Progressprogrammet här i parlamentet satte medlemsstaterna upp sina respektive mål och började arbeta.
Programmet fick mycket gott resultat, och det finns ingen anledning att tro att programmet därför inte kommer att pågå som planerat till 2013.
Programmet har varit och är ämnat för de grupper som befinner sig i en ogynnsam situation, och de har kunnat få hjälp genom detta program.
Nu håller den ekonomiska krisen på att utvecklas till en social kris.
Arbetslösheten ökar månad för månad, och Progress-åtgärderna behövs även nu.
Men på samma gång går kommissionen vidare med sitt önskemål om att minska medlen till dessa åtgärder som fortfarande är under genomförande.
Det är ett oansvarigt och oacceptabelt tillvägagångsätt.
Jag är säker på att vi i parlamentet inte kan godkänna mikrokreditinstrumentet förrän det står klart varifrån pengarna till dessa åtgärder ska tas, inte förrän det står klart att medlen ska komma från annat håll än från de planer som är ämnade för alla dem som har det svårt.
(LV) Fru talman! Effekterna av den globala ekonomiska krisen är fortfarande påtagliga i medlemsstaternas ekonomier, men det är unga entreprenörer och chefer för småföretag som drabbas hårdast av krisen.
Deras affärsidéer får för närvarande inget stöd från långivarna.
Den ekonomiska tillväxten sker i samband med att det skapas nya jobb. Nya jobb skapas när företagen får tillgång till finansiering för att förverkliga sina idéer.
I det här krisläget vill bankerna tyvärr inte låna ut pengar till företagen eftersom de är rädda för att ta risker.
Det privata kapitalet har alltså sinat.
Under sådana förhållanden brukar det vara mikroföretag och unga entreprenörer som drabbas hårdast.
De har idéer om utveckling men saknar finansiering, och det är uppenbart att om dessa företag inte kan utvecklas kommer inga nya jobb att skapas. Men det krävs nya jobb för att vi ska kunna resa oss ur den ekonomiska krisen.
En lösning på problemet är EU-instrumentet för mikrokrediter, som ska ge 100 miljoner euro till utveckling av mikroföretag och nya företag genom omfördelning av medel från befintliga finansieringskällor.
I motsats till de stora stimulanspaketen, som man under det senaste året har inrättat huvudsakligen för att rädda det finansiella systemet som sådant, är det här programmet riktat direkt till entreprenörerna och inte till bankerna.
Det innebär att man låter pengarna gå raka vägen för att hjälpa till att skapa nya jobb och stimulera realekonomin.
Jag uppmanar mina kolleger i parlamentet att inte tveka inför beslutet att inrätta det här mikrokreditprogrammet.
Medlemsstaterna befinner sig i kris nu.
Europa behöver nya jobb nu. Stödet till nya initiativ från entreprenörer behövs omedelbart.
(EL) Fru talman! Bara det faktum att alla politiska grupper samtycker till och är överens om EU-instrumentet för mikrokrediter för sysselsättning och social inkludering visar hur nödvändigt det är.
Det är mycket viktigt att den som har förlorat jobbet, eller riskerar att förlora det, och inte kan hitta en lösning på problemet på de vanliga bankmarknaderna får tillgång till ett mikrolån eller en mikrokredit.
Men för att idén om mikrokrediter ska fungera i praktiken måste den fungera korrekt och genomföras snart. Det innebär att vi på torsdag när vi röstar om budgeten för 2010 måste säga ja till de första 25 miljonerna som ska komma ur budgeten.
Men det räcker inte.
Jag anser att det behövs ytterligare 75 miljoner ur budgeten. Att ta pengar från Progressprogrammet vore som att ta från dem som är mindre fattiga och utsatta för att ge till dem som är fattigare och mer utsatta.
Det skulle innebära att instrumentet med mikrokrediter i grunden hade upphört som koncept.
Man bör ha i åtanke att Progress betyder framsteg med att utveckla Europas sociala dimension. Om det inte sker och pengarna tas från Progressprogrammet har vi tagit ett steg tillbaka.
Det är just därför som jag tycker att rådet ska anta Europaparlamentets ståndpunkt.
(BG) Fru talman, mina damer och herrar! EU har antagit ett antal olika åtgärder för att bekämpa den ekonomiska krisen i över ett år nu.
Till skillnad från övriga åtgärder syftar mikrokreditinstrumentet faktiskt till att hjälpa de mest utsatta grupperna i samhället, som har svårt att komma in på eller komma tillbaka till arbetsmarknaden.
Solidaritetstanken, som är en av EU:s grundprinciper, kräver att de ägnas särskild uppmärksamhet.
Det finns nu ett stort intresse för det här instrumentet, särskilt i Bulgarien, och jag antar att det är likadant i övriga länder också.
Jag har hållit mig informerad i frågan ända sedan debatterna inleddes, och många företrädare följer utvecklingen i medierna.
Det ligger i EU-institutionernas intresse att visa EU:s medborgare att det är vår omedelbara uppgift att se till dem som påverkas av krisen och till samhällets fattigaste medborgare.
Det kommer att göra medborgarna övertygade om att institutionerna är effektiva och står nära dem.
Det råder vissa tvivel om huruvida instrumentet kommer att nå ut till och vara till nytta för dem som det är avsett för.
Det råder en oerhört stor brist på kapital att låna, vilket har bidragit till den ökade arbetslösheten.
100 miljoner euro räcker inte för att hjälpa alla som saknar arbete att hantera risken för socialt utanförskap.
Det är trots allt inte alla som har förmåga att utöka ett företag. Det är inte alla som kan få utbildning.
Det viktiga är att beslutet fattas snabbare och att mikrokreditinstrumentet börjar verka i så stor omfattning som möjligt, så att de som har idéer och näsa för företagande kan sätta igång nu när det fortfarande råder en allvarlig kris.
Nästa år har utsetts till Europaåret för bekämpning av fattigdom och socialt utanförskap, så låt oss vidta lämpliga åtgärder och inte försena återhämtningen.
(DE) Fru talman, mina damer och herrar! Vi kan utan tvekan se lovande tecken på att ekonomin och finansmarknaderna kommer att stabiliseras under 2010, och jag vill också påminna er om att detta endast varit möjligt genom samordningen på EU-nivå.
Men vi ser naturligtvis stigande arbetslöshetstal och vi måste utgå ifrån att de fortsätter att stiga under nästa år. Därför välkomnar jag det nya finansieringsinstrumentet för personer som vill starta en egen verksamhet.
Det är ju allmänt känt att arbetstillfällen skapas i små och medelstora företag.
I många år har vi diskuterat ekonomiskt stöd till dessa företag.
Men varje år har vi upptäckt att medlen inte går till de ändamål de var avsedda för.
Jag hade möjlighet att ta del av ett slutfört pilotprojekt förra veckan, men jag hann inte ta med erfarenheterna av detta i det här betänkandet.
Därför vill jag berätta om det här.
Deltagarna i pilotprojektet var egenföretagare eller ville bli egenföretagare, och dessa fick vägledning i ett år på vägen mot en egen verksamhet.
Det var så framgångsrikt att jag uppmanar till det tas med i det här projektet, med andra ord att man inom projektet inte bara tillhandahåller finansiering för dem som ska starta eget företag, utan även för dem som stöder dessa personer.
Detta är nödvändigt eftersom bankerna, som ju inte ger några lån, ändå ser en viss risk i detta avseende.
Jag tror att man kan utjämna den risken med hjälp av detta stöd.
Det andra som nämndes gång på gång i diskussionerna om detta var att vi inte får sätta en undre gräns för lånen.
Hittills har man bara kunnat ta lån på minst 5 000 euro.
Personerna behöver inte alltid så mycket.
Då räcker det med mycket mindre belopp, och det bör vi ta hänsyn till i det här programmet.
(LT) Jag vill understryka att en av EU:s viktigaste uppgifter för närvarande är att hejda den massarbetslöshet som orsakats av den utdragna passiviteten och den sociala krisen.
Det är olyckligt att vi inte lyckades komma överens om mikrokrediter som finansieringsform under trepartssamtalen.
Under denna socialt och ekonomiskt sett svåra period skulle det vara en otillfredsställande att som i kommissionens förslag omfördela 100 miljoner euro från Progressprogrammets budget, eftersom man på så vis inte minskar det sociala utanförskapet för de mest utsatta grupperna.
Jag är övertygad om att mikrokreditinstrumentet blir mer effektivt och ändamålsenligt om man samordnar det med nationella, regionala och lokala program och avsätter tillräckliga resurser.
Det är också viktigt att ta hänsyn till att den sociala välfärden i EU är direkt kopplad till sysselsättningen och möjligheterna att hitta ett arbete.
Därför föreslår jag att kommissionen inte bara ska ta hänsyn till dem som riskerar att förlora sina jobb utan även till dem som har svårigheter att komma in på eller komma tillbaka till arbetsmarknaden.
Det fanns även före den ekonomiska recessionen många utbildade och hårt arbetande medborgare som inte hade några egentliga möjligheter att få anställning, och därför flyttade många av dem från EU.
När det gäller de socialt utsatta uppmanar jag kommissionen och rådet att tänka på att det finns fler socialt utsatta grupper än ungdomar, exempelvis kvinnor, personer med funktionsnedsättning och äldre, som behöver säkrad sysselsättning.
Det finns alltså inget annat sätt än att skaffa ytterligare medel till mikrokreditinstrumentet.
(Talaren godtog en fråga ställd i enlighet med blåkortsförfarandet i artikel 149.8 i arbetsordningen.)
(DE) Fru talman! Vi har nu lyssnat till tre eller fyra talare ur gruppen Progressiva förbundet av socialdemokrater och demokrater i Europaparlamentet.
Dessa har sagt att de inte vill ta några pengar från Progressprogrammet. Men enligt ändringsförslagen ska det kallas Progress-instrumentet och Pervenche Berès har även sagt att 60 miljoner euro ska tas från Progressprogrammet.
Det är två tredjedelar!
Jag skulle vilja veta hur socialdemokraterna egentligen ställer sig i frågan.
Ska instrumentet finansieras genom Progressprogrammet - ja eller nej?
(LT) Jag skulle vilja svara att den bästa lösningen vore att skaffa ytterligare medel, eftersom Progressprogrammet i grunden riktar sig till samma grupper och detta skulle innebära att effekten säkerligen uteblir om det inte tillkommer några resurser.
Låt oss därför sätta oss ner och tillsammans komma fram till en lösning, för arbetslösheten håller på att nå en smärtsam nivå och det drabbar verkligen många som redan har det svårt.
(EN) Fru talman! Tre och en halv miljon människor i EU blev av med sina jobb det senaste året.
Det går inte att förändra läget med 100 miljoner euro.
Om man ser till att hundra miljoner människor är sysselsatta i små och medelstora företag blir det bara en euro per anställd.
Men det är i alla fall en början som bör välkomnas, eftersom finansieringen för närvarande är det största problemet, som kommissionsledamot Vladimír Špidla påpekade.
Ett exempel på detta är en situation som jag fick kännedom om i helgen. Ett företag drabbades av att en betydande order försenades med tre månader och ansökte om ett brygglån i den bank som företaget hade gjort affärer med i 15 år.
Ansökan avslogs.
Företagets chef fick beskedet att lånet bara skulle beviljas om han använde sin egen privata bostad som säkerhet.
Det gjorde han, och en vecka senare fick han ett brev där man återkallade brygglånet med anledning av att de nu befann sig i en högrisksituation.
Följden blev att företaget fick läggas ned och ytterligare tio personer blev övertaliga.
Det får mig att hålla med min kollega Marian Harkin om att dessa medel så långt det är möjligt bör gå till icke-kommersiella banker som kreditföreningar, som åtminstone i mitt land finns i alla städer och gör ett enastående arbete, detta eftersom alla dessa berättelser tyder på att de kommersiella bankerna inte lånar ut ens de resurser som de fått från Europeiska investeringsbanken utan i stället behåller dem för att stärka sin egen ekonomi.
Av dessa två skäl tycker jag att vi bör vara mycket mer noggranna med var pengarna hamnar än med varifrån de kommer.
Om de hamnar hos rätt personer är det de mest välplacerade pengarna på länge här på EU-nivå.
Slutligen vill jag kommentera greve Dartmouths tämligen obetänksamma uttalande om den tiggande handen.
Det handlar inte om en tiggande hand.
Det handlar om att hjälpa dem som kan hjälpa andra att skapa sysselsättning och behålla sitt arbete.
Vi är mycket stolta och glada över att vi gick med i valutasamarbetet, och vi tänker stanna kvar.
(FR) Fru talman! Enligt klausulen om socialpolitik i Lissabonfördraget måste EU ta hänsyn till sysselsättningen, det sociala skyddet och kampen mot social utslagning.
Den ekonomiska och finansiella kris som drabbat Europa har lett till en mycket allvarlig kris för människorna och samhället, och det är omöjligt att bedöma konsekvenserna för tillfället.
Hittills har huvuddelen av insatserna syftat till att stabilisera bankerna och förhindra konkurser.
Förutom åtgärder för att förhindra arbetslöshet måste vi skapa ett instrument som ger ny stimulans till den ekonomiska tillväxten i EU.
Det instrument som kommissionen använder är utformat för att skapa en infrastruktur som i sin tur ska göra det möjligt för medborgarna att arbeta.
I praktiken är det möjligt att byta en tillfällig strategi mot en långsiktig strategi.
Detta instrument måste inrättas snabbt, i januari 2010.
Vår debatt i dag och våra beslut når fram till många människor som drabbats av ojämlikhet och många ungdomar som vill komma ut i arbetslivet och som vi bara borde ge en hjälpande hand.
Jag vill återigen nämna det förslag som redan lagts fram om att skapa en enskild budgetpost på 50 miljoner euro för det här instrumentet.
Det skulle ge cirka 6 000 europeiska entreprenörer möjlighet att starta företag, utveckla dem och på så vis skapa nya jobb.
Det viktigaste är dessutom att vi förbättrar tillgången till resurser och framför allt ger bättre information till medborgarna om alla de projekt som de kan ansöka om.
(PL) Fru talman! Hundratusentals européer har drabbats hårt av följderna av den ekonomiska krisen, för de har förlorat sina jobb.
Arbetslösheten har ökat i alla EU-länder och det är denna del av krisen som drabbar våra medborgare värst.
Den hjälp som behövs når fram till finansinstituten.
Olyckligtvis når hjälpen inte fram i tid till dem som riskerar att bli av med jobbet, och det är de som kommer att känna av den pågående krisen under längst tid.
Därför är även jag glad över inrättandet av EU-instrumentet för mikrokrediter för sysselsättning och social inkludering.
Det är särskilt värt att påpeka kombinationen av detta instrument med det allmänna målet om stöd till entreprenörskap.
De medel som tillförs genom detta instrument kommer att stimulera till nya företag.
Det är goda nyheter för vår ekonomi, eftersom den bygger på de små och medelstora företagen, och det är i de små och medelstora företagen som jobben skapas.
Instrumentet passar perfekt ihop med den idé om stöd till entreprenörskap som läggs fram i den europeiska stadgan för småföretag.
Det är viktigt att företagen även får hjälp i ett senare skede, och inte bara vid starten, eftersom de ekonomiska resurserna från instrumentet bara gör nytta för dem som använder dem och för ekonomin om de företag som startas överlever på marknaden.
Jag hoppas också att entreprenörskap, i synnerhet när det gäller små och medelstora företag, inte bara ska diskuteras under krisen.
Vi bör anta en övergripande strategi för entreprenörskap, eftersom de här företagen inte bara ger jobb till våra medborgare under krisen.
(IT) Fru talman, mina damer och herrar! Det skulle ha stor betydelse om vi med 2010, Europaåret för bekämpning av fattigdom och socialt utanförskap, kunde markera skapandet av nytt gemensamt finansieringsinstrument avsett för mikrokrediter till dem som inte får tillgång till bankernas system men som har planer på mikroföretag.
Som vi vet har mikrokrediter visat sig vara ett utmärkt redskap för att skapa tillfällen till eget företagande och sprida sociala värden i utvecklingsländerna, särskilt för kvinnor.
Det har blivit en ny strategi för FN och Världsbanken, men det har också använts i försök med positiva resultat i många länder, i många medlemsstater, bland andra Italien, särskilt för invandrare, kvinnor och ungdomar.
Genom att anta det här betänkandet ger parlamentet mitt i en allvarlig ekonomisk och finansiell kris inte bara en strategisk möjlighet till social inkludering utan även en positiv utmaning till bankernas system, eftersom man utvecklar en ny strategi och nya krafter i samarbete med icke-vinstbringande organ och med lokala och nationella institutioner.
Jag välkomnar antagandet av många ändringsförslag, som jag inte ska upprepa, men jag vill säga att vi i dag inte bara ber om resurser till mikrokrediter utan även begär att mikrokredit ...
(Talmannen avbröt talaren.)
(DE) Fru talman, herr kommissionsledamot, mina damer och herrar! Förra månaden lade kommissionen fram EU:s strategi 2020 som är en fortsättning på målen i Lissabonstrategin och där man bland annat uppmanar till ett mer socialt Europa.
Om vi strävar efter att säkra en varaktig sysselsättning för EU:s medborgare måste vi särskilt nu i detta svåra ekonomiska läge se till att människorna själva kan förverkliga sina egna goda idéer och skapa egen försörjning.
EU-instrumentet för mikrokrediter för sysselsättning syftar till att ge tillfälle till en ny start och underlätta vägen till entreprenörskap.
Övergången till egenföretagande sker ofta stegvis.
Det är lättare att klara av små investeringar i början än att ta på sig berg av skulder.
Särskilt kvinnor efterlyser en mer hanterbar risk när de ska starta eget företag, och de ansöker ofta om startkapital för att kunna etablera företaget och för att sedan när företaget går bra kunna expandera.
Kvinnor vill växa med sina företag.
Därför behöver medborgarna erbjudas lån på så små belopp som möjligt.
Med detta menar jag belopp som är väsentligt mindre än 25 000 euro, som är det belopp som i allmänhet tillhandahålls i form av en mikrokredit.
Det är särskilt under den ekonomiska krisen måste det finnas tillräckliga likvida medel för befolkningen som helhet.
Om det skulle hjälpa till att hålla nere de ofta höga räntorna och administrativa avgifterna för mikrokrediter, skulle vi få tillfälle att ge ny stimulans till ekonomin.
Jag välkomnar den idé som läggs fram i kommissionens förslag.
Parlamentets utskott är oeniga om finansieringen.
Det finns verkligen skäl att ifrågasätta befogenheterna i EU:s politik på detta område.
Medlemsstaterna bär det främsta ansvaret.
Men som jag ser det kan medel från EU:s program för sysselsättning och social solidaritet (Progress), särskilt enligt detta förslag, ge människor möjlighet att bli egenföretagare.
Vi talade tidigare om att utnyttja fonden för justering för globaliseringseffekter och förhoppningsvis ska vi diskutera Progressprogrammet de närmaste dagarna. Och de här EU-finansierade mikrokrediterna är ett idealiskt och nödvändigt instrument.
Jag tycker det är onödigt att upprepa att detta ska lösa eller vara ett försök att lösa problemen för de medborgare som har störst behov av hjälp.
Det enda sättet att ta sig ur detta är att lösa sysselsättningsproblemet, som är vårt sorgebarn, så vi borde försöka se till att det händer något så snart som möjligt och att det finns solida garantier när det gäller resurserna till det här instrumentet. Det behövs nämligen mycket mer resurser än dem vi har hört diskuteras i kväll, och vi borde verkligen inte föra över pengar från det ena instrument till det andra, eftersom pengarna behövs i alla tre programmen.
Enligt min mening ska man absolut inte ta 100 miljoner euro från Progressprogrammet, eftersom även det har samma mål, utan det bör finnas en fullt tydlig och separat budgetpost med garantier om mycket större resurser.
(FR) Fru talman, herr kommissionsledamot, mina damer och herrar! Först och främst vill jag tacka föredraganden för hennes arbete och våra kolleger i parlamentet för deras hårda arbete med att skapa det här nya mikrokreditinstrumentet.
Det här EU-instrumentet gör det möjligt att bevilja mikrokrediter till småföretagen och till personer som har förlorat jobbet och vill starta en egen verksamhet.
Det är de mest utsatta, särskilt arbetslösa och ungdomar, som har drabbats hårdast i dessa kristider.
I år har faktiskt mer än 3,5 miljoner förlorade arbetstillfällen registrerats i EU.
Antagandet av det nya instrumentet gör det lättare för dessa personer att få tillgång till det kapital de behöver för att starta eller utveckla ett företag och förverkliga sina drömmar om entreprenörskap.
Vi får inte glömma att mer än en tredjedel av mikroföretagen bildas av arbetslösa.
I min region blir jag ofta kontaktad av medborgare som skulle vilja ha stöd till att starta ett eget företag.
Jag är övertygad om att det här nya initiativet ska bära frukt när det gäller både att behålla och att skapa nya arbetstillfällen.
Förslaget underlättar för investeringar av små belopp och ger mikroföretagen tillfälle att växa.
Fru talman! Jag välkomnar det verkliga mervärdet av mikrokrediterna, som går hand i hand med nya stödåtgärder som utbildning och mentorskap, vilket ger ungdomar och arbetslösa möjlighet att få garantier och stöd till sina investeringsplaner.
Jag hoppas att det här nya instrumentet ska främja sysselsättningen och antas så snart som möjligt samt att parlamentet och rådet ska enas om att göra det till ett bestående instrument, vilket är mycket viktigt för våra medborgare och särskilt nu under krisen.
Mina damer och herrar! Vi får inte glömma att det är i de små och medelstora företagen som jobben skapas.
(IT) Fru talman, mina damer och herrar! Mikrokreditinstrumentet för sysselsättning ingår i ett paket med initiativ som har antagits på EU-nivå, och det erbjuder arbetslösa en ny start och öppnar dörren till egenföretagande för några av de mest utsatta grupperna i EU, bland annat ungdomar.
Detta nya instrument kommer att utvidga det riktade finansiella stödet till nya entreprenörer mot bakgrund av den nuvarande situationen med minskat kreditutbud.
Enskilda företagare och nyblivna mikroföretagare kommer också att stödjas genom mentorsprogram, utbildning, coachning och kapacitetsuppbyggnad, utöver det räntestöd som Europeiska socialfonden kan tillhandahålla.
Mot bakgrund av den nuvarande situationen med bankernas minskade utlåning och svårigheterna att få lån är det uppenbart att om de svagaste grupperna i samhället, arbetslösa och utsatta grupper, vill göra något, starta en egen verksamhet, måste detta stödjas kraftfullt. Det är ju ett av de instrument som kan bidra till att motverka den ekonomiska krisens givna epilog, nämligen en ändlös sysselsättningskris.
Även om vi nu ser tecken på ekonomisk återhämtning, ser det fortfarande mörkt ut när det gäller sysselsättningen.
Men det är nödvändigt att Progress-medlen betalas ut som planerat. Vi får inte verka för att resurser tas från Progressprogrammet.
Resurserna måste tas från andra källor och framför allt samordnas med andra EU-initiativ, så att vi visar oss starka och gör en kraftfull insats för att hjälpa de arbetslösa i Europa.
(FR) Fru talman, herr kommissionsledamot, mina damer och herrar! Jag vill göra er uppmärksamma på mikrokrediternas grundläggande betydelse för jobben i dessa kristider.
Mikrokrediter ger de arbetslösa tillfälle till en ny start tack vare riskspridning och finansieringsinstrument, som gör det möjligt för dem att ägna sig åt entreprenörskap.
Mot bakgrund av den ekonomiska krisen och den avsevärda minskningen av antalet beviljade lån stöder jag kommissionens förslag om att inrätta ett mikrokreditinstrument som riktar sig till de mest utsatta grupperna, i synnerhet kvinnor, ungdomar och arbetslösa.
Jag vill framföra mitt stöd till kollegerna i Europeiska folkpartiets grupp (kristdemokrater) som tillsammans med övriga grupper - socialdemokrater, liberaler och konservativa - har lagt fram kompromissförslag om ändringar för att mikrokreditinstrumentet ska kunna inrättas så snabbt som möjligt med början 2010.
(PL) Fru talman! Progressprogrammet är ett viktigt initiativ som syftar till att hjälpa medlemsstaterna att på ett effektivt sätt förverkliga målen på områdena sysselsättning och socialpolitik.
Förra veckan deltog jag i ett möte med medlemmarna i programkommittén om genomförandet av Progressprogrammet.
Jag drog följande slutsatser: Den annonskampanj som ska ge programmets potentiella förmånstagare information om programmets räckvidd genomförs för det första inte på ett tillräckligt synligt sätt.
För det andra finns merparten av informationen om anbud och uttagningsförfarande bara på tre språk, nämligen engelska, tyska och franska.
Det utgör ett funktionellt hinder för personer som inte behärskar något av dessa språk.
Jag tycker det finns skäl att se över principerna för reklamkampanjen.
Vi bör så snart som möjligt öka kännedomen om Progressprogrammet och sprida information om det i hela unionen.
(RO) För mikrokreditinstrumentet för sysselsättning och social inkludering eftersträvar man och måste man eftersträva enkla förfaranden, så att de berörda kan dra nytta av det på ett effektivt sätt.
Men jag anser att mikrokreditinstrumentet borde vara mer inriktat på personer som förlorat sina jobb, är missgynnade i förhållande till den traditionella kreditmarknaden och vill starta eller fortsätta att utveckla sina mikroföretag, bland annat som egen verksamhet.
Jag anser att man måste ägna särskild uppmärksamhet åt ungdomar som enligt den senaste EU-statistiken tyvärr står inför ännu längre perioder av arbetslöshet eller får tillfälliga anställningar.
Dessutom ska det inom en snar framtid bli möjligt att med hjälp av en årlig rapport om användningen av budgetmedel göra en grundlig analys och vid behov utöka budgeten.
Om vi överför belopp från det ena programmet till det andra riskerar vi att undergräva båda två.
(DE) Fru talman! I dag har vi diskuterat Europeiska fonden för justering för globaliseringseffekter och nu talar vi om mikrokrediter.
Båda instrumenten är absolut nödvändiga för att motverka den finansiella och ekonomiska krisens effekter i EU och stimulera arbetsmarknaden i Europa.
Vi behöver båda instrumenten, eftersom inte alla är ämnade att bli entreprenörer.
Vi bör inte heller ha som mål med sysselsättningspolitiken att enbart av företagsekonomiska skäl göra egenföretagare av tidigare anställda och förvärvsarbetande utan egen verksamhet.
En del av dem borde i så fall snarare benämnas ”skenbara egenföretagare”.
Medlemsstaterna måste även vidta förebyggande åtgärder när det gäller detta.
Men för alla dem som vill anta utmaningen att bli egenföretagare måste resurser göras tillgängliga så att de kan starta eller utöka sin verksamhet.
Men dessutom måste man se till att den vanliga socialförsäkringen fortsätter att gälla, och detta är Europaparlamentets och medlemsstaternas skyldighet.
Vi behöver nya pengar till nya idéer.
(LT) Jag tror att parlamentets ledamöter nu är helt eniga om att stödinstrumentet för mikrokrediter verkligen behövs.
Levnads- och arbetsförhållandena har förändrats väsentligt och arbetslöshetens gissel som drabbat nästan alla medlemsstater gör att vi måste lägga fram vissa förslag om att ändra vissa stödinstrument.
Hittills har huvuddelen av det ekonomiska stödet varit öronmärkt för storföretag och organisationer, och det har många gånger framhållits att vanliga EU-medborgare hittills knappast kunnat hoppas på något ekonomiskt stöd.
Jag anser att kommissionens framtida lösning att komma överens med parlamentet är absolut nödvändig.
100 miljoner är bara början.
Det är ett första försök, men jag är övertygad om att det kan bli framgångsrikt.
Av diskussionen framgår tydligt att parlamentet stöder mikrokreditinstrumentet och jag tror inte det råder någon större oenighet när det gäller kärnfrågan. Jag tror också att man ligger tämligen nära rådets ståndpunkt när det gäller kärnfrågan.
Det är frågan om finansiering som fortfarande är öppen.
Naturligtvis ingår finansieringsfrågan också i medbeslutandeförfarandet, vilket innebär att det är ytterst nödvändigt och önskvärt att försöka nå en kompromiss, och det gläder mig att debatten tyder på en stor vilja att utan dröjsmål återuppta förhandlingarna med rådet.
Debatten tyder också på att möjligheten att nå en kompromiss på vissa områden.
I debatten nämns och kritiseras ofta kommissionen när det gäller frågan användningen av Progressprogrammet inom ramen för det nya instrumentet.
Jag måste säga att det inte har varit någon enkel fråga för kommissionen, eftersom man varit tvungen att röra sig inom ramen för den befintliga budgeten eller inom ramen för det interinstitutionella avtalet.
Det går bara att använda de pengar som finns tillgängliga.
När vi gjorde bedömningen att använda Progressprogrammets resurser var vi mycket noggranna med att överväga följderna och kom till slutsatsen att det visserligen inte är någon optimal lösning men att det antagligen är en av de möjliga lösningarna.
Det nämndes upprepade gånger i debatten att detta handlade om nonchalans eller att flytta pengar från den ena skålen till den andra.
Det stämmer inte eftersom alla analyser visar tydligt att de resurser som används inom ramen för mikrokrediter beräknas ge en femfaldig effekt.
I det andra programmet skulle resurserna få index 1, men i mikrokreditprogrammet kan de teoretiskt sett nå upp till index 5.
Ur det perspektivet handlar det inte bara om att flytta pengar från den ena skålen till den andra utan om ett nytt sätt att använda resurserna.
Jag upprepar att det inte var något lätt beslut att fatta, och jag tror inte ens att det var det enda beslutet, och i debatten om en kompromiss kan vi säkert hitta en rimlig utgångspunkt, eller åtminstone hoppas jag det.
Idén om mikrokrediter bygger på att tydligt påstående om att det nuvarande finanssystemet inte ger tillräckliga resurser till små och mycket små företag i synnerhet. I systemet används med andra ord inte humankapitalet hos människor i de så kallade utsatta grupperna.
Jag ser det som bortkastade tillfällen i stor omfattning och det gläder mig därför att kommissionen har föreslagit det här instrumentet och att parlamentet sätter så stort värde på det.
Som jag redan har sagt är idén att använda humankapitalet hos de personer som vanligen inte har möjlighet att använda sitt kapital till entreprenörskap.
Men det är också mycket viktigt att utnyttja tiden.
Enligt min mening skulle en orimligt lång debatt motverka syftet med detta instrument som behövs särskilt i dessa kristider.
Jag tror också att det kommer att behövas när krisen är över och att det kommer att bli en bestående del av EU:s arbetsmarknad och ekonomiska politik.
Tack för de uppskattande anmärkningarna och kommentarerna.
Låt mig uttrycka mitt stöd till dem som har uttryckt sin besvikelse över kommissionens ovilja att kompromissa.
Jag måste också påpeka för kommissionsledamoten att en omfördelning av resurser som uteslutande hör till Progressprogrammet ger budskapet att när det gäller medel till social inkludering kan vi bara förvänta oss att stödja de mest utsatta om vi tar medlen ur källor med samma syfte.
Vi lyckas inte hitta någon annan sorts medel.
Jag tycker det är oacceptabelt.
Medbeslutandeförfarandet innebär också att alla, var och en av parterna, måste vidta åtgärder.
Parlamentet har utarbetat ett antal förslag i frågan, men det har inte kommit några sådana förslag från rådet eller kommissionen, vilket skulle ha hjälpt oss att komma överens.
Jag måste säga till Elisabeth Schroedter att vi genom att försvara Progressprogrammet här visar vår övertygelse om att detta program måste genomföras så snart som möjligt, och det är en utbredd övertygelse om att vi fortfarande vill nå en kompromiss om detta.
Det stöd som ges kommer bara att få effekt om instrumentet kan inrättas i början av 2010.
Om parlamentet faktiskt röstar i frågan den här veckan, har parlamentet från sin sida gjort vad det kan för att se till att programmet inrättas i början av 2010.
Eftersom parlamentet antagligen röstar för att ta 25 miljoner euro från sina egna resurser till nästa år, och om parlamentet röstar för hela beloppet, kommer det att vara tillräckligt för att kommissionen ska underteckna de avtal som kan underlätta inrättandet av programmet.
Jag tycker att detta speglar parlamentets konstruktiva ansats.
I alla fall anser jag att programmet är utomordentligt viktigt med tanke på social inkludering.
Jag vill också be de kolleger i parlamentet som stöder detta att gå med på att inte ta hela beloppet ur Progressprogrammet och att försöka skaffa resurser från de egna regeringarna, under förutsättning att dessa länders regeringar företräds av ledamöterna i kommissionen.
Debatten är härmed avslutad.
Omröstningen kommer att äga rum i morgon.
Skriftliga förklaringar (artikel 149)
Den ekonomiska krisen har blivit en överhängande påtaglig social kris som vi ännu inte har någon lösning på.
En av de faktorer som skulle kunna bidra till återhämtningen är långivningen, men den har tyvärr nått sin lägsta nivå sedan 1991 i euroområdet och har kollapsat som aldrig tidigare i de nya medlemsstaterna, såsom Rumänien.
Det är en av de faktorer som skapar ovisshet om utsikterna att övervinna recessionen.
Mot denna bakgrund välkomnar jag kommissionens förslag om att inrätta mikrokreditinstrumentet.
Men för att se till att åtgärderna för social inkludering blir effektiva måste man ge instrumentet en separat budgetpost.
Omfördelningen av medel från Progressprogrammet skulle påverka programmets specifika riktlinjer för unionens åtgärder och ge en varningssignal när det gäller den sociala öppenheten i EU:s verkställande organ, som hittills tyvärr har varit utomordentligt motvilliga när det gäller att visa tillräckligt mycket samhällsengagemang.
Krisen påverkar alla utsatta grupper, men vi får inte bortse från den omfattande ungdomsarbetslösheten.
En av fem ungdomar i Europa saknar jobb och det kan få åtskilliga återverkningar på ekonomisk och social nivå, och likaså när det gäller demografi och kriminalitet.
Därför anser jag att det är lämpligt att i högre grad inrikta sig på att förbättra möjligheterna för ungdomar att komma in på arbetsmarknaden.
Sedan i höstas har över 5 miljoner EU-medborgare förlorat sina arbeten, vilket har resulterat i sammanlagt 22,5 miljoner arbetslösa i Europa.
Mot denna bakgrund kan vi inte ignorera den allvarligt höga arbetslösheten bland ungdomar.
Det är djupt oroande att var femte ung människa i Europa står utan arbete, när det får återverkningar både på ekonomisk och social nivå, och sett ur en demografisk och brottsrelaterad synvinkel.
I vissa länder är procentandelen unga som saknar arbete dessutom högre jämfört med andelen arbetslösa i befolkningen i stort.
Till exempel är var tredje ung människa i Lettland arbetslös, medan ungefär 43 procent av Spaniens medborgare under 25 år är drabbade av problemet.
Jag anser att fokus måste riktas mer på ungdomarna.
Initiativet från kommissionen till EU-instrumentet för mikrokrediter, som ska finansieras med en särskild budgetpost, kommer i detta hänseende att hjälpa till att uppmuntra och motivera unga människor till att komma ut på arbetsmarknaden, och därigenom minska arbetslöshetstalen som har stigit i den här gruppen.
De ansträngningar som nu görs både på EU-nivå och nationell nivå måste ökas för att förbättra erbjudandet om mikrokrediter.
EU-instrumentet för mikrokrediter måste ge användbart stöd till de arbetslösa och utsatta människor som vill starta eller driva mikroföretag.
Jag anser att EU-instrumentet för mikrokrediter bör finansieras med särskild kreditgivning, eftersom målgruppen för detta stöd inte är samma som för Progressprogrammet.
Progressprogrammets anslag ska inte under några omständigheter minskas i dessa kristider, eftersom de riktar sig till de mest utsatta grupperna.
Jag anser även att EU-instrumentet för mikrokrediter bör få en tillräckligt stor budget för att på ett effektivt sätt kunna uppnå sina mål för arbete och social integration.
Medlemsstaterna och EU i stort måste fortsätta att effektivt genomföra Progressprogrammet i en tid av global ekonomisk kris.
Skriftliga förklaringar för införande i registret (artikel 123 i arbetsordningen): se protokollet
Inkomna dokument: se protokollet
15.
Nominering av en ledamot av revisionsrätten - Eoin O'Shea (IE) (
3.
Effekterna av den globala finansiella och ekonomiska krisen på utvecklingsländerna och utvecklingssamarbetet (
Före omröstningen:
Herr talman! Jag vill tacka alla som har deltagit i utarbetandet av detta betänkande.
Jag vill bara påpeka att det finns ett muntligt ändringsförslag till punkt 31.
Som vi kommit överens om ska jag nu läsa upp den andra delen av den engelska versionen.
(EN) ”Parlamentet anser därför att det är lämpligt att undersöka om det är möjligt att ingå en överenskommelse med långivarländerna om ett tillfälligt moratorium eller skuldavskrivning för de fattigaste länderna för att göra det möjligt för dem att genomföra konjunkturutjämnande ekonomiska strategier för att begränsa krisens allvarliga följder. Parlamentet föreslår att ansträngningar görs för att underlätta åtgärder för transparent tvistlösning i skuldfrågor.”
Herr Guerrero, om vi inte har fått fel information gäller det här muntliga ändringsförslaget punkt 34 och inte punkt 31.
(Enrique Guerrero Salom bekräftade att ändringsförslaget gällde den andra delen av punkt 34.)
Då var det klart.
(Omröstningen ägde rum.)
(Det muntliga ändringsförslaget beaktades.)
- Före omröstningen om punkt 22:
(FR) Herr talman! Vi har anmält ett muntligt ändringsförslag gällande punkt 22.
Jag vill påpeka att punkt 22 gäller global styrning och i synnerhet sammansättningen av G20-gruppen, vilken märkligt nog inte har någon företrädare från de minst utvecklade länderna.
Det muntliga ändringsförslaget syftar till att avhjälpa denna brist och den text jag föreslår parlamentet fyller detta behov.
(FR) Herr talman! För en stund sedan bad ni oss välkomna Tunisiens delegation.
Kan ni be den tunisiska delegationen att ingripa för ett frisläppande av Taoufik Ben Brik, en begäran från hela parlamentet?
(DE) Herr talman! Jag vill ta upp en ordningsfråga.
Jag är mycket nöjd med resultatet av omröstningen.
Men detta var till största delen ett initiativbetänkande och vi har enats om ett annat förfarande för sådana fall.
Nu har vi fått ha en enskild omröstning om ett initiativbetänkande.
Vi måste lösa detta för annars kommer vi att ha enskilda omröstningar om alla initiativbetänkanden i framtiden.
Skulle ni kunna be utskottet för konstitutionella frågor att klargöra saken?
I annat fall kan den tolkning som görs av parlamentets enheter rasera hela syftet med reformen.
Herr Swoboda, det kan ordnas.
Det är möjligt att begära delad omröstning, i enlighet med det förfarande som grupperna själva har begärt.
I alla händelser kan allt revideras. Det kan revideras i framtiden, men för närvarande är det som det är.
1.
Administrativt samarbete och kampen mot skatteundandragande i fråga om mervärdesskatt (omarbetning) (
37.
Befogenhet att delegera lagstiftning (
8.
Betänkande om kommissionens vitbok: Anpassning till klimatförändring: en europeisk handlingsram (
Herr talman, mina damer och herrar! Klimatförändringen är ett verkligt hot som vi måste vara redo att bemöta, trots att den kommer att påverka våra länder i varierande grad.
Ekosystemens nedbrytning kommer att utgöra ett hårt slag mot hälsan i våra ekonomier och hos de europeiska medborgarna.
Vi har redan tidigare efterlyst klimatdiplomati och rättvisa: vi är nu tvungna att skapa detta, genom att tala med enad röst.
Jag är övertygad om att EU bör behålla ledningen i kampen mot klimatförändringen och att varje försening med att genomföra dessa åtgärder kommer att öka de miljömässiga, sociala och ekonomiska kostnaderna på ett oproportionerligt sätt.
Vi måste först av allt erkänna de lokala och regionala myndigheternas centrala roll och behovet av att samarbeta med dem för att samordna de miljömässiga och ekonomiska innovationer som främjas genom tekniska framsteg.
Genom att anta vitboken uppmanar vi kommissionen och medlemsstaterna att främja offentlig-privata partnerskap för att hjälpa till att finansiera alla de initiativ som är knutna till anpassningspolitiken.
Varje kvadratmeter av vårt territorium måste tas om hand för att skydda jorden och behålla vattnet för att förhindra erosion och fylla på akviferer, däribland genom direkt återföring av ytvatten.
För att en anpassning ska vara möjligt krävs en systematisk strategi som omfattar förnybara energikällor.
Jag vill varmt tacka alla mina kolleger som har bidragit till framgången med detta betänkande.
(Applåder)
Sammansättningen på delegationen till parlamentarikerkommittén Cariforum-EU (tidsfrist för ingivande av ändringsförslag): se protokollet
Utskottens och delegationernas sammansättning: se protokollet
Avslutande av sammanträdet
Genomförda reformer och utvecklingen i Moldavien (debatt)
Den första punkten är kommissionens uttalande om genomförda reformer och utvecklingen i Moldavien.
ledamot av kommissionen. - (EN) Herr talman! När det gäller förbindelserna mellan EU och Moldavien råder det enighet om att vi har gjort stora framsteg på rekordtid, men inrikes står landet fortfarande inför många utmaningar.
Folkomröstningen den 5 september var avsedd att lösa det politiska dödläget genom att ändra reglerna för presidentvalet. Detta misslyckades.
Det är beklagligt. En annan viktig fråga var emellertid också huruvida folkomröstningen skulle uppfylla demokratiska standarder.
Att dessa standarder faktiskt efterlevdes har bekräftats av internationella observatörer. Det är ett uppmuntrande tecken.
Valet den 28 november är lika viktigt för att befästa demokratin i landet. Vi kommer att fortsätta att sända skarpa budskap i detta avseende till alla berörda parter.
Därefter är samtliga politiska aktörer tvungna att samarbeta, för att både välja en president och utse en regering som kan klara av att leda landet genom ett kritiskt reformarbete.
Samtidigt kommer vi att upprätthålla vårt orubbliga stöd till de strukturella reformer som genomförs av den moldaviska regeringen.
Jag vill belysa några viktiga aspekter.
EU är inte bara den ojämförligt största bidragsgivaren till Moldavien; i mars lyckades man också mobilisera mer än fyrtio bidragsgivare för att stödja Moldaviens reformer.
De utlovade ett imponerande belopp på 1,9 miljarder euro för åren 2010-2013, vilket även omfattade vårt eget åtagande på 550 miljoner euro.
Under de senaste månaderna har vi i god tid svarat på ett antal av regeringens särskilda behov genom att bereda policyförslag på en övergripande nivå till ministrar, stödja demokratiseringsinsatser på områden med anknytning till rättsstatsprincipen, hjälpa till att organisera samråd med väljarna, åtgärda akuta behov efter förra sommarens översvämningar och förbättra möjligheterna för den moldaviska vinexporten.
Tillsammans med den moldaviska regeringen har vi aktivt samarbetat med befolkningen i den transnistriska regionen genom småskaliga projekt, främst på det sociala området.
Under nästa år kommer vi att inleda genomförandet av det heltäckande programmet för institutionell uppbyggnad inom ramen för det östliga partnerskapet.
Programmet kommer att hjälpa Moldavien med förberedelserna för, och genomförandet av, de associeringsavtal som vi för närvarande förhandlar om.
Den senaste förhandlingsrundan i Chisinau den 13-14 oktober visade återigen att förhandlingarna går framåt i mycket snabb takt.
Vårt stöd har också utformats som direkta överföringar till den moldaviska budgeten.
Sedan sista kvartalet 2009 har 37 miljoner euro betalats ut som sektoriellt budgetstöd, och ytterligare 15 miljoner euro kommer att utbetalas inom kort.
Av dessa belopp har omkring 8,5 miljoner euro direkt avsatts för att hjälpa den fattigaste delen av befolkningen.
Nu när talman Jerzy Buzek har undertecknat det relevanta lagstiftningsbeslutet förväntar vi oss att inom kort kunna betala ut 40 miljoner av den första delen av ett makrofinansiellt stöd.
I samma anda kommer vi att fortsätta med vårt fulltecknade program av politiska kontakter och tekniskt utbyte.
Om några dagar kommer jag att träffa premiärminister Vlad Filat i Luxemburg.
I november kommer underkommittén EU-Moldavien för handel att undersöka hur Moldavien har svarat på kommissionens främsta rekommendationer i syfte att förbereda förhandlingar om ett djupgående och omfattande frihandelsområde.
Vi har också tillsammans med Moldavien inlett en särskild dialog om mänskliga rättigheter och en dialog om energi, och vi förhandlar om ett avtal om luftfartstjänster.
Vi har aktivt följt upp den viseringsdialog som inleddes i juni.
Nästa måndag förväntas rådet (utrikes frågor) tillkännage slutsatser om denna fråga utifrån resultatet av de informationsuppdrag som oberoende experter utförde i september.
Syftet med denna debatt är att vi ska diskutera de reformer som Moldavien genomförde under förra året och de framsteg som gjorts på vägen mot en europeisk integration.
Landet har funnits med på EU:s dagordning under ett års tid eftersom det har uppfyllt sina åtaganden.
Jag vill ta upp några av dessa åtaganden.
En plan har utarbetats över prioriterade åtgärder att vidta på väsentliga reformområden, utöver ytterligare en plan för en reform av rättsväsendet.
Genomförandet av båda planerna har påbörjats.
En dialog om mänskliga rättigheter har inletts.
Dessutom undertecknade det moldaviska parlamentet Internationella brottmålsdomstolens stadga i september.
Det förs intensiva förhandlingar om associeringsavtalet med utmärkta resultat så här långt.
Bara ett år har passerat, men de som deltagit under det inledande förfarandet garanterar att det kommer att fortsätta.
Moldavien är den stat som har gjort störst framsteg inom EU:s östliga partnerskap.
Därför uppmanar jag rådet att bedöma denna stat enskilt på egna meriter.
Framsteg tyder på politisk vilja, hårt arbete och engagemang, vilket bör belönas.
Vi belönade länderna på västra Balkan för de åtgärder som de vidtagit.
Låt oss gå vidare och göra likadant för Moldavien också.
I dialogen om viseringar har Moldavien gjort stora framsteg på samtliga fyra områden.
Därför ber jag rådet att vid nästa sammanträde den 25 oktober uppmana kommissionen att utarbeta en handlingsplan så att medborgare från Moldavien kan resa utan visum.
Direkta kontakter mellan människor är värt mer än deklarationer.
När det gäller Transnistrien är en lösning av avgörande betydelse för den politiska och ekonomiska stabiliteten i Moldavien och denna region.
EU bör spela en mer kraftfull roll på politisk nivå och vi bör delta genom gemensamma projekt som bidrar till förändringar som människor kan uppfatta.
Slutligen har den europeiska integrationsprocessen bidragit till att upprätta demokrati och frihet i en omfattning som aldrig tidigare skådats i Europas historia.
Se bara på hur situationen i Central- och Östeuropa har förändrats under de senaste tjugo åren.
Fred råder nu även i länderna på västra Balkan och reformer är på gång.
Låt oss göra vad som krävs för att också uppnå en sådan situation i Moldavien.
för S&D-gruppen. - (EN) Herr talman! Moldavien har ett val, dvs. valet mellan en ”transnistrisering” eller en ”europeisering”.
Med andra ord ett val mellan ett oligarkiskt förflutet av sovjetisk natur och en framtid av säkerhet, välgång och social rättvisa.
Moldaviens utveckling har hittills påverkats negativt av landets inhemska politiska instabilitet.
Landets grundläggande problem är inte knutet till de externa utmaningar som landet står inför, utan till en intern splittring bland de politiska aktörerna.
Denna inhemska politiska instabilitet har inneburit att den styrande koalitionen inte haft tillräckligt med tid för att genomföra sina proeuropeiska lösningar.
Moldavien står nu inför en vändpunkt.
Resultatet av detta tidiga val bör syfta till att leda landet mot en framtid av europeisk modernisering.
Vi uppmanar därför alla politiska aktörer i Moldavien som föreslår en framtid av europeisk modernisering för landet att undvika onödig protagonism eller konfrontationer, och att inrikta sig på att utveckla en allmän vision i syfte att hjälpa landet att uppnå sina europeiska mål.
för ALDE-gruppen. - (EN) Herr talman! För arton månader sedan upprördes parlamentet av de brutala händelserna i Chisinau.
Några veckor senare hade vi det stora nöjet att till vår åhörarläktare välkomna ledarna för landets demokratiska politiska partier, som slagit in på en ny bana.
Vi delade det moldaviska folkets entusiasm för en ny framtid.
Vi har sedan dess glatt oss över de framsteg som landet gjort.
Ytterligare framsteg återstår att göra - inte minst när det gäller att ställa förövarna för dessa brutala händelser inför rätta - men om Moldavien ger den nuvarande koalitionen förnyat mandat vid valet i nästa månad finns det, trots svårigheterna med den ekonomiska lågkonjunkturen, goda chanser att landet kan fortsätta sin omvandling.
Den brittiske författaren Francis Bacon konstaterade att hoppet är en bra frukost men en dålig middag.
Moldaviens styrande partier bör vara förvissade om att reformernas genomförande följer de rättsakter som möjliggör dessa reformer.
Tiden är inte på vår sida.
Mycket behöver åstadkommas på kort tid.
Min grupp berömmer kommissionsledamot Štefan Füle och hans tjänsteenheter för deras arbete med att bistå Moldavien.
Vi välkomnar bildandet av Moldaviens vänner och det storartade möte som hölls med europeiska länder i syfte att hjälpa Moldavien framåt.
Det görs stora insatser från EU:s sida för att hjälpa detta förtvivlat fattiga land att närma sig EU:s standarder.
Jag hoppas att rådet, när det i nästa vecka behandlar viseringsreglerna, hjälper oss att hitta en väg framåt i visumfrågan.
Som en av unionens fäder sade bestäms ett lands EU-strävanden inte av EU utan av den europeiska andan hos landets befolkning.
Vi uppmanar det moldaviska folket att visa denna europeiska anda vid valet i nästa månad.
Herr talman! Vi välkomnar de framsteg som Moldavien gjort och hoppas att den kommande valprocessen kan stärka de demokratiska institutionerna ytterligare och säkerställa att rättsstatsprincipen och de mänskliga rättigheterna respekteras i Moldavien.
Vi vet att det finns ett brett stöd i det moldaviska samhället för ett framtida moldaviskt medlemskap i EU - inte Nato.
Trots deras olika politiska plattformar har samtliga partier i det moldaviska parlamentet förklarat sig vara för ett europeiskt samarbete och en europeisk integration.
Men mot bakgrund av mitt eget hemland Lettlands erfarenheter av EU-medlemskapet har jag under mina samtal med moldaviska politiker försökt förklara att EU-medlemskapet inte kan vara ett mål i sig.
Det är mycket viktigt att påskynda försöken att genomföra djupgående och enhetliga ekonomiska och rättsliga reformer, i synnerhet genom att bekämpa korruptionen.
Det moldaviska samhället är multietniskt och flerspråkigt. Det finns dessutom väsentliga skillnader i hur man bedömer historiska händelser.
Därför är det mycket riskfyllt att skapa ytterligare skiljelinjer inom det moldaviska samhället.
Genom ett nyligen utfärdat dekret har den 28 juni fastställts som årsdag för den sovjetiska ockupationen, vilket utlöste en negativ reaktion hos en stor del av den moldaviska befolkningen. Snarare än att stärka samhället fick detta en motsatt effekt.
Det moldaviska samhället rymmer också flera olika nationaliteter bland befolkningen.
Det faktum att en stor del av de bofasta har dubbelt medborgarskap innebär också stora skillnader i fråga om rättigheter, och vi bör därför försöka avskaffa dessa skillnader och upprätta ett viseringsfritt system för samtliga moldaver.
Herr talman! Ingen bestrider att Moldavien har en lång väg att gå innan landet når sitt slutliga mål om anslutning till EU, som är ett mål som stöds av min grupp, ECR.
Moldavien är fortfarande ett av Europas fattigaste länder, trots att det är med i WTO, och är som sådant sårbart för organiserad brottslighet, människohandel och korruption.
Moldavien fortsätter att vara lamslaget av den pågående fastlåsta konflikten med den rysktalande och politiskt ryskdominerade utbrytarregionen Transnistrien.
Sedan kommunisterna drevs bort från makten för 15 månader sedan har Moldavien emellertid börjat göra väsentliga framsteg.
Partierna i Alliansen för europeisk integration, den koalition som i dagsläget styr landet, har visat en imponerande förmåga att samarbeta för att påskynda Moldaviens integrering i Europeiska unionen.
Unionen bör för egen del upprätthålla sina påtryckningar gentemot den moldaviska regeringen för ytterligare framsteg med de ekonomiska reformerna samt för en förbättrad rättsstatsprincip och ett gott styrelseskick.
Vi bör emellertid också belöna och samarbeta mer med regeringen i Chisinau.
Viseringsfrågan har nämnts, men jag vill också ta upp frågan om Euronest, som innebär möjligheter för politiker från både EU och Moldavien att diskutera gemensamma intressen.
Tyvärr har Euronest - som jag tog upp i ett betänkande under parlamentets förra mandatperiod - förblivit lamslaget till följd av tvisten om den vitryska representationen. Tvisten är en följd av att vårt parlament inte har erkänt det vitryska parlamentet, som inte har valts på demokratisk väg.
Jag hoppas att alla tydligt europeiska länder inom det östliga partnerskapet, nämligen Moldavien, Ukraina och ett framtida demokratiskt Vitryssland, en dag kommer att bli kandidatländer för anslutning till EU.
Herr talman! Denna debatt visar på EU:s engagemang för det splittrade Moldavien, vilket gläder mig innerligt.
I mitt hemland Nederländerna har medborgare under flera års tid åstadkommit vissa inspirerande sociala initiativ som ger unga människor från Moldavien goda framtidsutsikter.
I detta sammanhang vill jag också stolt nämna Orhei-stiftelsen i Bunschoten-Spakenburg, en by där man med stor entusiasm har hanterat liknande problem.
Jag kan se människorna från denna stiftelse i ögonen, eftersom vi också talar om denna fråga här, och visar vårt engagemang.
För övrigt strävar Moldavien efter ett djupgående, övergripande handelsavtal med EU.
Kommissionsledamot Štefan Füle nämnde också detta.
Herr kommissionsledamot, hur ser situationen ut på detta område och har det skett några påtagliga framsteg ännu?
Det är avgörande att försäljningsmöjligheterna för de moldaviska produkterna vidgas, i synnerhet när det gäller jordbruksprodukter och viner från Chisinau. Moldaviens främsta traditionella försäljningsmarknad Ryssland stänger nämligen regelbundet sina gränser eller begränsar införseln av politiska skäl.
Herr kommissionsledamot, du har redan nämnt detta, men finns det något sätt för EU att avhjälpa detta behov från Moldaviens sida?
Slutligen en fråga om den tyska förbundskanslern Angela Merkels ”Meseberg-initiativ”.
Finns det i dagsläget ett genuint engagemang från Rysslands sida för att nå en lösning i frågan om Transnistrien, i utbyte mot en förstärkt politisk dialog mellan EU och Ryssland?
Jag har hört det antydas att Kreml inte vidtar några åtgärder för närvarande.
Herr kommissionsledamot, jag vill särskilt önska dig framgång och uthållighet i försöken att föra Moldavien närmare EU.
(EN) Herr talman! Det finns gott om bevis på att Moldaviens åtagande om att efterleva europeiska värderingar och standarder är genuint och effektivt.
Bland våra grannländer i öst är Moldavien det land som lyckats bäst med att genomföra en proeuropeisk politik.
Moldavien har i själva verket lyckats uppfylla kriterierna för euron i överensstämmelse med länderna på västra Balkan.
Det positiva prejudikat som Moldavien skapat bör erkännas och uppmuntras.
De demokratiska institutionernas försämrade situation i grannlandet Ukraina ökar Moldaviens betydelse för EU:s politik mot Öst.
I detta sammanhang är det avgörande att det allmänna valet den 28 november bekräftar Moldaviens fortsatta strävan mot en europeisk integration.
Det är definitivt hög tid för EU att sända en positiv signal till Moldavien och moldaverna.
Tusentals moldaviska familjer är splittrade på grund av att de förnekas visum.
Viseringsdialogen mellan EU och Moldavien utgör en stor möjlighet för oss.
Denna dialog bör gå in i en operativ fas.
Låt oss hoppas att rådet (utrikes frågor) den 25 oktober kommer att uppmana kommissionen att utarbeta en handlingsplan för viseringsliberalisering.
Ett proeuropeiskt integrerat Moldavien skulle ha fördelaktiga effekter på EU:s östliga gräns, där svaga regeringar och olösta konflikter utgör ständiga hot mot den europeiska stabiliteten.
(BG) De utmaningar som Moldavien för närvarande står inför, och som också är en del av vårt allmänna mål, omfattar en förstärkning av den multietniska staten och dess identitet, en politisk lösning på problemet med Transnistrien och ett medlemskap i EU för Moldavien, som en autonom, självständig stat.
Processen med en viseringsliberalisering är särskilt viktig.
Vi har haft liknande fall i länderna från före detta Jugoslavien där viseringsliberaliseringen gett goda resultat.
Utvecklingen mot att tillämpa ett påskyndat förfarande för att simultant utfärda bulgariska och rumänska pass till moldaviska medborgare är ingen lösning på problemet utan medför istället vissa risker.
Samtidigt måste myndigheterna i Chisinau se till att de 90 miljoner euro i makrofinansiellt stöd som EU har beviljat blir kännbart för alla moldaviska medborgare, oavsett etniskt ursprung.
Detta är också särskilt viktigt för den bulgariska minoriteten i Moldavien, som lever i en av landets fattigaste ekonomiska regioner.
(RO) Som ledamot av den parlamentariska samarbetskommittén EU-Moldavien har det varit ett nöje för mig att följa Moldaviens positiva framsteg, och jag kan bekräfta att Moldaviens engagemang för det europeiska arbetet har varit tydligt under det senaste året.
Jag vill på den här punkten påminna om de reformer som gjorts på det ekonomiska området, samt inom rättsväsendet och den offentliga förvaltningen.
Samtidigt bör vi vara realistiska och erkänna att övergångsprocessen i Moldavien inte är okomplicerad, och att flera reformer fortfarande återstår att genomföra.
Det gläder mig att det görs framsteg i de diskussioner som syftar till en viseringsliberalisering.
Jag anser emellertid att kommissionen behöver utarbeta en tydlig färdplan för att uppnå detta mål, och för att kanske till och med avskaffa viseringskravet helt och hållet i framtiden.
Moldavien kommer att stå inför en avgörande prövning i samband med valet till parlamentet den 28 november, och jag hoppas att den europeiska väg som landet har valt att följa kommer att godkännas av befolkningen, och fortsätta.
Makrofinansiellt och politiskt stöd från EU:s institutioner och från vissa medlemsstater har varit av största betydelse.
Mot bakgrund av de positiva resultaten av vår politik uppmanar jag EU:s institutioner, dvs. parlamentet, rådet och kommissionen, att fortsätta sina åtgärder till stöd för Moldavien.
(PL) För tio dagar sedan hade jag möjlighet att besöka Moldavien som en del av en särskild delegation från utskottet för utrikesfrågor tillsammans med bland andra mina ledamotskolleger Monica Luisa Macovei och Graham Watson.
Vi var i Moldavien vid en ytterst viktig tidpunkt för landet - några veckor efter den misslyckade konstitutionella reformen den 5 september och några veckor före det mycket viktiga parlamentsvalet, som ni vet kommer att hållas den 28 november.
Vad vi framför allt upplevde var ett mycket starkt stöd från nationen och det moldaviska samhället för den europeiska integrationsprocessen.
Närmare tre fjärdedelar av moldaverna stöder denna process.
Vi såg också de väldiga framsteg som har gjorts av premiärminister Vlad Filats regering på vägen mot en europeisk integration och med det stora antalet reformer, däribland väsentliga framsteg med att bekämpa korruptionen som tidigare tärt hårt på landet.
Givetvis förekommer det problem, som både är en följd av finanskrisen och ett resultat av den ännu olösta situationen i Transnistrien.
För att reformprocessen ska fortsätta efter den 28 november behövs emellertid en tydlig signal från EU. Jag hoppas därför att man under det följande rådsmötet kommer att kunna driva igenom processen för en viseringsliberalisering.
(RO) Även jag vill tacka alla de som har möjliggjort denna debatt.
Det är vår plikt att betrakta Moldavien med stor ansvarskänsla, särskilt nu när valet närmar sig.
Den styrande Alliansen för europeisk integration har genom sina särskilda insatser visat att den är redo att inleda en omfattande process av politiska, ekonomiska och institutionella reformer, och därigenom går den i spetsen på detta område inom det östliga partnerskapet.
Detta sker efter åtta år av kommuniststyre, då grundläggande rättigheter såsom yttrandefrihet och rätten till rättvis behandling varit föremål för allvarliga kränkningar.
Moldaviens reformprocess måste fortsätta, framför allt inom rättsväsendet och på området för inrikes frågor.
Korruptionen måste bekämpas effektivt, och rättslig frihet garanteras.
Samtidigt måste man se till att frihetsberövande åtgärder utförs säkert och humant, så att grundläggande mänskliga rättigheter efterlevs.
Moldavien har nu haft en politisk kris under mer än 18 månader till följd av att presidentvalet och godkännandet av folkomröstningen misslyckades.
Jag anser att det kommande valet den 28 november är ett stort vågspel som äventyrar Moldaviens närmande till EU.
Demokratin utsätts återigen för en svår prövning.
Jag vill på ett ansvarsfullt sätt påstå att ett misslyckande för demokratin i Moldavien vid det kommande valet i viss utsträckning även kommer att beteckna ett misslyckande för EU:s politik i landet.
Vi behöver en partner i EU:s omedelbara närhet som antagit våra gemensamma värderingar.
Jag vill avsluta med att betona att det språk som talas av de moldaviska invånarna nu är ett officiellt språk i EU.
Detta är ytterligare ett skäl till att landet bör få vårt stöd.
(BG) Det gläder mig att parlamentet ägnar sin tid åt att diskutera situationen i Moldavien, ett land som i allt väsentligt är europeiskt.
I detta hänseende bör vi nämna att den styrande koalitionen för europeisk integration i själva verket bidragit en hel del till processen med att föra Moldavien närmare EU, och för detta bör den berömmas.
Samtidigt förväntar sig landets medborgare fler resultat på områdena för ekonomi och social utveckling.
Det är ingen slump att detta håller på att bli den nuvarande kampanjens viktigaste fråga.
Att upprätta förbindelser med EU är ingen engångsföreteelse.
Det är en långsiktig process, och Moldaviens tillnärmning måste bli oåterkallelig politik.
Misslyckandet med att ändra konstitutionen har lett till detta politiskt instabila tillstånd, som riskerar att upprepas efter det förestående valet.
Därför vädjar jag till de ledande politiska aktörerna, oavsett skillnader och valresultat, att göra vad som krävs för att garantera politisk stabilitet i Moldavien. Detta kommer att ge dem möjlighet att agera i medborgarnas intresse och främja landets europeiska framtid.
(RO) När parlamentsledamöter i Rumänien visar intresse för, och uttalar sig om, situationen i Chisinau beskrivs detta som rumänsk imperialism av moldaviska kommunister, oavsett om det är president Traian Băsescu eller ledamöter av Europaparlamentet som yttrar sig.
Kommunisterna i Chisinau vill med andra ord att regeringen i Bukarest ska tiga.
Jag anser inte att de kan förvänta sig något sådant.
Tvärtemot är det vår plikt att säga vår mening.
Den främsta orsaken till detta är att ett stort antal ursprungligen europeiska, rumänska, bulgariska och andra medborgare lever i Moldavien.
Jag anser att de boende i Moldavien, i likhet med alla övriga europeiska medborgare, ska kunna åtnjuta de rättigheter som deras politiska ställning ger dem.
För det andra bör vi rikta vår uppmärksamhet mot Chisinau, eftersom landets koalitionsregering nu har agerat under mer än ett års tid för en europeisk integration.
Det handlar inte bara om koalitionens benämning.
Om den hade hetat Alliansen för Ryssland hade vi förvisso inte visat så mycket intresse för den.
Den benämns som Alliansen för europeisk integration, men det är inte bara namnet som räknas, utan det är denna regerings mycket modiga åtgärder.
Monica Luisa Macovei och kommissionsledamot Štefan Füle har förklarat vad dessa modiga åtgärder inneburit.
I förra veckan besökte jag Chisinau och Tiraspol och lade märke till att landets europeiska strävanden också står på spel i valkampanjen, som ska inledas inför valet i november.
De moldaviska medborgarna ska i själva verket inte bara välja mellan olika politiska företrädare utan också mellan ett fortsatt eller avbrutet närmande mot EU.
Låt oss inte lura oss själva.
Jag såg att till och med ledaren för EU:s delegation i Chisinau började bedra sig.
Kommunisterna vill inte ha någon integration.
Kommunisterna demonstrerade sin önskan för drygt ett år sedan.
Demonstrationerna i april var ett mycket tydligt bevis på var kommunisterna i Chisinau har sina intressen.
Därför hoppas jag att medborgarna kommer att förstå partiernas budskap och inställning, och att politikerna själva också förstår de önskningar som folket uttrycker vid valurnorna.
(PL) Vi bör fråga oss varför vi ägnar så mycket uppmärksamhet åt ett sådant litet land som ligger i närheten av Svarta havet, men som saknar tillgång till samma hav.
Orsaken till att vi talar om Moldavien är kanske att det är ett litet land där två världar möts.
En av dessa världar, som en gång symboliserade Sovjetunionen, håller med stora svårigheter på att förpassas till det förgångna.
Moldavien är ett delat land.
En del av landet är under ockupation och stöds av externa aktörer.
Jag anser att landet förtjänar vårt stöd.
Det är ett litet land som bebos av ett mycket modigt folk som vill närma sig EU och upprätta demokrati.
Herr kommissionsledamot, situationen i Moldavien påminner om en idé inom fysiken som säger att det inte är styrkan i sig som är viktig utan den punkt mot vilken den riktas.
Dessa miljontals euro som ni talade om är inte särskilt imponerande.
Det är bara ett marginellt belopp, men om det riktas rätt vid rätt tidpunkt kan det åstadkomma de positiva effekter som vi önskar.
Jag lyckönskar alla dem som vill upprätta demokrati i Moldavien.
Jag är inte intresserad av partitillhörighet, men jag skulle vilja att Moldavien stärks och att landet kan bygga en bättre framtid för sitt folk och bli vår partner inom en nära framtid.
(SK) De framsteg som Moldavien hittills har gjort tyder på att landet skulle kunna bli ett exempel på en framgångssaga bland deltagarländerna i EU:s östliga partnerskap.
Den nuvarande proeuropeiska regering som leds av Alliansen för europeisk integration har gett de moldaviska medborgarna ett tydligt och viktigt politiskt perspektiv för framtida framsteg när det gäller att bygga upp landets demokrati.
Det är emellertid också sant att den interna politiska situationen har påverkats negativt av den utdragna tvisten om en konstitutionell reform.
Efter den misslyckade folkomröstningen borde det kommande valet överbrygga dödläget i de politiska förhandlingarna mellan partierna.
Jag anser att EU uttryckligen bör erkänna de viktiga framsteg som den nuvarande regeringen har uppnått när det gällt att stärka förbindelserna med unionen.
På måndag den 25 oktober förväntas rådet (utrikes frågor) utfärda sina slutsatser om Moldavien.
Rådet borde uttrycka sitt stöd för de proeuropeiska åtgärder som den nuvarande regeringen hittills har vidtagit och, vad viktigare är, rådet skulle kunna uppmana kommissionen att utarbeta en handlingsplan avseende viseringsliberaliseringen.
Detta är en viktig fråga för Moldaviens medborgare.
Givetvis kommer det slutliga resultatet främst att bero på valresultatet.
Vad beträffar Europaparlamentet anser jag att vår hållning gentemot Moldavien borde vara mer positiv.
Vi borde på ett tydligare sätt visa vårt stöd för landets proeuropeiska aktörer och även visa dem att vi är angelägna om att Moldavien ska bli en framtida medlem i ett förenat Europa.
Vi bör övertyga dem om att en sådan framtid även ligger i deras bästa intresse.
(EN) Herr talman! Moldavien har kommit en bra bit på vägen sedan Molotov-Ribbentroppakten delade upp Europa i maktsfärer, och Moldavien blev en del av dåvarande Sovjetunionen.
Moldavien är i dag en självständig stat.
Det är sant att landet har många problem.
Samtidigt är det ett demokratiskt land på väg mot en europeisk integration, så i dag vill jag uppmuntra alla politiska klasser i det landet, alla demokratiska politiska aktörer och alla etniska samfund att undvika onödiga konfrontationer. I stället bör man satsa på att utveckla en bred vision för Moldavien i syfte att hjälpa landet att uppnå sina europeiska mål.
Sist men inte minst gäller det frågan om Transnistrien.
Transnistrien borde prioriteras högt på vår dagordning, och jag välkomnar initiativet från Tysklands förbundskansler Angela Merkel och några andra länders politiska ledare för att lösa denna fastlåsta konflikt.
(EN) Herr talman! Moldavien är en sista rest av ”den latinska kulturen” utanför EU.
Historien har haft en stor roll i detta.
Grannskapspolitiken och det östliga partnerskapet har förbättrat Moldaviens utsikter att först närma sig och sedan anslutas till EU, efter att landet har uppfyllt de nödvändiga villkoren.
Trots att valet närmar sig har den nuvarande koalitionen ökat reformtakten, vilket EU har bemött på vederbörligt sätt.
De ansvariga på båda sidor bör gratuleras.
Både takten för de inhemska reformerna och EU:s svar bör snarare förr än senare nå den punkt där det inte finns någon återvändo.
Moldaviens förändring är givetvis beroende av en lösning på Transnistrienkonflikten.
I detta avseende uppmuntrades vi av de senaste diskussionerna om denna fråga som tillkännagavs vid toppmötet mellan Tyskland och Ryssland i Potsdam. Diskussionerna återupptogs vid det senaste trepartsmötet i Deauville, då man förmodligen drog fördel av Rysslands uppenbara villighet att nå en lösning.
Låt oss hålla våra löften och samarbeta för att denna sista rest av den ”latinska kulturen” ska föras in i EU.
(DE) Herr talman! När vi vid tidigare tillfällen har behandlat Balkanländerna, t.ex. när vi betonade problemen i Kosovo eller Bosnien, har vi tenderat att förbise Moldavien.
EU borde för länge sedan har iklätt sig rollen som medlare i de konflikter som berör Moldavien och dess grannländer.
Det är beklagligt att Moldavien nu har förkastat EU:s erbjudande att medla i Transnistrienkonflikten.
Det är ingen slump att Moldavien är den europeiska familjens styvbarn.
Det beror på landets kaotiska, före detta socialistiska ekonomi.
Som vi vet har det främsta industriområdet i östra Moldavien förklarat sin självständighet med stöd av Ryssland, och därigenom har regionen sanktionerat landets ekonomiska nedgång, eftersom ekonomin baseras uteslutande på jordbruket.
När Moldaviens medborgare går till valurnorna i slutet av november för att utse en ny regering är det viktigt att se till att valet avlöper väl för att förhindra ytterligare oro och en intensifiering av konflikten med t.ex. Rumänien.
(PL) Herr kommissionsledamot! Jag hade möjligheten att följa det förra valet i Moldavien.
När vi talade med företrädarna för de dåvarande oppositionspartierna uttryckte de en stor önskan om förändring.
Denna förändring har ägt rum.
Den nuvarande premiärministern Vlad Filat, som tidigare yttrade sig som företrädare för oppositionen, har tydligt förklarat sina europeiska strävanden.
Vi välkomnade effekterna av hans arbete när han besökte oss här i parlamentet.
Effekterna av hans arbete bekräftades också av delegationen från utskottet för utrikesfrågor som nyligen besökte Moldavien.
De inhemska problemen, i synnerhet frågan om Transnistrien, samt landets splittring och söndring, som är en symbol för landets förflutna och för dess delning, är mycket svåra frågor.
Vi måste stödja den process som kan möjliggöra att Transnistrien införlivas i Moldavien.
Här finns ett antal problem, däribland migrationsfrågan.
Herr kommissionsledamot, varje form av stöd till Moldavien, och här instämmer jag med min ledamotskollega...
(Talmannen avbröt talaren.)
(IT) Herr talman! Förra helgen reste jag till Chisinau i Moldavien.
Jag närvarade vid ett konvent som anordnats av kulturministern om Moldaviens integration i Europa med särskild hänvisning till kulturen.
Jag uppskattade väldigt mycket den stora önskan om tillväxt, framför allt genom en rad initiativ, som omfattade allt från byggandet av infrastruktur och vägar, elnät och andra typer av nät till yrkesutbildning för alla branscher och repetitionskurser för andra yrken.
Moldaviens befolkning är mycket intresserad av att anslutas till EU.
Regeringen strävar efter att Moldavien verkligen ska integreras i EU inom den närmaste framtiden, och man arbetar för detta.
Det är bra att EU för närvarande betonar ...
(Talmannen avbröt talaren.)
(EN) Herr talman! Antalet naturliga mottagare av EU-medel är för närvarande knappt hälften av det totala antalet medlemsstater.
I och med att vi utvidgar unionen till att omfatta alltfler, och till och med fattigare, öststater kommer andelen nettomottagare att öka till möjligen två tredjedelar.
Detta kommer självfallet att ske på bekostnad av nuvarande nettobetalare, men även på bekostnad av de medlemsstater som för närvarande är nettomottagare.
Vi får ofta höra att viseringslättnader inte kommer an på migrationen, och då åsyftas givetvis laglig migration.
Däremot finns ett klart samband mellan viseringslättnader och olaglig migration, dvs. smuggling av människor som arbetar för lägre ersättning än minimilöner och under arbetsförhållanden som inte uppfyller minimikrav.
Migrationen kommer också att leda till att landet töms på människor i arbetsför ålder som skulle kunna föra landet ut ur fattigdomen.
Slutligen vill jag säga att Moldavien förklarade sig självständigt från Sovjetunionen 1991.
Vill landet verkligen avstå från sin självständighet för EU, oavsett hur mycket det får motta i silvermynt?
ledamot av kommissionen. - (EN) Herr talman! Jag uppskattar verkligen den här diskussionen.
Jag uppskattar diskussionens läglighet och framför allt detta framstående parlaments tydligt enhetliga budskap och stöd.
Moldavien befinner sig vid en vändpunkt i landets historia.
Kommissionen har agerat aktivt för att hjälpa den moldaviska regeringen att uppnå så mycket som möjligt av sitt ambitiösa reformprogram under det senaste året.
De reformer som vi stöder återspeglar utan undantag de åtskilliga mål som finns med i handlingsplanen EU-Moldavien.
Det är avgörande för Moldaviens framtid att dessa reformer lyckas.
Vi har uttryckt vårt stöd för visionen om ett modernt och blomstrande Moldavien med en försonad befolkning. Vi stöder också landets territoriella integritet som har återupprättats vid så många tillfällen och inte bara den 30 september när den så kallade gruppen av vänner som Graham Watson hänvisade till besökte Chisinau.
Det råder inga tvivel om att vi genom EU:s historia har lärdomar att dela med oss av.
Moldavien är på god väg.
Jag är övertygad om att landet kommer att kunna nå den politiska kompromiss som krävs för att upprätthålla löftet om reformer.
Vi kommer i största möjliga utsträckning att fortsätta att stödja Moldaviens medborgare och tillhandahålla det externa stöd som krävs för reformerna.
Vi kommer att fortsätta att stödja dem för att de ska visa bärkraft vid det kommande parlamentsvalet.
Även jag hoppas uppriktigt att vi efter detta val kommer att få se en inkluderande politisk process i Moldavien som är inriktad på en proeuropeisk agenda, och att omvandlingsprocessen fortsätter till fördel för de moldaviska medborgarna och EU.
För att avsluta debatten har jag mottagit sex resolutionsförslag som ingetts i enlighet med artikel 110.2 i arbetsordningen.
Debatten är härmed avslutad.
Omröstningen kommer att äga rum i dag, torsdagen den 21 oktober 2010, kl. 12.00.
Skriftliga förklaringar (artikel 149)
Även jag välkomnar de framsteg som EU har gjort under det senaste året i förhållande till Moldavien.
Jag vill gratulera mina ledamotskolleger som har lagt fram detta resolutionsförslag.
Rumänien har allt sedan landets anslutning till EU engagerat sig för Moldaviens sak i EU.
Jag anser att ett konkret bevis på detta engagemang framgår av det antal rumänska parlamentsledamöter från olika politiska grupper som har gett sitt stöd till resolutionen.
De 90 miljoner euro som beviljats Moldavien i makroekonomiskt stöd har varit, och är fortfarande, den livlina som landet och dess medborgare behövt för att göra framsteg, och i synnerhet uppfylla de åtaganden som landet har gjort på området för reformer, rättsstatsprincipen och bekämpandet av korruptionen.
Moldavien har två huvudsakliga problem som måste få en lösning.
Det första gäller Transnistrien, där EU:s regeringar är tvungna att bidra på ett mer specifikt och beslutsamt sätt, samtidigt som förhandlingar måste återupptas.
Det andra problemet, som uppenbarligen kommer an på de demokratiska politiska aktörerna i Moldavien som vi bör uppmuntra, är det sätt på vilket valet kommer att genomföras den 28 november.
Vi måste garantera att medborgare både inom och utanför landet faktiskt har rätt att rösta fram en central regering.
Tack.
Avslutande av sammanträdet
(Sammanträdet avslutades kl. 23.40.)
1.
Användning av EU:s solidaritetsfond: Irland, översvämningar i november 2009 (
Avslutande av sammanträdet
(Sammanträdet avslutades kl. 23.40.)
Utökning av räckvidden för direktiv 2003/109/EG till att omfatta även personer som beviljats internationellt skydd (debatt)
Nästa punkt är ett betänkande av Claude Moraes, för utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor, om utökning av räckvidden för direktiv 2003/109/EG till att omfatta även personer som beviljats internationellt skydd - C6-0196/2007 -.
föredragande. - (EN) Herr talman! När jag nu inleder mitt inlägg är jag rädd att det bara kommer att vara jag själv, PPE-samordnaren och kommissionsledamoten kvar i kammaren.
Jag beundrar din uthållighet, Cecilia Malmström.
Jag borde inte ta av min talartid för att säga detta, men jag kunde inte låta bli.
Tack även till PPE-gruppen för att ni finns här vid denna sena timme.
Kommissionsledamot Cecilia Malmström! Du och rådet har gjort en enorm arbetsinsats för att rädda detta förslag som innebär att de som aldrig borde ha uteslutits från det ursprungliga direktivet om varaktigt bosatta tredjelandsmedborgares ställning nu garanteras sina rättigheter.
En ny chans att inkludera dessa medborgare gavs 2008, men tyvärr gick denna chans om intet eftersom rådet inte lyckades nå enhällighet i frågan.
Det är därför en glädjens dag i dag då man lyckats enas om ett förslag som lagts fram av en av mina föregångare som samordnare för min grupp, Martine Roure.
Jag känner även stor tacksamhet gentemot rådet.
I debatten tidigare, då rådet inte var närvarande, framhöll jag att om rådet varit närvarande här i dag skulle jag ha tackat rådet också, eftersom vi under Belgiens ordförandeskap gjort betydande framsteg.
Det är något jag är mycket tacksam för.
Förslaget kommer att få direkta positiva följder för alla som beviljats internationellt skydd och som har bott i EU i mer än fem år men inte kan få permanent uppehållstillstånd.
Det innebär ett slutgiltigt stopp för den särbehandling som dessa personer utsatts för i förhållande till andra tredjelandsmedborgare och ger dem ökad trygghet i EU.
Den centrala frågan i förhandlingarna har rört hur man ska beräkna den tidsperiod som en person uppehållit sig lagligt inom EU och som ska uppgå till fem år.
Vi stödde kommissionens uppfattning att även den tid då förfarandet pågått bör räknas med.
Men detta var något som rådet kraftigt motsatte sig.
Detta var en fråga som vi såg som mycket viktig, med tanke på att asylförfarandet i vissa medlemsstater kan ta många år.
Den kompromiss som vi har nått fram till i förhandlingarna innebär att åtminstone halva tiden för asylförfarandet kommer att räknas med. Om ett förfarande tar mer än 18 månader kommer tiden för hela förfarandet att räknas med.
Jag drar mig för att gå in på frågan om jämförelsetabeller, men jag är förpliktad att säga någonting om dem, även om jag helst skulle slippa.
Jag vill dock be institutionerna att försöka nå en överenskommelse sinsemellan i denna fråga.
Jag vill särskilt be rådet att tänka på hur viktigt det är med jämförelsetabeller för att kunna övervaka lagstiftningens genomförande.
Vi befann oss i en mycket besvärlig situation eftersom denna fråga kunde ha försenat många av de ärenden som olika grupper inom detta parlament ser som mycket viktiga.
Jag ser även mycket positivt på att förslaget innebär att såväl flyktingar som personer som beviljats subsidiärt skydd omfattas.
Vi måste se till att utvecklingen fortsätter när det gäller att sammanjämka skyddsnormerna med de rättigheter som båda dessa grupper har, som i det s.k. skyddsdirektivet.
Förslaget innehåller även många garantier mot ”refoulement” (dvs. utvisning eller avvisning av en person till ett land där denne riskerar att utsättas för trakasserier).
Med tanke på att flyktingar som beviljats skydd nu kan röra sig mellan olika medlemsstater är det viktigt att deras behov av skydd aldrig glöms bort.
Medlemsstaterna kommer därför att bli tvungna att göra en kommentar om detta i ett permanent uppehållstillstånd och måste i samband med en eventuell avvisning samråda med den medlemsstat som beviljade skyddet.
I förslaget tas även frågan om överföring av skyddsansvaret till en annan medlemsstat upp, något som regleras på nationell nivå.
Personens permanenta uppehållstillstånd måste då ändras så att det skyddar mot ”refoulement”.
Vi har också sett till att principen om att familjer ska hållas samman respekteras vid en avvisning till en annan medlemsstat, men att denna princip inte ska tillämpas per automatik om det inte kan anses ligga i övriga familjemedlemmars intresse att följa med den person som ska avvisas.
Den överenskommelse som vi nått i denna fråga är ett exempel på den nya typ av samarbete som kan ske mellan de tre institutionerna när det gäller asylfrågor och laglig migration tack vare de nya förutsättningar som Lissabonfördraget gett.
Det visar att vi kan nå en överenskommelse med medlemsstaterna om en progressiv lagstiftning på asylområdet.
Jag vill återigen tacka de olika gruppernas skuggföredragande samt Marya Nedelcheva, Cecilia Wikström och övriga kolleger som bidrog till att detta blev vad jag, paradoxalt nog, vill kalla en trevlig trepartsdiskussion.
Jag vill tacka alla de som bidragit till att detta blev möjligt.
Herr talman! Jag vill börja med att tacka Europaparlamentets föredragande Claude Moraes.
Han har gjort ett fantastiskt arbete tillsammans med sitt team av skuggföredragande.
Parlamentet, kommissionen och rådet har verkligen kunnat enas.
Även ministern har varit till stor hjälp.
Den kompromiss som har nåtts är välbalanserad och ligger i linje med förslaget från 2007.
Att personer som beviljats internationellt skydd kan få status som varaktigt bosatta i ett EU-land kommer att ge en högre skyddsnivå och ökad rättssäkerhet för flyktingar i Europa och kommer att underlätta deras integration i våra samhällen.
Detta utgör även den första byggstenen i vårt asylpolitiska paket - den första delen av ett lagstiftningspaket i sex delar - och det första steget mot vårt gemensamma mål att senast 2012 ha nått fram till ett gemensamt europeiskt asylsystem.
Det kommer att skicka en stark politisk signal om att vi kan nå enighet, att vi är beredda att slå in på denna svåra men nödvändiga väg och göra framsteg och att vi kan agera förnuftigt och konstruktivt i denna fråga.
Jag vill verkligen tacka er för detta.
När det gäller de så omtalade jämförelsetabellerna har kommissionen avgett en förklaring till rådet om detta.
Jag vill gärna läsa upp den för er: ”Kommissionen erinrar om sitt åtagande att se till att medlemsstaterna upprättar jämförelsetabeller som beskriver kopplingen mellan medlemsstaternas införlivandeåtgärder och EU-direktivet och att de översänder dem till kommissionen inom ramen för införlivandet av EU-lagstiftningen.
I kommissionens förslag från 2007 om ändring av direktivet om varaktigt bosatta tredjelandsmedborgares ställning framfördes kravet att det bör vara obligatoriskt med sådana jämförelsetabeller. Kommissionen beklagar att ett sådant krav inte fick något stöd.
Som en kompromiss och för att säkerställa att förslaget om ändring av direktivet om varaktigt bosatta tredjelandsmedborgares ställning kan antas utan dröjsmål kan kommissionen gå med på att kravet på att det ska vara obligatoriskt med jämförelsetabeller ersätts med en formulering där medlemsstaterna anmodas att se till att sådana tabeller upprättas.
Kommissionens hållning i detta ärende ska dock inte ses som prejudicerande.
Kommissionen kommer att fortsätta sina ansträngningar för att tillsammans med Europaparlamentet och rådet nå fram till en lämplig lösning i denna institutionsövergripande fråga.”
Jag tror vi kan enas om detta.
Det är viktigt att denna förklaring har förts fram och tas till protokollet.
Som jag sade tidigare i debatten står kommissionen fast vid denna ståndpunkt.
Men när det gäller just detta betänkande är det mycket viktigt att vi har nått en överenskommelse.
Jag vill återigen tacka er alla för era bidrag.
Herr talman, fru kommissionsledamot, Claude Moraes, mina damer och herrar! Först av allt vill jag ge föredraganden Claude Moraes en eloge för en utmärkt arbetsinsats och för ett exemplariskt samarbete med skuggföredragandena, kommissionen och rådet.
Med detta betänkande har vi tagit ett stort steg framåt mot ett samordnat europeiskt asylsystem.
Överenskommelsen med rådet var nödvändig och jag ser mycket positivt på att vi har lyckats nå framsteg i denna fråga.
Det asylpolitiska paketet omfattar dock mycket mer, och det finns också mycket kvar att uträtta här.
Vi får därför inte luta oss tillbaka och tro att man inom rådet kommer att vara lika samarbetsvillig vid framtida förhandlingar.
Detta vill jag ha sagt som en inledning.
När det gäller det innehållsmässiga vill jag, utan att upprepa vad föredraganden sagt, återkomma till två punkter.
Först och främst vill jag betona hur viktigt det är att tredjelandsmedborgare integreras i våra samhällen.
Invandrare som kommer till våra länder utgör en stor tillgång för våra ekonomier.
Men vi kan inte ta emot alla och på vilka villkor som helst.
Flera regeringar har under de senaste månaderna insett att deras integrationsmodell har varit ett misslyckande.
(Talmannen avbröt talaren.)
för ALDE-gruppen. - Herr talman! Låt mig först tacka vår föredragande Claude Moraes, som på ett för honom sedvanligt högkvalitativt sätt och med en uppriktig vilja att framhålla humanitära och medmänskliga principer har utarbetat det betänkande som vi har att ta ställning till.
Människor som har beviljats internationellt skydd i ett medlemsland kommer ofta att stanna där under mycket lång tid, kanske resten av sitt liv, eftersom utsatthet och förföljelse i det land de flytt från tenderar att bestå under mycket lång tid.
Många som har beviljats internationellt skydd befinner sig alltså i samma situation som dem som räknas som flyktingar.
Rimligen bör man också räknas som bofast i ett land när man har levt där i fem år. Det var också inriktningen hos både kommissionen och parlamentet.
Rådet ville annorlunda, vilket jag beklagar.
Jag vill också lyfta fram att familjemedlemmar till den person som har beviljats internationellt skydd måste ha egna möjligheter att gestalta sina liv.
Till exempel vid en utvisning så måste familjen få välja om man följer med eller stannar kvar.
Jag är glad över att parlamentet nu kommer att anta detta betänkande.
Jag beklagar att rådet inte har gått med på de så kallade correlation tables (jämförelsetabellerna) men jag välkomnar att vi går framåt med de betänkanden som ska ingå i det gemensamma europeiska asylpaketet.
Förhoppningen är att rådet nu ska inta en mer lyssnande hållning.
Vi har alla samma deadline att möta, och det är 2012.
Nu gäller det att lämna invanda positioner och se till den alleuropeiska hållningen och det gemensamma bästa när det gäller asyl- och migrationsfrågor.
Annars kommer ordet solidaritet snart att förlora sin betydelse.
Jag vill ånyo tacka föredraganden Claude Moraes för hans goda arbete och för ett mycket fint, för att inte säga excellent, samarbete med detta betänkande.
Herr talman! Förra veckan besökte jag Aten med utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor, och när jag var där talade jag med Mamuth.
Mamuth är 26 år gammal och kommer från Eritrea.
Han kom till Europa via Grekland och reste sedan vidare till Nederländerna där han hade velat stanna eftersom han har en del kontakter där, men han skickades tillbaka till Grekland.
Mamuth berättade att om han till slut får flyktingstatus i Grekland kommer han inte att kunna resa fritt och att det skulle ta evigheter att få grekiskt medborgarskap.
Det finns många fler som Mamuth som har rätt till ett nytt liv och inte förtjänar att bli skickade fram och tillbaka över gränserna, och det är för deras skull som jag gläder mig åt att detta parlament nu kommer att se till att denna situation ändras samt åt att Claude Moraes har lyckats ta det första steget mot ett asylpolitiskt paket.
Det är också viktigt att Mamuth, som alltså skulle föredra att leva sitt nya liv i Nederländerna, ges möjlighet att jämföra olika länder, för denne unge man har rätt att få veta hur olika frågor hanteras i Grekland respektive Nederländerna, eller var han nu skulle vilja bygga upp sitt nya liv.
Tack Claude Moraes, tack för ett gott samarbete. Nu får vi se hur lång tid processen tar för Mamuth.
(MT) Herr talman! Jag vill börja med att tacka Claude Moraes och ge honom en eloge för hans betänkande.
Jag stöder betänkandet och välkomnar det eftersom det kommer att innebära nya rättigheter för personer som ansöker om internationellt skydd, däribland flyktingar.
Det kommer att ge dessa personer vissa rättigheter som faktiskt redan ges till tredjelandsmedborgare som har bott lagligt i EU i fem år.
Men det finns några problem med detta betänkande.
Jag kommer från ett land som drabbats av det problem jag talar om, dvs. att fem år är en alldeles för lång tid för att få de rättigheter som denna lagstiftning avser.
Detta gäller i synnerhet i de länder som tar emot en enorm mängd människor som sedan blir kvar eftersom de fastnar i det land de först anlände till.
Förutom mitt eget land finns det även andra som under den senaste tiden drabbats av liknande problem, t.ex.
Grekland. Dessa länder tar emot ett stort antal människor som måste vänta fem år på att få de rättigheter som denna lag föreskriver.
Till slut kommer de förstås att få status som varaktigt bosatta och kommer då även att kunna flytta till andra EU-länder, vilket kan vara till stor hjälp för länder som Grekland, Malta, Cypern m.fl.
Jag anser således att denna lag visserligen är bra, men att den kunde ha gjorts bättre genom att den föreskrivna väntetiden på fem år hade kortats ned.
Jag vill avsluta med att tacka föredraganden Claude Moraes för att han uppmärksammat detta problem och gjort vad han kunnat genom att i slutet av motiveringsdelen införa en, må vara symbolisk, hänvisning till denna problematik.
(RO) Herr talman! Även jag vill börja med att ge min kollega Claude Moraes en eloge för detta betänkande.
Dessutom vill jag tacka honom för hans enastående insatser som samordnare inom utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor.
Jag tycker att det är alldeles förträffligt att detta nya direktiv äntligen kan fylla det rättsliga vakuum som rått när det gäller det problem med uppehållstillstånd som personer som beviljats internationellt skydd ställs inför inom EU.
Dessa människor som har bosatt sig i en EU-medlemsstat befinner sig i dagsläget i en vansklig situation när det gäller rättssäkerheten eftersom de under nuvarande förhållanden inte kan söka permanent uppehållstillstånd, till skillnad från andra tredjelandsmedborgare.
De ska inte diskrimineras, utan måste precis som andra tredjelandsmedborgare ha rätt till permanent uppehållstillstånd, med tidigare laglig bosättning som enda villkor.
Jag menar att det vid beräkningen av vistelsetiden hade varit bättre om man beaktat den totala tid som personen uppehållit sig lagligt inom EU, räknat från det datum då ansökan om internationellt skydd lämnades in.
Samtidigt måste man beakta att dessa människor alltid kommer att vara sårbara utanför EU, varför varje ansats till att dra in deras internationella skydd eller uppehållstillstånd måste ske med fullständig respekt för deras grundläggande rättigheter och i enlighet med principen om ”non-refoulement”.
Direktivet innehåller även bestämmelser för vilka förfaranden som ska tillämpas om det blir aktuellt med en avvisning eller ett upphävande av det internationella skyddet.
Jag anser att vi måste rösta för Claude Moraes betänkande, med tanke på att det utgör en del av ett större lagstiftningspaket för EU:s asyl- och migrationssystem.
(DE) Herr talman!
Jag betraktar inte detta betänkande genom ett rosenrött skimmer, utan jag väljer att se det utifrån ett perspektiv som omfattas av de medborgare i våra medlemsstater som oroas inför tanken att flyktingar som bott fem år i en medlemsstat ska beviljas permanent uppehållstillstånd.
Denna regel ska tillämpas inom hela EU:s territorium.
Detta innebär att när en flykting väl har bosatt sig i en medlemsstat som har relativt slapp asyllagstiftning kan denne efter fem år välja att bosätta sig i vilken annan medlemsstat som helst - och förstås kommer flyktingen att som första asylland välja det land som har den mjukaste lagstiftningen eller en lagstiftning med flest kryphål i för att sedan välja att bosätta sig permanent i ett land med hög social standard.
Detta kommer att resultera i sekundär migration och missbruk av reglerna.
Även ackumuleringen av fem års vistelse är en problematisk del av asylsystemet eftersom de administrativa förfarandena ofta fördröjs med avsikt och blir föremål för olika utredningar.
En utvidgning av direktivets räckvidd skulle innebära att en ännu större börda läggs på medlemsstater med hög social standard och som redan har enorma problem att brottas med utan att dessutom behöva försöka integrera flyktingar.
Jag kommer att ställa mig mycket kritisk till detta betänkande.
ledamot av kommissionen. - (EN) Herr talman! Jag har inte så mycket mer att tillägga.
Det råder stort samförstånd här för ett stöd för Claude Moraes insats när det gäller detta så viktiga direktiv.
Jag vill bara än en gång framhålla för Claude Moraes m.fl. vilken viktig byggsten detta utgör.
Jag tror att förslaget kommer att få ett starkt stöd vid omröstningen i morgon.
Det här är ett första steg på vår gemensamma väg mot 2012 och vårt asylpolitiska paket.
Jag hoppas bara att denna anda av konstruktivt samarbete kommer att fortsätta, eftersom jag behöver och även räknar med ert stöd i samband med övriga direktiv.
Herr talman! Jag vill uttryckligen tacka kommissionsledamoten för hennes arbete i denna fråga.
Vi hoppas att det första steget i asylfrågan kan fullbordas vid omröstningen i morgon - som jag hoppas innebär en överlägsen seger för förslaget - och ett av skälen till att vi hoppas på detta är att även om asylpolitiken kommer att fortsätta att vara en av de mycket känsliga frågorna i detta parlament, och framför allt för de mindre länderna, som Simon Busuttil också klargjort, kan varje liten del av asyllagstiftningen få oproportionerliga konsekvenser inte bara för de mindre länderna, utan även för t.ex. en konflikthärd som Grekland.
Vi bör alla gå fram med försiktighet, precis som vi gjort i detta betänkande. Det finns några punkter i motiveringsdelen som bör säkerställa att medlemsstaternas synpunkter tas på mycket stort allvar, inte minst när de kommer från medlemsstater som tar denna fråga på allvar.
Jag anser t.ex. att vi lyckats få med såväl Marya Nedelchevas synpunkter om integration som Cecilia Wikströms invändningar angående familjemedlemmar och avvisningar, samt även frågor rörande våld i hemmet och andra frågor.
Det är när vi har ett sådant samarbete som förhandlingarna går så bra på de högre nivåerna inom kommissionen och rådet, tack vare det arbete som vi utför här i parlamentet tillsammans med våra kolleger.
Och, Judith Sargentini, avslutningsvis har jag försökt komma på ett nytt sätt att uttrycka hur ytterst viktigt det är med jämförelsetabeller.
Att säga att de asylsökande nu väntar på att jämförelsetabeller ska införas är förmodligen det mest uppfinningsrika och kreativa sättet att lobba för en resolution om jämförelsetabeller, så jag hoppas att rådet lyssnade nu.
Jag vill återigen tacka alla mina kolleger för det stöd de gett detta betänkande efter så lång tid.
Debatten är härmed avslutad.
Omröstningen kommer att äga rum tisdagen den 14 december 2010.
Inkomna dokument: se protokollet
Frågestund (frågor till kommissionen)
Nästa punkt är frågestunden (B7-0001/2011).
Följande frågor har ställts till kommissionen:
Del I
Angående: Användning av EU-medel
Enligt en artikel nyligen i Financial Times har EU endast använt 10 procent av de 347 miljarder euro som anslagits för utveckling av fattiga regioner för perioden fram till 2013.
I artikeln sägs också att den finansiering som öronmärkts för små och medelstora företag har kommit att användas av multinationella bolag (Coca-Cola, IBM, Nokia Siemens) samtidigt som andra stora företag (Twining, Valeo) använder EU-medel för att flytta sina verksamheter till länder där arbetskraften är billigare och därigenom bryter mot bestämmelserna som uttryckligen förbjuder sådana metoder.
Vad anser kommissionen om uppgifterna i den artikeln och vilka åtgärder övervägs för att förhindra att liknande situationer uppkommer i framtiden?
Herr talman! Kommissionen välkomnar Financial Times granskning eftersom den ger ett viktigt bidrag till att inleda och bredda en allmän diskussion om sammanhållningspolitikens effektivitet och ändamålsenlighet.
Kommissionen är medveten om att användningen av medlen brukar vara långsammare i början på en programperiod.
De senaste uppgifterna visar dock att kommissionen har gjort fler betalningar inom ramen för sammanhållningspolitiken under det fjärde kvartalet 2010 än någonsin tidigare.
De allra flesta betalningarna var mellanliggande betalningar, dvs. ersättningar för utgifter som redan uppkommit och verifierats i medlemsstaterna.
Det är alltså säkert att takten i utnyttjandet av medlen för sammanhållningspolitiken ökar.
Utnyttjandenivåerna i form av EU-betalningar till medlemsstaterna är nu 21 procent för Sammanhållningsfonden, 22 procent för Europeiska regionala utvecklingsfonden och 23 procent för Europeiska socialfonden.
När det gäller stöd till multinationella och stora företag betonar kommissionen att ett primärt mål för sammanhållningspolitiken är tillväxt och skapandet av nya arbetstillfällen i vissa regioner och medlemsstater.
Allt stöd till produktiv investering måste ses i det sammanhanget.
Främjandet av arbetstillfällen och ekonomisk tillväxt kan uppnås på många sätt, från etablering av småföretag till att stödja större företag.
Insatserna inom sammanhållningspolitiken stöder produktiva investeringar som främst är inriktade på små och medelstora företag, i enlighet med föreskrifterna i förordningarna om Europeiska regionala utvecklingsfonden och Europeiska socialfonden.
Kommissionen betonar också den roll som små och medelstora företag spelade under förhandlingarna om de nuvarande programdokumenten.
De allra flesta produktiva investeringar och investeringar i utvecklingen av den inneboende potentialen är inriktade på små och medelstora företag.
Det kan dock förekomma fall då man i överensstämmelse med förordningarna beviljar medfinansiering till större företag under förutsättning att målen för de berörda fonderna och programmen respekteras.
Sammanlagt har 55 miljarder euro i företagsstöd beviljats mellan 2007 och 2013 inom ramen för sammanhållningspolitiken, varav en stor del utgörs av innovationsstöd till små och medelstora företag.
Kommissionen vill påpeka att multinationella företag inte är mottagare av stöd från Europeiska socialfonden.
Arbetstagare får samfinansierad utbildning.
Europeiska socialfonden stöder människor.
Det handlar om att tillhandahålla utbildning och omskolning samt att förbättra människors kompetens för att förbereda och hjälpa dem att hitta ett arbete.
En arbetstagare som anställs i ett visst företag kan mycket väl sedan bli anställd av ett annat företag.
Det viktiga är det kompetenskapital som arbetstagarna förvärvar så att de kan stanna kvar på arbetsmarknaden, inte vilken typ av företag som tillhandahåller utbildningen.
Från politisk synpunkt anser kommissionen att företag inte bör få EU-finansiering för investeringar som leder till förlust av arbetstillfällen i samma företag i en annan region i EU, eftersom nettoeffekten av ESF-investeringen då kan bli noll eller negativ.
I de fall då ett företag som har fått stöd från sammanhållningspolitiken lägger ned verksamheten eller slutar att stödja ett projekt inom fem år - eller tre år när det gäller små och medelstora företag - måste finansieringen betalas tillbaka.
Min sista - men viktiga - punkt är att även om det självklart finns utrymme för förbättringar bör och får inte detta överskugga de stora positiva effekter som sammanhållningspolitiken har.
Jag försäkrar er att kommissionen inte ryggar tillbaka inför problemen.
Vi har faktiskt tidigare föreslagit ändringar, varav en del fick gehör, och vi kommer att fortsätta att driva på för förbättringar av sammanhållningspolitiken.
Sammanhållningspolitiken ger klara fördelar för de fattigare regionerna i Europeiska unionen, men även klara fördelar för övriga Europa.
(RO) Jag vill tacka kommissionsledamoten även för kvaliteten på de upplysningar som har lämnats.
Jag vill dock göra ytterligare en kommentar.
I en debatt som denna om ett sådant ämne anser jag att vi snarare bör inrikta oss på framtida åtgärder för att se till att vi undviker liknande situationer och, om jag får lov att säga det, kanske det är ännu viktigare för oss att fråga oss själva om det inte är troligt att medborgarnas förtroende för EU-institutionernas arbete kommer att minska när dessa siffror blir allmänt uppmärksammade.
(DE) Herr talman, herr kommissionsledamot! Jag vill särskilt tacka för klargörandet eftersom det ger förutsättningar för en förnuftig diskussion och ett klart åtagande för våra små och medelstora företag.
Trots allt står de för två tredjedelar av Europas arbetstillfällen och betalar 80 procent av skatterna.
Min fråga är därför om du tror att vi i framtiden kan stärka ramförutsättningarna för forskning och forskningsinfrastrukturen en aning mer.
(LT) Herr talman! Jag har följande fråga.
Pengar från strukturfonderna och i synnerhet pengar från Europeiska socialfonden är mycket viktiga.
Medlen är avsedda att förbättra arbetstagarnas kvalifikationer och bevara arbeten så att de utförs av kvalificerade personer.
Anser du att det råder lika villkor för rika internationella företag, eftersom de själva måste ge ett bidrag för att kunna få medel från strukturfonderna eller Europeiska socialfonden, och små och medelstora företag, som också vill utbilda sitt folk och vill ha kvalificerade anställda?
Planerar du inte någon form av förslag här, eftersom villkoren inte är lika för stora företag och för små och medelstora företag?
Herr talman! Tack för era frågor.
När det gäller forskningens infrastruktur får små och medelstora företag redan betydande resurser från Europeiska regionala utvecklingsfonden, särskilt för att främja innovation - där de får innovationsstöd i storleksordningen tiotals miljarder euro.
Under perioden 2000-2006 inriktade sig över 30 000 företag på detta område på ett fokuserat sätt.
Vi funderar över att stor vikt också bör fästas vid forskningsinfrastrukturen, särskilt i framtiden - inte bara på det ekonomiska området, utan även inom grundforskningen.
Det är möjligt att vi även under den innevarande perioden kommer att stödja forskningsinfrastrukturprojekt som också ingår i färdplanen för Esfri - Europeiska strategiska forumet för forskningsinfrastruktur - med sådana medel för första gången, eftersom undersökningar av projektet har visat att det har en mycket varaktig effekt i en region utöver själva projektet genom de arbetstillfällen som kommer att skapas, inte bara forskningsarbeten, utan även i leverantörsföretag eftersom även grundforskningsinfrastruktur behöver tjänster och förnödenheter.
Med andra ord kan det bli ett verkligt nav i ett visst område i en region - i detta fall en region i Ungern.
Detta ska också skicka ut en signal inför den kommande programperioden, kanske till universiteten, vilket till sist också kommer att få konkreta effekter.
Redan i dag sker nästan en tredjedel av universitetsforskningen inom tillämpad forskning, vilket till sist är till godo för ekonomin och skapar varaktiga arbetstillfällen.
Om jag får lov går jag nu över till damens fråga. Inom ramen för Europeiska socialfonden är det i allmänhet anställda eller tillfälligt arbetslösa som får stöd till utbildning för att förbättra sina förutsättningar på arbetsmarknaden.
Detta kan ske inom det företag där de är anställda. Om de inte är anställda kan det vara för att förbättra deras färdigheter eller helt enkelt göra dem generellt bättre kvalificerade för andra tänkbara typer av arbeten.
Jag kan ge ett exempel - eftersom det kanske var detta som du syftade på och eftersom det har utsatts för mycket kritik - och det är anställda hos McDonald's som har erbjudits vidareutbildning.
Här måste vi göra en klar åtskillnad: det rörde sig om utbildningsåtgärder för McDonald's anställda för att göra dem bättre kvalificerade på arbetsmarknaden och i arbetslivet.
Som ni vet - det har faktiskt fått en del kritik - är arbeten hos McDonald's, eller med ett engelskt slanguttryck McJobs, i allmänhet deltidsanställningar som inte kräver några större kvalifikationer. Dessa arbeten utförs ofta av studerande.
Det handlar om att höja deras kompetens.
När det gäller intern fortbildning, som i det här projektet, bar exempelvis McDonald's alla kostnader själv.
Med andra ord försöker och strävar vi efter att se till att den fortbildning de anställda får koncentreras på deras personliga kvalifikationer.
Därför anser jag att det inte bör göra någon skillnad om personerna är anställda eller inte. Vårt mål måste i stället vara att ytterligare förbättra kvaliteten på varje persons färdigheter så att de blir mer lämpade för en alltmer rörlig arbetsmarknad och därmed att så långt möjligt undvika arbetslöshet.
Angående: Europeiska instrumentet Progress för mikrokrediter
Genomförandet av det europeiska instrumentet Progress för mikrokrediter för sysselsättning och social delaktighet förfaller gå långsammare än väntat, vilket kan äventyra dess syfte och står i stark kontrast till den hastighet med vilken instrumentet antogs i mars 2010.
Vad tänker kommissionen göra för att påskynda processen och se till att instrumentet når ut till de mest sårbara människorna samtidigt som den rätta geografiska balansen tryggas?
Vad tänker kommissionen göra för att få medlemsstaterna att finansiera mentors- och utbildningsprogram och för att även säkerställa att räntebetalningar subventioneras med medel från Europeiska socialfonden så som man kommit överens om?
Hur kommer kommissionen att se till att informationen om Progress-instrumentet för mikrokrediter når ut till målgrupperna?
Kära kolleger! Jag är glad över att kunna rapportera att båda delarna av europeiska instrumentet Progress för mikrokrediter - garantidelen och kontantdelen - nu är helt operativa.
Endast tre månader efter ikraftträdandet av beslutet har kommissionen färdigställt mandatet för Europeiska investeringsfonden att starta garantiinsatser för tillhandahållare av mikrofinansiering.
I november inrättade kommissionen en särskild investeringsfond.
Det gör att de första mikrolånen kommer att börja tillhandahållas den här månaden.
Jag är också glad över att rapportera att kommissionen har lyckats säkerställa ytterligare medel för mikroföretagare i Europa.
Europeiska investeringsbanken kommer att svara för EU:s bidrag på 100 miljoner euro, och fler bidragsgivare kan förväntas.
Det gör att den totala lånevolymen inom ramen för instrumentet Progress för mikrokrediter som väntat kommer att uppgå till cirka 500 miljoner euro.
Dessa pengar kommer att vara till nytta för arbetslösa, för människor som riskerar social utestängning och för utsatta människor som har svårt att få tillgång till den vanliga kreditmarknaden.
Två viktiga punkter i kommissionens uppdrag till Europeiska investeringsfonden är att säkerställa att instrumentet når ut till målgrupperna och att främja den geografiska balansen.
De åtgärder som hittills har godkänts eller håller på att förberedas tyder på att båda målen kommer att uppnås.
Från och med början av 2011 kommer mikrolån att tillhandahållas genom en inledande mikrofinansieringsinstitution i Belgien som är inriktad på missgynnade stadssamhällen, och genom en stiftelse i Nederländerna som är inriktad på enskilda personer som saknar tillgång till vanlig finansiering.
Europeiska investeringsfonden har tillkännagett att de åtgärder som håller på att förberedas även kommer att få en balanserad geografisk täckning.
Cirka 40 procent förväntas involvera förmedlare som investerar i Europa och cirka 60 procent i Central- och Östeuropa.
Det är välkänt att mikrofinansiering är mest effektivt om nyföretagare och mikroföretag ledsagas genom stödtjänster för företag.
Kommissionen kommer därför att vidta åtgärder för att stödja de myndigheter som förvaltar medlen från Europeiska socialfonden och förmedlande organ för att intensifiera främjandet av egenföretagande och mikroföretag.
Under den innevarande programperioden för Europeiska socialfonden har medlemsstaterna öronmärkt över 2,7 miljarder euro för att främja företagande.
Företagare kan också stödjas genom räntesubventioner.
Det är de enskilda medlemsstaterna som bestämmer om räntor ska subventioneras via Europeiska socialfonden eller inte.
För närvarande har endast en medlemsstat, Litauen, meddelat att den utnyttjar denna möjlighet.
Slutligen kommer kommissionen att främja information om instrumentet Progress för mikrokrediter.
De som tillhandahåller mikrokrediter och befinner sig närmast de tilltänkta mottagarna kommer att informera om att mikrolån är tillgängliga.
Kommissionen kommer att använda de befintliga nätverken av arbetsförmedlingar, Europeiska socialfondens förvaltningsmyndigheter och icke-statliga organisationer och informera om framstegen inom instrumentet Progress för mikrokrediter.
Sist men inte minst kommer man inom kampanjen Unga på väg att ägna särskild uppmärksamhet åt möjligheterna för unga från olika bakgrunder att starta egna företag och få mikrolån.
(HU) Herr talman! Det gläder mig att höra kommissionsledamotens rapport, och jag vill klargöra en del.
När vi fick rapporten från kommissionen och Europeiska investeringsfonden för ett par veckor sedan nämndes en totalsumma på ungefär 200 miljoner euro.
En av mina frågor gällde just detta att det ursprungliga löftet eller planen var 500 miljoner euro.
Jag skulle vilja veta var dessa ytterligare medel kom ifrån.
Jag anser att det är mycket viktigt eftersom detta är ett högprioriterat program för att begränsa effekterna av krisen, och det var delvis därför som vi skyndade på med antagandet.
Den andra viktiga frågan var om medlemsstaterna stöder subventioner av räntebetalningar samt utbildnings- och mentorinslagen från socialfonden.
Detta ingick också i den ursprungliga planen, och sedan tycktes kommissionen försumma frågan.
Det är mycket viktigt att lämna information och att se till att informationen når ut till människor.
(PL) Herr talman, herr kommissionsledamot! Jag vill tacka dig för den här informationen.
Jag håller helt med om att det instrument som vi diskuterar i dag är mycket viktigt.
Det är dock värt att nämna att vi också bör svara på frågan om vilka stater som utnyttjar instrumentet Progress för mikrokrediter.
Det oroade mig att du sade i ditt svar att vi bör sörja för olika fördelningsnivåer efter stat och geografiskt område.
Har några stater hittills använt instrumentet?
(RO) Herr talman! De unga är de som helt klart har drabbats hårdast av den ekonomiska och finansiella krisen, men vi får inte heller glömma arbetslösa människor som är äldre än 45 år.
Jag vill ställa följande fråga till kommissionsledamoten, eftersom du nämnde att 60 procent av det europeiska instrumentet Progress för mikrokrediter kommer att gå till Central- och Östeuropa: Har du tagit reda på vad det är som hittills har förhindrat att länderna i denna del av Europa utnyttjar instrumentet tillräckligt?
Tack för ert intresse och era kommentarer.
Ämnet mikrokrediter täcks faktiskt av flera generaldirektorat, och László Andor har en viss ledande roll när det gäller innehållet.
Det är dock också något som vi är berörda av på det regionalpolitiska området.
När det gäller räntenivåer finns det vissa medlemsstater som har bestämt ett tak - som ett villkor så att säga - som ligger på ungefär 8 till 9,5 procent.
Det som också måste beaktas är dock naturligtvis - och detta har redan diskuteras, bland annat under förberedelserna för allt detta - att omkostnaderna är relativt höga i förhållande till de faktiska lånen och därmed de kostnader som måste täckas.
En förnuftig medelväg måste hittas, vilket jag anser att vi har lyckats med.
Jag går nu över till den andra frågan och kan berätta för er att instrumentet Jasmin - som är avsett att stödja lämpliga förberedelser för mikrokrediter och bana väg för förmedlarna att etablera och utbilda sig - för närvarande används för att förbereda 15 institutioner i 15 olika länder, vara elva finns i Central- och Östeuropa och fyra i Västeuropa.
Jag kan inte plocka fram alla länderna direkt från minnet, men det handlar framför allt om de nya anslutningsländerna, och vi förväntar oss att ytterligare 20 förmedlare kommer att förberedas enligt Jasminprogrammet under de kommande åren.
När det gäller den sista frågan måste jag be er ursäkta att jag inte kan ge er ett svar direkt.
Ni kommer att få ett skriftligt svar med utförliga förklaringar av det begränsade tillträdet.
Jag antar dock att det säkerligen ofta är kommunikationsproblem här och att det också ofta finns hinder eftersom många av de potentiella låntagarna är personer som inte längre kan få lån från vanliga banker, och det finns därför ofta en viss oro eller tveksamhet när det gäller att närma sig sådana inrättningar.
Om så är fallet och det blir en ingrodd och etablerad uppfattning är det dock nödvändigt att genomföra lämpliga informationsverksamheter på området.
Angående: Ytterligare stödåtgärder för små och medelstora företag inom ramen för turismpolitiken
Världskonkurrensens effekter är kännbara inom turismen precis som inom andra delar av ekonomin.
För att Europeiska unionen ska förbli konkurrenskraftig inom sektorn har EU i Lissabonfördraget uppställt som mål att främja konkurrenskraften och skapa en miljö som är gynnsam för affärsutveckling.
För detta ändamål har följande mål antagits: främja innovation inom turism, förbättra den allmänna kvaliteten på turisttjänster och utveckla personalens yrkeskunskaper.
Företag inom turismsektorn - varav många är små och medelstora företag - klarar inte alltid att uppnå dessa mål genom sina egna insatser utan stöd.
Detta beror på flera faktorer, till exempel begränsade ekonomiska resurser, brist på utbildad personal och oförmåga att snabbt reagera på förändring: därav behovet av ytterligare finansiering.
Anser inte kommissionen att det skulle vara önskvärt att utforma en samordnad strategi och en detaljerad handlingsplan som innefattar stödåtgärder för små och medelstora företag samt finansieringsåtgärder som skulle kunna bidra till att övervinna svårigheterna inom sektorn?
Herr talman, mina damer och herrar! Den europeiska turistbranschen möter liksom många andra ekonomiska sektorer den allt större utmaningen från globaliseringen.
Detta är en utmaning som kommissionen redan har betonat och tagit itu med vid flera tillfällen, särskilt i meddelandet ”En integrerad industripolitik för en globaliserad tid”.
Den 30 juni förra året antog kommissionen ett särskilt meddelande om turismen, med förslag - i enlighet med Lissabonfördraget och den nya Europa 2020-strategin - till ett konsoliderat politiskt ramverk för att förstärka konkurrenskraften inom sektorn för att göra europeisk turism till en verklig konkurrenskraftig, modern, hållbar och ansvarsfull bransch.
Skapandet av en miljö som befordrar utvecklingen av mikroföretag, små och medelstora företag inom turismsektorn är den princip som denna konsoliderade ram grundas på.
För att uppnå detta mål föreslog vi tre särskilda mål: för det första att stimulera konkurrenskraften inom den europeiska turismsektorn, för det andra att främja utvecklingen av hållbar, ansvarsfull turism av hög kvalitet och för det tredje att konsolidera Europas anseende och profil som en samling av hållbara turistmål och naturligtvis att maximera EU:s ekonomiska politik och instrument för att utveckla turism.
De initiativ som främjas bör ge sektorn de nödvändiga instrumenten för anpassning till de utmaningar som dess näringsidkare står inför och arbeta mot en hållbar utveckling av sektorn i fråga om konkurrenskraft.
Särskilda åtgärder kommer naturligtvis att vidtas för att främja innovation inom turismsektorn, förstärka kvaliteten på de anställdas yrkeskunskaper, eftersom vi inte längre får betrakta turism som en sektor som enbart består av familjeföretag. Vi måste också beakta hur vi kan göra den mer modern och konkurrenskraftig.
Jag ska ge ett par exempel på utbildning och yrkeskunskaper: en IKT- och turismplattform kommer att lanseras för att underlätta sektorns och dess företags anpassning till utvecklingen inom marknaden för nya informationstekniker och förbättra deras konkurrenskraft.
Alla dessa förslag och idéer finns med i kommissionens meddelande, som har godkänts av rådet och som vi debatterar i parlamentet - föredraganden är närvarande i kammaren.
Branschens företagare kommer att uppmuntras att utnyttja unionens olika program, till exempel Leonardo, ramprogrammet för konkurrenskraft och innovation, Erasmus för unga entreprenörer, Europeiska socialfonden och andra program.
En strategi för att främja diversifiering av turisttjänster och tillkomsten av ett elektroniskt observatorium för europeisk turism kommer också att bidra till att skapa en gynnsam miljö för sektorns aktörer.
Dessutom måste jag påpeka att små och medelstora företag kan dra nytta av andra generella initiativ för att få tillgång till finansiering.
Jag vill nämna kommissionens gemensamma initiativ Jeremie, Europeiska investeringsfonden och Europeiska investeringsbanken, som syftar till att förbättra tillgången till medel särskilt för mikroföretag, små och medelstora företag genom kanalisering av riskkapital, lån, säkerheter, mikrokrediter och andra former av återbetalningspliktigt stöd.
Till sist vill jag påpeka att små och medelstora företag inom turistsektorn helt täcks av de åtgärder som föreslås inom ramen för småföretagsakten, vars syfte är att främja affärsklimatet för just dessa företag.
Parlamentet kommer att få den uppdaterade texten om ett par veckor.
Småföretagsakten kommer alltså att bli ett instrument för att skydda små och medelstora företag som erbjuder en stor potential för utvecklingen av en sektor som jag hoppas ska kunna förstärkas under det närmaste året, eftersom jag är absolut övertygad om att en europeisk politik i enlighet med fördraget kan ge mervärde åt det utmärkta arbete som redan utförs av Europas regioner och medlemsstaterna.
Jag kan därför försäkra ledamoten som ställde frågan att kommissionen och jag själv har åtagit oss att se till att alla små och medelstora företag inom sektorn får stöd och hjälp i sina försök att få tillgång till EU:s ekonomiska instrument som ett led i en politisk strategi för att göra turismen till en av våra viktigaste näringslivssektorer.
(LT) Herr talman! Förmodligen hoppas alla vi som är här i parlamentet i dag att den prognos som kommissionsledamoten gav om turismens framtida utveckling faktiskt kommer att bli verklighet och att området inte bara kommer att utvecklas utan att även vara gynnsamt för investeringar.
Som ni vet är turismen hittills ojämnt utvecklad inom Europeiska unionen, och det finns objektiva och subjektiva skäl till det.
Jag har en fråga.
I Östersjöstrategin anges Östersjöregionen som ett av huvudmålen.
Vad har egentligen uppnåtts på detta område under året?
(IT) Herr talman, herr kommissionsledamot, mina damer och herrar! Jag vill tacka Zigmantas Balčytis för denna fråga som sätter i centrum för vår diskussion att parlamentet vill få möjlighet att inom de närmaste månaderna återigen behandla det parlamentsbetänkande som jag är ansvarig för.
Först och främst måste vi ge kommissionens vice ordförande Antonio Tajani en eloge för att ha gett ett mycket starkt stöd till den nya europeiska turismpolitik som föreskrivs i Lissabonfördraget med det meddelande som antogs i juni och den genomförandeplan som lades fram för ett par veckor sedan.
Dessa två dokument är särskilt inriktade på små och medelstora företag och på konkurrenskraften inom sektorn, med särskild betoning av innovations- och utbildningsfrågor.
I fråga om finansiering måste vi agera på två fronter: För det första måste vi öka medvetenheten om att fonderna finns och se till att de utnyttjas mer, och för det andra måste parlamentet starkt förespråka - herr talman, jag avslutar här - införlivandet av budgetrubrikerna för turismpolitiken i budgetramen för perioden 2014-2020.
(RO) Det finns vissa länder som till exempel använder det regionala programmet för konkurrenskraft och innovation eller det operativa programmet för att utveckla turism och när det gäller Grekland det operativa programmet för regional utveckling.
Jag vill fråga dig om du tänker inrätta en europeisk ram för att öka de små och medelstora företagens utnyttjande av EU-medel för utveckling av turismen.
Jag vill tacka Zigmantas Balčytis eftersom han har gett mig möjlighet att tala om den fråga som av alla dem som jag ansvarar för som kommissionsledamot ligger mig närmast om hjärtat. Som den första kommissionsledamoten för turism anser jag att turismpolitiken tillsammans med industri- och rymdpolitiken är prioriterade.
För att ge ett konkret svar är den centrala frågan förutom de politiska initiativ som jag har försökt att genomföra sedan jag blev kommissionsledamot den som Carlo Fidanza tog upp i sitt inlägg: eftersom EU inte ansvarade för turismpolitiken före Lissabonfördragets ikraftträdande ingår inte de medel som behövs för EU ska kunna bidra till en stark insats för turismen i den aktuella budgetramen.
Vi har intressanta program som exempelvis Kalypso, som i Spanien har förstärkt med ett antal i mina ögon mycket positiva initiativ.
Jag förstår dock klart den poäng som Carlo Fidanza gör i det betänkande som parlamentet är på väg att lägga fram, men det kommer att finnas stöd eftersom de medel som är öronmärkta för turismpolitiken kommer att ökas i nästa budgetram.
De kan ökas i det åttonde ramprogrammet eller genom införande av särskilda budgetposter.
Det viktiga är dock att parlamentet tar fram problemet i ljuset eftersom det är svårt att ge konkreta svar om de ekonomiska instrumenten inte finns på plats.
Detta innebär dock inte att vi inte kommer att agera mycket bestämt.
Som ni vet har ett otal initiativ tagits, det belgiska ordförandeskapet arrangerade ett stort evenemang på Malta och det ungerska ordförandeskapet har redan tillkännagett att det kommer att arrangera ett särskilt evenemang för turism - detta var ämnet för vårt första möte, som hölls i Budapest för ett par dagar sedan.
Jag är glad över att Zigmantas Balčytis tog upp frågan om turism i Östersjöområdet: turism är inte en fråga som enbart rör ekonomierna i Medelhavsländerna - Spanien, Frankrike, Italien, Grekland och Malta.
Det är en ytterst viktig resurs för hela Europeiska unionen, inklusive länderna i Central- och Östeuropa, som har egna turistorter och en egen potential att utveckla.
När det gäller Östersjöstaterna anser jag att en av frågorna - som för övrigt tas upp i den text som godkändes den 30 juni förra året - är relationen till de nya framväxande klasserna, till den nya medelklassen i Ryssland.
Miljontals ryssar planerar att turista och alltså att resa utanför sitt eget land.
Vi har ett problem när det gäller viseringar.
Samma problem finns i fråga om Kina, misstänker jag. Kommissionen och turismministrarna är beredda att försöka lösa problemet med potentiella besökare från både Ryssland och Kina.
Vi vill skynda på det hela och göra det enklare för dem att få komma till våra länder.
Dessutom är Östersjöstaterna närmare Ryssland och kan skörda de potentiella ekonomiska fördelarna av att ta emot turister även från den växande medelklassen.
Detta är centralt för vårt arbete att främja turismpolitiken, och jag är också uppmuntrad av att många ministrar från olika medlemsstater, inklusive Storbritannien - jag träffade den nya brittiska turismministern för ett par veckor sedan i London - och Frankrike är positiva till att stödja EU:s turismpolitik.
Det är viktigt att identifiera ett antal ingångsportar, eftersom Europa måste representera ett mervärde.
Jag är glad över att kommissionsledamot Androulla Vassiliou i den text om idrott som antogs i dag har försökt ta in synpunkten att stora idrottsevenemang, som den kommande olympiaden i London, är ett utmärkt tillfälle för hela Europeiska unionen.
Kort sagt måste vi se till att varje land i EU kan agera som en ingångsport för turister som besöker det landet men sedan reser vidare och besöker andra europeiska länder när de är klara.
Detta är den ytterligare åtgärd som kommissionen kan vidta, och jag anser att parlamentets stöd är viktigt.
Får jag lov att tacka er nu för era framtida insatser, bland annat i diskussionen om turismpolitiken men även i alla diskussioner om de kommande budgetverksamheterna.
Del II
Angående: Program och initiativ för att modernisera den högre utbildningen
Studier har genomförts i vissa medlemsstater för att ta reda på hur högskoleinstitutioner har anpassats till de nya kraven på arbetsmarknaden och vilka utsikter de studerande har att hitta ett arbete när de är klara med sin examensutbildning.
Forskningen har tyvärr visat att många universitet utbildar specialister för en marknad som redan är mättad.
Högskolornas studieplaner tar inte alltid hänsyn till arbetsmarknadens behov och de som drabbas mest av detta är därför de nyutexaminerade.
I sitt arbetsprogram för 2011 nämner kommissionen modernisering av den högre utbildningen och anger att förslag kan komma att läggas fram om det system som ska tillämpas för att bedöma och öka insynen i högskoleinstitutionernas verksamheter.
Eftersom så är fallet, vilka särskilda program- och modellinitiativ kommer kommissionen att anta för att modernisera den högre utbildningen i Europa?
Kommer kommissionen att utarbeta en särskild strategi för den högre utbildningen för att se till att unga nyutexaminerade kan hitta ett arbete så snart som möjligt?
Hur mycket är kommissionen redo att satsa i framtida program och initiativ av detta slag för ungdomar?
Herr talman! Utbildning är bara en av de viktiga faktorer som bestämmer anställbarheten.
Risken att bli arbetslös är 40 procent lägre för personer med examen från högre utbildning än för sådana som endast har gymnasieutbildning.
Arbetslösheten och undersysselsättningen bland ungdomar är dock oacceptabelt hög i dag.
Alltför många utexaminerade kämpar för att klara steget ut på arbetsmarknaden och få ett kvalitetsarbete som motsvarar deras utbildningsbakgrund.
Insatserna för att förbättra anställbarheten börjar naturligtvis långt före den högre utbildningen.
Kommissionen arbetar med medlemsstaterna för att identifiera de färdigheter eller nyckelkompetenser som ungdomar behöver för att lära sig i skolan.
I dag behöver unga ett bredare spektrum av färdigheter än tidigare för att kunna leva och verka i en globaliserad ekonomi.
Många kommer att bli verksamma i arbeten som ännu inte finns.
Många kommer att behöva avancerade färdigheter i språk, interkulturella förbindelser och företagande.
Tekniken kommer att fortsätta att förändra världen på sätt som vi inte kan föreställa oss så att förmågan att fortsätta att lära sig och vara innovativ kommer att bli viktiga faktorer för anställbarheten.
Vägledning är också viktigt.
Unga människor möter ett allt större utbud av utbildningsalternativ.
De behöver kunna fatta informerade beslut.
För detta krävs bättre information om utbildningsvägar, bland annat en klar bild av möjligheterna att få arbete.
Vi behöver utveckla en yrkesmässig vägledning av kvalitet och en yrkesutbildning med ett starkt engagemang av arbetsmarknadens institutioner.
Om vi går över till högre utbildning har kommissionen som ni vet nyligen lanserat Ungdom på väg - ett flaggskeppsinitiativ inom Europa 2020-strategin för att göra utbildningen mer relevant för unga människors behov.
Vi börjar nu genomföra olika delar av den strategin.
Senare under året planerar kommissionen ett nytt meddelande om modernisering av den högre utbildningen.
Vi kommer att mäta framstegen i att göra den högre utbildningen mer relevant för behoven i det kunskapsbaserade samhället, inklusive frågan om anställbarhet.
Vi kommer att identifiera de viktigaste utmaningarna för framtiden och ge vårt svar.
Som ett led i dessa ansträngningar kommer kommissionen att förstärka den europeiska plattformen för dialog mellan universitet och företag för att öka de studerandes anställbarhet och utveckla utbildningens roll i kunskapstriangeln.
I en mer global och rörlig värld kan öppenhet om högskoleinstitutionernas resultat stimulera både konkurrens och samarbete och bli ett incitament för fortsatta förbättringar och modernisering.
Befintliga internationella rangordningar kan dock ge en ofullständig bild av universitetens resultat.
I år kommer kommissionen att lägga fram resultaten av en förstudie för att utveckla ett alternativt och flerdimensionellt rangordningssystem som avspeglar högskoleinstitutionernas mångfald.
Europa behöver bli bättre på att förutse morgondagens behov av kompetens.
Därför har kommissionen lanserat En agenda för ny kompetens och nya arbetstillfällen, som går hand i hand med vårt initiativ Unga på väg.
Genom En agenda för ny kompetens och nya arbetstillfällen tittar vi på hur vi kan hjälpa våra ungdomar att bli mer anställbara.
Framför allt behöver vi ge människor rätt kombination av färdigheter så att de kan anpassa sig till vårt snabbföränderliga samhälle.
Vår nya kompetenskarta för EU, som blir operativ 2012, kommer att hjälpa till att prognostisera inte bara de färdigheter som arbetsgivarna behöver i dag, utan också de färdigheter som behövs i framtiden.
I vår tänker kommissionen föreslå nya europeiska riktmärken för rörlighet i utbildningssyfte och om utbildningens roll för att göra människor anställbara på den kunskapsbaserade arbetsmarknaden.
EU-programmen för att stödja utbildning och ungdomar, inklusive program för rörlighet som Erasmus, kan hjälpa ungdomar att förbättra sina chanser på arbetsmarknaden genom att tillägna sig värdefull internationell erfarenhet och utveckla sin intellektuella förståelse.
(LT) Herr talman, fru kommissionsledamot! Tack för ditt verkligt utförliga svar.
Jag skulle dock vilja ställa en följdfråga.
Europeiska unionen måste garantera alla medborgare rätt till högre utbildning av god kvalitet.
I medlemsstaterna finns det dock många skillnader mellan utbildningssystemen, kostnaderna för högre utbildning och tillhandahållandet av lån för att betala studierna.
Hög ränta på lån som tagits för att betala studierna och ogynnsamma villkor för återbetalning av lånen avskräcker ofta ungdomar från att bedriva högre utbildning i sitt eget land och främjar en kompetensflykt till andra länder.
Tänker kommissionen publicera en vägledning om önskade villkor för tillhandahållande av studielån?
(PL) Herr talman! Jag vill ställa en enda fråga till kommissionsledamoten, även om vi diskuterar olika saker just nu.
Jag vill fråga kommissionsledamoten om något arbete sker för att öka medlen för utbytesprogram för studerande i Europa.
Jag har intrycket att den finansieringspool som vi har för Erasmus och andra program har varit oförändrad i flera år.
För närvarande är dessa stipendier verkligen mycket låga.
(EL) Fru kommissionsledamot! Det är riktigt att denna särskilda fråga omfattas av subsidiaritet.
Medlemsstaterna finansieras dock av medel från EU för att modernisera utbildningsplanerna i medlemsstaterna.
Under exempelvis den tidigare och tredje stödramen från gemenskapen utnyttjade många medlemsstater gemenskapsmedel för detta ändamål.
Jag har en mycket konkret fråga: Har kommissionen uppgifter om effektiviteten av de medel som gavs och kommer att ges till medlemsstaterna?
För det första om frågan om skillnader mellan högskoleinstitutioner: Det stämmer exakt!
Det är därför som vi vill ha insyn i universitetens resultat.
Det är därför som vi nu slutför förstudien på vars grund vi ska våga titta på rangordningen av universitet, kartläggning av universiteten och deras standarder för att ge de studerande bättre informerade alternativ.
Målet är att de ska veta var de ska studera, vad de ska studera och vilken standard universitetet har som de söker sig till.
I fråga om avgifter håller jag nog med om att höga avgifter kräver rättvisa lån, men ni vet säkert att detta är medlemsstaternas ansvar.
Vi vet att det enda som ekonomerna är överens om är att investering i utbildning ger långsiktiga resultat, tillväxt och arbeten. Jag uppmanar därför alltid regeringarna att inte skära ned universitetsinvesteringarna eller utbildningsinvesteringarna i allmänhet.
Jag håller dock med ledamoten som ställde frågan om otillräckligheten av rörlighetsstöd som Erasmus.
Det är därför vi återigen genomför en förstudie - som utförs av London School of Economics, som jag hoppas kommer att vara klar om ett par månader - på grundval av vilken vi tillsammans med Europeiska investeringsbanken ska undersöka möjligheterna att skapa ett europeiskt studielån för rörlighet.
Jag är säker på att detta kommer att ge alla studerande, oavsett om de är fattiga eller rika, möjlighet att utnyttja dessa förträffliga rörlighetsbidrag.
När det gäller Georgios Papanikolaous fråga talade han om strukturutvecklingsmedel som regeringarna kan använda till att bygga upp sin utbildningsinfrastruktur.
Tyvärr är strukturfonderna inte mitt ansvar, men jag ska ta reda på av kommissionsledamot Johannes Hahn om det finns några rapporter från medlemsstaterna om resultatet av dessa bidrag, och i så fall ska ni förstås få veta det.
Angående: Skolresultat för elever i EU-medlemsstaterna
De nyligen offentliggjorda resultaten av den internationella undersökningen om 15-åriga skolelevers prestationer (Pisa-undersökningen 2009) visar att EU:s konkurrenskraft är allvarligt hotad eftersom endast två EU-länder hör till de tio bästa på området läsförmåga (nivåerna5-6).
Inom matematik var endast tre EU-länder bland de tio bästa och ingen av dem tillhörde de fem bästa.
År 2020 kommer både dessa ungdomar och de yngre eleverna att vara aktiva på arbetsmarknaden eller på väg att bli det och det är därför nödvändigt att vidta omedelbara och effektiva åtgärder i medlemsstaterna om vi vill förbättra kvaliteten på elevernas undervisning betydligt.
Kommer kommissionen att göra en grundlig utvärdering av ovanstående undersökning och lämna uttryckliga rekommendationer om förfaranden med bevisad effektivitet?
Finns det några planer för att sammanställa ett program för att sprida sådana beprövade och testade förfaranden eller inrätta ett forum för att diskutera utmaningarna som måste mötas?
Bör diskussioner föras med medlemsstaterna för att bestämma vilka åtgärder som behöver vidtas för att förbättra deras resultat?
Som ni vet bestämmer varje enskild medlemsstat hur det egna utbildningssystemet ska utformas.
Det överensstämmer med artikel 165 i fördraget om Europeiska unionens funktionssätt.
Trots det samarbetar kommissionen med medlemsstaterna för att främja ömsesidigt lärande och utbyte av god praxis.
Som vi anger i Europa 2020-strategin är det avgörande för EU:s framtid som ett kunskapsbaserat och integrerat samhälle att utbildningssystemen reformeras och moderniseras så att de ligger i nivå med de bästa i världen.
OECD:s PISA-undersökning är en viktig resurs för sådant utbyte.
Den senaste PISA-undersökningen, som offentliggjordes i december 2010, ger EU:s medlemsstater ett blandat intryck.
Det finns tecken som tyder på betydande förbättringar i vissa system, men som helhet återstår det mycket att göra.
Resultaten blir en viktig grund för de framtida diskussionerna mellan kommissionen och medlemsstaterna.
Den referensram för EU som antogs av rådet i maj 2009 syftar till att föra de grundläggande färdigheterna i läsning, matematik och naturvetenskap till en adekvat nivå genom att sänka andelen icke godkända femtonåringar till under 15 procent till år 2020.
Låt mig nu läsa upp något ur PISA-rapporten som är mycket viktigt.
Andelen elever som inte var godkända i läsning ökade från 21 procent 2000 till 24 procent 2006, men sjönk till 20 procent 2009.
OECD:s mål för 2010, att minska andelen från 20 till 17 procent år 2000, uppnåddes emellertid inte.
Andelen underkända elever i matematik och naturvetenskap har minskat sedan 2006.
Det gjordes större framsteg inom naturvetenskap än inom matematik och andelen underkända är i dag lägre inom naturvetenskap än inom matematik.
Med 2006 som utgångspunkt ligger EU bra till vad gäller framstegen mot målet 2020 för andelen underkända.
I genomsnitt, och för de tre discipliner i de 25 EU-staterna för vilka det finns uppgifter tillgängliga, var 22,5 procent underkända 2006.
År 2009 hade den andelen minskat till 19,6 procent Som vi kan se har alltså EU som helhet gjort vissa framsteg.
Kommissionen kommer naturligtvis att analysera PISA-resultaten och offentliggöra sina slutsatser i nästa årliga lägesrapport om referensramen, 2011.
I november 2010 uppmanade rådet kommissionen och medlemsstaterna att fokusera det gemensamma arbetet på följande områden: utformning av läroplaner, motivation till läsning, läs- och skrivfärdigheter, matematik, naturvetenskap och teknik, den nya teknikens påverkan på grundfärdigheterna och möjligheterna att utnyttja den för att hjälpa studenterna till självständighet och att hålla motivationen uppe, könsskillnader i prestanda och attityder, kopplingen mellan studenternas bakgrund och deras basfärdigheter och, slutligen, frågor som gäller lärare och lärarutbildare samt skolornas etik och egenskaper.
I sina slutsatser uppmanade rådet också kommissionen att inrätta en högnivågrupp om läs-och skrivfärdigheter och en temainriktad arbetsgrupp för matematik, naturvetenskap och teknik.
Jag tänker starta upp högnivågruppen om läs- och skrivfärdigheter den 1 februari.
Denna grupp ska föreslå politiska åtgärder som bygger på bästa praxis och forskning, vilket kommer att hjälpa medlemsstaterna att förbättra konsekvensen och effektiviteten när det gäller att tillhandahålla grundläggande färdigheter inom ramen för strategierna för livslångt lärande. Gruppen kommer att slutföra sitt arbete och offentliggöra sin rapport till halvårsskiftet 2012.
Den tematiska arbetsgruppen för matematik, naturvetenskap och teknik har dessutom redan inrättats.
Den består av nationella beslutsfattare och experter och arbetar utifrån ömsesidigt lärande och utbyte av bästa praxis.
Den temainriktade arbetsgruppen kommer att ange och sprida politiska åtgärder för att förbättra läget för personer med svaga grundläggande färdigheter på nationell nivå.
Jag vill också understryka att Comeniusåtgärderna för programmet för livslångt lärande bland annat prioriterar ökad motivation inom naturvetenskap och matematik och förbättrade läs- och skrivfärdigheter.
(LT) Herr talman! Jag vill fråga om det kanske har gjorts undersökningar i vissa länder som kan förklara studenternas svaga resultat och framsteg?
Handlar det om finansiering eller är det strukturbetingat?
Vad anser ni om primärutbildningen?
Forskning har genomförts på studenter i högre årsklasser, men hur är det med de yngre som har för avsikt att fortsätta sina studier?
Jag kan redovisa alla de uppgifter vi har om de olika medlemsstaterna. Vi har inte analyserat dem.
Det är inte vår uppgift att ta reda på varför vissa medlemsstater klarar sig sämre än andra, men under arbetets gång har vi utbytt exempel på bästa praxis.
Det gläder mig verkligen att kunna säga att vissa länder som har följt exemplen på bästa praxis har gjort väldigt goda framsteg sedan 2006 när det gäller de flesta av dessa indikatorer.
När det gäller grundskolans tidigare del har vi dessvärre inte några undersökningar liknande PISA.
Det finns ingen sådan undersökning.
Angående: Uppsplittring av de digitala marknaderna och konsekvenser för utbildningssystemet och investeringarna i geografiskt isolerade områden
Enligt kommissionens meddelande om en digital agenda för Europa är Europa alltjämt ett lapptäcke av nationella Internetmarknader, och européerna kan inte dra nytta av fördelarna med en digital inre marknad på grund av problem som faktiskt går att lösa, exempelvis bristande nätinvesteringar.
Detta får till resultat att utbildningen i många isolerade regioner (bergs- och öregioner) släpar efter tekniskt, och likaså påverkas investeringarna på flera håll.
Jag vill fråga kommissionen följande::
Informations- och kommunikationsteknik (IKT) står med sitt årliga marknadsvärde på 660 miljarder euro för 5 procent av EU:s BNP, och lämnar ett ännu mycket större bidrag till den totala produktivitetsökningen (20 procent direkt från IKT-sektorn och 30 procent från IKT-investeringar).
Är det på gång några gemensamma åtgärder för att ta tag i problemet med knappa nationella nätinvesteringar, särskilt i geografiskt isolerade regioner?
I kommissionens meddelande om Europa 2020 och i meddelandet om den digitala agendan för Europa angavs målet att alla EU:s medborgare ska ha tillgång till grundläggande bredbandstjänster senast 2013 och att alla medborgare ska få tillgång till betydligt högre Internethastigheter på över 30 megabyte per sekund till 2020, samt att minst 50 procent av alla EU:s hushåll ska ha Internetanslutningar på över 100 megabyte per sekund.
Kommissionen är medveten om att det utan ett kraftfullt offentligt ingripande finns risk för att bredbandstjänsterna inte introduceras optimalt, att de snabba, beprövade nätverken koncentreras till tättbebyggda områden och att isolerade landsbygdsområden släpar efter.
Det skulle dessutom få negativa effekter på utbildningssystemen och möjligheterna att integrera informations- och kommunikationsteknik i utbildningen.
Enligt färska uppgifter har bara 67 procent av skolorna i EU tillgång till bredband och det råder stora skillnader mellan olika medlemsstater och mellan tätt och glest befolkade områden, 73,7 respektive 60,6 procent.
För att undvika risken att introduktionen inte blir optimal har kommissionen antagit ett bredbandspaket som omfattar en gemensam ram för både den nationella och den regionala politiken, som bör utvecklas för att man ska kunna uppfylla målen.
Sådana politiska åtgärder bör framför allt sänka kostnaden för bredbandsutbyggnad inom hela EU:s territorium genom att garantera en god planering och samordning och genom att minska de administrativa bördorna.
Kommissionen har redan agerat för att öka investeringarna i avlägsna områden och regioner inom ramen för EU:s sammanhållningspolitik genom att avsätta cirka 2,3 miljarder euro för perioden 2007-2013.
Genom kommissionens meddelande om en ekonomisk återhämtningsplan för Europa blev det också möjligt att avsätta 360 miljoner euro till bredbandsinsatser för landsbygdsområden genom Europeiska jordbruksfonden för landsbygdsutveckling.
I programpaketet meddelade kommissionen att den kommer att förstärka och rationalisera finansieringen av höghastighetsbredband genom EU:s instrument till 2014 och undersöka hur man kan få fram kapital för bredbandsinvesteringar genom kreditförstärkningar som backas upp av Europeiska investeringsbanken (EIB) och EU:s fonder.
Ett förslag från kommissionen och EIB i frågan väntas under 2011.
En annan pelare i den digitala agendan gäller digitala färdigheter.
Här föreslår vi bland annat att man ska betrakta digitala kunskaper och kompetenser som ett prioriterat område för förordningen om Europeiska socialfonden under nästa programperiod och ange digital kompetens som ett komplement till Europass för att garantera insyn.
Som ni vet är utbildning helt avgörande för att utveckla digital kompetens i vårt samhälle och vi håller med om att vissa regioner kan komma att släpa efter utan lämpliga investeringar.
Enligt färska EU-data - de avser 2006 - hade bara 67 procent av skolorna tillgång till bredband, och det förelåg stora skillnader mellan olika medlemsstater och mellan tätt och glest befolkade områden.
Vi ska just påbörja en ny undersökning om skolorna och resultaten kommer att bli tillgängliga i slutet av året.
(EL) Jag vill tacka kommissionsledamoten, för ett mycket detaljerat svar.
Jag vill gärna lägga till följande fråga: I EU:s 2020-strategi anges att vårt mål är en digital inre marknad för hushåll och företag, vilket betyder lika möjligheter i fråga om tillträde, men det betyder också lika möjligheter i fråga om utveckling.
Du har själv sagt i samband med utfrågningar i de behöriga utskotten, till exempel utskottet för kultur och utbildning, att det kommer att behövas cirka 500 000 nya jobb inom de här sektorerna under de kommande fem åren.
Jag har en mycket specifik fråga: Vidtar vi alla de åtgärder som krävs för att se till att de här nya jobben fördelas rättvist, utan att man utesluter geografiskt avlägsna områden?
Herr talman! Svaret är ja.
Det låter väldigt bra.
Tack så hemskt mycket!
Angående: 116 000 - Hotline för saknade barn
Kommissionen har nyligen riktat en sista uppmaning till medlemsstaterna att så snart som möjligt aktivera EU:s hotline 116 000 för saknade barn.
Via detta telefonnummer skulle barn som befinner sig i utsatt läge kunna få den hjälp och det stöd som de behöver.
För närvarande är hotlinenumret 116 000 fullt funktionsdugligt endast i 12 medlemsstater.
Anser kommissionen att det faktum att denna service inte fungerar ordentligt i hela EU kan medföra att barn utsätts för risker?
Kommer människor att informeras om att denna service saknas i deras land eller i det land som de besöker?
Måste varje medlemsstat införa denna service i sin helhet på ett korrekt sätt?
Stämmer det inte att misslyckandet med att tillhandahålla en adekvat service i alla medlemsstater när det gäller detta nummer, kan utsätta barn för risker?
Herr talman! Kommissionen håller med Liam Aylward om att det krävs större insatser i många medlemsstater för att aktivera EU:s journummer 116 000 för saknade barn.
Enligt de reviderade telekomreglerna, och då tänker jag i första hand på artikel 27a i direktivet om samhällsomfattande tjänster, ska medlemsstaterna göra allt de kan för att se till att medborgarna har tillgång till tjänsten som driver ett journummer för att rapportera fall av saknade barn.
Kommissionen övervakar noggrant medlemsstaterna och hjälper dem att införliva den nya bestämmelsen i sin nationella lagstiftning, något som ska vara genomfört till den 25 maj 2011.
Den 17 november förra året antog kommissionen meddelandet ”Ring 116 000: det europeiska journumret för försvunna barn”.
Syftet med meddelandet är att förnya kommissionens uppmaning till medlemsstaterna att snarast aktivera EU:s journummer och att se till att tjänsten håller samma höga kvalitet i hela EU för att ge medlemsstaterna praktiskt stöd.
I meddelandet framhålls nuvarande bästa praxis i de olika medlemsstaterna för att ta itu med de viktigaste problemen i samband med driftskostnader och telekomkostnader för journumret 116 000.
Kommissionen tänker använda dessa exempel på bästa praxis till att utarbeta en uppsättning gemensamma miniminormer som kan garantera en tjänst av hög kvalitet inom hela EU, så att föräldrar och barn kan räkna med samma hjälp oavsett var de befinner sig.
Detta omfattande arbete går utöver de frågor som gäller elektronisk kommunikation och som jag har ansvaret för, och samordnas därför av min kollega Viviane Reding.
(EN) Fru kommissionsledamot! Tidigare har ni nämnt kostnader och bristen på information som hinder för att aktivera detta journummer i vissa medlemsstater.
Vilka åtgärder tänker ni vidta för att ta itu med dessa hinder och tänker ni er dessutom att denna tjänst ska aktiveras fullt ut i samtliga medlemsstater?
Slutligen undrar jag vilka alternativ som står till förfogande för de medlemsstater som har svårt att finansiera journumret, för att se till att det verkligen aktiveras i hela EU?
Självklart gör vi vad vi kan.
Den ärade ledamotens resonemang verkar förnuftigt.
Som jag nämnde tidigare är kostnaden en viktig fråga i sammanhanget.
Själva journumret är det minst problematiska i detta avseende.
Problemet är uppföljningen.
Den fråga vi bör fokusera på är inte bara själva journumret, utan uppföljningen.
Vi övervakar och stöder medlemsstaterna vad gäller aktiveringen, och vi är medvetna om att det är de som ska ta initiativet vad gäller den nationella lagstiftningen.
Vi är också medvetna om att det i samband med den nuvarande finansiella krisen är ännu svårare för medlemsstaterna att hitta resurser för att finansiera uppföljningen.
Några organisationer har erhållit EU-finansiering för vissa projekt.
Den tillgängliga EU-finansieringen är inte till för att täcka hela driftskostnaden för tjänsterna, utan syftar till att hjälpa till att utveckla 116 000-tjänsterna genom konkreta projekt.
Naturligtvis måste vi vara kreativa.
De som är engagerade i sådana här projekt och de nationella regeringarna bör också vara kreativa när det gäller att utnyttja budgetresurser, företagens sociala ansvar och privata donationer för att hitta resurser så att man till slut kan göra det som vi alla skulle vilja göra.
Angående: Alpin järnvägskorridor
Hur ser kommissionen på det nuvarande läget vad gäller bygget av Brennertunneln och det faktum att det krävs järnvägsanslutning till tunneln på båda sidor samt att järnvägssträckan München-Mühldorf-Freilassing-Salzburg måste byggas ut?
Herr talman! Frågan om trafiken genom alperna är extremt allvarlig, men läget ser ganska ljust ut för närvarande.
Trots en svår finansiell miljö gör man framsteg med Brennertunneln och dess norra och södra tillfarter.
Det här projektet har högsta prioritet och kommissionen beslutade att avsätta en budget på närmare en miljard euro för ändamålet.
För det första, när det gäller själva Brennertunneln nådde man viktiga framsteg under den österrikisk-italienska mellanstatliga kommissionens möte den 19 november 2010 i närvaro av EU:s samordnare Pat Cox.
Österrike och Italien skrev under ett avtal om den totala kostnaden för Brennertunneln på åtta miljarder euro.
Österrike godkände en optimerad arbetsplan som gör att förberedande arbeten för huvudtunneln kan påbörjas 2011.
Den italienska regeringen godkände att arbetena påbörjas genom ett åtagande som garanterar att kostnaderna är täckta under hela byggperioden.
För det andra kan jag rapportera om goda framsteg när det gäller tillfarterna på båda sidor.
Italien har godkänt att arbetet påbörjas på den södra tillfartsleden och att man börjar med den första sektionen, Fortezza-Ponte Gardena.
Österrike har också gjort goda framsteg vad gäller den norra tillfartsleden.
Österrike har ett avsnitt i nedre Inndalen som kommer att stå färdigt 2013, eller ännu tidigare.
När det slutligen gäller de gränsöverskridande förbindelserna mellan Österrike och Tyskland kommer man inte att kunna nå det ursprungliga målet att arbetet ska slutföras senast 2012.
På den tyska sidan kommer arbetet inte att påbörjas förrän 2012 och det kommer att ta cirka tre år.
I november 2010 offentliggjorde Tyskland emellertid sin nationella investeringsplan, som inkluderar avsättningar för positiv utveckling av den norra tillfartsleden mellan München och den österrikiska gränsen.
Sektionen med ett enda spår kommer att uppgraderas och hela avsnittet kommer att elektrifieras.
Nästa steg blir ett samförståndsavtal mellan Tyskland och Österrike om detta avsnitt och sedan måste planeringsprocessen för infrastrukturförvaltningen påbörjas.
(DE) Tack, Siim Kallas, för det vänliga svaret..
Men du besvarade inte den andra delen av frågan, där jag nämnde München-Mühldorf-Freilassing, som är en del av huvudlinjen från Paris till Budapest och som är särskilt viktig om man tänker på den bayerska kemiska triangeln och på att avlasta tillfartsleden till Brenner.
Om Brennertunneln genomförs kommer Rosenheim-sektionen att bli överbelastad och det blir då viktigt att utveckla München-Mühldorf-Freilassing-Salzburg, som också är ett projekt med högsta prioritet för kommissionen.
Jag måste fråga dig om du anser att det är möjligt att ställa ytterligare finansiering till förfogande för detta i nästa budgetplan. Det handlar trots allt om en gränsöverskridande fråga.
Det som händer i alperna är säkert bra, men på grund av detta memorandum gör den grekiska regeringen nedskärningar och minskar antalet tjänster, vilket isolerar Grekland från järnvägsnäten i Europa och på Balkan. Som skäl anger regeringen, på samma sätt som kommissionen, de grekiska järnvägarnas stora skulder.
Min fråga är därför följande: Vad anser du om denna utveckling, dvs. nedskärningarna i järnvägstjänsterna?
För det andra, omfattar de grekiska järnvägarnas skulder pengar för att medfinansiera infrastrukturarbeten tillsammans med EU?
När det gäller Grekland kan jag inte svara, eftersom jag inte känner till detaljerna.
Jag har inte fått någon information om de här problemen.
När det gäller det prioriterade projektet nummer 17, München-Mühldorf-Freilassing-Salzburg, så pågår det.
Det inledande arbetet påbörjades 2007.
En del av arbetet är avklarat.
Den 19 april 2010 påbörjades arbetet med den nya tvåspåriga järnvägsbron över floden i Mühldorf och det kommer att slutföras.
Denna bro finansieras helt av den tyska återhämtningsplanen.
Den kostar 11,7 miljoner euro, så det går framåt och vi anser inte att detta är ett viktigt problem i nuläget.
Angående: Att skicka sms samtidigt som man kör - trafiksäkerhet
En förare som skickar sms löper 23 gånger större risk att vara med om en olycka.
Sms:ande i samband med körning kräver årligen flera tusen dödsoffer i trafiken, och antalet personskador ökar i en oroväckande takt för varje år.
Trots att kommissionen erkänner behovet av att öka trafiksäkerheten och se till att trafiksäkerhetsreglerna genomförs finns det ingen EU-täckande lagstiftning som förbjuder användning av sms, e-post eller Internet vid körning av ett motorfordon över en viss, på förhand fastställd, hastighetsgräns.
Tekniken för att förhindra användning av sms, e-post och Internet samtidigt som man kör finns redan. Avser kommissionen att lägga fram någon EU-lagstiftning för att råda bot på denna livsfarliga vana?
Kommissionen håller med om att det är extremt farligt att skicka sms eller att ägna sig åt några andra ovidkommande aktiviteter samtidigt som man kör.
Under 2009 släppte kommissionen en rapport om användningen av mobiltelefoner samtidigt som man kör.
Den rapporten finns publicerad på Europa-webbsidan för trafiksäkerhet.
Vi har emellertid ingen statistik om antalet olyckor som beror på detta.
Samtliga medlemsstater har lagar som åtminstone indirekt förbjuder användning av sms, e-post och Internet samtidigt som man kör.
Även om man inte direkt nämner användningen av mobiltelefoner, så finns det krav i den nationella lagstiftningen på att förarna måste vara helt koncentrerade på sitt bilkörande.
Mot den bakgrunden tänker kommissionen inte införa ett ytterligare skikt av EU-lagstiftning för att förbjuda användning av sms, e-post och Internet vid körning av ett motorfordon.
Vi hoppas att medlemsstaterna ska ta hand om den här frågan på lämpligt sätt.
(GA) Herr talman! Jag är besviken på svaret jag fick från kommissionsledamot Siim Kallas.
Det är oerhört viktigt att de olika medlemsstaterna samarbetar.
Vi måste göra allt vi kan för att minska antalet dödsfall och allvarliga skador på vägarna.
Ett nytt fenomen på Europas vägar är att folk skickar sms samtidigt som de kör. Medlemsstaterna har olika regler.
Vi måste öka samarbetet.
Jag är besviken på att kommissionsledamoten inte kan lova oss mer i samband med detta.
(EN) Jag vill gratulera min kollega Jim Higgins till att ha tagit upp denna oerhört viktiga fråga.
Jag delar hans oro över den brist på entusiasm som kommissionsledamoten visade när det gäller att se till att bästa praxis tillämpas i hela EU.
Jag vill fråga honom varför kommissionen inte åtminstone kunde försöka uppmuntra medlemsstaterna till att införa samma regler i hela EU och se till att de följs för att främja säkerheten och skydda liv?
(ES) Herr talman! Jag har bara begärt ordet för att informera er, mina damer och herrar, om att jag är föredragande för frågan om gränsöverskridande påföljder, där rådet har fått möjlighet att öppna upp förteckningen över överträdelser - som faktiskt förekom i kommissionens inledande förslag - och där frågan om användningen av mobiltelefoner förekom.
Dessvärre deltar varken Storbritannien eller Irland i den förändring av rättslig grund som tillhandahålls genom rådets avtal eftersom de har valt att inte vara med.
Detta är ett av de problem vi har och som vi i parlamentet kanske kunde åtgärda.
Jag hoppas att de här länderna i diskussionerna med rådet ska förtydliga sina intressen, även om vi inte vet något om dem.
Det verkar som om Storbritannien nu tänker ansluta sig.
En bred handlingsplan för säkerheten och genomförandet av den planen har haft extremt hög prioritet för kommissionen, och vi har verkligen gjort enorma framsteg. Vi har kraftigt minskat antalet olyckor i Europa.
Jag kan berätta att dödstalet i mitt eget land var 400 i början av 1990-talet, medan det var nere på 78 förra året. Och detta naturligtvis med en tiofaldig ökning av antalet fordon på vägarna.
Det är en kraftig förändring.
Detta är viktigt, och tack så mycket Inés Ayala Sender för att du påminner oss om gränsöverskridande verkställighet av trafikpåföljder, vilket är ett extremt viktigt steg mot en bättre trafiksäkerhet.
Det beslutet togs av rådet i december och vi kommer nu att genomföra det.
Jag tror inte att ett ökat antal lagar på EU-nivå är något universalmedel. Att vi, oavsett problem, måste ha EU-lagstiftning.
Samtidigt som alla kritiserar att vi har för mycket EU-lagstiftning är detta, som jag ser det, emellertid en fråga där medlemsstaterna är lika oroliga som den europeiska allmänheten, och om gränsöverskridande verkställighet av trafikpåföljder kan skapa ett europeiskt område för trafiksäkerhet, så är detta mycket viktigt.
De frågor som på grund av tidsbrist inte hade besvarats skulle erhålla skriftliga svar (se bilagan).
Frågestunden är härmed avslutad.
(Sammanträdet avbröts kl. 20.15 och återupptogs kl. 21.00.)
Föredragningslista för nästa sammanträde: se protokollet
Avslutande av sammanträdet
Utsläppsnormer för nya lätta lastfordon (debatt)
Nästa punkt är ett betänkande av Martin Callanan, för utskottet för miljö, folkhälsa och livsmedelssäkerhet, om förslaget till Europaparlamentets och rådets förordning om utsläppsnormer för nya lätta nyttofordon som ett led i gemenskapens samordnade strategi för att minska koldioxidutsläppen från lätta fordon - C7-0271/2009 - 2009/0173 (COD)).
föredragande. - (EN) Herr talman! Det gläder mig att få inleda dagens debatt med betänkandet om utsläpp från lätta nyttofordon.
Innan jag går in på detaljerna i texten vill jag rikta några tackord till först och främst skuggföredragandena från alla politiska grupper, till föredragandena och ledamöterna i utskottet för transport och turism och utskottet för industrifrågor, forskning och energi för deras åsikter, och slutligen till kommissionsledamoten och hennes team - vi har haft ett antal mycket konstruktiva möten om detta.
Jag vill också tacka det belgiska ordförandeskapet för dess mycket hårda arbete under trepartsförhandlingarna och, slutligen, ett stort tack till Jos Vervloet och Isobel Findlay från miljöutskottets sekretariat, som har varit ett fantastiskt stöd under hela processen.
Jag har särskilt uppskattat Isobels hjälp i de komplexa frågorna kring kommittéförfarandet.
Vi har väntat på den lagstiftning som nu föreslås ända sedan liknande lagstiftning infördes för personbilar.
Personligen var jag inte helt övertygad om behovet av denna lagstiftning, eftersom de flesta lätta lastbilar köps av företag, både stora och små, som redan är mycket medvetna om behovet av ekonomiska och bränsleeffektiva fordon.
Jag har därför under hela processen framhållit betydelsen av att ha ett ambitiöst men realistiskt långsiktigt mål och ett lämpligt kortsiktigt mål som tar hänsyn till dels vad som krävs för industrins produktionscykel, dels behovet av miljöförbättringar.
Huvudfokus i vår debatt har hela tiden legat på det långsiktiga målet.
Kommissionens ursprungliga förslag till gränsvärde var 135 g CO2/km, vilket av många ansågs vara helt omöjligt att uppnå.
Utvecklings- och produktionscyklerna är längre för lätta nyttofordon än för personbilar.
Lätta nyttofordon används också, som namnet antyder, främst för nyttoändamål. Jämfört med personbilar finns det mycket lite utrymme att laborera med fordonens form och vikt för att minska utsläppen.
De huvudsakliga sätten att åstadkomma detta hos lätta nyttofordon är ändringar av fordonens motorer och mekanik - vilket tar betydligt längre tid och är betydligt kostsammare än att bara ändra karosseriet eller minska vikten.
Dessutom används redan dieselmotorer i de lätta nyttofordonen i betydligt högre utsträckning än i personbilar.
När kommissionen offentliggjorde sitt ursprungliga förslag klargjorde många av tillverkarna att de inte kunde gå lägre än 160 g CO2/km, en siffra som i sin tur framstod som alltför oambitiös för de flesta av oss i parlamentet.
I det paket som vi slutligen enats om, och som ligger framför er i dag, har vi en ganska rimlig kompromiss på 147 g CO2/km.
Med beaktande av de högre kostnaderna för att minska koldioxidutsläppen från lätta nyttofordon, jämfört med personbilar, och de längre utvecklings- och produktionscyklerna, anser jag personligen att detta ger en bra balans mellan strävan efter att förbättra miljönormerna och fastställandet av realistiska och genomförbara mål för fordonsindustrin.
Det faktum att vi på grund av denna kompromiss från ena hållet anklagas för att vara alltför eftergivna mot industrin, och från andra hållet får höra att vi är alltför miljömedvetna, tycker jag tyder på att vi faktiskt hittat den rätta balansen.
En avsnitt i kommissionens förslag som enligt alla grupper var ogenomförbart gällde den mycket komplicerade frågan om etappvis färdigbyggda fordon.
Det är självklart orättvist att straffa den som tillverkat grundfordonet när denne inte är ansvarig för vad som händer med fordonet i ett senare skede av produktionen.
I paketet som ni har framför er i dag finns ett mycket klokt förslag om att kommissionen ska se över frågan före årets slut. Här anges också grunderna för hur denna översyn bör gå till.
Jag anser att det paket som vi har förhandlat fram och som läggs fram för parlamentet i dag som ändringsförslag 58 är det bästa möjliga resultatet.
Jag gläder mig åt det stöd som jag förhoppningsvis har hos de flesta av de största politiska grupperna.
Det balanserar behovet av bättre miljönormer med realistiska och uppnåeliga mål som inte kommer att skada industrin eller utgöra en risk för arbetstillfällena i unionen.
Generellt är jag inte positiv till överenskommelser vid första behandlingen, utan anser att man helst ska undvika dem så långt möjligt.
I det här fallet bringar dock en överenskommelse vid första behandlingen klarhet och säkerhet till en sektor som fortfarande lider av den globala ekonomiska krisens efterverkningar, samtidigt som vi lägger ribban för hårda men rättvisa miljönormer som vi alla vill se.
Jag hoppas att kollegerna kommer att stödja paket tillsammans med mig i dag.
Herr talman! Jag vill först och främst gratulera föredraganden Martin Callanan och skuggföredragandena till deras ansträngningar för att nå en överenskommelse om kommissionens förslag om lätta nyttofordon.
Som Martin Callahan påpekat var dessa diskussioner verkligen svåra så här i efterdyningarna av den ekonomiska nedgången.
Jag vill inte sticka under stol med att det kompromisspaket som de interinstitutionella diskussionerna har resulterat i är mindre ambitiöst än kommissionens förslag på flera punkter.
De viktigaste av dessa är att uppfyllandet av det kortsiktiga målet skjuts upp med ett år, sanktionerna för överträdelser - ”avgifter för extra utsläpp” - sänks, och ambitionen för det långsiktiga målet minskas.
Det förvånar nog ingen att om jag säger att jag skulle ha föredragit ett mer ambitiöst resultat, och många av er delar säkert den uppfattningen.
Men den här kompromissen är ändå ett viktigt steg framåt.
Den innebär att vi fram till 2020 minskar de genomsnittliga koldioxidutsläppen från lätta nyttofordon från baslinjen 2007 på 203 gram koldioxid per kilometer till 147 gram per kilometer.
Det är en genomsnittlig minskning av utsläppen från de lätta nyttofordonen på 28 procent på 13 år.
Med tanke på att efterfrågan på lätta nyttofordon förväntas öka kommer ökad bränsleeffektivitet att vara en viktig faktor för att minska utsläppen från transporter.
Kompromissen kommer också att generera en nettobesparing under fordonets livstid på över 2 200 euro per fordon för konsumenterna, som främst är små och medelstora företag.
Dessutom kommer målen att stimulera innovation inom industrin och göra det möjligt för tillverkarna att utnyttja övergången till en koldioxidsnål ekonomi och därmed öka sin konkurrenskraft på lång sikt.
Kom ihåg att denna förordning bör ge tillverkarna ett försprång på världsmarknaden där liknande normer för koldioxidutsläpp sannolikt kommer att följa och efterfrågan på energieffektiva fordon förväntas öka.
Förordningen täpper dessutom till en stor lucka i lagstiftningen mellan personbilar och lätta lastbilar och minimerar därmed potentialen för snedvridande effekter av förordningen om koldioxidutsläpp från personbilar.
Man kommer inte att kunna kringgå koldioxidnormerna genom att registrera om stora bilar som lätta lastbilar.
Som ni alla vet släpper transportsektorn ut mer i dag än 1990, vilket i hög grad uppväger de minskningar som gjorts inom andra sektorer.
Detta är naturligtvis inte hållbart.
Transportsektorn måste i mycket högre omfattning bidra till EU:s övergripande koldioxidmål.
Denna förordning är ännu ett instrument som ska hjälpa medlemsstaterna att uppfylla sina åtaganden att fram till 2020 minska koldioxidutsläppen från de sektorer som inte omfattas av utsläppshandeln.
Jag ser denna överenskommelse som ännu ett bevis för Europeiska unionens beslutsamhet att uppnå klimatmålen och jag hoppas att ni kommer att ge ert stöd till kompromisspaketet vid omröstningen senare i dag.
Herr talman! Antagande vid första behandlingen bör vara ett undantag.
I detta fall var det möjligt eftersom vi på de mest kontroversiella punkterna kunde komma fram en kompromiss mellan kommissionens förslag och förslagen från utskottet för miljö, folkhälsa och livsmedelssäkerhet och utskottet för industrifrågor, forskning och energi.
Detta resultat kunde uppnås enbart tack vare att vi gick in i förhandlingarna med ett gemensamt förhandlingsmandat från alla grupper.
Jag vill särskilt tacka Martin Callanan för det engagemang han har visat.
Vi kan vara stolta över resultatet.
Det är på många områden identiskt med industriutskottets förslag.
Projektet vi nu har inlett är ambitiöst, men genomförbart för industrin och framför allt kommer det att ge användarna möjlighet att köpa prisvärda, moderna fordon med lägre koldioxidutsläpp.
Detta gäller särskilt små och medelstora företag, hantverkare, detaljhandlare och mikroföretag som använder denna typ av fordon.
(Talmannen avbröt talaren.)
Bland mina handlingar finns en punkt från industriutskottet som inte togs med, men som ändå antogs med knapp majoritet.
Det gäller förslaget om hastighetsbegränsare.
Detta blir nu en fråga för medlemsstaterna, som måste fastställa sina egna regler.
På det stora hela är vi därför nöjda med kompromissen.
Utskottet för industrifrågor, forskning och energi är berett att stödja hela paketet.
Herr talman! Det stämmer att transportsektorn är en av de sektorer där utsläppen måste minskas.
Vår brådska att minska utsläppen får dock inte undergräva konkurrenskraften hos EU:s biltillverkare.
Detta krav är särskilt angeläget med tanke på den rådande ekonomiska krisen, som redan har fått allvarliga konsekvenser för EU:s bilindustri.
Ur det perspektivet anser jag att målet 147 g CO2/km i genomsnittligt utsläpp från nya lätta nyttofordon är väl ambitiöst, och jag är mycket nyfiken på den genomförbarhetsstudie som kommissionen ska göra på grundval av de uppdaterade resultaten.
Samtidigt följer jag med stor uppmärksamhet de upprepade ansträngningarna från kommissionen och vissa andra parter, som verkar anse att det föreslagna målet tvärtom inte är tillräckligt ambitiöst, och som vill återuppta debatten kring denna fråga och försöka ändra förordningen för att fastställa strängare mål.
Jag anser att de ekonomiska aktörerna behöver garantier för att lagstiftningen inte kommer att ändras hela tiden.
Det är dags att ge biltillverkarna arbetsro och låta dem utveckla nya motorer så att de kan anpassa sig till reglerna och de nya målen.
I detta sammanhang bör vi också hålla ögonen på skäl 24, där man överväger möjligheten att utvidga användningen av hastighetsbegränsande anordningar till lätta nyttofordon.
Jag är glad över att denna fråga ska behandlas särskilt och att den debatten kommer att handla om affärsmässiga beslut och inte om ideologier.
Mina damer och herrar, vi måste hålla fast vid våra tider, eftersom vi har ett fullt program och omröstningen är klockan 12.
Herr talman! I dag företräder jag Anja Weisgerber, vår skuggföredragande för utskottet för miljö, folkhälsa och livsmedelssäkerhet, som är mammaledig.
Vi skickar henne våra varmaste lyckönskningar.
Hon har gjort ett utmärkt arbete med detta ärende.
På det stora hela är vi alla nöjda med kompromissen.
Den var inte lika svår att uppnå som i fallet med personbilar, eftersom nyttofordonen inte är en lika känslomässig fråga.
Ändå stod vi inför stora miljömässiga och ekonomiska utmaningar.
Ur ett klimatpolitiskt perspektiv är det viktigt att bördan fördelas jämnt längs alla länkar i kedjan, och även denna länk måste bidra med sin del.
Vi måste dock se till att inte slipa så mycket på länken att den riskerar att brytas.
Vad menar jag med det?
Kostnaderna för åtgärder av detta slag som berör små och medelstora företag innebär naturligtvis en betydande utmaning för dem.
Småföretagen kommer att fundera mycket noga över om det är värt att ersätta sina gamla fordon och investera i nya.
Därför var vi tvungna att fokusera mindre på de tekniska aspekterna och mer på de ekonomiska.
Om det bara gällt tekniken kunde vi ha uppnått mycket mer, men kostnaderna för detta hade definitivt överförts på de små och medelstora företagen och det hade inte gett det önskade resultatet.
Nu får vi vänta några år för att få reda på om den här förordningen är bra, det vill säga om vi verkligen lyckas uppnå de önskade utsläppsnivåerna.
Om förordningen bara att leder till att vi får driva in straffavgifter är inte målet nått.
Vi måste noga övervaka hur situationen utvecklas.
Herr talman, mina damer och herrar! Jag vill börja med att tacka för ett gott och konstruktivt samarbete.
Vi har uppnått en bra kompromiss, ur både miljömässigt och ekonomiskt perspektiv.
Även om vi enligt min mening kunde har gått längre när det gäller gränsvärdet, så är den lagstiftning som vi antar i dag fortfarande den strängaste i världen för lätta nyttofordon.
Det får vi inte glömma.
Som Connie Hedegaard påpekade är dessa särskilda rättsakter som vi inför för de mindre sektorer som ligger utanför utsläppshandeln mycket viktiga för att vi ska nå de mål vi har satt upp.
Fordon som drar mindre bränsle ger ett mervärde inte bara för klimatet utan också för luftkvaliteten.
Med en gräns på 147 g CO2/km, vilket motsvarar 5,6 liter diesel, kommer att fordonen att producera mindre luftföroreningar.
Det innebär att luftkvaliteten i våra städer kommer att förbättras.
Det är ett viktigt steg framåt vi tar i dag.
Min grupp röstar för detta kompromisspaket eftersom det innehåller en viktig punkt där det anges att vi senast 2014 måste utvärdera om de mål som vi antar i dag har uppfyllts eller överskridits och om vi behöver göra några justeringar på området.
Detta var ett grundläggande krav från vår grupp.
Jag har haft långa diskussioner med min kollega Mario Pirillo om kompromissen och detta var en av de grundläggande förutsättningarna för hela paketet.
Några har redan kommenterat den första behandlingen.
Vi bör i framtiden se till att vi antar färre texter i första behandlingen.
I det här fallet är det godtagbart, eftersom förhandlingarna i slutändan endast gällde två gram.
Det fanns inget behov av att ta det i andra behandlingen.
Men om parlamentet antar alla texter under första behandlingen berövar vi oss själva en del av våra rättigheter.
Jag vill också ta upp frågan om testcykeln.
Det kommer att bli mycket viktigt för oss att ha en standardiserad testcykel i framtiden som förhoppningsvis vid någon tidpunkt kommer att gälla i hela världen och som kommer att visa de verkliga värdena.
De nuvarande testcyklerna är inte realistiska och det krävs förbättringar på detta område.
Internationella förhandlingar pågår och jag hoppas att de kan slutföras med framgång, eftersom det skulle innebära att lagstiftningen kommer att återspegla den faktiska körcykeln.
Jag vill än en gång tacka alla berörda.
I dag är en bra dag för Europeiska unionens klimat- och miljöpolitik.
Herr talman! När det gäller huruvida det är klokt att nå en överenskommelse under första behandlingen bör vi inte hålla så hårt på våra principer som vissa ledamöter har rekommenderat.
Det bör alltid bero på ärendet.
Hur går diskussionerna?
Hur kontroversiellt är ämnet?
I fråga om regleringen av koldioxidutsläpp från lätta nyttofordon var det uppenbart att institutionernas ståndpunkter inte var särskilt långt ifrån varandra.
Därför skulle det inte ha varit mödan värt att inleda den andra behandlingen, utom möjligen i den fråga som är föremål för hetare diskussioner, det vill säga det långsiktiga målet.
Kommissionen har aldrig helt klargjort, och det framgår heller inte av konsekvensbedömningen, hur en minskning av utsläppen från dagens 203 gram till 135 gram inom 10 år - det är de siffror som nyss nämndes av Connie Hedegaard - ska kunna genomföras på ett ekonomiskt hållbart sätt.
Det motsvarar en nedskärning med 34 procent, något som går långt utöver våra andra klimatmål.
Parlamentets viktigaste uppgift var att göra detta mål mer realistiskt och genomförbart i ekonomiska termer.
Det är vad vi har gjort.
Jag är glad över att Matthias Groote tog upp mina argument, eftersom ett genomsnitt för hela fordonsflottan på 147 gram är långt ifrån vad kommissionen ursprungligen föreslog, men det är samtidigt det i särklass mest ambitiösa målet i världen.
Vi ska dock inte försöka inbilla oss att en gräns för koldioxidutsläpp från lätta nyttofordon kommer att rädda världens klimat.
Jag vill tacka alla, däribland föredragandena för deras hårda arbete.
Det gläder mig att vi har fått en stor majoritet för denna kompromiss.
för Verts/ALE-gruppen. - Herr talman! Tack föredragande Martin Callanan, du har varit väldigt professionell och inkluderande i genomförandet av förhandlingarna.
Däremot kommer jag inte att tacka för uppgörelsen.
Vi i Verts/ALE anser att kommissionens ursprungliga förslag var realistiskt och bra, men tyvärr är uppgörelsen alldeles för svag.
Den gör inte bilindustrins konkurrenskraft någon nytta, för var kommer man att sälja bilar år 2020?
Jo, det kommer man att göra i Asien, och där kommer man att efterfråga extremt energisnåla fordon.
Så vill vi gynna industrins konkurrenskraft bör vi fastställa mycket högre mål.
Uppgörelsen kommer inte heller att gynna miljön, för även om varje lastbil släpper ut 28 procent mindre så är det ingen som tror att trafiken inte kommer att öka fram till 2020.
Därmed kommer utsläppsmålen om en minskning på 30 procent, som vi antagligen kommer att uppnå genom förhandlingar i Durban i Sydafrika, inte heller att nås.
Dessutom tjänar inte ens ekonomin på det, eftersom ingen väl räknar med att bensinpriset 2020 kommer vara runt 13 kronor eller 1,30 euro per liter, utan det kommer givetvis att vara mycket högre.
Därmed var de kalkyler som låg till grund för kommissionens ursprungliga förslag mycket mer realistiska och till och med då låg de nästan för högt om man ska räkna ekonomiskt effektivt.
Så tyvärr vinner inte konkurrenskraften, ekonomin eller miljön på den här uppgörelsen.
Tvärtom tror jag att den naturliga tekniska utvecklingen faktiskt kommer att nå längre än den här uppgörelsen säger.
Det blir en sämre planeringshorisont för industrin, eftersom konsumenterna år 2020 med all säkerhet kommer att efterfråga bilar som drar högst 120 g CO2/km.
Det är också tråkigt att vi sänkte böterna för dem som inte uppnår målen.
Då kommer vi inte heller att uppnå lagstiftningens mål - om det nu inte blir som jag tror: att vi kommer att nå det här ändå med naturlig utveckling.
Det är samma sak med superkrediter: Det lurar oss att tro att utsläppen är mindre än vad de är om man räknar en elbil trippelt.
Så tyvärr vi kan inte stödja den här uppgörelsen, men jag vill ändå tacka alla inblandade.
Herr talman! Jag vill tacka för att du modererar den här debatten delvis på tjeckiska.
Främst vill jag dock tacka föredragandena och huvudföredraganden Martin Callanan för det arbete de har utfört.
Lagen som vi diskuterar är kopplad till den klimatpolitik som förs här i Europaparlamentet, och det här är inte rätt plats att kritisera den politiken och hela konceptet.
Vi måste inse att detta huvudsakligen handlar om ensidiga åtgärder från parlamentets sida, som inte har någon motsvarighet i resten av världen, utanför EU.
Vi måste överväga vad som skulle vara en bra motivation och vad som skulle vara en orimlig börda för EU:s företag, och jag är säker på att detta betänkande närmar sig en bra motivation.
I det avseendet håller jag verkligen inte med Carl Schlyter.
EU:s konkurrenskraft är inte och kommer inte att vara betjänt av att man hämmar EU:s industri.
Alla fakta pekar på att EU:s industri är på nedgång och flyttar utanför våra gränser.
Åtgärder på området för lätta nyttofordon är långt mer komplicerade än för personbilar, och lägger en mycket större börda på de små företagen, vilket redan har påpekats här.
Jag vill avsluta med att tacka alla föredragandena. Jag ser den uppnådda kompromissen som ett enastående arbete.
Herr talman, mina damer och herrar! Innan jag börjar diskutera lätta nyttofordon vill jag påminna om att EU:s biltillverkare har uppnått EU:s produktmål vad gäller koldioxidutsläpp från personbilar, flera år innan tidsfristen 2015, genom att vidta lämpliga tekniska åtgärder.
Det är nu uppenbart att tillverkarna allvarligt överdrev under förhandlingarna om tidsfristen och målen för åtgärderna för koldioxidutsläpp från personbilar, vilket ledde till att kraven urvattnades.
Tillverkarna använder samma strategi i sin lobbyverksamhet när det gäller målen för minskning av koldioxidutsläppen från lätta nyttofordon.
Jag undrar hur en majoritet här i parlamentet medvetet kan upprepa detta misstag och än en gång ge efter för bilindustrins krav.
Så här i klimatförändringens tid menar jag att det viktiga är att skydda miljön och trygga mänsklighetens framtid.
Om parlamentet åtminstone kunde stödja kommissionens förslag så skulle detta placera EU:s bilindustri i spetsen för den tekniska utvecklingen och därmed trygga dess konkurrenskraft.
Kommissionen har föreslagit ett mål på 135 g CO2/km.
Tack vare en övergångsperiod skulle tillverkarna inte ha varit tvungna att uppnå den gränsen förrän 2020.
Detta menar jag skulle ha varit möjligt.
I stället har en klen kompromiss tvingats fram under påtryckningar från rådet, bakom stängda dörrar, som innebär att biltillverkarna nu bara måste minska koldioxidutsläppen från lätta nyttofordon till 197 g CO2/km fram till 2020.
Denna svaga kompromiss är en gåva till industrin.
Superkrediter, övergångsperioder och poolning kommer att vattna ur den redan svaga gränssättningen ännu mer.
Tillverkarnas lobbyverksamhet bland ledamöterna här i parlamentet och påtryckningar i rådet från de fordonstillverkande länderna Tyskland, Frankrike och Italien har lett till detta dåliga resultat, som innehåller en mängd kryphål.
Betänkandet är oacceptabelt.
Det strider mot EU:s klimatmål och det kommer att bromsa upp den tekniska innovationen.
Gruppen Europeiska enade vänstern/Nordisk grön vänster kommer att rösta emot detta betänkande.
Herr talman! Min far är småföretagare.
Han har en elfirma och den enda anledningen till att han fick chansen att starta sitt företag var de skattelättnader och möjligheter som skapades av den konservativa premiärministern och sanna euroskeptikern Margaret Thatcher på 1980-talet.
Liksom alla småföretagare brottas han med byråkrati och reglering - varav en hel del kommer härifrån, från Europaparlamentet.
Min fars företag kommer att förbli litet.
Men det är den här typen av företag som är grundvalen för den brittiska ekonomin och de utgör svindlande 73 procent av alla företag i Storbritannien.
Min far kör en lätt lastbil, och som så många andra småföretagare får han kämpa på grund av lågkonjunkturen.
Jag är mycket orolig för att denna lagstiftning kommer att sätta småföretag som min fars i konkurs för alltid, eftersom vi fått veta att lagstiftningen kommer att medföra prishöjningar på lätta nyttofordon på upp till 5 000 euro.
Småföretagare har inte råd med denna kostnad nu när de kämpar med ekonomin.
Min kollega från den socialdemokratiska gruppen sade att detta är en bra dag för Europeiska unionens klimat- och miljöpolitik.
Men om detta går igenom kan jag garantera att det blir en dålig dag för småföretagare över hela kontinenten.
(Talaren godtog att besvara en fråga (blått kort) i enlighet med artikel 149.8 i arbetsordningen)
(EN) Herr talman! Varför kan inte du, Paul Nutall, förstå att den här åtgärden syftar till att förbättra bränsleeffektiviteten hos lätta nyttofordon?
Det innebär minskade kostnader för att köra dem, mil efter mil, i en tid då bränslepriserna är rekordhöga.
Detta hjälper företagen, det stjälper dem inte.
(EN) Herr talman! Än en gång visar parlamentet att man inte har en aning om vad som händer i den verkliga världen.
Människor kämpar där ute, och vad denna lagstiftning gör - och det har vi fått helt klart för oss - är att öka kostnaden för lätta lastbilar som körs av många småföretagare över hela kontinenten.
Priset kommer att öka med minst 5 000 euro.
Det är helt och hållet fel, och det är något som vi inte har råd med under en lågkonjunktur.
(EN) Herr talman! När jag lyssnar till diskussionerna om hur man ska kunna krama mer pengar ur småfolket med klimatförändringarna som förevändning, slås jag av två saker.
Den första är att ingen talar om global uppvärmning längre.
Även de mest världsfrånvända bland parlamentsledamöterna har fått klart för sig att avslöjandena av bedräglig pseudovetenskap och rekordkalla vintrar över hela världen har gjort allmänheten mycket skeptisk, och det med rätta, till all den falska propagandan om drunknande isbjörnar.
Det andra som slår mig är fordonsflottan på parkeringen nedanför oss - Porche, Mercedes, BMW, stadsjeepar - en parad av bensinslukande lyx som körs av de människor som ogillande pekar finger åt de många vita skåpbilarna och gör upp planer för att försvåra arbetslivet ytterligare med hastighetsbegränsare och straffavgifter, allt detta för en dogm baserad på kritiserad statistik som förts fram av en klick köpta akademiker, finansierad och höjd till skyarna av superrika med egna intressen i det gröna industriella komplexet - Al Gore, prins Charles, Shell och Goldman Sachs - som alla nu är i färd med att stjäla en förmögenhet ur de skatter som skördats genom subventioner till vindkraftverk och handel med utsläppsrätter.
Även om jag uppskattar de ansträngningar som vissa parlamentsledamöter gjort för att mildra de värsta överdrifterna i denna koldioxidhysteri, är den enkla sanningen den att alla som sätter någon tro till den genomskinliga bluffen om en global uppvärmning orsakad av människan är delaktig i historiens mest dödliga bedrägeri.
Ja, jag säger dödliga, för det handlar inte bara om att råna vanliga människor och avindustrialisera västvärlden, det handlar också om att hundratusentals av världens fattigaste barn just nu svälter ihjäl på grund av att livsmedelsgrödor ersätts av biobränsle som subventioneras av skattebetalarna.
Men det ökar vinsterna för Monsanto och det ger parlamentsledamöterna resor med alla utgifter betalda till oljepalmsplantagerna i Malaysia, så då måste det väl vara okej?
Nej, det är inte okej, särskilt som det avleder uppmärksamheten från den verkliga krisen - som inte gäller utsläpp av koldioxid från fossila bränslen, utan att vi börjar få slut på oljan som driver vår civilisation.
Varje dag som slösas på tal om att begränsa utsläppen av naturens viktigaste gödningsmedel är en förlorad dag i kampen för att försörja fler och fler människor med mindre och mindre energi.
Om det inte vore en sådan tragedi skulle det vara en fars.
(Talaren godtog att besvara en fråga (blått kort) i enlighet med artikel 149.8 i arbetsordningen)
(EN) Herr talman! Du har fel, Nick Griffin, när du säger att detta har varit en kall vinter över hela världen.
Det var faktiskt bara i vissa delar av norra Europa och vissa centrala delar av USA som det var kallt.
Globalt sett var 2010 ett av de två varmaste åren i historien.
Det faktum att det blir kallare här nu var också ganska förutsägbart, för om Golfströmmen trycks ned av smältvatten från Arktis, så är det en förklarlig effekt.
Så nej, 2010 var en mycket varmt år, klimatförändringen är verklig och de åtgärder vi vidtar är bra för ekonomin.
(EN) Herr talman! Jag vet inte om man här i kammaren noterade att gårdagens snöfall i Korea slog ett 100-årigt rekord, så det rör sig alltså inte om ett fåtal platser.
Precis som för två år sedan i Köpenhamn, när klimatkonferensen hölls där, var det kallare än på årtionden i Cancùn när klimatkonferensen hölls där.
För det andra finns det inga som helst bevis för att smältvatten från Arktis skulle hindra Golfströmmen.
Den har inte förändrats alls.
För det tredje skulle dina argument vara effektivare om datormodellerna för klimatförändringarna hade förutsett detta för ett par år sedan.
Det gjorde de inte.
För ett par år sedan fick vi höra att våra barn inte skulle veta vad snö var.
Det var verkligen rena rappakaljan.
När det slutligen gäller den statistik som påvisar global uppvärmning är faktiskt den viktigaste faktorn, som alla ignorerar, att 65 procent av världens väderstationer finns inom 10 meter från en artificiell värmekälla.
Praktiskt taget alla finns i städer.
Sovjetunionens sammanbrott har medfört att de flesta väderstationerna i naturligt kalla områden har lagts ned.
Det är detta som har snedvridit statistiken, som är en fundamental bluff skapad av människor som påhejade av FN letat efter tecken på en global uppvärmning orsakad av människor för att kunna införa de lösningar som de vill ha.
(FR) Herr talman, fru kommissionsledamot! Jag vill börja med att gratulera föredraganden till denna överenskommelse.
Som våra debatter visat har överenskommelsen varit svår att nå.
Jag tror att alla kan hålla med om vad som sagts.
Ja, klimatförändringarna existerar naturligtvis, men lätta nyttofordon är inte bilar som folk köper för att det är roligt att köra dem eller för att de är passionerat intresserade av dem.
Det är fordon som människor använder som ett arbetsredskap, vilket innebär att målet 147 g CO2/km år 2020 ger en bra balans.
Jag skulle ha föredragit en något högre gräns, men detta är åtminstone ett förslag som jag tycker är mer balanserat än kommissionens ursprungliga.
Det förslaget skulle ha lett till att tillverkarna påtvingades tekniska mål med tillhörande innovationskostnader som skulle fått stora ekonomiska konsekvenser för slutkonsumenterna som vi inte vill lägga mer börda på, eftersom de genomgår en exceptionell krisperiod.
Ändå välkomnar jag införandet av incitament för tillverkning av bränsleeffektivare fordon och straffavgifter för biltillverkare som inte uppfyller målen.
Allt detta är därför verkligen ett steg i rätt riktning.
Jag välkomnar också straffavgifterna.
Det är bra att vi har kunnat hitta en gemensam grund för straffavgifterna som är desamma som de som gäller för personbilar.
Därför röstar jag gärna för detta betänkande.
(IT) Herr talman, mina damer och herrar! För att klara övergången till en koldioxidsnål ekonomi och nå de mål som anges i klimatpaketet måste vi reglera koldioxidutsläppen inom olika sektorer, bland annat inom fordonsindustrin.
Jag är mycket nöjd med förhandlingarna som lett till en överenskommelse med rådet om att begränsa utsläppen till 147 g CO2/km fram till 2020.
Detta är en realistisk gräns som utgör en bra balans mellan miljömässiga, sociala och industriella regler.
Jag hoppas att jag också gjort min del i detta som skuggföredragande för utskottet för industrifrågor, forskning och energi.
Överenskommelsen tar hänsyn till den ekonomiska kris som sektorn genomgår och gör även rimliga eftergifter för skillnaderna mellan personbilssektorn och sektorn för lätta nyttofordon.
Precis som vi sett hända efter förordningen om personbilar, kommer EU:s bilindustrin att också lyckas med att utveckla grön, konkurrenskraftig och miljövänlig teknik för de lätta nyttofordonen.
Jag hoppas att även industrin kommer att kunna utnyttja den miljömässiga utmaningen och investera ännu mer i innovation och forskning.
(EN) Herr talman! Frågan är om vi kunde ha uppnått mer om denna åtgärd hade införts för att förbättra bränsleeffektiviteten hos nyttofordon snarare än att minska koldioxidutsläppen.
I praktiken är det naturligtvis samma sak, men det ena ses som en kostnad för företagen, och det andra ses som en besparing.
Paul Nuttall säger att åtgärden kommer att leda till prishöjningar på 5 000 euro per fordon.
Jag tror inte att åtgärden kommer att höja fordonspriset alls.
Låt oss ha denna debatt om tre år igen och se vem som får rätt.
Faktum är att oljepriset nu ligger på 100 US-dollar per fat.
Det är mer än vad kommissionen räknade med när den gjorde sin bedömning.
De potentiella besparingarna för företagen är större, och jag önskar att PPE-gruppen kunde erkänna detta.
PPE har uttalat sig på uppdrag av de stora tillverkningsföretagen, i stället för på uppdrag av alla de företag som använder lätta nyttofordon och som behöver mer bränsleeffektiv teknik för att kunna sänka kostnaderna.
Tillverkarna har gjort stora tekniska framsteg under de senaste åren.
Vi bör driva på den ambitionen.
Jag hoppas att kommissionen återkommer med en översyn om ett par år och ser till att dessa ambitioner får en reell chans att förverkligas.
(Talaren godtog att besvara en fråga (blått kort) i enlighet med artikel 149.8 i arbetsordningen)
(EN) Herr talman! Anser du verkligen, Chris Davies, att det är rätt att rösta för en lagstiftning som i praktiken kommer att leda till att kostnaderna för ett fordon ökar?
Både du och jag vet att det kommer bli så.
Det som detta kommer att leda till är att man sätter små företag i Liverpool och Manchester - i din egen valkrets - i konkurs.
Tycker du detta är rättvist?
Tycker du detta är moraliskt rätt?
Är du beredd att stå på denna plattform vid valet om tre år?
(EN) Herr talman! Den brittiska regeringen, närmare bestämt transportdepartementet, har faktiskt gjort en bedömning av effekterna av denna åtgärd.
Man fann att den sannolikt skulle bli mer fördelaktig för företagen än vad kommissionen hade uppskattat.
Nettobesparingen för att köra ett fordon, då bränslepriserna ligger på rekordnivåer, är större än den eventuella ökningen av kostnaden för fordonet - en nettobesparing för företagen och lägre priser för konsumenterna.
Detta är vad UK Independence Party är så fast beslutna att kämpa mot.
Därmed arbetar partiet för att få företagen att betala mer än de behöver.
(IT) Herr talman, mina damer och herrar! I förslaget fastställdes ursprungligen ett gränsvärde för utsläpp på 135 g CO2/km för lätta nyttofordon på lång sikt, dvs. detta skulle uppnås senast 2020.
Tillverkarnas enhälliga uppfattning var dock att det var tekniskt omöjligt att respektera denna gräns.
Om betänkandet hade godkänts som det var skulle koldioxidhalten på global nivå ha minskat med 0,00014 procent, att jämföra med den extremt stora ekonomiska effekten på mer än 45 miljarder euro bara för EU, vilket oundvikligen skulle ha lett till en genomsnittlig prisökning på omkring 3 800 euro per fordon.
Trots dessa problematiska frågor nåddes en överenskommelse med rådet vid första behandlingen som sätter gränsvärdena för utsläpp på 147 g CO2/km fram till 2020, med förbehåll för genomförbarheten, vilken måste bedömas av kommissionen före januari 2013.
Detta beslut är hur som helst enbart politiskt och har absolut ingenting att göra med de verkliga villkoren för industrin eller marknaden, eller konsumenternas intressen.
Vi kommer att rösta emot betänkandet, eftersom vi anser att de ekonomiska effekterna är för stora i förhållande till den obetydliga minskningen av koldioxidhalterna globalt.
(ES) Herr talman! Jag vill först gratulera föredraganden Martin Callanan, som har arbetat mycket hårt och, framför allt, fått ett bra resultat.
Det var inte alls lätt att nå en överenskommelse vid första behandlingen om en så här pass komplicerad förordning.
Bilindustrin är av avgörande betydelse i Europeiska unionen.
Det är dessutom en bransch som är engagerad i EU:s utsläppsminskningsmål och i teknisk innovation.
Den här överenskommelsen är en stabil ram som ger våra fordonstillverkare rättssäkerhet.
Jag anser att utsläppsmålen är både ambitiösa och realistiska.
Tillverkarna kommer att behöva minska utsläppen till 147 g CO2/km till 2020.
Jag är säker på att de kommer att lyckas, och därmed bidra till EU:s mål att minska utsläppen med 20 procent fram till 2020.
Men det finns också annat av intresse i den nya förordningen, som superkrediter och satsning på alternativa bränslen.
Biodrivmedel förespråkas tydligt i linje med EU:s mål för förnybara bränslen för 2020.
Jag framhåller detta uppenbara faktum, för om kommissionen fortsätter med sina tvekande förslag om biodrivmedel så kommer vi inte att uppnå målen för 2020.
Jag vill avsluta med att gratulera skuggföredraganden för Europeiska folkpartiets grupp (kristdemokrater), som just blivit mamma och som har arbetat mycket hårt och bidragit till att göra överenskommelsen till en framgång.
Herr talman! Jag vill börja med att tacka föredragande Martin Callanan, skuggföredraganden och alla andra som har varit inblandade i arbetet med detta direktiv.
Vi får nu äntligen en reglering av utsläppen också från lättare nyttofordon och det är viktigt.
Direktivet behöver nu införas så snart som möjligt.
Samtidigt nådde vi inte så långt som många av oss ville, och det tycker jag att vi ska tala ärligt och öppet om.
Vad vi ser är ett miljö- och industripolitiskt beslut som tydligt har påverkats av den ekonomiska krisen och av det faktum att så många europeiska regeringar, konservativa högerregeringar, har valt att möta denna ekonomiska kris med enbart nedskärningar och inga investeringar.
Detta resulterar i hög arbetslöshet och låg efterfrågan och påverkar både personbilsindustrin och industrin för lätta nyttofordon.
Visst kan man kalla det här för realism, men vad det handlar om är en påtvingad anpassning till den ekonomiska krisen och nedskärningspolitiken.
Kommissionen har alltså varit ambitiösare än till och med parlamentets miljöutskott, och det är inte vanligt.
Jag är tacksam för att det här beslutet ändå innehåller en översyn av utsläppsmålen år 2014.
Då hoppas jag att vi får en andra chans att visa att vi menar allvar med att konkurrenskraft och höga klimatpolitiska ambitioner inte står i konflikt med varandra, utan tvärtom kan hjälpa varandra framåt.
(FR) Herr talman, fru kommissionsledamot! Det är motvilligt som jag kommer att rösta för den slutliga kompromissen.
Förhandlingarna var förfärliga och enligt min mening är denna omröstning ett beslut som tvingats på oss genom ett maktspel inom parlamentet och rådet.
De största producentländerna har, med stöd av en majoritet av ledamöterna som är känsliga för branschens argument, lyckats hindra oss från att fastställa ett ambitiöst utsläppsminskningsmål.
Jag vill framhålla att kommissionen hade föreslagit ett mål på 135 g CO2/km till 2020.
Parlamentet visar alltså här mindre ambitioner än kommissionen, och det är beklagligt.
Bilindustrin, som har kämpat emot denna förordning - och det har vi just sett ytterligare exempel på - har uppenbarligen inte insett att den har allt att vinna på att gå i bräschen för utsläppsminskningen, särskilt eftersom en undersökning från Europeiska federationen för transport och miljö som gjordes i november förra året har visat att tekniska lösningar finns.
Undersökningen visade att EU:s biltillverkare har minskat koldioxidutsläppen från personbilar med 2-10 procent under 2009, och att en japansk tillverkare så gott som nått sitt mål sex år i förtid.
Jag kommer att rösta för kompromissen eftersom vi annars riskerar att förstöra denna bedrift, hur liten den än må vara, i en andra behandling.
Jag vill dock understryka att vi gör tillverkarna en björntjänst genom att försvara status quo och att de berörda statliga myndigheterna underlåter att fullgöra sitt uppdrag genom att inte uppmuntra innovation.
(IT) Herr talman, mina damer och herrar! Vi har uppnåt ett mycket ambitiöst resultat.
Koldioxidutsläppen från dessa fordon ligger för närvarande på 200 g per kvadratkilometer.
Att minska detta till 147 g sänker därför tröskeln med över 25 procent.
Jag vill dessutom betona att marginella minskningar är de dyraste och vi bör därför vara försiktiga.
Jag anser också att denna särskilda kategori av fordon inte kan jämföras med personbilar vilket ofta har hänt här i kammaren.
Produktionscyklerna är mycket längre och det skulle bara ha en 1,5-procentig inverkan på koldioxidutsläppen inom hela transportsektorn.
Om vi inte fastställer vårt centrala mål kommer det att leda till att vi bestraffar en sektor som redan har lidit av en abrupt minskning på över 30 procent, något som framför allt har skadat små och medelstora företag, och alla vi här i kammaren bekräftade för bara 12 timmar sedan att vi ville stödja dessa företag, på grund av den viktiga ekonomiska och sociala roll de spelar som det enda verkliga redskapet för sysselsättning i Europa.
Vi måste därför vara mycket noggranna.
Jag välkomnar det arbete som har utförts, men vi behöver definitivt övervaka det hela noggrant.
(NL) Herr talman! Den text vi har framför oss är verkligen en kompromiss och vi skulle ha önskat att vi hade varit lite mer ambitiösa här och där, särskilt när det gäller val av tidpunkt och nivån på straffen.
Å andra sidan är det viktigt att utsläppsnormer fastställs för denna kategori av fordon - något som tycks ha slunkit igenom nätet lite, med tanke på att det redan finns ett antal regler för både person- och lastbilar.
Utvecklingen går i rätt riktning, men som ni själv sade har antalet nyttofordon ökat enormt de senaste åren och det ser ut som om de kommer att fortsätta att öka under kommande år.
Som ledamot i utskottet för transport och turism skulle jag kort vilja återkomma till hastighetsbegräsningarna.
Vi har i utskottet föreslagit att hastighetsbegränsningen ska fastställas till 120 km i timmen från 2018, vilket verkligen inte är orimligt.
Som ni vet finns det redan en gräns för lastbilar och jag tror att det skulle vara klokt att lagstifta om detta, både av miljö- och av trafiksäkerhetsskäl.
Jag tror det måste ske på europeisk nivå eftersom det inte är så mycket mening med att överlämna detta till medlemsstaterna.
Fru kommissionsledamot! Jag skulle vilja uppmana dig att ta upp frågan igen med din kollega Siim Kallas - han är här i kammaren med oss - studera den och lägga fram ett förslag.
Jag tror att det skulle vara positivt för era respektive ansvarsområden: miljön och trafiksäkerheten.
(DE) Herr talman, kommissionsledamot Hedegaard, mina damer och herrar! Vi är inte här i dag för att diskutera klimatet.
Vi behöver bara göra det som är möjligt.
Jag välkomnar den kompromiss som har uppnåtts.
Genom att begränsa utsläppen till 147 gram per kilometer från 2020 fastställer vi mycket tydliga normer.
Det kommer att skapa incitament för att utveckla ny teknik som kan öka energieffektiviteten och bekämpa klimatförändringarna.
Fordonsanvändarna kommer också att ha nytta av dessa innovationer som kommer att spara bränsle och därmed pengar.
Små transportbilar används huvudsakligen av handelsidkare, små och medelstora företag, jordbrukare och vinodlare.
De körs vanligtvis endast korta sträckor och används ofta i många år, till dess att företaget lämnas över till nästa ägare.
Kostnaden för dessa fordon måste därför vara hanterliga.
Högre investeringskostnader måste finansieras på grundval av energieffektivitet och energibesparingar.
Det långsiktiga målet med 2020 ger oss tillräckligt med tid för övergångsperioder så att forskningsorganisationer och industrin kan utveckla och tillverka nya motorer.
Det mål vi har satt upp är realistiskt, nåbart och fortfarande effektivt.
Jag hoppas att det får ett brett stöd.
(PL) Herr talman! Alla inom vägtransportsektorn, både tillverkare av personbilar och tillverkare av lätta nyttofordon, bör bidra till att begränsa de totala koldioxidutsläppen.
Jag välkomnar därför den kompromiss som utarbetats av Europaparlamentet, rådet och kommissionen, där det fastställs gränser för utsläpp och straff om dessa gränser inte respekteras.
Att fastställa obligatoriska och ambitiösa gränser som också är realistiska kommer att innebära en utmaning för den europeiska bilindustrins möjligheter till innovation.
Den kommer att fungera som ett incitament för att öka forsknings- och utvecklingssatsningar som syftar till att finna nya designlösningar som kan användas för att tillverka mer miljövänliga fordon.
Vi måste ha våra egna gröna tekniker så att vi kan undvika att importera fordon, vilket har varit fallet med hybridtekniken.
Jag anser att de lagstiftningsbeslut vi har fattat kommer att fungera som en lämplig stimulans för att mobilisera europeiska tillverkare som kommer att inse att grön teknik utgör ett tillfälle till utveckling.
(FR) Herr talman!
Jag skulle vilja börja med att gratulera föredraganden till hans ståndpunkt och jag noterar att parlamentet trängts in mellan en kommission som är mycket ambitiös och ett råd som, precis som vanligt, är försiktigt mellan klimatskeptiker och klimatkritiker och mellan dem som stöder industrin och miljövänner.
Detta är därför en balanserad ståndpunkt som förblir ambitiös eftersom målet på 147 gram år 2020 ger branschen tid att åstadkomma det tekniska språnget och samtidigt uppmuntrar den att verkligen bli effektiv.
Förlängningen av ändringsperioden till 2018 är positiv och kommer att göra forskning inom, och tillverkning av, icke miljöförstörande bilar attraktivare.
Jag har avslutningsvis två kommentarer.
Jag välkomnar självfallet att förslaget har godkänts vid den första behandlingen och jag förstod inte fullt ut kommentarerna från vår kollega nyss när han sade att han föredrog en andra behandling.
För det andra beklagar jag, i likhet med Saïd El Khadraoui, avsaknaden av anordningar för hastighetsbegränsning, eftersom det innebär att vi kommer att fortsätta att bli omkörda på motorvägen av de enda fordon som ännu inte håller hastighetsbegränsningarna, nämligen lätta nyttofordon.
(RO) Herr talman! Den här förordningen innebär ett framsteg när det gäller att successivt uppnå målen att minska koldioxidutsläppen från lätta nyttofordon i Europa.
Det blir möjligt genom att det skapas incitamentsystem som gör bilarna effektivare och genom att det införs straff för tillverkare som inte uppfyller dessa mål.
Jag tror emellertid inte att den nya lagstiftningen om minskning av koldioxidutsläppen kommer att äventyra situationen för vare sig biltillverkare eller kunder.
De nya bestämmelserna måste ta hänsyn till oron bland små och medelstora och europeiska biltillverkare som begär att det successiva införandet av utsläppsgränser ska inledas efter 2015, eftersom de bilar som ska säljas under 2014 redan befinner sig på utvecklings- och produktionsstadiet.
Siffran 147 gram är en acceptabel kompromiss jämfört med de siffror som har nämnts.
Kommissionen måste emellertid noga övervaka förhållandet mellan bilindustrin och användarna för att bedöma hur åtgärden påverkar priserna och därmed verksamheten för små företag.
(PL) Herr talman! Tillverkningen av lätta nyttofordon och tillhörande tekniska frågor kräver mycket stora investeringar och en långsiktigare strategisk plan och tillverkningscykel än vad som gäller för passagerarfordon.
Att godkänna ett sådant långsiktigt mål var grundläggande för att garantera industrin tillverkningssäkerhet.
Å andra sidan bör vi inte bortse från den gräns på 147 g som ska uppnås senast 2020.
Det inledande kortfristiga målet, dvs. gränsen på 175 g, som infördes i syfte att uppnå målet på 147 g senast 2020, kommer att avsevärt öka kostnaden för att tillverka lätta nyttofordon, vilket gör dem dyrare för många små företag som använder dem i sitt dagliga arbete.
Jag hoppas att detta inte leder till en påtaglig nedgång i försäljningen av nya fordon, vilket i sin tur skulle innebära att tekniskt äldre fordon som orsakar mycket högre utsläppsnivåer skulle finnas kvar längre på vägarna.
(IT) Herr talman, fru kommissionsledamot, mina damer och herrar! Den kompromiss som uppnåtts med rådet förefaller definitivt mer balanserad och realistisk än kommissionens ursprungliga förslag som var så ambitiöst att det föreföll delvis utopiskt, eftersom det inte tog vederbörlig hänsyn till industrins villkor och inverkan på marknaden.
Alltför mycket ideologiskt miljökämpande innebär alltid en riske för att sannolikheten för nåbara resultat minskar, och leder till att miljön skadas.
Enligt min uppfattning kan det, trots att det långsiktiga målet på 147 g koldioxid/km senast 2020 ännu inte är optimalt, visa sig vara mer rimligt och realistiskt än det som ursprungligen föreslogs.
Jag välkomnar även de planerade incitamenten för ekologiska innovationer men enligt min uppfattning återstår en kritisk fråga: beslutet om utsläpp från så kallade färdigbyggda fordon, det vill säga de som byggs i flera steg.
Jag hoppas att kommissionen respekterar sitt åtagande att lämna ett specifikt lagstiftningsförslag om detta före årets slut.
(RO) Herr talman! Jag välkomnar det utmärkta arbete som föredraganden Martin Callanan och min kollega Matthias Groote har utfört genom detta betänkande.
Bestämmelsen kommer att tvinga tillverkare att utveckla ny grön teknik och även om detta till synes innebär en ny börda för dem kan det öka bilindustrins konkurrenskraft på den globala marknaden.
Samtidigt kommer det att bidra till att uppfylla åtagandena när det gäller minskning av koldioxidutsläppen, i linje med EU:s strategi.
Kompromissändringsförslagen ger tillverkarna tillräckligt med tid för att förbereda genomförandet av ny teknik, och kommissionen får tid att utveckla ett effektivt system för att övervaka överträdelser av bestämmelserna på området.
(PT) Herr talman! Hanteringen av innovation, med andra ord forskning och utveckling av ny teknik och nya produktionsprocesser, deras genomförande i stor skala och valet av lämplig tidpunkt för att genomföra dem, bör som sina vägledande kriterier först och främst ha skyddet av det allmänna intresset, förbättring av livskvalitet för allmänheten och skyddet av miljön.
Dessa principer, snarare än smala kommersiella intressen hos industri och företag, bör i första hand styra ansträngningarna i riktning mot innovation och hanteringen av deras genomförande.
Detta gäller även utsläpp från fordon.
Med tanke på att transportsektorn står för en avsevärd andel av koldioxidutsläppen bör en lämplig del av ansträngningarna för att minska dessa vara inriktade på detta område.
Det är därför viktigt att fortsätta att förbättra fordonens energieffektivitet, minska bränsleförbrukningen och rent allmänt utveckla teknik för låga koldioxidutsläpp.
Detta har nu blivit möjligt genom vetenskaplig och teknisk utveckling som tar hänsyn till den successiva och ofrånkomliga bristen på fossila bränslen redan från första början, något som redan är mycket viktigt att ta hänsyn till.
(FR) Herr talman, fru kommissionsledamot! Jag ska fatta mig kort.
Jag kommer att rösta för den här texten eftersom jag anser att kompromissen är ett steg i rätt riktning.
Samtidigt beklagar jag att den inte har gått så långt som förslaget från Connie Hedegaard.
Jag skulle därför nu vilja att ni berättade för oss, efter debatten och före omröstningen om några timmar, vad det förfarande som ni kommer att anta för de närmaste två åren består av, eftersom det ska göras en översyn 2013, vilket gör det möjligt för oss att utan dröjsmål, såsom vår grupps föredragande Matthias Groote ville, driva kampen vidare för att minska utsläppen från dessa lätta nyttofordon.
Det är min fråga till dig, Connie Hedegaard, och jag vet att du kommer att vara orubblig så att vi kan göra framsteg trots branschens lobbyverksamhet, som jag, i likhet med ett antal av mina kolleger som har talat i ärendet, anser är olämplig.
(DE) Herr talman, kommissionsledamot Hedegaard! Jag kan inte dölja att jag är en av dem som mycket hellre skulle ha antagit ett mål på 135 gram i dag.
Jag anser emellertid att den här kompromissen återspeglar verkligheten och visar att vi är beredda att göra en allvarlig gemensam ansträngning för att begränsa och minska koldioxidutsläppen.
EU har nyligen lyckats minska de totala kolidioxidutsläppen med 9 procent.
Utsläppen inom transportsektorn har däremot ökat med närmare 30 procent.
Enbart ur detta perspektiv anser jag att det steg vi i dag tar är ytterligare ett i rätt riktning.
Vi bör emellertid inte tillåta oss att distraheras av att de verkliga problemen inom transportsektorn ligger någon annanstans, med tanke på den totala ökningen på 29 procent.
Vi behöver med andra ord starkt fokusera på att utveckla kollektivtrafiken.
Vi får inte öka bördorna för de små och medelstora företagen utan ska i stället underlätta för pendlare och skynda på järnvägsbyggandet.
Vi kommer att uppnå mycket mer genom att gå från individuella transporter till kollektiva.
Jag anser att vi tar det första steget i rätt riktning eftersom vi när allt kommer omkring talar om en minskning på 25 procent.
(NL) Herr talman! Jag vill gratulera samtliga men jag skulle ha velat se ett mer ambitiöst resultat.
Mycket mer ambitiöst.
Och varför?
Jag ska ge er fem skäl: Mer innovation, större konkurrenskraft för Europa, miljön, självfallet, eftersom detta kunde ha bidragit till att vi sparar råvaror, och det skulle också ha varit billigare för konsumenten.
I Europa är vi starkt beroende av import av råvaror för energi.
Med renare teknik skulle vi ha gjort många fler besparingar och vi skulle också ha gett en enorm impuls till vår starka bilindustri att ta fram ren, intelligent teknik som skulle kunna säljas var som helst i övriga världen och som kunde ha gett oss ett försprång.
Det skulle ha varit billigare och effektivare, just för att vi är så beroende av import.
Det skulle också ha resulterat i besparingar för konsumenten.
Inköpspriset kanske hade varit högre, men det skulle till slut ha blivit billigare per kilometer.
Det skulle framför allt ha varit av stort intresse för små och medelstora företag.
För nederländarna är uttrycket ”ta hand om dina cent så kommer euron att ta hand som sig själv” fortfarande mycket intressant!
(ES) Herr talman! Jag skulle också vilja tacka föredragandena och särskilt vår skuggföredragande, Matthias Groote, för ett förslag som kommer att uppmuntra vår industri att bli grönare.
Jag tycker dock att det är högst beklagligt att vi har förlorat ett gyllene tillfälle att införa hastighetsbegränsare som är avgörande för att bidra till att förbättra luftkvaliteten.
Jag vill påpeka att direktivet redan har varit obligatoriskt i över en och en halv månad, vilket har märkts i städer som Barcelona, där den socialistiska ledningen har satt hastighetsgränsen till 80 km i timmen. Det är skillnad mot andra städer såsom Madrid eller Valencia som har konservativa ledningar, och där befolkningen löper stor risk att drabbas av allergier och andningssjukdomar.
Hastighetsbegränsare skulle ha hjälpt oss att minska dessa problem, och även att förbättra vägsäkerheten och minska antalet omkomna.
Det är därför beklagligt och vi hoppas att vi kommer att kunna uppnå detta i framtida lagstiftning.
Herr talman! Först en kort kommentar till Gilles Pargneaux som undrade vilka planerna var för de närmaste åren.
För det första måste naturligtvis kommissionen, precis som vi har kommit överens om, bedöma de framsteg som gjorts och förvissa sig om att saker och ting är genomförbara.
Det är vad vi alla har kommit överens om, men vi har självfallet skäl att anta att det är genomförbart eftersom vår konsekvensanalys redan har visat detta.
Vi är medvetna om kostnaden och konsekvenserna av det vi gör, och den nivå vi väljer att införa.
Vi tror därför att det kommer att bli genomförbart, men vi tittar självfallet på allt detta.
Jag skulle bara vilja säga att om vi inleder debatten på nytt om målet för 2020 kan det leda till osäkerhet i planeringen så vi bör därför nu naturligtvis betona att ett långsiktigt mål har fastställts.
Många tillverkare uppskattar detta eftersom det ger dem den långsiktiga planering och den förutsägbarhet som de verkligen behöver.
När allt kommer omkring uppskattar de det.
Det var också ett svar till Oldřich Vlasák och hans oro.
Bara en kort kommentar till Paul Nuttall - jag vet inte om han fortfarande är här - eller snarare till hans far eftersom han absolut inte behöver oroa sig över något, med undantag för att hans son använder siffror från en källa som jag inte är bekant med.
Faktum är att kostnaden för detta är mycket lägre än vad Paul Nuttall påstår och man sparar mer pengar i form av bränslekostnader än vad själva kostnaden är.
Så när allt kommer omkring kommer inte Paul Nuttalls far att endast spara pengar - han kommer att göra en nettovinst.
Han kan också förklara att hans barn och barnbarn kommer att få renare luft.
Det vi försöker göra här är att öka innovationen inom en mycket viktig industrisektor för Europa.
Det är vad vi försöker göra.
Jag ska avsluta debatten med att bara säga att vi har fördelen att ha skaffat oss bred erfarenhet av lagstiftning när det gäller bilar.
I samtliga fall visade det sig att tillverkarna kunde uppfylla lagstiftningen snabbare och till lägre kostnader än de påstått.
Jag skulle inte bli förvånad om samma sak händer med dessa transportbilar.
Regler för personbilar finns nu.
Nu är det dags för transportbilar.
Jag uppskattar det mycket breda stöd som denna lagstiftning fått.
Nästa sak vi behöver titta på inom detta område blir tunga nyttofordon och där ser jag självfallet fram emot att samarbeta med Europaparlamentet.
Herr talman! Låt mig kort besvara flera av de kommentarer som framförts här.
Carl Schlyter sade att han ansåg att det var dåligt för europeisk industri och att det skulle leda till att fler lätta nyttofordon tillverkas i Asien.
Jag måste säga att jag helt enkelt inte förstår den kommentaren.
Vi fastställer de ojämförligt mest utmanande målen i världen, mycket strängare än reglerna i staterna eller någonting som finns i Kina eller Fjärran östern.
Sabine Wils jämförde förordningen med förordningen för personbilar.
Jag tycker att det är en felaktig jämförelse.
Möjligheterna att minska utsläppen från personbilar är mycket större på grund av lägre vikt och byte av bränslemix.
Dieseln är redan mycket vanligare på marknaden för transportbilar.
Transportbilar är naturligtvis mycket mer ett nyttofordon och köps av affärskunder.
Jag är rädd att Paul Nuttall inte är kvar till slutet på den här debatten, men han har fel i de siffror som han har lämnat.
Det kommer att leda till totala kostnadsbesparingar för många företag.
Jag måste säga att jag skulle ha lite mer respekt för kommentarerna han lämnade om EFD-koncernen verkligen hade brytt sig om att sända en enda företrädare till något av våra trepartsmöten eller till något av våra skuggmöten för att framföra att de gillar att tala för småföretagens räkning.
(Applåder)
Sammanfattningsvis tycker jag detta är ett bra resultat.
Det ger den bästa balansen för det första beträffande företagens kostnader, men även när det gäller miljöförbättringar.
Oavsett vilken uppfattning man har om klimatförändringarna måste bränsleeffektivitet - att använda dyrbara resurser effektivare - vara en god sak.
Debatten är avslutad.
Omröstningen kommer att äga rum vid middagstid i dag (15 februari 2011).
Skriftliga förklaringar (Artikel 149)
Överenskommelsen med rådet är resultatet av tuffa förhandlingar ansikte mot ansikte med intensiv lobbying från branschen.
Genom hela förfarandet har vi stått emot tillverkarnas massiva påtryckningar för att försvaga förordningen och framför allt sänka ambitionen med de långsiktiga målen för att minska koldioxidutsläppen.
Det var ett svårt dilemma eftersom många av oss har bilindustrier som redan har det kämpigt på grund av den ekonomiska situationen.
Men vi visste av erfarenheterna från förordningen om personbilar att bilindustrin har gjort enorma framsteg när det gäller innovation och utveckling av renare teknik eftersom lagstiftningsramen uppmuntrade dem i rätt riktning.
Vi ville upprepa denna framgång med lagstiftning för transportbilar - inte bara av miljöskäl, utan för att större bränsleeffektivitet i slutändan kommer att minska kostnaderna för många företag.
Vi har en kompromisstext som, även om den inte är lika ambitiös som vi skulle ha velat, kommer att leda till en betydande minskning av koldioxidutsläppen från transportbilar och bidra till EU:s ambitioner att minska utsläppen till 2020 och därefter.
Jag vill gratulera föredraganden och skuggföredragandena till deras framgångsrika förhandlingar med rådet.
Vägtransportsektorn är den näst största källan till utsläpp av växthusgaser i EU och utsläppen fortsätter att öka.
Alla typer av fordon, inbegripet lätta nyttofordon, bör därför omfattas av förordningar som syftar till att minska dessa utsläpp.
Målsättningen att minska utsläppen av växthusgaser kommer att uppnås lättare om det finns en lagstiftning som täcker hela EU, snarare än nationell lagstiftning med olika målsättningar.
Vi behöver därför kombinera ambition med realism och förnuft.
Med tanke på att små och medelstora företag sannolikt är de som mest använder lätta nyttofordon och att dessa står för 99,8 procent av företagen och 67,4 procent av arbetstillfällena i EU bör vi därför inte ha mål som kan äventyra dem.
Jag instämmer därför i målet med 147 g koldioxidutsläpp per kilometer för nya lätta nyttofordon i EU om det är bekräftat att detta är genomförbart.
Jag välkomnar också det faktum att en gemensam hastighetsgräns för denna typ av fordon inte har införts på EU-nivå.
Jag välkomnar denna åtgärd och det är mycket viktigt att en balans upprätthålls mellan skydd av miljön och skydd av arbetstillfällen och små och medelstora företags konkurrenskraft i EU.
1.
Avtalet EG/Sydafrika om handel, utveckling och samarbete (
1.
Medielagen i Ungern (
- Före omröstningen:
Herr talman! Innan den planerade omröstningen om resolutionen om medielagen i Ungern vill jag uppmärksamma mina ledamotskolleger om den senaste utvecklingen av situationen och lägga fram ett konkret förslag.
För fyra dagar sedan antog Ungerns parlament de ändringar - alla ändringar - som kommissionen krävde trots att ledamöter från Ungerns socialistiska parti och gröna parti röstade nej.
Kommissionsledamot Neelie Kroes deltog vid omröstningen, och hon meddelade att den ändrade versionen av lagen följde europeisk lagstiftning och i synnerhet stadgan om de grundläggande rättigheterna.
Ändå ignoreras dessa fakta helt i vänstergruppernas resolution som vi ska rösta om vid lunchtid idag.
Texten är i princip samma som för tre veckor sedan, och inget nämns om omröstningen i det ungerska parlamentet.
Min fråga är denna: lever detta parlament i verkligheten eller i en låtsasvärld?
Är denna resolution riktad mot den ungerska regeringen, eller mot Europeiska kommissionen, som inte längre har några invändningar mot lagen?
(Applåder)
Jag vill framför allt fråga ordföranden för den liberala gruppen: har du eller har du inte förtroende för kommissionsledamot Neelie Kroes?
Europeiska folkpartiets grupp (kristdemokrater) anser att parlamentet förlorar sin trovärdighet om den antar texter som inte motsvarar verkligheten.
Måste vi bli en arena för att samla nationella politiska poäng?
(Applåder)
Mot bakgrund av detta drar PPE-gruppen tillbaka sin egen resolution och uppmanar övriga grupper att göra samma sak.
Parlamentets trovärdighet står på spel.
Mina damer och herrar! Förslaget är helt tydligt.
Som jag förstår det har Europeiska folkpartiets grupp (kristdemokrater) dragit tillbaka sin resolution.
Vi har därför endast en resolution, som har ingivits av flera av de politiska grupperna.
Jag vill be företrädarna för de politiska grupperna att kommentera detta.
Herr talman, mina damer och herrar! Joseph Daul talade om verklighet.
Verkligheten är att den ungerska regeringen eller det ungerska parlamentet har ändrat lagen, och det är bra, för jag kommer ihåg den debatt i denna kammare där vissa personer - inklusive du själv, herr Daul - sade att inget behövde ändras utan att allt var bra.
Nu måste det plötsligt ändras.
(Applåder från vänster)
Men det är också verklighet - och även detta kan man läsa - att både OSSE:s representant för mediefrihet och företrädaren från Europarådet säger att ändringarna är bristfälliga.
Det är verkligheten, herr Daul.
Det är verkligheten.
(Applåder från vänster)
Vid vår grupps sammanträde igår, där jag var ordförande, diskuterade vi lagen och ändringarna. Precis som OSSE och Europarådet kom vi fram till att ändringarna är bristfälliga.
Vilket beslut som än tas idag, om du vinner, herr Daul, eller om vi vinner, så kommer vi inte att ge upp kampen för mediefrihet, herr Lange.
Om du gör så är det din sak.
(Applåder från vänster)
Mediefrihet är ett oantastligt element i en demokrati.
Vi vill ha demokrati och vi vill ha mediefrihet.
Vi ber er därför att rösta därefter idag.
Vi vet att det även finns vissa ledamöter i er grupp som håller med oss.
Vi måste kämpa för mediefrihet, både i Ungern och på andra ställen.
(Applåder från vänster)
Mina damer och herrar, ledamotskolleger! Som jag förstår det drar de fyra politiska grupperna inte tillbaka sin förklaring.
Vi skulle kunna avsluta debatten här och gå vidare till omröstningen, men om jag förstår rätt så vill även Gruppen Alliansen liberaler och demokrater för Europa i Europaparlamentet göra ett uttalande.
Varsågod.
Herr talman! Man vände sig specifikt till oss här.
Naturligtvis har vi förtroende för kommissionsledamot Neelie Kroes arbete.
Hennes utredning av sekundärlagstiftningen var exemplarisk.
Vi önskar att kommissionsledamoten som utredde primärlagstiftningen hade gjort sitt jobb på samma sätt, eftersom det är där problemet ligger.
(Applåder från vänster)
I verkligheten omfattar situationen de saker som Hannes Swoboda just nämnt, nämligen att både Europarådet och OSSE anser att ändringarna är bristfälliga.
Ungerns vice premiär- och justitieminister Tibor Navracsics har själv erkänt att detta inte var någon betydande ändring av medielagen.
Jag kan nämna skyddet för journalistiska källor, som ännu inte är reglerat, eller mediemyndighetens sammansättning och makt.
Alla dessa frågor kvarstår att diskutera.
Jag vill därför, på Gruppen Alliansen liberaler och demokrater för Europas vägnar, meddela att vi inte kommer att dra tillbaka resolutionsförslaget utan istället kräva att omröstningen äger rum.
Mina damer och herrar! Vi ska nu rösta om de fyra politiska gruppernas resolution.
Muntliga frågor och skriftliga förklaringar (ingivande): se protokollet
Datum för nästa sammanträdesperiod: se protokollet
7.
Statsstödda exportkrediter (
för GUE/NGL-gruppen. - (EN) Herr talman! Jag vill meddela att GUE/NGL-gruppen vill stryka omröstningen med namnupprop om båda delarna av ändringsförslag 10.
Liksom vid den förra omröstningen har de skuggföredragande och jag själv beslutat att inte låta lagstiftningsresolutionen gå till omröstning i parlamentet. Vi fortsätter förhandlingarna med rådet i hopp om att man tar hänsyn till parlamentets omröstning i dag.
2.
Ansvarsfrihet 2009: EU:s allmänna budget, Europeiska ombudsmannen (
1.
Ansvarsfrihet för 2009: EU:s allmänna budget, Avsnitt III, Kommissionen (
Interinstitutionellt avtal om ett gemensamt öppenhetsregister - Ändring av arbetsordningen efter upprättandet av ett gemensamt öppenhetsregister
Nästa punkt är en gemensam debatt om
betänkandet av Carlo Casini, för utskottet för konstitutionella frågor, om ingående av ett interinstitutionellt avtal mellan parlamentet och kommissionen om ett gemensamt öppenhetsregister, och
betänkandet av Carlo Casini, för utskottet för konstitutionella frågor, om att ändra Europaparlamentets arbetsordning till följd av inrättandet av ett gemensamt öppenhetsregister för Europaparlamentet och kommissionen.
föredragande. - (IT) Fru talman, fru minister, herr kommissionsledamot, mina damer och herrar! Jag kommer att behandla båda betänkandena i mitt inlägg eftersom de handlar om samma fråga.
I och med den här debatten och den efterföljande omröstningen kommer vi att avsluta arbetet och förhandlingarna i den arbetsgrupp som leddes av Diana Wallis och bestod av kolleger från samtliga politiska grupper samt en kommissionsdelegation ledd av Maroš Šefčovič, och som har lett till att vi har kunnat utarbeta ett avtal om inrättande av ett gemensamt öppenhetsregister.
Utskottet för konstitutionella frågor har utarbetat detta betänkande på bara några månader och har också slutfört betänkandet om ändringen av parlamentets arbetsordning.
Personligen blev jag väldigt förvånad över den offentliga uppmärksamhet som detta öppenhetsavtal har fått.
Jag är rädd för att folk tror att resultaten kommer att ha större effekt än vad som faktiskt var meningen.
Insyn och öppenhet är en garanti för att de rätta politiska åtgärderna vidtas, men är inte rätt instrument för att komma åt korruptionen.
Händelserna nyligen där journalister har försökt korrumpera några parlamentsledamöter kan ske även utanför parlamentet.
Dessutom skulle de som eventuellt skulle låta sig korrumperas veta hur de kan undvika att bli identifierade och registren är därför ingen garanti.
Det rätta verktyget för den uppgiften är straffrätten.
Men om medlemsstaternas straffrätt inte räcker till måste vi se över artiklarna 82-86 i Lissabonfördraget, överväga om korruption av Europaparlamentsledamöter kan anses vara ett gränsöverskridande brott eller en handling som på annat sätt skadar unionens finansiella intressen, och bestämma oss för om vi bör inrätta en europeisk offentlig åklagare eller ej, vilket dessutom skulle vara ett stort steg på vägen mot enighet.
Öppenhetsregistret har en mer blygsam uppgift.
I en del länder har begreppet lobbyist en negativ mening, medan lobbyverksamhet i andra länder närmast ses som en offentlig tjänst eftersom lobbyisterna informerar beslutsfattarna om frågor som de kanske inte skulle känna till annars.
Detta är särskilt viktigt för Europaparlamentet, eftersom de frågor som ledamöterna arbetar med ofta är mycket komplexa och tekniska och vi nästan alltid måste finna en lämplig avvägning mellan företag och länder med olika intressen.
Det är här lobbyisterna gör stor nytta.
Vi bör alltså inte kalla dem lobbyister längre, utan intressenter.
Det kan naturligtvis finnas motstridiga intressen, och det är helt i sin ordning.
Jag har arbetat som domare och jag kan säga att korsförhör av motsatta sidor anses vara ett villkor för att få fram sanningen och skapa rättvisa.
Därför är det bra att vi har lobbyister eller intressenter med motstridiga intressen: det viktiga för en domare - och därmed även för Europaparlamentets ledamöter i det här fallet - är att man behåller sin tankefrihet, sitt oberoende och ärligt söker efter sanningen.
Därför har vi inrättat öppenhetsregistret i en ömsesidig överenskommelse mellan parlamentet och kommissionen med förhoppningen om att rådet snart kommer att ansluta sig till avtalet.
De som vill företräda sina intressen har fritt tillträde till våra lokaler, men de måste vara inskrivna i registret, där alla upplysningar som behövs för att identifiera deras rättsliga och finansiella status kommer att registreras.
Registret är offentligt.
Det finns även organisationer som inte har själviska intressen, utan som vill samarbeta i utformningen av EU-politiken på grund av allmänna värderingar, som kyrkor, politiska partier och regioner.
De behöver inte skrivas in i registret, men om de har separata kontor som uteslutande har uppgiften att hålla kontakt med EU-institutionerna måste de skrivas in i registret. De omfattas dock av ett annat rättsligt system än intressenterna.
Såsom redan har angetts innebär det nya registret även en ändring av arbetsordningen.
Därför har två betänkanden utarbetats, men detta är hur som helst bara ett första steg mot fullständig insyn.
Vissa hypoteser har redan utforskats och kan omvandlas till regler efter ytterligare övervägande. I punkt 9 i betänkandet om ingående av avtalet anges därför möjligheten att registret ska omfatta uppgifter om de lobbyister som har beviljats ett möte med en berörd ledamot angående en viss rättsakt.
Det lämnas stort utrymme för möjliga ändringsförslag, vilket gör att jag måste uttrycka en negativ åsikt om ändringsförslag som skulle innebära en begränsning av sådana framtida överläggningar.
Jag hoppas dock att rådet kommer att ansluta sig till avtalet inom kort och att vi också når ett omedelbart och brett samförstånd här i parlamentet, vilket skulle utgöra ett starkt budskap när det gäller insynskravet och även en uppmaning att agera.
Jag hoppas att omröstningsresultatet blir närmast enhälligt.
rådets ordförande. - (HU) Fru talman, herr kommissionsledamot, mina damer och herrar! Insyn och öppenhet är en särskilt viktig princip för demokratiska institutioner.
Detta gäller särskilt EU-institutionerna eftersom de - och det är allmänt känt - ofta anklagas för att inte låta människorna vara delaktiga och för att verka i det fördolda.
Rådet vill garantera största möjliga insyn och öppenhet mellan EU:s institutioner och organ.
Rådet är också medvetet om att medborgarna förväntar sig att de personer som de har utsett att styra dem arbetar efter strängast möjliga normer, och därför välkomnar vi Europaparlamentets och rådets initiativ att inrätta ett öppenhetsregister.
Jag välkomnar särskilt Carlo Casinis betänkanden.
Om parlamentet antar dem kommer det att bli möjligt att inrätta öppenhetsregistret under de närmaste månaderna, på grundval av betänkandena.
På så sätt kan vi återigen visa att EU är engagerat i insyn och öppenhet, inte bara i ord, utan även i handling.
Jag vill passa på att betona att jag är medveten om att rådet har inbjudits att delta i öppenhetsregistret.
Rådet tänker för närvarande inte delta fullt ut i processen eftersom rådet, till skillnad från parlamentet och kommissionen, till sin karaktär inte påverkas av intressenters verksamhet.
Dessa personer och organisationer kontaktar i allmänhet inte rådet som institution, utan inriktar sitt arbete på medlemsstaterna.
Men jag har redan sagt att rådet är berett att delta i registret och följa den här verksamheten.
Vi är också beredda att diskutera aspekter av rådets eventuella roll i detta med parlamentet och kommissionen, naturligtvis utan att fördröja ikraftträdandet av avtalet mellan de två institutionerna.
På grundval av rådets beslut nyligen överväger vi nu möjligheten att utfärda en politisk förklaring så att registret kan inrättas i juni.
kommissionens vice ordförande. - (EN) Fru talman! Insyn och öppenhet är en fråga som både intresserar och oroar medborgarna och det är viktigt att öka EU:s demokratiska legitimitet.
Jag är mycket glad över att kunna informera er om att vi redan i dag har över 3 800 poster i kommissionens register.
Därför är jag fullständigt övertygad om att införandet av ett gemensamt öppenhetsregister kommer att utgöra ytterligare ett stort steg framåt i arbetet med att öka insynen i EU:s beslutsprocess och direkt bemöta medborgarnas oro i det här sammanhanget.
Jag vill berömma det mycket konstruktiva arbete som vår gemensamma arbetsgrupp har utfört.
I det sammanhanget vill jag även berömma Diana Wallis, vår talman för i dag, vår föredragande Carlos Casini, och även Jo Leinen och Isabelle Durant.
Det var en fantastisk grupp och det var ett verkligt nöje att arbeta med er.
Resultatet av vårt arbete är ett mycket välavvägt och praktiskt utkast till interinstitutionellt avtal, som vi lägger fram för parlamentet för behandling och debatt i dag.
Om det blir ett positivt omröstningsresultat i morgon kommer våra två institutioner att gemensamt kunna inrätta registret i juni.
Detta kommer helt klart att sända en stark politisk signal som bekräftar att vi är fast beslutna att arbeta på ett öppet och etiskt sätt på EU-nivå.
Syftet med registret är att öka insynen för medborgarna när det gäller organisationer och egenanställda personer som är engagerade i EU:s politiska arbete eller försöker påverka EU:s beslutsprocess.
Jag har förstått att det har uppstått en viss oro över regionala offentliga organ, så det är bäst att jag klargör det.
Frågan var om de ska registrera sig.
Om vi läser texten noggrant inser vi att ett registreringskrav inte skulle avspegla deras verkliga identitet och inte heller avspegla att de representerar sina medborgare direkt enligt respektive författningssystem.
Vid en noggrann genomläsning av avtalsinnehållet framgår det dock att det finns fullständiga garantier i det här avseendet.
Faktum är att det uttryckligen anges i texten att lokala, regionala och kommunala myndigheter inte behöver registrera sig.
Detta synsätt förstärks även genom bilaga I, där det anges att offentliga myndigheter inte behöver registrera sig.
Lokala, regionala och kommunala myndigheter, inbegripet de representationer som ingår i förvaltningen av dessa och som har institutionella eller konstitutionella arbetsuppgifter behöver inte heller registrera sig.
Jag hoppas att detta klargör de frågetecken som jag har märkt av under de senaste dagarna.
Några sista ord om den interinstitutionella dimensionen.
Jag tror att vi alla är överens om att det gemensamma samarbetet mellan kommissionen och parlamentet skulle förstärkas ytterligare om rådet också deltog.
Därför är jag mycket glad över och tackar varmt det ungerska ordförandeskapet för att det har lyckats ändra ståndpunkten i rådet och för att det har skapat en positiv anda och inställning när det gäller att se hur vi bäst kan organisera förbindelserna mellan rådet, kommissionen och parlamentet i driften av registret. Det är nämligen en mycket viktig politisk signal att våra tre institutioner tar den här frågan på så stort allvar och att vi kommer att hantera insynsfrågan tillsammans.
Med ett sådant starkt politiskt stöd från samtliga tre institutioner är jag säker på att vi mycket snart kommer att nå gränsen 4 000 registreringar.
för PPE-gruppen. - (DE) Fru talman, fru minister, herr kommissionsledamot! Insyn och öppenhet är en hörnsten i demokratin, som garanterar att man vet vem som utövar inflytande och hur besluten fattas.
Sedan Lissabonfördragets ikraftträdande har Europaparlamentet fått avsevärt utökade befogenheter.
Därför är det också helt rätt att våra arbetsmetoder alltid ska vara öppna för diskussion och att vi även bör ifrågasätta det vi själva gör.
Förhandlingarna mellan Europaparlamentet och kommissionen om öppenhetsregistret har varit en framgång och vi har nått ett utmärkt resultat.
Jag vill återigen understryka att det är bra att vi har lyckats utforma tydliga regler för lokala och regionala myndigheter, och även för kyrkor, som avspeglar deras intressen.
Jag vill också påpeka att vi inte ser lobbyverksamhet som något negativt i sig.
Vi behöver expertåsikter och vi måste kunna anlita experter för vårt arbete.
Det viktiga är ju trots allt att vi, som parlamentariker, fritt kan överväga frågor och fatta oberoende beslut.
Jag anser att vi parlamentariker har mycket att vara stolta över.
Om vi gör en nationell jämförelse ser vi att endast ett fåtal EU-medlemsstater har inrättat öppenhetsregister på denna nivå.
I Berlin, huvudstaden i mitt land, där jag också råkar bo, finns inget öppenhetsregister och vi bör alltså vara medvetna om att detta är ett verkligt viktigt steg framåt.
Till rådet vill jag säga att om den här frågan inte är ett problem för dem eftersom lobbyisterna har mycket lite inflytande i rådet, borde det i så fall betyda att det är ännu lättare för dem att ansluta sig till öppenhetsregistret.
Rådet bör därför kunna övervinna det interna motståndet.
Avslutningsvis vill jag påpeka att om vi i parlamentet vill slippa undan lobbyisternas inflytande mer i framtiden kommer vi att behöva ytterligare stödresurser och mer personal, så att vi kan åstadkomma mer för EU-medborgarna.
för S&D-gruppen. - (DE) Fru talman, mina damer och herrar! För det första vill jag tacka föredraganden och alla som har arbetat med den här frågan eftersom en lång tid av hårt arbete äntligen kommer att avslutas efter morgondagens omröstning.
Det är en bra dag för EU, för Europaparlamentet som institution och för kommissionen, eftersom vi har lyckats inrätta ett gemensamt öppenhetsregister.
Det är ett viktigt steg på vägen, men vi behöver göra mer.
Jag vill ta upp två punkter.
För det första är registret egentligen inte obligatoriskt.
Det måste klargöras i det här läget.
Jag har en fråga till kommissionen om detta: kommissionen har alltid hävdat att det inte finns någon lämplig rättslig ram för detta.
Är kommissionen beredd att inrätta en sådan rättslig ram, så att vi får ett obligatoriskt register efter översynen?
Det var glädjande att höra rådets uttalande om att det inte ser några svårigheter med att ansluta sig till vårt register, som Manfred Weber nyss påpekade.
Jag hoppas att rådet kommer att följa upp detta, eftersom registret faktiskt bara kan bli fullständigt om samtliga tre EU-institutioner har ett gemensamt och även obligatoriskt register.
Vår grupp är för det ändringsförslag som lagts fram av en av de andra grupperna med ett krav på att de pengar som läggs på lobbyverksamhet även ska anges i öppenhetsregistret, och vi kommer att stödja det ändringsförslaget.
När det gäller de olika nationella lobbygrupperna har det klargjorts att de inte kommer att tas med i registret.
Jag vill tacka alla mina kolleger för deras kompromissvilja i den här frågan.
Det skulle verkligen ha varit en plump i avtalet om nationella lobbygrupper ska behandlas på samma sätt som branschlobbyister eller andra yrkesorganisationer.
Fru talman! Den senaste tidens skandaler har verkligen visat vilken makt lobbyister kan ha över parlamentet, så den liberala gruppen välkomnar varmt rationaliseringen av lobbyistregistret, som effektivt skapar ett öppet och direkt system som ska medföra ökad insyn och förbättrade samrådsprocesser.
Jag välkomnar särskilt punkt 9 i betänkandet, där presidiet uppmanas att inrätta ett system med vägledande förteckningar varigenom föredragandena kan registrera de lobbyister som har bidragit under utarbetandet av en rättsakt.
Det är en känslig fråga, men jag anser att det skulle vara ett ytterligare steg framåt för att öka parlamentets folkliga legitimitet och kvaliteten på vårt lagstiftningsarbete.
Systemet blir först fullständigt när rådet - som är den andra kammaren i vår lagstiftande församling - ansluter sig, men jag välkomnar de trevande stegen framåt och tackar ordförandeskapet för dess uttalande här i eftermiddag.
(Talaren godtog att besvara en fråga (blått kort) i enlighet med artikel 149.8 i arbetsordningen.)
(DE) Fru talman! Jag vill tacka Andrew Duff för att han tar upp frågan om vägledande förteckningar.
Anser du att de vägledande förteckningarna, vars räckvidd inte har fastställts ännu, kan leda till att Europaparlamentets arbete begränsas?
En annan fråga: hur stor inverkan tror du att de vägledande förteckningarna kommer att få?
(EN) Fru talman! Jag anser att de vägledande förteckningarna bör vara ett experiment.
Precis som med alla experiment skulle användningen spridas om det slår väl ut.
Jag anser dock att detta bör begränsas till föredragande som är ansvariga för att utarbeta ett förslag till en rättsakt för parlamentets räkning.
De bör offentliggöra namnen på de personer som de har haft offentliga sammanträffanden med under arbetets gång.
Dessutom anser jag att detta skulle uppmuntra en intelligent och välgrundad lobbyverksamhet i parlamentet.
Vi vet alla att vi är beroende av branschspecialister och experter för att utarbeta förslag av hög kvalitet.
Fru talman! Jag vill börja med att tacka Carlo Casini för hans arbete med detta interinstitutionella avtal.
Ledamöterna av utskottet för konstitutionella frågor och kommissionen har gjort ett bra arbete och tagit fram ett meningsfullt och praktiskt inriktat betänkande som kommer att leda till ökad insyn och öppenhet i lagstiftningsprocessen.
Fru talman, det är bra att det är du som har ordförandeskapet i dag eftersom jag vill tacka dig för dina insatser i förhandlingarna mellan parlamentet och kommissionen.
Betänkandet är proportionellt och användbart och jag är övertygad om att det kommer att göra nytta.
Man bekräftar den viktiga roll som regionala och lokala myndigheter spelar i utformningen av EU-lagstiftningen, och gör därför en tydlig åtskillnad mellan lobbyister och lokala och regionala myndighetstjänstemän.
Även om betänkandet är ett steg i rätt riktning återstår fortfarande arbete att göra.
Jag hoppas att öppenhetsregistret - om det faller väl ut - kommer att utvecklas till ett obligatoriskt register för lobbyister.
Jag instämmer i Andrew Duffs förslag om att föredragandena bör ange namnen på de lobbyister som de har haft kontakt med under utarbetandet av en rättsakt.
Det råder inget tvivel om att våra väljare ser på oss parlamentsledamöter med en viss misstänksamhet.
Ju mer insyn och öppenhet desto bättre.
Med tanke på detta vill jag bara påpeka att ett problem med det här avtalet är att det saknas en institution.
Det är en besvikelse att rådet inte har anslutit sig.
Som medlagstiftare bör medlemsstaterna enas och ansluta sig till registret så vi får en verkligt öppen lagstiftningsprocess.
för Verts/ALE-gruppen. - (DE) Fru talman, mina damer och herrar! Politik bygger på förtroende.
Parlamentets ledamöter har valts i ett fritt och hemligt val av medborgarna i våra medlemsstater, som med all rätt förväntar sig att vi respekterar deras intressen, det vill säga det allmänna bästa, i allt vi säger och gör och att vi inte agerar i eget intresse eller tredje parters intresse, vare sig de är företag eller andra intressegrupper.
Men vi är också medvetna om att vi till exempel i Bryssel är omgivna av över 10 000 yrkeslobbyister, som gör exakt vad deras arbetsbeskrivning antyder, nämligen att försöka utöva inflytande över parlamentets och kommissionens ledamöter.
Det kan man inte stoppa eftersom det är fullständigt normalt - vi lever i ett fritt och öppet samhälle - men vi måste göra våra röster hörda inom denna struktur och upprätthålla vårt oberoende.
Vi har inte alltid lyckats med det och det har funnits ledamöter som har brutit mot dessa regler, vilket är ett av de främsta skälen till att vi vill ändra våra regler.
Insyn och öppenhet är en av de viktigaste förutsättningarna för förtroende, och det är exakt vad vi arbetar med för närvarande.
Efter ytterst långdragna förhandlingar har vi lyckats enas med kommissionen om ett öppenhetsregister.
Jag skulle visserligen ha föredragit att rådet också hade varit med ombord.
Gruppen De gröna/Europeiska fria alliansen har kämpat länge för öppenhetsregistret.
Vi gläder oss över att vi äntligen har lyckats inrätta det och är också stolta över resultatet, men jag måste säga att vi inte är nöjda med alla aspekter.
Vi skulle ha föredragit att registret hade varit obligatoriskt, inte bara för dem som arbetar inom kommissionens och parlamentets byggnader, utan även för dem som arbetar på annat håll, till exempel över ett glas vin i en av Bryssels många barer.
Vi vill inte att registret endast ska gälla för parlamentet och kommissionen, utan även för rådet.
Vi vill att den ekonomiska information som lämnas ska vara mer exakt och meningsfull.
Vi anser vidare att de belopp som är involverade ska mätas på samma sätt i stället för den metod som föreslås nu, enligt vilken mindre transaktioner mäts i storleksintervaller på 50 000 euro, medan större transaktioner mäts i större intervaller, vilket gör det svårt att veta exakt hur mycket pengar det handlar om.
Vi är också för regelbundna kontroller som utförs av ett gemensamt sekretariat.
Icke desto mindre är detta en bra dag för EU eftersom vi får mer insyn och öppenhet.
Jag vill tacka alla som har varit med och arbetat med detta för de goda resultaten.
för GUE/NGL-gruppen. - (DA) Fru talman! Detta betänkande är ett steg i rätt riktning mot ökad öppenhet och ett obligatoriskt lobbyistregister för alla som försöker påverka EU.
Men vi har fortfarande långt kvar innan vi når vårt mål.
Dessutom måste vi se om vårt eget hus, vilket fallen med de korrumperade parlamentsledamöterna har visat.
Vi måste klargöra att det inte är godtagbart att Europaparlamentets ledamöter har någon form av betalt arbete vid sidan om som kan ifrågasätta vår integritet.
Dessutom måste vi ha effektiva kontrollmetoder och regler för att fastställa följderna om någon bryter mot reglerna.
Vi måste också skapa tydliga regler för skydd av visslare, för att förhindra att budbäraren blir skjuten.
Vi ser fram emot arbetsgruppens rapport och hoppas på en snabb översyn av det avtal vi diskuterar i dag och av parlamentets arbetsordning.
(Talaren godtog att besvara en fråga (blått kort) i enlighet med artikel 149.8 i arbetsordningen.)
(DE) Fru talman! Søren Bo Søndergaard, jag ville fråga dig vad du anser om förslaget om vägledande förteckningar och om att öppenhetsregistret fortfarande inte kommer att vara obligatoriskt, vilket innebär att det kommer att finnas stora kryphål även i framtiden.
(DA) Tack för din fråga.
Den ger mig möjligheten att upprepa en sak jag redan sagt, nämligen att vi fortfarande har långt kvar innan vi når vårt mål.
Vi anser inte att vi redan har gjort det, utan att det fortfarande saknas något.
Det står klart att det är absolut nödvändigt att registret blir obligatoriskt.
Vi anser att förslaget om ett digitalt ”fotavtryck”, dvs. vägledande förteckningar för rättsakter, är bra och att vi bör använda oss av det, men vi anser naturligtvis att även detta måste vara obligatoriskt för att det ska fungera.
Men som jag sade, det vi har nu är ett steg i rätt riktning, och när vi får rapporten från arbetsgruppen och texten ska ses över - den ska nämligen ses över inom två år - hoppas vi att vi kan uppnå vårt mål fullständigt, eftersom det är viktigt inom det här området.
(EN) Fru talman! Nu får vi äntligen ett öppenhetsregister!
Det är inte förvånande att det enda skälet till att vi har kunnat åstadkomma detta är att driftiga brittiska journalister lyckades bevisa hur lätt vissa Europaparlamentsledamöter föll för lockelsen att tjäna extra pengar.
Vid den tidpunkten bekände Europaparlamentet, inte helt olikt polischefen i filmen Casablanca, att det var chockerat - chockerat - över att upptäcka att korrupt lobbyverksamhet hade skett mitt framför näsan på oss.
Registret är hur som helst exakt samma sak som att stänga stalldörren efter det att hästen har sprungit ut.
Det är inte mycket som kommer att förändras med registret, lobbyisterna kommer alltid att ta sig igenom.
Ett frivilligt registreringssystem infördes, men det var ineffektivt.
Nu kommer vi att sprida lite ljus över vad som pågår, men det mesta kommer i alla fall att döljas i den stillastående dunkla dammen, affärerna kommer att pågå som vanligt.
Som vanligt kommer de som följer reglerna också att få bära den största byråkratiska bördan, och de som bryter mot bestämmelserna hittar sätt att fortsätta.
Så länge som så stora belopp av skattebetalarnas pengar flyter omkring i Bryssel kommer det alltid att finnas skrupelfria lobbyister, precis som att det alltid finns hyenor där det finns kadaver.
(Talaren godtog att besvara en fråga (blått kort) i enlighet med artikel 149.8 i arbetsordningen.)
(DE) Herr talman! John Stuart Agnew, jag tycker att det är positivt med välorganiserade åsiktsutbyten under debatterna, men jag tycker däremot att det är mindre trevligt när fakta förvrängs.
Därför vill jag be dig att korrigera ditt senaste uttalande.
Du har just hävdat att parlamentet bara diskuterar öppenhetsregistret för att ett antal brittiska dagstidningar uppmärksammade allmänheten på en viss historia.
Jag uppmanar dig att förklara för parlamentet och för allmänheten i stort att vi redan hade börjat diskutera den här frågan och parterna redan hade enats om öppenhetsregistret när den nyhet som du talar om ens hade skett.
(EN) Herr talman! Det verkar vara den utlösande orsaken till allt detta.
Jag vill inte att några brittiska ledamöter ska vara här i alla fall.
Jag förstår inte varför vi ska behöva stå ut med att utländska institutioner som denna sköter våra affärer.
Ju längre vi rör oss mot söder, desto värre blir korruptionskulturen.
Jag tycker inte om det, och jag vill inte att mitt land ska ha någon del i det.
(DE) Herr talman! Vi är alla väl medvetna om att inte bara Europaparlamentet utan hela EU lider av ett enormt trovärdighetsproblem.
Jag är säker på att det är något som Gerald Häfner inte vill höra talas om, men även om parlamentet äntligen har kunnat enas om öppenhetsregistret, utan tvivel genom att ge efter för påtryckningarna till följd av lobbyskandalen nyligen, kommer det i alla fall att vara tandlöst.
Jag anser att ett frivilligt register helt enkelt är hyckleri och att det inte kommer att bidra till ökad öppenhet eller att ministerrådet kommer att vara berett att delta i det, så vi har inte ens alla lagstiftande organ ombord.
Även om rådet skulle ansluta sig kommer det ändå att finnas en hel massa kryphål.
Uppenbarligen finns det hundratals expertgrupper som arbetar med de officiella rapporter som offentliggörs av kommissionen, men namnen på de medlemmar i de rådgivande kommittéer som sammanträder bakom stängda dörrar förblir en välbevakad hemlighet.
Enligt min åsikt behöver vi inte bara ett register över allt arbete som utförs av företag eller i internationella frågor, utan även för allt betalt lobbyarbete som utförs av intressegrupper som yrkesorganisationer och fackförbund.
Våra medborgare har rätt att förvänta sig verklig insyn även i det här fallet.
(EL) Herr talman! Jag gratulerar Carlo Casini till hans betänkande, som är mycket lyckat.
Insynsfrågan berör även parlamentarikernas värdighet, det råder det inget tvivel om.
Men ju fler åtgärder vi vidtar desto mer främjar vi insyn och öppenhet och fungerande förbindelser mellan EU-institutionerna, arbetsmarknadens parter och intressegrupper.
Enligt förslaget till nytt register garanteras insyn och öppenhet i hela det breda spektrumet av institutionella kontakter och registret samlar speciella intressegrupper, företrädare för det civila samhället och för offentliga myndigheter i olika kapitel, vilket innebär att man gör åtskillnad mellan intressegruppers och officiella institutionella talesmäns roller.
Registreringen skyddar identiteten för intressegrupper genom att ange dem separat och ger dem en ställning där de kan tala direkt och omedelbart med EU-institutionerna.
Efter ratificeringen av Lissabonfördraget har Europaparlamentets befogenheter utökats, vilket innebär att fler företrädare för olika intressegrupper vill göra sina röster hörda.
Avslutningsvis är det främsta syftet med öppenhetsregistret att bidra till insyn och en demokratisk pluralistisk samverkan mellan arbetsmarknadens parter, de medborgare som röstade fram oss parlamentsledamöter och EU-institutionerna.
Det är självklart att samtliga EU-institutioner och överordnade tjänstemän måste delta i registret.
(ES) Herr talman! Jag vill tacka Carlo Casini för hans betänkanden om öppenhetsregistret.
Vi upplever en kris av oerhörd omfattning som vi har dragits med länge vid det här laget, och som hotar att pågå ännu längre.
En kris som denna förvärrar människornas levnadsvillkor och försämrar deras framtidsförväntningar.
När vi på grund av en ekonomisk kris inte kan få igenom politiska åtgärder med positiva resultat för allmänheten måste vi kämpa för att få igenom politiken med en obetingad respekt för de politiska värderingar som vi förespråkar: åtstramning, ärlighet, närhet till allmänheten och öppenhet.
Öppenhetsregistret är ett steg framåt mot insyn, men det är bara ett steg.
Jag håller med mina kolleger som sagt att registret måste vara obligatoriskt, att rådet måste ansluta sig och att oegentligt uppförande måste bestraffas hårdare.
(DE) Herr talman, mina damer och herrar! När vi röstar om öppenhetsregistret i morgon kommer vi att ta ett viktigt steg i rätt riktning, men det står klart att sista ordet inte är sagt i den här frågan.
För det första gläder det mig att vi har valt ett nytt namn för Europaparlamentets lobbyregister, som härrör från 1996 och som från och med nu kommer att benämnas ”öppenhetsregistret”.
Jag tycker dock att det är beklagligt att se vilka personer och organisationer som måste registrera sig för att få ett ettårigt passerkort till parlamentets byggnader - listan omfattar offentliga institutioner och organ.
Som jag har sagt tidigare kan jag förstå varför en advokatfirma måste registrera sig, men jag har däremot svårare att först varför offentliga organ som aldrig har varit aktiva på partipolitisk nivå, och aldrig kommer att vara det, måste registrera sig.
Oavsett all insyn vi har skapat handlar det ändå om varje ledamots moraliska kompass, eftersom den anger om de tänker rätt, vem de beslutar att inte träffa och vem de väljer att lyssna eller inte lyssna till.
De personer som kontaktar oss använder ju också många olika kommunikationskanaler.
(DE) Herr talman! Att följa vår moraliska kompass kan vara svårt.
Jag anser att det handlar om vårt oberoende som parlamentsledamöter.
Lobbyarbete blir naturligtvis ett problem om någon försöker ändra på våra övertygelser genom att använda alla argument de kan, särskilt om argumenten är oärliga.
Faktum är att lobbyregistret nu bara omfattar 2 800 av de 20 000 lobbyisterna i Bryssel.
Här i parlamentet har vi också alldeles för få möjligheter att utveckla tillräckligt kvalificerad expertis, men det kan vi snabbt ändra på genom att rikta om finansieringen och det skulle jag verkligen stödja.
Öppenhetsregistret kanske bara är en liten seger, men det kan ses som ett steg i samma riktning som Washington, där lagen om offentliggörande av lobbyverksamhet har funnits en tid.
Det fungerar bättre än något vi har här.
För min del anser jag att vi inte bara bör införa ett ”rättsligt fotavtryck” dvs. vägledande förteckningar vid utarbetande av rättsakter, så snart som möjligt, utan även ett rättsligt ”fingeravtryck”, dvs. att vi bör offentliggöra namnen på alla lobbyister som vi kommer i kontakt med och vad vi diskuterar med dem.
Gå gärna in på min webbsida, där jag har installerat en lobbyisträknare, som registrerar alla kontakter med lobbyister, vare sig jag arbetar med en rättsakt eller inte.
(GA) Herr talman! Betänkandet är viktigt eftersom det handlar om själva kärnan i vårt arbete här i parlamentet, dvs. att utarbeta och genomföra regler och lagar.
(EN) Precis som Carlo Cassini sade är begreppet ”lobbyist” lite missriktat eftersom det skapar ett intryck av en privilegierad ställning eller korruption eller båda, medan dessa personer i verkligheten är experter på sina respektive områden som hjälper till att informera oss om detaljer och nyanser av de olika rättsakter som vi utarbetar förslag om.
Själv arbetar jag just nu med ett yttrande över dataskydd och det är förvånande att se hur många grupper som har kommit till mig med sina åsikter.
Om vi driver fram ett register skulle jag vilja registrera även dem som kontaktade mig, för då skulle vi ha verklig öppenhet.
Ett officiellt register över lobbyister, men även ett register över dem som vill påverka oss.
Det skulle skapa verklig insyn, ökad trovärdighet och i slutändan ökat förtroende.
(EN) Herr talman! Det har ofta sagts att våra medborgare inte vet att parlamentet har fått större befogenheter sedan Lissabonfördraget.
Det kan mycket väl vara sant och är i så fall mycket olyckligt eftersom ni kan vara säkra på att lobbyisterna - eller de som utger sig för att vara lobbyister, vilket har visat sig nyligen - är mycket medvetna om vilka befogenheter parlamentet har.
Vi medbeslutar om nästan all viktig lagstiftning i EU, och det är bra eftersom vi företräder folket i EU.
Vi är den enda direktvalda institutionen.
Men även om parlamentet är och kommer att fortsätta vara en av de mest öppna institutionerna i EU anser jag fortfarande att ökade befogenheter medför större ansvar, och det är just detta vi måste sträva efter under de kommande månaderna.
Dagens avtal med kommissionen är inte dåligt, men lobbyisterna måste bli skyldiga att ange sina namn och verkliga intressen i ett register.
Det är också vad parlamentet redan kräver av lobbyister som kommer till oss.
Jag hoppas att de andra institutionerna kommer att följa vårt exempel.
Jag avslutar med följande kommentar.
Som ni nämnde är jag medordförande för den arbetsgrupp som vi har inrättat.
Jag kan inte säga så mycket om vad vi diskuterar i detalj, men jag försäkrar er om att parlamentets uppförandekod kommer att bli en av de öppnaste, med regler som gör våra medborgare stolta och som får oss själva att känna oss hedrade över att vara ledamöter av denna utomordentliga institution.
- (SK) Herr talman! Jag vill börja med att välkomna att det framlagda avtalet kommer att bidra till att förbättra öppenheten och insynen i EU, men ärligt sagt är det fortfarande långt ifrån idealiskt.
Det är dock bra att lobbyisterna nu har större anledning att ansluta sig till registret, eftersom de inte kommer in i Europaparlamentet annars.
Tillgången till information om lobbyister, inklusive deras namn, har också förbättrats, och vi bör även välkomna att de lobbyister som inte följer reglerna kommer att bestraffas på olika sätt, de kan t.ex. strykas från registret, vilket innebär att de blir svartlistade.
Frågan är bara om dessa åtgärder är tillräckliga.
Jag kan inte hålla med om att registreringen faktiskt är obligatorisk när endast registrerade lobbyister har tillträde till parlamentet.
För att skapa ökad insyn måste registreringen vara rättsligt obligatorisk, och jag hoppas att vi kommer att åstadkomma det under den nuvarande mandatperioden.
Vi måste också förbättra reglerna för rapporterna från lobbysammanslutningar när det gäller deras utlägg för lobbyverksamhet.
Enligt det nuvarande systemet kan lobbyisterna rapportera mycket mindre belopp än de egentligen har lagt ut.
Det är lika viktigt att det råder insyn i de finansiella källor som lobbyister och konsultfirmor får sina intäkter från.
Avslutningsvis vill jag tillägga att jag verkligen skulle uppskatta om ledamöterna inte blandade ihop frågan om öppenhetsregistret med uppförandekoden, eftersom den är en helt annan fråga.
Ledamöter som på något sätt har fallit offer för falska lobbyfirmor - även om det är deras eget fel - bör inte motiveras på det sättet när reglerna för öppenhetsregistret fastställs.
Herr talman! Mycket är redan sagt men förtjänar att upprepas.
Det är bra att vi nu äntligen är överens om ett lobbyistregister.
Vi är många som har kämpat länge för det.
Men fortfarande är det ett mycket försiktigt förslag.
Jag väljer ändå att se det som ett första steg som kan utvecklas till en bred offentlighetsprincip i EU:s samtliga institutioner.
Det är väldigt bra med dagens markeringar från rådet och från kommissionsledamot Maroš Šefčovič.
Offentlighet och öppenhet är ett av få riktigt effektiva instrument för att minimera riskerna för övertramp och fusk.
Det är också en viktig väg för att öka förtroendet för oss som verkar i detta politiska system och för politik i största allmänhet.
Nästa steg bör vara att alla institutioner omfattas, att registret görs obligatoriskt och att det, i likhet med vad som görs i en del skandinaviska länder, kompletteras med ett meddelarskydd för ”visslarna”, som också är kolossalt viktiga för verklig öppenhet och transparens.
Tack.
- (SK) Herr talman! Jag välkomnar och stöder fullständigt inrättandet av ett öppenhetsregister och en förteckning över lobbyister, både för organisationer och de oberoende lobbyister som deltar i utarbetandet och genomförandet av EU-politiken, eftersom en skärpning av normerna för att garantera stabiliteten och integriteten hos EU:s offentliga förvaltning och stärka institutionsreglerna är en garanti för EU:s demokratiska fungerande.
Men registret får naturligtvis inte hindra ledamöterna från att fullgöra de arbetsuppgifter de har tilldelats enligt sitt mandat och sammanträffa med sina väljare eller företrädare för offentliga organ som agerar för EU-medlemsstaternas räkning i Europaparlamentet.
Det måste dock finnas tydliga regler för företrädare för speciella intressegrupper för att säkra en öppen, insynsvänlig och lämplig dialog med de personer och organisationer som på något sätt vill delta i utarbetandet av EU-lagstiftning och påverka den processen.
(EN) Herr talman!
Jag talar som föredragande för betänkandet om förordning (EG) nr 1049/2001 om allmänhetens tillgång till offentliga handlingar. Jag välkomnar detta avtal, som överensstämmer med andan av insyn och öppenhet i den förordningen.
Det är ännu ett steg i rätt riktning eftersom insyn och öppenhet står i centrum för den demokratiska beslutsprocessen och vi bör vara medvetna om alla som påverkar och ibland har ett olämpligt inflytande på politiken, förfarandena och resultaten.
Men vi måste göra mer, vi måste se till att insynen och integriteten i det arbete som utförs av lobbyister på EU-nivå är av hösta nivå.
Dessutom måste det nya registret tas i drift så snabbt som möjligt, och så snart vi har gjort det måste alla personer och organisationer som omfattas av det lämna korrekt och aktuell information så vi kan se vem som påverkar vad.
Avslutningsvis vill jag citera Jana Mittermaier från organisationen Transparency International: ”Det nya registret kommer att bli ett test för alla lobbyisters åtagande för ökad insyn.”
Tydligare kan det inte sägas.
(ES) Herr talman! Jag vill påpeka att 2000-talet är webbens, WikiLeaks och den institutionella insynens århundrade.
Detta innebär att det krävs öppenhet och deltagande för allmänheten, och allmänheten måste ges ett visst medansvar i beslutsprocessen.
Vi måste besluta tillsammans och därför måste vårt arbete också vara proaktivt.
Vi kan inte bara vänta på att lobby- och intressegrupper ska pressa oss, vi måste göra oss besväret att närma oss allmänheten och lyssna till människorna.
Jag anser därför att öppenhetsregistret och de vägledande förteckningarna kommer att bli effektiva.
Syftet är absolut inte att begränsa arbetet och orsaka rädsla, detta är i stället en möjlighet att förbättra våra betänkanden och mäta våra resultat.
Jag anser att det är det enda sättet för oss att utvecklas och bli ett modernt parlament.
Jag har haft ansvaret för ett betänkande, och när jag skrev motiveringen lyssnade jag till alla aktörer som jag arbetade med. Vi måste göra en tydlig åtskillnad mellan våra arbetsmetoder och de oansvariga handlingar som vi har sett tidigare.
(FR) Herr talman! Även jag är nöjd med texten, som jag gärna röstar för i morgon.
Jag vill bara påpeka att de skandaler vi har sett den senaste tiden är försök till mutor, inget annat.
Detta är en allvarlig fråga och det har hänt saker på sistone.
Vi inledde dock vårt arbete långt före den senaste tidens allvarliga händelser, som behandlas i ett annat betänkande.
De är isolerade fall, och även i det fallet har vi gjort ett bra arbete.
Vi kan emellertid se att ett antal grupper använder betydande resurser och gör allt de kan för att påverka beslutprocessen i så hög utsträckning som möjligt.
Registret är därför ett steg i rätt riktning.
Jag medverkade i arbetet med det och jag är också oerhört nöjd med allt arbete som har utförts.
Men det krävs ytterligare åtgärder.
Registret måste bli ett dynamiskt instrument som ses över årligen.
Det bör vara allt annat än strikt.
Jag anser faktiskt att den tekniska utvecklingen och de hjälpmedel som används av lobbyisterna kommer att tvinga oss att kontinuerligt se över instrumentet för att se till att det är effektivt och genom riktlinjer kartlägga vem som arbetar med lobbyverksamhet, för hur mycket pengar och på vilket sätt.
Jag är också absolut för rättsliga fotavtryck - jag menar de vägledande förteckningarna - som kan innehålla uppgifter om antalet lobbyister och namnen på de personer som de har sammanträffat med, och jag tycker att det är bra om vi kan få reda på exakt vem som sade vad och vem som påverkade vem.
Avslutningsvis är det en sak att offentliggöra registret och en helt annan att förklara hur det fungerar.
Medborgarna måste också få tillgång till registret så att de kan använda informationen på ett meningsfullt sätt när de vill sätta sig in i vår beslutsprocess.
Därför kommer vår grupp att oreserverat rösta för den här texten.
(DE) Herr talman! Lobbyverksamhet är ett centralt instrument för medborgarnas deltagande i det politiska livet, och därför är det viktigt att förhindra missbruk.
Det är också därför som det snabbt krävs ett öppenhetsregister för samtliga institutioner, inte bara för parlamentet och kommissionen utan även för rådet, eftersom det faktiskt är där som alla beslut fattas.
Jag vill upprepa att registreringen måste vara obligatorisk, inte bara för tillträde till parlamentet eftersom alla lobbyister ju inte hittar sina kontakter i parlamentets byggnad, utan även och oftare i restauranger, vid cocktailmottagningar eller på gymmet.
Jag vill även säga ett par ord om insyn i politiska partier.
Även om de är enmanspartier som agerar självständigt och försöker framställa sig själva som ärligast i världen, måste dessa partier och personer uppfylla insynskraven.
De måste garantera insyn när det gäller deras tillgångar, hur stora offentliga medel de beviljas och hur stora ersättningar de får för kampanjkostnader, med andra ord de verkliga belopp som de fått från offentliga organ i sina egna länder under valkampanjerna.
Dessa kostnader måste dokumenteras på ett öppet sätt.
(PL) Herr talman! Tack för att jag får ordet.
Precis som majoriteten här i parlamentet håller jag med om att registret utgör ett framsteg när det gäller insynen i lagstiftningsförfarandet, men enligt min mening är det bara ett första steg.
Vi bör allvarligt överväga andra åtgärder och lösningar.
Enligt min mening är den viktigaste frågan vad Europaparlamentsledamöterna får eller inte får göra.
Får de endast arbeta som parlamentsledamöter här i parlamentet eller får de också syssla med annat vid sidan av sitt arbete här?
Personligen anser jag att dessa andra verksamheter bör fastställas noggrant och att de bör vara begränsade till vetenskapligt arbete och publikationer.
Allt annat arbete i olika styrelser kommer alltid att ge upphov till frågetecken och tvivel.
Herr talman! Europaparlamentet har genom Lissabonfördraget fått ökade maktbefogenheter och det innebär också ett större ansvar.
Transparensen i vårt arbete är därför oerhört viktig, med tanke på att vi arbetar med lagstiftning för 500 miljoner människor och ofta väldigt stora ekonomiska värden.
Den lista för lobbyister som nu beslutats i kompromissen är naturligtvis väldigt värdefull, och jag hoppas att vi kan gå vidare med ett meddelarskydd för visslare.
Jag hoppas vidare att vi kan gå vidare och se till att uppgifterna i registret för ekonomiska ansvarsförbindelser eller ägande blir obligatoriska, och inte frivilliga som i dag är fallet.
Jag hoppas också att vi får en diskussion om vilka sidouppdrag som ur etisk synvinkel är lämpliga när man har ett uppdrag som EU-parlamentariker.
Jag uppskattar kompromissen och ser den som en väg framåt, men det finns många fler steg att ta på den väg som leder mot transparens, öppenhet och större demokratiskt förtroende.
Tack.
kommissionens vice ordförande. - (EN) Herr talman! Jag anser att Manfred Weber har helt rätt när han säger att vi ska vara stolta över att öppenhetsregistret drivs gemensamt eftersom jag, med undantag för Förenta staterna och Kanada, inte känner till något annat land utanför EU där ett öppenhetsregister som det vi kommer att inrätta fungerar.
Här avser jag också medlemsstaternas huvudstäder.
Frågan om huruvida registret ska vara obligatoriskt togs upp av flera talare, först Matthias Groote och därefter Gerald Häfner.
I arbetsgruppen diskuterar vi denna fråga mycket ingående.
Problemet är att vi för närvarande inte har någon rättslig grund för att tvinga företag, medborgare eller intressegrupper att registrera sig för att utöva sitt yrke.
Som EU-förvaltning kan vi inte vägra att ha kontakt med sådana personer eller organisationer på den grunden.
Därför har vi funderat över hur vi på ett positivt sätt kan motivera företag, organisationer och lobbyister att registrera sig. Jag anser att vi har åstadkommit en hel del, eftersom vi med parlamentets samtycke faktiskt håller på att göra detta register obligatoriskt.
Med våra gemensamma insatser, tillsammans med rådet, kommer vi att öka registrets anseende och pressa på så mycket vi kan. Under de närmaste åren kommer vi att se hur det fungerar och detta kommer att ge oss ytterligare erfarenhet för att kunna göra en bra översyn, där vi ser hur vi kan förbättra systemets funktionssätt ännu mer.
När det gäller kraven på lämpliga kontroller av finansieringen av verksamheten för dem som registrerar sig kan jag försäkra er om att kommissionen redan utför stickkontroller av alla som finns i registret och jag är säker på att dessa kontroller till och med kommer att öka när vi väl driver registret gemensamt.
Alla som är med i registret kan vara säkra på att om det finns något olämpligt så kommer vi att upptäcka det, påtala det och försöka rätta till det, och vi kommer inte att vara rädda för att namnge de ansvariga.
Jag blev väldigt glad över att höra - jag kommer tillbaka till den frågan eftersom flera talare påpekade att den är viktig - att samtliga tre institutioner gör framsteg i detta arbete.
Efter det att det ungerska ordförandeskapet nu har inlett arbetet är jag säker på att vi inte kommer att slösa bort en enda minut och vi kommer att försöka inleda de interinstitutionella samtalen med rådet så snart som möjligt så att vi, och det är jag säker på, kan finna ett lämpligt sätt att driva registret tillsammans, och att de tre institutionerna arbetar mot samma mål i den här frågan, dvs. ökad insyn i EU:s lagstiftning.
Den sista punkten jag vill nämna togs upp av flera talare och beskrevs av Carlo Casini. Öppenhetsregistret är definitivt ingen silverkula eller en magisk lösning för att bekämpa korruption.
Vi vet mycket väl att höga moraliska standarder, etik, värdighet och tydliga regler är avgörande i det här sammanhanget.
Men registret kommer däremot att vara ett mycket bra instrument och en bra indikator på att de som registrerar sig är beredda att följa reglerna och arbeta på ett öppet sätt, att de inte har något att dölja och - vilket bör vara en viktig ledstjärna för oss alla - att de kommer att arbeta med oss i ett verkligt partnerskap och utbyta information med oss, och att de slutligen har förtroende för vår framtida kommunikation.
rådets ordförande. - (HU) Herr talman, herr kommissionsledamot, mina damer och herrar! Som företrädare för en medlemsstat som har en lagstiftning om lobbyverksamhet sedan 2006, välkomnar jag dagens debatt samt att parlamentet och kommissionen kan komma överens i frågan om ett öppenhetsregister.
Öppenhet har alltid varit en viktig fråga för rådet.
Under 2008 och 2009 lyckades vi inte göra några genombrott i förhandlingarna, men jag är väldigt glad över att vi nu under det ungerska ordförandeskapet fick ett genombrott. Rådet är redo att garantera insyn i processerna och delta i verksamheten såtillvida det kan göra det - vi får se i vilken omfattning det blir.
Vi är redo att förhandla om vårt deltagande och, som jag angav i mitt inledande anförande, vi tror att vi kan offentliggöra vår avsikt i en politisk förklaring i juni.
Men detta betyder inte att vi skulle ansluta oss till det interinstitutionella avtalet.
Anledningen till att medlemsstaterna nu kan anta formuleringen - som jag än en gång måste betona utgör stora framsteg i jämförelse med tidigare år - är att lobbyisterna inte kontaktar rådet som europeisk institution, det finns ytterst få exempel på det.
De inriktar sig snarare mot medlemsstaterna, deras regeringar och statliga organ.
Rådet är därför inte utsatt för lobbyverksamhet i samma utsträckning som kommissionen eller parlamentet.
Herr talman, herr kommissionsledamot, jag hoppas att samarbetet blir effektivt och att vi kommer att kunna komma fram till den politiska förklaringen efter förhandlingarna.
föredragande. - (IT) Herr talman, mina damer och herrar! Jag vill förtydliga några punkter.
Jag vill också kraftfullt betona att avtalet var klart långt innan historien med de brittiska journalisterna bröt ut.
Tyvärr är detta ett sätt att sprida falsk information via media.
Den stora italienska tidningen Corriere della Sera har till exempel i dag skojat med EU och skrivit att vi agerade alltför sent och först efter händelserna med journalisterna.
Det är inte sant.
Det föranleder en omotiverad misstro mot EU.
Avtalet ingicks långt tidigare.
Diskussionen uppstod först något senare, för när skandalen väl var ett faktum funderade vi på om vi kunde stärka avtalet ytterligare.
Men texten förblev oförändrad.
Det är det första förtydligandet.
Den andra punkten avser frågan om skyldighet.
Registret är redan obligatoriskt.
De som vill utöva lobbyverksamhet måste skriva in sig i registret.
Jag förstår inte vad ”obligatoriskt” betyder. Det kan inte betyda att alla bolag, alla företag eller alla medborgare måste skrivas in i registret.
Det är omöjligt.
Det är upp till varje parlamentsledamot att uppmana dem som vill utöva lobbyverksamhet att registrera sig innan de tar kontakt.
Den tredje punkten avser möjliga framtida ändringsförslag.
En arbetsgrupp är tillsatt i detta syfte och jag anser att den behöver ha så stor handlingsfrihet som möjligt.
Jag instämmer i att vi bör identifiera lobbyisterna som vi möter under förhandlingarnas gång, men jag vet inte om den uppgiften tillkommer föredraganden eller om den bör tillkomma ordföranden.
Arbetsgruppen är fri att lägga fram alla nödvändiga rekommendationer.
Jag vill slutligen tacka både Maroš Šefčovič, som har gjort mycket stora insatser för att genomföra avtalet, och företrädaren för den ungerska regeringen för bland annat försäkran om att rådet inom kort ska ansluta sig till avtalet, något som utan tvekan var osäkert eftersom rådet företräder den andra kammaren i det här fallet.
Om rådet också inrättar registret skulle det betonas mer effektivt att EU:s struktur består av en regering - kommissionen - och ett lagstiftande organ, som består av både medborgarnas och medlemsstaternas företrädare.
Men jag inser att det finns fler frågor som måste besvaras, eftersom ministerrådet företräder medlemsstaterna.
Jag är ändå övertygad om att vi kommer att uppnå ett positivt resultat.
Debatten är härmed avslutad.
Omröstningen kommer att äga rum onsdagen den 11 maj 2011.
Skriftliga förklaringar (artikel 149 i arbetsordningen)
, skriftlig. - (EN) Vi är alltid stolta över att vara den mest öppna europeiska institutionen.
Men under de senaste åren har det visat sig att oavsett vilka fördelar detta medför, har systemet även sina nackdelar.
Vi är alla medvetna om hur europeiska medborgare har förlorat och fortfarande förlorar tilltro till EU och - låt oss vara ärliga - till oss parlamentsledamöter.
Ett viktigt sätt för att få tillbaka förtroendet är att öppet redogöra för det vi gör och hur vi påverkas i vårt arbete.
Det gemensamma öppenhetsregistret som vi ska anta i dag genom att rösta ja till bägge betänkandena som lagts fram, utgör ett första steg i den riktningen.
Det är ett ”första steg” eftersom det inte kommer att lösa alla våra problem.
Även om det är svårt att genomföra i dag, ska vi i framtiden sträva efter obligatorisk registrering av lobbyister.
Jag vill också understryka att ett sådant register inte ersätter våra enskilda försök till öppenhet och behovet av att se över vårt arbete i det avseendet.
Jag välkomnar kommissionens och Europaparlamentets gemensamma öppenhetsregister.
Men det bör utgöra endast ett av flera mycket viktiga steg mot ökad insyn i lagstiftningsprocessen, som bör gälla samtliga tre europeiska institutioner.
Europaparlamentet är villigt att föra en allvarlig debatt om lobbyverksamhet och bestämmelserna om lobbyverksamhet.
Det statuerar också ett exempel för de medlemsstater som fortfarande måste ta steget.
Jag anser att öppenhetsregistret också kommer att bidra till ökad tilltro till den politiska verksamheten.
Men dess verkliga inverkan kommer främst att bero på hur var och en följer de strängaste reglerna.
, skriftlig. - (NL) Jag kan bara välkomna kommissionens och parlamentets gemensamma arbete för att inrätta ett gemensamt öppenhetsregister för lobbyister, tankesmedjor och andra intresseorganisationer.
I varje fråga på vår agenda måste vi helt öppet kunna lyssna till olika intressegrupper.
Det finns förresten inget fel i det att organisationer försvarar sina egna intressen, om det sker öppet och väl balanserat.
Principen om ”legislative footprint” (vägledande förteckning), enligt vilken föredragandena måste ange vem de har varit i kontakt med i samband med utarbetandet av förslagen, är en bra åtgärd.
Jag har redan tagit upp det i mitt betänkande om leksakers säkerhet.
Tydliga anvisningar för en allmän tillämpning av principen kommer att öka insynen.
Det är också ett lämpligt instrument för att slå hål på de myter om lobbyverksamhet som sprids bland allmänheten, vars gemensamma intressen vi parlamentsledamöter ska främja.
Att rådet också angav att det är redo att ansluta sig till registret innebär att vi kommer att ha ett enda register för alla EU-lobbyister. Det är något som vi tillsammans med Europaparlamentet har arbetat för under flera år.
Jag stöder därför systemet.
18.
Handelsförbindelserna EU-Japan (omröstning)
(PL) Herr talman! I detta ändringsförslag skulle PPE-gruppen vilja stryka ordet ”starkt” i punkt 2.
Jag hoppas att det inte finns några invändningar.
Öppnande av sammanträdet
1.
Sri Lanka: uppföljning av FN-rapporten (debatt)
Nästa punkt är debatten om sex förslag till resolutioner om Sri Lanka.
(EN) - Herr talman! I Sri Lankas regerings brutala krig mot den tamilska minoriteten dödades åtminstone 40 000 tamiler inom loppet av några veckor och hundratusentals internerades i fångläger ute i det fria.
FN-rapporten erkände långt om länge officiellt de brott som hade begåtts mot det tamilska folket.
Tyvärr bör man inte göra sig några illusioner om att rapporten kommer att ändra tamilernas situation i Sri Lanka.
Dagen efter rapportens publicering rapporterade man att FN:s generalsekreterare endast skulle starta en internationell undersökning om Sri Lankas regering samtycker eller om ett internationellt forum, såsom FN:s säkerhetsråd, kräver en undersökning.
Mot bakgrund av karaktären på Sri Lankas regering är det uppenbart att den inte kommer att tillåta någon internationell undersökning.
Det belyser än en gång behovet av att genomföra en kampanj för en verkligt oberoende undersökning om krigsbrotten och för att Rajapaksa-regimen ska hållas ansvarig för dem.
Den 18 maj kommer protester att genomföras i hela världen, vilka anordnas av många grupper, däribland kampanjen för solidaritet med tamilerna, för att uppmärksamma den andra årsdagen av detta blodiga krig.
En förenad kamp från singaleser och tamiler behövs fortfarande för att besegra denna regim och kämpa för rätten till självbestämmande för det tamiltalande folket.
Herr talman! Vi behöver bara höra dessa inledande kommentarer för att förstå varför jag djupt beklagar att vi har denna debatt i dag.
Den stöds av extremistelement i den tamilska diasporan, samma individer som har hjälpt till att upprätthålla LTTE:s terroristkampanj under många år genom politisk verksamhet och ofta genom brott.
Naturligtvis var de sista skedena av LTTE-kampanjen förfärliga.
I FN:s Darusman-rapport, som är den omedelbara förevändningen för denna debatt, konstateras tydligt och klart att under slutfaserna använde LTTE civilbefolkningen som mänskliga sköldar, intensifierade tvångsrekryteringen av civila, inklusive barn, till sina led, avrättade civila som försökte fly från konfliktzonen och utplacerade artilleri i närheten av fördrivna civilpersoner och civila inrättningar, såsom sjukhus.
Detta ursäktar inte beskjutningen av civila mål, men den sätts i ett sammanhang och visar var skulden ligger.
I stället för att försöka föra samman Sri Lankas folk finns det de som försöker fortsätta en kampanj av hat och splittring.
De ser Darusman-rapporten som ett vapen i denna kampanj och vill bara sätta Sri Lankas regering på de anklagades bänk.
Denna taktik är ondskefull och kontraproduktiv.
Sri Lankas regering och kommissionen har inrättat en kommission för dragande av lärdomar och åstadkommande av försoning (LLRC) för att undersöka anklagelser om kränkning av de mänskliga rättigheterna.
Låt oss göra allt vi kan för att stödja dem och Sri Lankas folk i stället för att gå till angrepp mot dem.
Herr talman! Från de allra första orden har ni alla förstått att debatten skulle bli mycket livlig och att det skulle finnas två åsikter.
Jag skulle vilja säga att min grupp inte lierar sig med vare sig med den eller med den andra sidan, utan helt enkelt stöder rättvisa och försoning.
Jag tror inte att det kan bli någon försoning om inte rättvisa skipas i dessa länder, som Sri Lanka, men det finns säkert många andra som har upplevt ohyggliga krig.
Vad gör nu denna FN-rapport som Geoffrey Van Orden refererar till?
Den upprepar helt enkelt fakta och kräver en mekanism för internationell rättvisa, som man vet måste godkännas av regeringen.
Det är det allra minsta.
Hur skulle ni vilja att ett folk försonades?
Det gäller båda sidor, Geoffrey Van Orden.
Det är inte bara på tamilsidan.
Det har förekommit brott på båda sidorna.
Båda sidorna är ansvariga.
Rättvisa måste skipas av båda sidorna.
I rapporten konstateras också, och jag ber om ursäkt för detta, att den försoningskommission som just nämnts inte hade ett utredningselement av tillräckligt hög standard.
Till sist är jag rädd för att ett nationellt rättviseorgan inte kommer att slutgiltigt resultera i ett klargörande av fakta.
Därför säger jag helt enkelt och i alla deras namn som har lidit på båda sidor, att denna kammare bara kan stödja detta betänkande för att sprida mer ljus och åstadkomma mer rättvisa.
Det är det enda budskap som jag skulle vilja vidarebefordra i dag.
Jag kommer inte att ha använt all min tilldelade tid men detta är det väsentliga budskapet för denna kammare.
Herr talman! I februari åkte jag till Sri Lanka med delegationen för förbindelserna med Sydasien.
Medan vi var där blev vi vittne till de enorma insatserna för att komma över följderna av ett 25-årigt inbördeskrig.
EU, FN och frivilligorganisationerna hjälper till, från att röja undan landminor genom HALO Trust till tamilernas återflyttning till sina tidigare hem.
Vi uppmanar regeringen där att svara positivt på FN:s expertpanels rekommendationer som uppmärksammade krigsbrott och brott mot mänskligheten från både singalesernas och LTTE:s sida.
Det är uppmuntrande att regeringen har tillsatt en kommission för att åstadkomma försoning, införa rättsskipning, lösa språkproblem och hantera problemet med tidigare soldater i frontlinjen.
Den konsekventa beredvilligheten att samarbeta, viljan att integrera minoriteter och försäkran om att upprätthålla internationella rättsliga normer bildar basen för utvecklingen av ett land som utan våld och terror har en verklig framtid.
Vi uppmanar med eftertryck EU:s höga representant att stödja insatser av detta slag.
Herr talman! Konflikten i Sri Lanka är visserligen slut men många frågor återstår att besvara.
Ett slut på en konflikt innebär inte nödvändigtvis att konflikten är över i människors sinnen.
Seger är inte samma sak som fred.
Det krävs tid, ansträngning och speciellt engagemang och stark vilja för att komma över ärren efter en konflikt.
Försoning är absolut nödvändigt.
Rättvisa är centralt för en ny start.
Därför borde Sri Lankas regering omedelbart inleda undersökningar om brotten mot internationell humanitär rätt och de mänskliga rättigheterna.
Båda sidor måste undersökas.
Internationella konventioner som Sri Lanka deltar i kräver utredningar om de påstådda kränkningarna och åtal mot dem som är ansvariga.
Bara genom en öppen och ärlig undersökning och genom rättvisa kan Sri Lankas befolkning läka såren efter en lång och svår konflikt och fortsätta sitt liv i fred.
ALDE-gruppen applåderar FN:s generalsekreterare Ban Ki-moons rapport och initiativ om Sri Lanka.
Vi stöder helt och fullt FN:s rekommendationer.
Herr talman! Den 23 maj 2009 undertecknade FN:s generalsekreterare Ban Ki-moon och Sri Lankas president Rajapaksa ett gemensamt uttalande där Sri Lanka samtyckte till att garantera ansvarsskyldighet för påstådda krigsbrott och brott mot mänskligheten under det krig som slutade i maj 2009.
Eftersom denna överenskommelse inte hade infriats av Sri Lankas regering tillsatte FN:s generalsekreterare en expertpanel för att ge honom råd om modaliteter för en ansvarsskyldighetsprocess.
I rapporten som publicerades helt nyligen gjorde man trovärdiga påståenden om att både regeringsstyrkorna och Tamilska befrielsetigrarna underlät att respektera normerna för internationell rätt.
I rapporten betonades behovet av ansvarsskyldighet på båda sidor.
Sri Lankas regering har avvisat panelens rapport och kallar den olaglig och vinklad.
Jag anser att det är ett objektivt skäl för ytterligare undersökningar.
I en tid när det förtjänstfulla och berättigade arbete som internationella organisationer för mänskliga rättigheter utför missaktas är det viktigt att parlamentet träder fram och försvarar internationell rätt.
Krigsbrott får aldrig förbli ostraffade var de än inträffar.
Herr talman! Inbördeskriget i Sri Lanka varade i 25 år och slutade med ett nederlag för de tamilska tigrarna.
De sista skedena av kriget var särskilt blodiga och tusentals dog under krigets sista månader.
Enligt den nya rapporten från FN är det mycket troligt att de tamilska tigrarna och regeringstrupperna kommer att befinnas skyldiga till de allvarliga brott mot internationell humanitär rätt och mänskliga rättigheter som begicks i konfliktens slutskeden.
De tamilska tigrarna misstänks för att ha skjutit civila som försökte fly.
Regeringen dödade civila med bomber.
Båda dessa är allvarliga brott och får inte nonchaleras.
Därför är det viktigt att FN kan genomföra en opartisk och öppen undersökning om denna fråga.
Tyvärr har Sri Lankas regering varit obenägen att tillåta att undersökningarna fortsätter utan dess godkännande om inte FN:s medlemsstater enhälligt insisterar på det.
Det är ytterst viktigt att Sri Lanka intar en konstruktiv hållning och är villigt att samarbeta.
En känsla av ansvar är nödvändig för försoningsprocessen.
EU måste stödja insatser för att stärka Sri Lankas ansvarskänsla.
I slutsatserna i Darusman-rapporten från FN konstateras att massakrer på tiotusentals civila, krigsbrott och brott mot mänskligheten liksom andra hemska kränkningar av humanitär rätt har begåtts både av Tamilska befrielsetigrarna (LTTE) och Sri Lankas regering.
Att genomföra en oberoende undersökning och ställa de ansvariga inför rätta är inte ett politiskt val utan en skyldighet enligt internationell rätt.
Den försoningskommission som har inrättats av regeringen uppfyller inte grundläggande krav på oberoende.
Därför måste det internationella samfundet - särskilt EU och FN:s säkerhetsråd - erbjuda sitt ovillkorliga stöd för rapportens rekommendationer och vidta brådskande åtgärder för att skapa en oberoende internationell mekanism för att övervaka Sri Lankas regerings åtgärder, garantera att brott som begåtts på båda sidor undersöks och söka rättvisa för Sri Lankas folk.
Herr talman! Jag vill stödja denna resolution om kränkningar av de mänskliga rättigheterna och krigsbrott som begåtts i Sri Lanka.
Det är ytterst viktigt att vi, förutom att uttrycka vår solidaritet med offren och fördöma våldet mot bakgrund av problemen beträffande rättsväsendets brist på oberoende, stöder att en seriös, opartisk öppen undersökning företas av en oberoende organisation så att de personer som är ansvariga på båda sidor av konflikten kan identifieras och straffas.
Straffrihet för krigsbrott måste upphöra om vi vill förhindra att de upprepas i framtiden.
I Sri Lanka bombades civilbefolkningen bland andra illgärningar.
För sjuttiofyra år sedan bombade Francos trupper staden Guernica i mitt eget land och dödade mer än hälften av befolkningen, en händelse som har avbildats utmärkt av Picasso.
Alltsedan dess har Guernica varit en universell symbol för fred och motstånd.
Det är emellertid allas önskan att göra framsteg och nå försoning.
Vi måste därför uppmuntra, hjälpa och också driva på Sri Lankas regering för att den ska fortsätta dessa åtal så att verklig fred och rättvisa kan åstadkommas.
Herr talman! FN-rapporten som publicerades den 11 april belyser de krigsbrott och brott mot mänskligheten vilka begicks i Sri Lanka under konflikten mellan Mahinda Rajapaksas regeringsstyrkor och de tamilska tigrarnas separatiströrelse.
Striderna i maj och juni 2009 ledde till krigsbrott och brott mot mänskligheten och tusentals civila miste livet.
Vi kan inte acceptera straffriheten för de ansvariga och för upphovsmännen till dessa brott.
Rajapaksas regering har gjort allt som står i dess makt för att förhindra publiceringen av FN-rapporten och bestrider till och med dess slutsatser.
I Sri Lanka är pressen försedd med munkavle och journalisterna utsätts för hotelser och godtyckligt frihetsberövande.
Oppositionens viktigaste informationsplats på nätet har fått sitt tillträde blockerat av de rättsliga myndigheterna samtidigt som tillträde till flyktinglägren för tillfället fortfarande är ytterst begränsat, också för FN.
Den tamilska minoriteten är offer för ett folkmord som man inte får nämna namnet på.
Vi måste skyndsamt skicka observatörer från parlamentet till norra Sri Lanka för att se vad som verkligen händer där och åter hävda principen om folkens självbestämmanderätt.
(Talaren godtog att besvara två frågor (blå kort) i enlighet med artikel 149.8 i arbetsordningen.
(EN) Herr talman! Jag hörde det direkt på franska och det ord som användes var 'génocide', vilket betyder folkmord och det har en särskild betydelse i internationell rätt.
Om något sådant var avsikten från Sri Lankas regering hur kommer det sig då att de just har släppt 200 000 tamiler som var fångar?
Det är absurt att anklaga Sri Lankas regering för folkmord.
Jag hoppas att ledamoten tar tillbaka det uttalandet.
(FR) Herr Tannock! Jag använde det ordet som en metafor, framför allt för att beteckna företeelsen.
Jag har emellertid klargjort att det inte var namnet.
Fakta måste fastslås.
Hur som helst det som händer den tamilska minoriteten kan man inte avfärda med ett enkelt smärtstillande medel.
(EN) Herr talman! Föregående talare nämnde att hon efterlyser någon slags kommission som ska resa till Sri Lanka för att se vad som försiggår på ort och ställe där.
Skulle jag kunna få påminna henne om att delegationen för förbindelserna med Sydasien just har varit i Sri Lanka - och jag ser flera medlemmar av den delegationen i kammaren.
Och min kollega, Thoman Mann, refererade faktiskt till besöket där: den föregående talaren lyssnar uppenbart inte på vad som pågår i denna debatt.
Människor har varit i Sri Lanka.
De känner till Sri Lanka och de vet vad som pågår.
Jag vet inte var Karima Delli får allt detta nonsens ifrån.
(FR) Du har rätt, vi har redan skickat en delegation dit och jag inser att den delegationen var av formidabel karaktär när jag förstår att du arbetade på den.
Men vi kan också utöva påtryckningar vilket innebär att vi absolut måste upprepa detta förfaringssätt.
Herr talman! Sri Lanka är ett härjat land.
Inbördeskriget slutade officiellt för nästan två år sedan och vi vet under vilka förhållanden det ägde rum.
I det landet misslyckades FN kapitalt.
Rapporterna från icke-statliga organisationer är fördömande.
Tusentals civila dödades mellan januari och maj 2009.
Illdåd begicks av båda lägren men det förefaller som om man accepterar att pro-regeringsstyrkor medvetet bombade zoner där de hade uppmanat civilbefolkningen att ta skydd.
Sedan dess har Sri Lankas regering manövrerat för att rentvå sig och hindra tillgång till rättvisa för dem som åtminstone måste kallas offer för krigsbrott.
Regeringen har inte upphört med att försöka underskatta antalet civila som var närvarande i krigszonen samtidigt som den till och med har berövat dem humanitärt bistånd, inklusive livsmedel, vatten och hälsovård.
De tamilska tigrarna har sin del i ansvaret för dessa fasor.
De tvångsinkallade barnsoldater och använde civilbefolkningen som mänskliga sköldar men det minskar på intet sätt regeringsmyndigheternas ansvar på ort och ställe.
Det rättfärdigar inget.
FN väntade länge innan det kritiserade situationen i landet.
Vad som är värre är att Sri Lankas regering har mångdubblat sina intriger för att förhindra publiceringen av särskilt den senaste rapporten och för att få dess slutsatser förkastade.
Vi kan bara välkomna rapporten av den 11 april.
Resolutionen framför oss i dag går i rätt riktning.
För min del skulle jag ha velat att den gick ännu längre.
Det är hög tid att internationell rättvisa gör vad den ska i Sri Lanka lika väl som annanstans.
Herr talman! Den långvariga militära konflikten mellan regeringsstyrkorna och Tamilska befrielsetigrarnas väpnade grupper, vilken har haft mycket blodiga konsekvenser för civilbefolkningen som bor i konfliktzonerna, upphörde 2009.
Efter krigets slut lovade Sri Lankas president Mahinda Rajapaksa att undersöka alla misstänkta brott mot militärlagarna och internationell humanitär rätt under den militära konflikten.
I FN-rapporten som publicerades i april i år konstateras att båda sidorna i konflikten utförde militära operationer utan att vidta åtgärder för att skydda civilbefolkningens rättigheter och liv.
Trots detta har ansvariga myndigheter i Sri Lanka två år efter krigets slut inte ställt de personer som är ansvariga för allvarliga kränkningar av humanitär rätt till svars.
De rättsliga myndigheterna är i många fall passiva och vi måste därför genom vår resolution stödja FN-insatser för att upprätthålla lagen och utkräva ansvar för dödandet och tortyren av tusentals civila under de brutala striderna mellan Tamilska befrielsetigrarna och regeringsstyrkorna i Sri Lanka.
(PL) Herr talman! De dramatiska händelserna i Sri Lanka som beskrivs i FN-rapporten visar vilka slags problem som kan orsakas av väpnade konflikter.
Det som inträffade där är ytterligare bevis på att försök att lösa meningsskiljaktigheter genom våld och vapenmakt skapar andra mycket stora problem.
I Europa har man i århundraden reflekterat över begreppet ett rättfärdigt krig.
Vad som är särskilt smärtsamt är att i den moderna världen medför även ett krig, som teoretiskt är rättfärdigt, oundvikligen lidande för oskyldiga och oberättigade offer.
Detta händer oberoende av hur vi definierar ett rättfärdigt krig.
I fallet Sri Lanka visar allt fler uppgifter på att kriget inte var rättfärdigt för någondera sidan.
Segraren har inte alltid rätt även om de alltid försöker bevisa att de har rätt.
Om det verkligen ska bli en försoning, såsom Sri Lankas regering har deklarerat, måste grunden för en sådan försoning vara sanningen om vad som hände under kampen mot de tamilska tigrarna.
Det kommer inte att bli en äkta försoning utan att man avslöjar de krigsbrott som begicks oberoende av vilken sida det var som begick dem.
Det kommer inte att bli någon försoning om båda sidor anser att deras egna synder är tabu och inte tillåter att de nämns.
(EN) Herr talman! Många i denna kammare har varit inblandade i Sri Lankas politik och självklart i Sri Lankas diasporas och det tamilska samfundets politik.
Det vi diskuterar i dag är en rapport av generalsekreterarens expertpanel om ansvarsskyldighet i Sri Lanka.
Jag har inte hört någon i kammaren hittills som ifrågasatt den rapportens reella kvalitet.
Jag har läst rapporten och jag har talat med många om rapporten på båda sidor.
Om vi nu säger att vi borde bordlägga rapporten, och inte göra undersökningar om vad som hände mellan januari och maj och verkligen inte öppna en möjlighet för att undersöka många anklagelser på båda sidor, vad är då meningen med en rapport av detta slag?
Jag tycker faktiskt att det är oavvisligt att en diasporaorganisation för det tamilska samfundet, det globala tamilska forumet, har sagt att trovärdiga anklagelser mot LTTE - och de har markerat detta mycket tydligt - också ska undersökas.
Vi har en rapport som borde få en uppföljning och jag talar varmt för behovet av ett riktigt förfarande för undersökning av ansvarsskyldighet, vilket skulle leda till sanning, rättvisa och försoning för Sri Lanka efter vad som kommer att bli en plågsam undersökning, men en undersökning som måste ske.
(EN) Herr talman! Det är skrämmande att nästan 100 000 människor dödades under den långdragna militära konflikten i Sri Lanka som slutade 2009, däribland tiotusentals civila, av vilka de flesta dog i slutskedet av konflikten.
Det internationella samfundet borde kräva en kraftfull internationell undersökning av trovärdiga rapporter om illdåd som begåtts på båda sidor.
Det är synd att länder som Kina och Ryssland motsatte sig diskussion om ämnet i FN:s säkerhetsråd och att FN:s generalsekreterare skulle vidta kraftfullare åtgärder för att undersöka de brott som begåtts.
FN:s expertpanel visade tydligt att både Sri Lankas regering och de tamilska rebellerna begick allvarliga brott mot internationell humanitär rätt och de mänskliga rättigheterna, eventuellt var de i vissa fall krigsbrott och brott mot mänskligheten.
Därför stöder jag helt och fullt att man omedelbart inrättar en internationell rättvisemekanism, såsom föreslås i FN-rapporten.
(FI) Herr talman, herr kommissionsledamot! Av FN-rapporten framgår tydligt att tusentals civila dog i artillerield från regeringstrupperna under de sista blodiga månaderna av inbördeskriget i Sri Lanka, vilket pågick i 25 år.
FN sade också att de tamilska rebellerna hade använt mer än 300 000 civila som mänskliga sköldar och skjutit civila som försökte fly.
Båda sidor begick därför allvarliga överträdelser mot de mänskliga rättigheterna och internationell rätt i en krigssituation.
Det är viktigt att försoningssamtal nu kommer igång, så att FN kan genomföra en opartisk och oberoende undersökning om krigsbrott.
Parlamentets resolution är välbalanserad i ordvalet och kommer att uppmuntra parterna att nå försoning och åstadkomma fred.
(RO) Herr talman! I slutsatserna från FN-rapporten som publicerades den 25 april 2011 framförs allvarliga anklagelser om de flertaliga brotten mot de mänskliga rättigheterna och normerna för internationell rätt, både av Sri Lankas regering och de rebellstyrkor som besegrades i inbördeskriget vilket varade gott och väl 28 år.
I rapporten konstateras faktiskt att regeringsstyrkorna dödade tiotusentals civila genom att bomba befolkade områden, sjukhus och till och med centrum för humanitärt bistånd som tillhörde FN.
Å andra sidan använde rebellstyrkorna många civila som mänskliga sköldar och de som försökte fly från konfliktzonen sköts på plats.
I likhet med andra talare före mig anser jag att en oberoende internationell mekanism behöver inrättas för att undersöka krigsbrotten i detta land men också de andra allvarliga brotten mot de mänskliga rättigheterna.
En opartisk öppen undersökning krävs som kan utröna vem som är ansvarig för dessa brott som har chockat det internationella samfundet.
(EN) Herr talman! Denna rapport som grundas på väl genomförda efterforskningar visar oss - förutom alla sina slutsatser - att än en gång är det sanningen som är det första offret för kriget.
Vad den inte lyckas göra är att dra upp riktlinjerna för den politik som behövs för att läka nationens sår.
Alltför många länder blundade alltför länge för vad som pågick.
Den rätta politiken behövs nu i form av en samlad insats av det internationella samfundet för att söka frigörelse och rättvisa för alla dem som har blivit så fruktansvärt drabbade.
(EN) Herr talman! Graham Watson har alldeles rätt när han säger att det första offret i alla krig, och särskilt i detta, är sanningen.
Givetvis måste vi också medge att civilbefolkningen är offer i detta slags konflikt och FN-panelen har klart visat att båda sidor är ansvariga: huvudsakligen regeringen men också Tamilska befrielsetigrarna och båda måste undersökas.
Det vi säger är att en ordentlig utredning inte är särskilt trolig om utredningskommissionen tillsätts av regeringen.
Det vi begär är att en oberoende kommission ska undersöka dessa anklagelser om krigsbrott och brott mot mänskligheten, som identifierats av FN-panelen.
Om vi inte inser behovet av detta kommer vi inte att få en lösning, för det kan bara bli fred om det blir rättvisa; rättvisa är endast möjlig med sanningen som grund; och sanningen kommer bara fram om vi får en oberoende undersökning.
(EN) Herr talman! Sri Lanka har äntligen fått fred efter ett kvarts århundrade av terroristuppror och FN-rapporten om Sri Lankas armés seger över de tamilska tigrarna är full av kritik men innehåller få väsentliga bevisade fakta.
Den strategi man valt i rapporten förefaller att undergräva de ansträngningar som nu görs av Sri Lankas regering för att främja sanning och förståelse, inte minst genom kommissionen för dragande av lärdomar och åstadkommande av försoning (LLRC), och att regeringen faktiskt har släppt mer än 200 000 internerade tamilska fångar.
Naturligtvis måste alla avsiktliga illgärningar mot civila av militären straffas.
Jag håller med om det, men det finns inga klara bevis på att detta var en avsiktlig regeringspolitik.
Jag skulle vilja påminna kammaren om att LTTE vägrade ett övervakat internationellt erbjudande om kapitulation och i stället föredrog att välja blodbad som sin exitstrategi, vilket var skrämmande.
Konsekvenserna nu av det internationella samfundets ambivalens gentemot Sri Lanka är tydliga: minskat inflytande och en oförmåga att forma en utveckling.
Under tiden har Kina ryckt in och blivit Sri Lankas närmaste vän och försvarare i FN.
Jag behöver knappast påminna kollegerna i kammaren om Kinas inställning till de mänskliga rättigheterna.
Herr talman! Den 25 april 2011 offentliggjorde FN den rådgivande rapporten från den expertpanel som utsetts av FN:s generalsekreterare om ansvar i samband med den väpnade konflikten i Sri Lanka.
Panelen fann trovärdiga anklagelser som om de kunde bevisas skulle vittna om att allvarliga brott mot internationell humanitär rätt och de mänskliga rättigheterna hade begåtts av Sri Lankas militär och LTTE, av vilka några skulle innebära krigsbrott och brott mot mänskligheten.
Panelen ger också en rad rekommendationer till FN:s generalsekreterare och Sri Lankas regering, vilka med panelens ord skulle kunna tjäna som ram för ett pågående och konstruktivt samtal mellan generalsekreteraren och Sri Lankas regering om ansvarsskyldighet.
Rekommendationerna innebär att Sri Lankas regering inleder reella undersökningar och att generalsekreteraren inrättar en oberoende internationell mekanism.
FN har fastslagit att FN:s generalsekreterare noggrant granskar rapporterna, slutsatserna och rekommendationerna och FN:s högkommissarie för mänskliga rättigheter har uppmanat Sri Lankas regering att snabbt vidta de åtgärder som föreslås av panelen och säkerställa rättvisa.
Sri Lankas regering har å sin sida förkastat rapporten i starkaste ordalag.
Tidigare i veckan publicerade den höga representanten Catherine Ashton ett uttalande på EU:s vägnar som återupprepade EU:s åsikt att en oberoende process för att ta itu med dessa ytterst allvarliga anklagelser borde bidra till att stärka försoningsprocessen och trygga varaktig fred och säkerhet i Sri Lanka.
Den höga representanten har betonat att frågan om ansvarsskyldighet bör ses som en väsentlig del av den nationella försoningsprocessen.
EU hoppas därför att Sri Lankas regering ska värdesätta rapportens konstruktiva mål och uppmanar den att inleda samtal med FN:s generalsekreterare om dess innehåll.
Debatten är härmed avslutad.
Omröstningen kommer strax att äga rum.
Skriftliga röstförklaringar (artikel 149)
Konflikten mellan Sri Lankas regering och Tamilska befrielsetigrarna (LTTE) upphörde i maj 2009 och resulterade i mer än 90 000 dödsfall.
Flera lankeser som hade varit tvungna att flytta på grund av våldet i sitt land har återvänt till sina hem efter våldshandlingarnas slut.
Det finns emellertid fortfarande 75 000 flyktingar som fortsätter att tillbringa ett hårt liv i läger i Tamil Nadu, Indien.
Sri Lanka ställs inför en dubbel utmaning.
Landet måste återhämta sig efter en långvarig kris.
FN:s expertrapport, som offentliggjordes den 25 april, fann anklagelserna om brott mot internationell humanitär rätt och de mänskliga rättigheterna trovärdiga.
I rättvisans och försoningens intresse i Sri Lanka är det nödvändigt att starta en opartisk, öppen och oberoende utredning.
Sri Lanka måste också förbereda sig för olika naturkatastrofer, såsom översvämningar, jordskred, cykloner och också torka vilka landet är utsatt för.
Undertecknande av rättsakter som antagits i enlighet med det ordinarie lagstiftningsförfarandet: se protokollet
Meddelande från ordförandeskapet
Mina damer och herrar!
Jag vill meddela följande: På grund av den utrymningsövning som genomfördes under omröstningen i dag kommer vi att höra alla röstförklaringar som sammanhänger med dagens omröstning i morgon, tillsammans med morgondagens röstförklaringar.
I morgon genomför vi också de omröstningar som skulle ha genomförts i dag, men inte kunde genomföras.
Det gäller också den omröstning som pågick när vi fick avbryta. Vi kommer att fortsätta från exakt samma punkt som vi hade kommit till, så att vi har en fullständig kontinuitet.
Välkomsthälsning
Jag har just fått veta att FN:s undergeneralsekreterare Muhammad Shaaban befinner sig på besöksläktaren.
Jag vill välkomna företrädaren för FN.
En ny flerårig budgetram för ett konkurrenskraftigt och hållbart Europa för alla (fortsättning på debatten)
Vi fortsätter nu med debatten om betänkandet av Salvador Garriga Polledo om en ny flerårig budgetram för ett konkurrenskraftigt och hållbart Europa för alla.
(FR) Herr talman! Salvador Garriga Polledos betänkande är en ambitiös, framåtblickande sammanfattning, och jag tackar honom och gratulerar honom till hans arbete.
Hans betänkande innehåller krav på ökade medel för att unionen bättre ska kunna genomföra sina målsättningar enligt Lissabonfördraget.
Med kraft väcks frågan om egna medel och därmed också frågan om huruvida vår institution är fri i sitt grundläggande politiska agerande när den röstar om sin budget.
Det föreslås att gemensamma politikområden ska utökas och utvidgas, framför allt sammanhållningspolitiken, som i det förflutna i hög grad bidragit till att göra EU till en modell för samarbete och förståelse mellan folk, och som kan fortsätta att göra det i framtiden.
Med den kommande fleråriga budgetramen kommer sammanhållningspolitiken, enligt Europaparlamentets mening, att kunna gå in i en ny fas genom att en mellankategori skapas för regionerna.
Vi föreslår alltså ett nytt paket för denna fond, som stärker de lika möjligheterna för alla våra europeiska territorier, oavsett deras ekonomiska förflutna, oavsett deras handikapp jämfört med mer utvecklade regioner och oavsett hur sårbara de är för den ekonomiska kris som vi just nu upplever eller en kris som vi kan komma att ställas inför i framtiden.
Sammanhållning mellan EU:s olika territorier är ett centralt, strategiskt mål som EU:s hela framtid är beroende av.
De förslag som lagts fram är steg i rätt riktning, och om de följs av handling kommer goda grunder att läggas för framtiden.
Omröstningen om Salvador Garriga Polledos betänkande blir ett enkelt val - det handlar om att välja ett Europa som går framåt, ett val som görs av dem som bortser från politisk tillhörighet och tror på Europas framtid.
(PT) Herr talman! I denna tid av allvarlig ekonomisk kris i euroområdet, till följd av nyliberal politik och bristande solidaritet och ekonomisk och social sammanhållning, är det oacceptabelt att man inte förespråkar ett avståndstagande från och en förändring av EU:s politik och dess finansiella resurser.
När vi genomgår en ekonomisk och social kris är en av våra största utmaningar att komma fram till en ny flerårig budgetram där EU-budgeten för ekonomisk och social sammanhållning ökas avsevärt, samtidigt som de obligatoriska nationella bidragen minskas till som mest 10 procent av vad som föreslås, särskilt för länderna med de största ekonomiska svårigheterna. Det måste vara en ram som innefattar ett åtagande om investeringar, om offentliga tjänster, om produktionsstöd, om skapande av arbete med rättigheter och om utrotning av fattigdom, sociala orättvisor och all slags diskriminering, särskilt på grund av kön.
Vi måste också främja fred, samarbete och utvecklingsstöd och kraftigt dra ned på utgifterna för militären och utlandsrepresentationen.
Av alla dessa skäl anser vi att detta betänkande inte alls är vad som behövs för en bättre, rättvisare framtid för EU och dess medborgare.
Mina damer och herrar! När jag tar över ordförandeskapet för det här sammanträdet förstår ni säkert alla att jag vill uttrycka min sorg och bestörtning över Jorge Semprúns bortgång för några timmar sedan, vid 87 års ålder.
Vi hyllar Jorge Semprún som en person som satt fängslad i koncentrations- och utrotningslägret Buchenwald och som kämpade mot nazisternas styrkor i Frankrike och mot Francos diktatur i mitt land Spanien.
Vi hyllar också den framstående politiskt engagerade författaren, som bl.a. medverkade i vårt program för det europeiska bokpriset, och den övertygade Europavänliga politikern.
Jag sörjer hans död både som kollega och som vän, och jag tänker be talman Jerzy Buzek att sända hans familj och den spanska regeringen ett budskap om uppriktigt deltagande och stöd, som jag är säker på att alla här står bakom.
(Applåder)
(IT) Herr talman! Det är ingen tvekan om att vi står inför ett av de mest kritiska ögonblicken i EU:s ekonomiska historia.
Just av det skälet har det utskott som vi lyckats inrätta under detta år definitivt haft en väsentlig roll.
Vi har inga förutfattade meningar mot en ökning av budgeten, men vi anser att vi måste undersöka var nedskärningar kan göras.
Det står klart att vi måste skära i EU-budgeten, för det händer tyvärr att EU-medel inte används på rätt sätt.
Och kanske är det just det sätt på vilket dessa medel används som gör att många EU-medborgare inte längre är så övertygade om att EU är värdefullt.
För att nämna ett exempel vill vi fästa er uppmärksamhet på de medel som går till utvidgningspolitiken - ibland vet vi inte var de hamnar.
Vad kan sägas om de oändliga belopp som spenderas på integration och som åstadkommit så lite?
Vissa skötsamma regioner får heller inte tillgång till medlen, som sedan beviljas andra regioner som antingen inte utnyttjar dem alls eller utnyttjar dem på ett bristfälligt sätt eller för syften som inte är helt legitima.
Vi vill att denna fråga ska ägnas största möjliga uppmärksamhet och att åtgärder - även hårda sådana - ska vidtas så att EU kan återupprätta sin trovärdighet.
(NL) Herr talman! Jag får givetvis begränsa mig till några grundläggande kommentarer.
För det första kan jag inte någonstans i betänkandet, trots dess omfattning, hitta ett enda seriöst försök att lägga fram förslag till strukturella besparingar, exempelvis avskaffande av vad som enligt min mening är fullständigt överflödiga EU-institutioner, t.ex. Europeiska ekonomiska och sociala kommittén, Regionkommittén och en hel del europeiska byråer av olika slag.
Inte heller har det gjorts något som helst försök att ställa frågan om huruvida det inte vore klokare av EU att begränsa sig till ett antal noggrant definierade kärnuppgifter.
Tvärtom.
För det andra bävar jag verkligen inför de upprepade förslagen om att EU bör införa sina egna skatter, eller utfärda europeiska statsobligationer, som förr eller senare måste återbetalas av någon.
I betänkandet antyds att åtgärder av det slaget inte skulle öka det totala skattetrycket på medborgarna, vilket givetvis är lögn och bedrägeri av värsta slag.
För övrigt skulle det ytterligare underminera det sista spår av tillsyn och kontroll som medlemsstaterna utövar över EU-institutionernas utgiftsdiarré.
Det är de viktigaste skälen till att jag verkligen inte kan stödja detta betänkande.
(RO) Herr talman! De utmaningar som EU står inför i dag kräver ett bestämt och konsekvent gensvar på EU-nivå.
Det gensvaret utgörs av 2020-strategin, ett instrument som skapats för att EU ska kunna återhämta sig och få tillbaka sin styrka.
I det betänkande som presenteras i dag placeras 2020-strategin i centrum för nästa fleråriga budgetram som är under utarbetande, tillsammans med den nya situation som är resultatet av de behörighets- och politikområden som föreskrivs i Lissabonfördraget.
Vid en tidpunkt när många medlemsstater står inför besvärliga skattemässiga justeringar måste EU-budgeten, varav 95 procent går till investeringar, ge ett mycket högt europeiskt mervärde.
I betänkandet krävs att två oerhört viktiga områden av EU-politiken - den gemensamma jordbrukspolitiken och sammanhållningspolitiken - ska ligga kvar på åtminstone dagens nivåer.
Anslagen inom dessa politikområden måste baseras på nya kriterier som säkrar ett korrekt utnyttjande av medlen för att åstadkomma största möjliga effektivitet och överensstämmelse med konvergens- och sammanhållningskriterier.
Transport- och energipolitiken måste stärkas.
Anslagen till forskning och utveckling, både på EU-nivå och på nationell nivå, måste bidra till framsteg inom all EU-politik.
Sjuårsperioden, den nya struktur som föreslås och ökad flexibilitet ger större trygghet när det gäller att genomföra och anpassa sig till förändrade prioriteringar.
För stabilitetens skull måste systemet med EU:s budgetmedel tas under nytt övervägande, så att dagens nationella bidrag ersätts med EU-medel.
Europeiska rådet antog nyligen ambitiösa mål för EU:s utveckling.
Rådet måste också godta att den femprocentiga budgetökning som föreslås i betänkandet är minimivillkoret för att dessa mål ska kunna nås.
Den kommande fleråriga budgetramen måste genomföras med hjälp av ett system för ekonomisk styrning som säkrar den finansiella stabilitet som krävs för genomförandet av EU-politiken.
Jag vill gratulera föredraganden Salvador Garriga Polledo.
(ES) Herr talman! Jag vill inleda mitt anförande med att berömma det arbete som utförts av föredraganden och alla ledamöter i det särskilda utskottet för de politiska utmaningarna och budgetmedlen för en hållbar Europeisk union efter 2013.
Framför allt måste jag berömma deras beslutsamhet under det gångna året att sträva efter att nå en majoritetsöverenskommelse och majoritetsstöd i parlamentet för ett betänkande som det som läggs fram i dag.
Betänkandet är den färdplan som EU måste följa om vi vill nå de politiska, ekonomiska och sociala mål vi har satt upp, och också om vi vill klara de utmaningar vi kommer att ställas inför under kommande år.
Det här är det manus vi måste följa för att ta oss ur krisen och se till att vår tillväxt är intelligent, hållbar och integrerad, såsom anges i Europa 2020-strategin.
Om vi håller med om att EU:s värde är mycket större än summan av de 27 medlemsstater det innefattar, om vi vill ha ett ansvarsfullt jordbruk av hög kvalitet, om vi vill nå millennieutvecklingsmålen, om vi vill hjälpa våra grannar i Medelhavsområdet med deras övergång till demokrati, om vi vill fortsätta att satsa på forskning och innovation, om vi vill fortsätta att bekämpa klimatförändringar och satsa på utbildning och Erasmusstipendier, om vi fortfarande tror på sammanhållningspolitiken som ett verktyg för hållbar utveckling och solidaritet mellan våra länder, och om vi fortfarande stöder t.ex. transeuropeiska energi- och transportnät - kort sagt, om vi vill ha mer Europa - då måste vi kräva en större budget för EU.
Därför varnar vi i detta betänkande för att vi utan tillräckliga medel inte kommer att kunna nå de mål vi har satt upp.
Vi vet att en del rådsmedlemmar inte vill öka budgeten - det har vi sett här.
Det har de inte velat under konjunkturuppgångar heller.
Nu säger de att det beror på krisen, men de ville ha nedskärningar även under förhandlingarna om den gällande budgetramen.
Det är därför vi ber rådet att, om det inte vill ha denna budgetökning, tala om för oss vilka mål det vill att vi inte ska nå.
I det här betänkandet beskriver vi inte bara den politik vi vill föra på olika områden.
Vi visar också hur den ska finansieras, och vi för en diskussion om egna medel.
Den diskussionen, som syftar till att få slut på den falska debatten om nettobetalare, handlar om att få till stånd finansiering utan allmosor och utan undantag - finansiering som är rättvis.
Vi har lagt fram flera förslag om hur det ska gå till, men jag föredrar ett av dem, och Janusz Lewandowski vet mycket väl vilket det är: skatten på finansiella transaktioner eller Robin Hood-skatten, som den kallas i många av våra länder.
En sådan skatt skulle göra det möjligt att få in mellan 200 och 300 miljarder euro.
Det är en skatt som bestraffar spekulanter och skulle tvinga alla som har skott sig på att spela hasard med våra pengar att betala.
Det är en skatt som skulle öka öppenheten och minska finansspekulationen och, framför allt, en skatt som inte skulle drabba medborgarna, eftersom den skulle tvinga dem som direkt bär ansvar för krisen att betala för sina utsvävningar.
Det är egentligen bara en sak vi ber er om: att sikta högre.
Vi ber er att sikta högre för att se till att det europeiska projektet kan gå vidare och inte kör fast, för det skulle kosta oss vår framtid.
(DE) Herr talman! Jag föddes i EU 1975, och det har präglat mitt politiska liv.
Därför smärtar det mig desto mer att tvingas leverera en kalldusch i denna fråga.
När det talas om ökningar måste diskussionerna leda till ett övervägande kring det korrekta utnyttjandet av medlen.
Betänkandet är visserligen ambitiöst i sin strävan att få stöd från en så stor majoritet som möjligt i parlamentet, men jag anser att det i sin nuvarande form saknar ambitioner när det gäller de mål och syften som eftersträvas.
Jordbruks- och strukturbudgetarna lämnas orörda.
Man vill däremot ha mer pengar till forskning och utveckling.
Den enda lösning som parlamentet kan komma på är mer pengar, vilket också framgår av betänkandet, men det anges inte tydligt var pengarna ska komma från.
Vi hör tal om unionens ”egna medel”, men det har inte definierats vad det egentligen rör sig om för medel.
Om folk verkligen på allvar ville ha strukturreformer kunde de t.ex. ha anammat förslaget från David Cameron om att gå till rådet och säga: Finansieringen ska frysas, men vi kräver att outnyttjade medel ska kunna överföras till nästa budgetår, så att vi kan fortsätta att spendera dem på livskraftiga projekt och spara pengar.
EU:s livskraft i framtiden bör inte mätas i decimaler.
I det avseendet är jag inte bara lite besviken på det här betänkandet.
(EN) Herr talman! I morse kom Joseph Daul rusande för att tala här i plenum om behovet av en större EU-budget, men han sprang så fort att han tappade andan och måste sluta tala.
Det åskådliggör på ett utmärkt sätt debatten om den fleråriga budgeten.
EU-budgeten är fastställd till omkring 1 procent av EU:s BNP, men kommissionen och parlamentet säger att det inte är tillräckligt och vill ha mer pengar.
Men EU kan inte göra slut på de pengar som finns; miljardtals euro i regionala sammanhållningsfonder går inte åt.
En del pengar måste betalas tillbaka till medlemsstaterna.
Så varför behöver ni mer pengar om ni inte kan göra slut på de pengar ni har?
Men så har vi några ”Pavlov” här i parlamentet: Martin Schulz, Joseph Daul och Guy Verhofstadt, som alla är frånvarande nu - de har försvunnit i stället för att vara här och tala om att inrikta budgeten på kvalitet i stället för kvantitet, exempelvis genom att begränsa regional- och sammanhållningsfonder till de fattigare medlemsstaterna och därmed spara 30 procent på dessa fonder, pengar som kan satsas på innovations- och framtidsorienterad politik.
Men jag är säker på att alla Pavlov i EU på nytt kommer att springa in i Europeiska rådets tegelvägg senare i år.
(FR) Herr talman! Som redan har sagts står det klart att de nationella budgetarna har svårigheter av olika skäl - både samma och olika skäl, men i samtliga fall förvärrade av krisen.
Budgetsituationen måste ses över i vart och ett av våra länder, oavsett hur regeringsmajoriteten ser ut.
Vi har två alternativ.
Det ena är att agera på egen hand och försöka få ihop utgifter och inkomster, varvid i vissa fall - enligt vad jag har hört - åtstramningar hyllas som ett självändamål och kännbara nedskärningar görs i de offentliga utgifterna och sociala förmånerna. Därigenom förvärras situationen för medborgarna.
Jag skulle förespråka det andra alternativet, nämligen att förena våra budgetansträngningar och se till att budgetsolidariteten fungerar genom att spela ut kortet med de egna medlen, främst genom en skatt på finansiella transaktioner.
Det är syftet med den budgetsamordning vi vill åstadkomma genom denna konventliknande konferens, ett förslag som vi lagt fram för rådet under förlikningsförfarandet och som vi har upprepat i detta betänkande.
Vi måste samarbeta - EU, nationella parlament och regeringar - för att komma fram till en gemensam hållning i utgifts- och budgetfrågor.
Vi kan inte både ha kvar kakan och äta upp den - vi kan inte göra nedskärningar och samtidigt satsa på infrastruktur.
Det går inte att bidra mindre men få mer.
Jag anser att denna konventliknande modell för dialog mellan regeringar, EU, nationella parlament och Europaparlamentet är det rätta sättet att på nytt bygga upp förtroendet för EU, både nu och på längre sikt.
(NL) Herr talman! Det här är ett mycket dåligt betänkande som förtjänar att omedelbart kastas i papperskorgen.
Just nu, när människor överallt står inför oerhört smärtsamma åtstramningsåtgärder, är det för galet för att vara sant att vi i EU föreslår att ännu mer pengar ska spenderas.
Tänk att vi agerar så när det skulle kunna se ut på ett helt annat sätt: inget mer slöseri med pengar, ingen finansiering till cykelbanor och crêperier i ett land som Nederländerna.
Vi bör koncentrera våra strukturfonder på de fattigaste länderna och bara på innovativa projekt av Europaomfattande betydelse i övriga medlemsstater.
Enligt betänkandet bör allt förbli som det är: mer pengar har begärts för Europeiska jordbruksfonden för landsbygdsutveckling, inga reformer av strukturfonderna har föreslagits, det finns inga konkreta förslag för ökad effektivitet.
Parlamentet borde skämmas, särskilt gruppen Alliansen liberaler och demokrater för Europa och Europeiska folkpartiets grupp (kristdemokrater).
Medan - märk väl - Mark Ruttes regering i Nederländerna lämnar de sjuka och funktionshindrade ute i kylan har samma grupper här i parlamentet ett glödande hål i fickorna.
Åtstramningsmästare hemma, storslösare i Bryssel.
Detta är skandal!
(IT) Herr talman, mina damer och herrar! Jag vill framhålla flera saker i detta viktiga betänkande, till att börja med EU:s inkomstsystem.
Vid det här laget står det klart att dagens mekanism har för många motsägelser, varav den mest kända är Storbritanniens korrigeringsmekanism.
Flera andra korrigeringar och kompensationer har därefter lagts till, vilket gör EU:s inkomstmekanism helt och hållet orättvis och allt annat än tydlig.
I det här skedet vore det bättre att övergå till ett direktinkomstsystem baserat uteslutande på medlemsstaternas bruttonationalprodukt, eller till en gemensam och enhetlig inkomstform, t.ex. mervärdesskatt.
EU-medborgarna får givetvis inte utsättas för ytterligare bördor, och EU bör inte heller ersätta medlemsstaternas skattepolitik, som måste förbli självständig och helt och hållet suverän på det här området.
I betänkandet fastställs olika prioriteringar, varav några är viktiga och andra mindre viktiga, men de är i samtliga fall mycket kostsamma.
Vi kan skaffa fram medel med hjälp av instrument som projektobligationer och euroobligationer, men de måste omfattas av oerhört stränga villkor så att det inte riskerar att uppstå ytterligare skulder, vilket vore farligt.
Som ledamöter av Europaparlamentet kan vi omedelbart bidra till att förbättra EU:s finanser.
Vi måste äntligen välja en enda plats för parlamentets arbete, vilket skulle ge besparingar på tiotals miljoner euro varje år.
Det här är inte demagogi utan bara ...
(Talmannen avbröt talaren.)
(EN) Herr talman! Guy Verhofstadts förlöjligande av den brittiska regeringen när han lät oss ta del av sin logik i frågan om varför Storbritannien bör överlåta mer pengar och mer makt till EU var ytterligare ett bevis för det uppenbara förakt som vissa här i kammaren känner för Storbritannien, dess nationella regering och dess medborgare.
Vad Guy Verhofstadt glömde att nämna är att det finns andra besparingar att göra för Storbritannien.
Företag som tvingas lägga 30 miljoner brittiska pund på att rätta sig efter EU-föreskrifter skulle kunna spara de pengarna genom att återta kontrollen från EU.
Brittiska fiskare skulle hemskt gärna vilja ha de 3,3 miljarder punden i sina fickor - värdet av den fångst som går förlorad när EU låter andra länder fiska på deras territorialvatten.
Janusz Lewandowski, du säger att EU-budgeten inte handlar om att duplicera en nationell budget.
Men den kan inte skiljas från medborgarnas verklighet.
I dag är det brittiska bidraget 6,4 miljarder brittiska pund, vilket stiger till över 10 miljarder brittiska pund om rabatten försvinner.
De pengarna kan bara fås fram genom högre skatter, nedskärningar i fråga om tjänster, skolor ...
(Talmannen avbröt talaren.)
(DE) Herr talman, mina damer och herrar! Vi måste ställa oss själva fem frågor:
För det första: Vilken budget behövs för 2020-strategin för tillväxt och sysselsättning?
För det andra: Vilken budget krävs i en valutaunion?
För det tredje: Vilka möjligheter har vi att göra besparingar?
För det fjärde: Vilken budget behövs för Europas förenta stater?
För det femte: Vilken roll ska Europa 2020-strategin spela?
Vill vi spela någon roll över huvud taget?
Vi i Europaparlamentet tar vårt ansvar på allvar.
Vi talar klarspråk.
I Österrike har vi ett talesätt: Om du inte betalar kommer orkestern inte att spela.
Vi vill nå våra mål, fullgöra våra skyldigheter, anta utmaningarna och hålla våra löften.
Fler funktioner, bättre konkurrenskraft, mer hållbar tillväxt, fler arbetstillfällen, mer forskning och ytterligare integration kan inte åstadkommas med mindre pengar och utan en finansiell översyn, utan en utvärdering av hur medel betalas ut i dag och utan egna medel.
Mer Europa kommer också att ge möjligheter till besparingar i medlemsstaterna.
Mer Europa kommer också att ge ökad effektivitet och är vår lösning med avseende på globaliseringen, framtiden och utlandsskulden.
Vad är det vi vill?
Vi vill inte frysa budgeten.
Den som försöker frysa budgeten kommer att skada EU och försämra vår förmåga att fullgöra våra skyldigheter gentemot medborgarna.
Vi vill införa en transaktionsskatt som utgör våra egna medel, anta utmaningarna och rätta oss efter fördraget i stället för att stoppa huvudet i sanden.
Det är vår strategi.
Låt oss sätta bollen i rullning och rösta för det här betänkandet.
(BG) Herr talman, herr kommissionsledamot, mina damer och herrar! Huvudtemat i Salvador Garriga Polledos betänkande är inte finanser utan politik.
Jag vill tacka honom och Jutta Haug, liksom alla kolleger i utskottet, för att de haft detta som sin huvudsakliga utgångspunkt under det arbete som pågått under hela året.
Ekonomiska medel är bara ett sätt att nå målen.
Politiken är det viktiga och det som måste betonas när nästa budgetram diskuteras.
Vi vet alla att det görs budgetnedskärningar i alla EU:s medlemsstater.
Det kommer att fortsätta under kommande år.
Nedskärningarna ingår i insatserna för att ta oss ur krisen.
Men vi får inte glömma att detta även har EU-aspekter: planen för ekonomisk utveckling, finansmarknadsregleringarna för att förhindra en ny kris, de åtgärder som för närvarande diskuteras när det gäller ekonomisk styrning i EU och EU-åtgärder som bara gör de nationella åtgärderna effektivare.
Därför är det olämpligt att nationella åtgärder som syftar till att åtgärda krisen och dess konsekvenser kolliderar med EU-åtgärder.
Att ingå i EU ger mervärde.
Mervärde och solidaritet är inte bara tomma ord.
Att förklara för nederländska skattebetalare att deras avgifter till EU ökar är inte detsamma som att förklara för bulgariska eller polska jordbrukare att det bidrag de får är tre gånger mindre och att de tvingas konkurrera på samma konkurrensutsatta marknad.
Det är inte lätt att rikta anklagelser mot grekiska skattebetalare, som genomgår en oerhört svår tid just nu därför att det europeiska finanssystemet fick en enorm summa pengar från Grekland för bara några år sedan.
Solidaritet har särskilda aspekter. De aspekterna hänger också samman med de prioriteringar som EU fastställt för de kommande åren.
Inget genombrott kan nås i fråga om forskning, energi, transport, ekonomisk styrning eller digital teknik om inte dessa sektorer får stöd av gemensam EU-politik.
Vi måste definitivt också överväga hur dagens EU-budget kan förändras.
Den innehåller ju reserver som måste begäras.
Men jag ska ge er ett exempel.
Reserverna kan inte ställas till förfogande genom att exempelvis all politik eller alla mål som rör energieffektivitet, transport och så vidare införlivas med sammanhållningspolitiken.
Att ta medel från befintliga program tillgodoser inte behovet av nya resurser om vi vill sätta upp nya mål för EU och om vi vill att den europeiska integrationen ska ge ett verkligt mervärde, även för skattebetalarna, som med rätta håller uppsikt över vartenda öre som går till EU-budgeten.
Därför måste vi också se EU-budgeten som en del av ett system, både för ekonomisk styrning och för förvaltning av den gemensamma valutan.
Minimiökningen på 5 procent, som ifrågasätts, är inte tillräcklig för att alla dessa frågor ska kunna lösas.
Därför måste vi också ställa frågor om europeiska projektobligationer, euroobligationer och andra finansieringsmetoder.
Herr talman! Jag måste säga att under alla mina år i det här parlamentet så är SURE-utskottets arbete det roligaste, det mest visionära, kort sagt det roligaste: det är roligt, det är vackert.
Allt det nödvändiga och allt det goda för Europas framtid finns med.
Dock är jag själv personligen oerhört oroad över det vi inte gjorde, och det är att göra prioriteringar.
Man har tagit till sig alla nya utmaningar, men man har också bibehållit allt det gamla.
Det kanske inte är möjligt att göra både och.
Vi borde ha prioriterat, vi borde ha prioriterat väldigt mycket hårdare, men det som är allra mest oroande i sammanhanget är att vi har överlåtit prioriteringarna åt ministerrådet.
Det är inget arv för framtiden, mina vänner.
(EN) Herr talman! Allmänheten, de hårt arbetande skattebetalare över hela Europa som faktiskt tjänar de pengar som så många här är så ivriga att få spendera, vill att EU ska göra mindre och göra det bättre.
De vill ha en liten EU-budget som tar hänsyn till att vi, oavsett vad vi tycker om det, lever i åtstramningstider.
De vill att EU ska fokusera på de mycket få områden där det faktiskt kan ge ett mervärde och lämna den övriga verksamheten till våra medlemsstater.
Tyvärr föreslås inget av detta i det här betänkandet.
Låt oss tala klarspråk: förslaget om en femprocentig ökning är fullständigt oacceptabelt, och detsamma gäller tanken på så kallade egna medel - det är bara ett försök från EU:s sida att få mer makt.
Budgeten bör moderniseras, och medel bör omfördelas till program som faktiskt ger fördelar i framtiden och inte syftar till att dölja tidigare misslyckanden.
Finansieringen av insatser för att rädda euron bör överlåtas till de länder som faktiskt ville ansluta sig till euron från början.
De av oss som varnade för att det var ett misstag bör inte tvingas att bidra.
Utskottet hade chansen att föra fram många av dessa konstruktiva och framtidssäkrade förslag, men man tog den inte.
Inget av detta har blivit av, och parlamentet bör förkasta betänkandet.
(HU) Herr talman! Det betänkande vi har framför oss är kanske det viktigaste under den här perioden.
Europaparlamentet är först av institutionerna att sammanställa sina tankar om de kommande sju åren, men utan att det påverkar kommissionens rätt att lägga fram förslag.
Det här är emellertid den enda möjligheten att undvika en skandal gällande vår rätt till samtycke som skulle tvinga oss att förkasta rådets förslag.
Alla våra partner vet alltså vad Europaparlamentet vill, och de kan ta intryck av det i möjligaste mån.
Jag vill rekommendera mina kolleger två dokument som är värda att läsa innan ni börjar tänka på ren kritik: Lissabonfördraget och själva betänkandet.
Stödet för egna medel är varken mer eller mindre än vad som föreskrivs i Lissabonfördraget.
Budskapet om att EU-budgeten behöver ökas en aning ser jag som mycket viktigt.
En aning betyder i det här sammanhanget att de 5 procent som föreslås även kommer att justeras för inflationen, vilket betyder att det inte är någon abnorm ökning vi talar om.
Det handlar inte om att utgifterna för jordbruk eller sammanhållning ska öka utan om att de inte får minska.
Miklós Zrínyi, en kroatisk-ungersk författare som levde på 1600-talet, sade - vid den tiden med avseende på turkarna - ”skada inte ungrarna!”.
Jag citerar honom och säger: Skada inte jordbrukspolitiken och skada inte sammanhållningspolitiken, för de som skadar dessa politikområden skadar inte bara ungrarna, rumänerna och slovakerna utan alla medborgare i de europeiska nationerna.
Ju mindre väljarstöd en politiker har, desto mer hänvisar han till medborgarna.
Jag menar att vi, som har stöd från en större politisk kraft, även företräder medborgarnas intressen, och det är därför vi säger: Skada inte jordbrukspolitiken och sammanhållningen!
(EN) Herr talman! Jag vill tacka föredraganden och ordföranden för deras arbete med det här betänkandet.
Det framgår av dagens debatt om betänkandet att det kommer att bli strid i rådet om ett antal frågor, bl.a. den generella ökningen, den brittiska rabatten och de egna medlen.
Ärligt talat tror jag att parlamentet har försökt komma fram till en del kompromisser, utom i frågan om den brittiska rabatten där ledamöterna från Storbritannien kommer att vara ensamma om sin åsikt.
I samband med långa, komplicerade och viktiga betänkanden som det här är det nästan oundvikligt med kompromisser, men jag välkomnar faktiskt en del av dem.
Jag välkomnar kompromissen om varaktigheten och strukturen för nästa budgetram.
Jag välkomnar också kompromissen om sammanhållningspolitiken.
Jag anser att sammanhållningspolitiken är nödvändig om vi ska lyckas få till stånd arbetstillfällen och tillväxt i EU efter 2013.
Därför behöver vi inför framtiden tillräcklig finansiering av sammanhållningspolitiken, åtminstone på samma nivå som i dag, om inte mer.
För att vara relevant för medborgarna måste nästa budgetram handla om sysselsättning och tillväxt.
Därför behöver vi, vid sidan av en stark sammanhållningspolitik, även strategier för finansiering av forskning och utveckling på våra universitet och i våra små och medelstora företag.
Åttonde ramprogrammet behöver därför tillräcklig finansiering för framtiden.
Vi måste också satsa på vår infrastruktur i EU - det gäller t.ex. transport, energi och bättre bredband i många landsbygdsområden - och vi får inte glömma just våra landsbygdsområden.
För att kunna genomföra alla dessa strategier för sysselsättning och tillväxt behöver vi genomförandemekanismer.
Dessutom behöver vi partner.
(Talmannen avbröt talaren.)
(FI) Herr talman, herr kommissionsledamot! Först och främst vill jag gratulera föredraganden till ett utmärkt betänkande och till hans utomordentliga arbete i det särskilda utskottet för de politiska utmaningarna och budgetmedlen för en hållbar Europeisk union efter 2013.
Ett av de främsta målen för framtida budgetramar är att införa instrument för att genomföra Europa 2020-strategin på gräsrotsnivå.
I detta betänkande finns en insikt om att det inte kommer att lyckas utan en sammanhållningspolitik och en jordbrukspolitik som är stabila och starka i budgethänseende.
Sammanhållningspolitiken, exempelvis, är inte det enda faktiska instrument som ger oss möjlighet att utveckla innovationer och skapa arbetstillfällen och tillväxt.
Reformer behövs, men vi kan också genomföra dem inom dessa politiska sektorer.
Jag vädjar därför till dig, Janusz Lewandowski, att se till att både regionalpolitiken och jordbrukspolitiken får behålla dagens budgetnivåer under den kommande budgetperioden, som parlamentet vill.
Det gläder mig dessutom att man i betänkandet också tar hänsyn till regioner där förhållandena är särskilt svåra, t.ex. de glesbefolkade områdena i norr.
De kommer också att behöva egna tilläggsbudgetar under den kommande budgetperioden.
(NL) Herr talman! Nyckelordet för EU är ”förtroende”.
EU-institutionerna i allmänhet, och Europaparlamentet i synnerhet, måste få tillbaka medborgarnas förtroende.
Hur kan det åstadkommas?
För det första, inte med mer Europa eller mer pengar för Europa, utan med ett bättre Europa, ett Europa med ett mervärde. EU bör inte lägga sig i frågor som idrott eller turism som medlemsstaterna mycket väl kan ta hand om själva.
För det andra, låt sammanhållningsfondens medel gå till de verkligt fattiga regionerna i EU.
Än i dag går 50 procent till rika medlemsstater som Tyskland och Frankrike.
Det är oacceptabelt.
Om vi får ordning på det här kommer vi att kunna tygla det onödiga slöseriet med pengar och fortfarande göra en nettovinst.
För det tredje, investeringar i framtidssäkrat jordbruk och industri.
Garriga Polledo-betänkandet blev ett misslyckande.
Allt och mer därtill har slängts i en stor gryta, och medborgarna förväntas smälta denna sörja.
Smaklig måltid, men se upp så ni inte sätter i halsen.
(PT) Herr talman, mina damer och herrar!
Jag vill gratulera föredraganden till hans utmärkta arbete, som har resulterat i ett betänkande som ger oss möjlighet till en bra start vid utformningen av en flerårig budgetram - en utmaning för kommissionen och rådet.
Det här är ett ambitiöst och samtidigt realistiskt betänkande.
Jag hoppas att alla institutioner har dragit rätt slutsatser av den finansiella, ekonomiska och sociala kris som bara långsamt släpper sitt grepp om oss.
En slutsats är tydlig för mig: bara ett enat EU som uppvisar solidaritet och en stärkt, harmoniserad och konsekvent ekonomisk styrning kan klara uppgiften att framgångsrikt möta de politiska utmaningar vi har framför oss.
Vi behöver mer och bättre Europa.
Vi måste prioritera unionsmetoden i stället för den mellanstatliga metoden.
Vi måste öka budgeten.
Vi har enats om Europa 2020-strategin; dess prioriteringar är tydliga och dess mål mätbara.
Den kommer att vara vägledande för kommande budgetramar.
Denna strategi kan dock bli framgångsrik bara om det finns en budget som motsvarar verksamheten inom dess ramar - dess målsättningar.
Den fleråriga budgetramen måste därför få den ekonomiska uppbackning som krävs för att nå upp till den ambition och det åtagande som präglar Europa 2020-strategin.
Sammanhållningspolitiken är också ett resultat av solidaritetsprincipen.
Det är viktigt att denna sammanhållning är ekonomisk, social och territoriell, och att den ger de fattigare regionerna ett uppsving.
Jag anser därför att det är väsentligt att finansieringen för sammanhållningspolitiken ligger kvar på åtminstone samma nivåer, vilket även gäller finansieringen för den gemensamma jordbrukspolitiken.
Det är också viktigt att gå mot en flerårig budgetram där mer än 80 procent av medlen inte kommer från nationella budgetar.
(HU) Herr talman! Krisen tvingar oss att se över både nationella budgetar och EU-budgetar i effektivitetshänseende och titta på hur de tjänar våra syften och hur stort mervärde, europeiskt mervärde, de bidrar med.
Jag vill tala om ett område som inte har nämnts hittills i dag, nämligen samarbetet i rättsliga och inrikes frågor, som genom Lissabonfördraget lyfts från medlemsstaternas behörighet till EU-nivå.
Vår önskan att åstadkomma stora förbättringar på det här området måste återspeglas under den kommande budgetperioden.
Vi måste definitivt tillhandahålla medel för Stockholmsprogrammet, som är ganska ambitiöst.
EU behöver välutbildade invandrare som kommer hit i enlighet med reglerna, och en gemensam migrationspolitik med tillräckliga resurser.
Händelserna i Nordafrika har på nytt fäst uppmärksamheten på vikten av en gemensam europeisk invandringspolitik och har visat behovet av integration som stöds med resurser, och behovet av europeisk solidaritet.
De senaste månaderna har det också blivit tydligt att försvaret av våra gemensamma värderingar, icke-diskriminering och mänskliga rättigheter också behöver skydd och resurser, och att vi måste förenkla utnyttjandet av medel för hantering av extraordinära situationer, samt att vi behöver egna medel för att skapa ett bättre, starkare och mer omfattande EU under den kommande perioden.
(EN) Herr talman! Jag vill gratulera föredraganden till allt hans arbete.
Det har varit oerhört omfattande sett till insatsen för att försöka nå samförstånd.
Det finns tre områden där jag skulle vilja se ändringar.
För det första behöver vi på längre sikt en femårig budgetram.
Om 2020 är ett sjuårsperspektiv bör vi ha som absolut villkor att nästa budgetram ska gälla en femårsperiod.
För det andra har inte tillräckligt mycket arbete ägnats åt att titta på hur vi får en revisionsförklaring för utgifterna.
De som förespråkar mer pengar på EU-nivå skulle ha bättre möjligheter att få gensvar om vi visste att vi kunde vara helt säkra på vart pengarna faktiskt går.
För att svara Guy Verhofstadt vill jag sist men inte minst säga att det är oklokt att peka ut en viss medlemsstat när ett antal medlemsstater är nettobetalare till budgeten.
Jag förespråkar starkt att vi sätter en gräns för medlemsstaternas nettobidrag i procent av BNP, för om vi ser framåt är det orealistiskt att tro att man kan få medlemsstaternas godkännande när deras nettobidrag fördubblas i tider av stora åtstramningar.
(DE) Herr talman! Den femprocentiga budgetökningen förklaras av utgifterna för Europeiska utrikestjänsten, gränsskydd, kriget mot terrorism, en ökning av utvecklingsbiståndet samt stöd för forskning och gränsöverskridande infrastruktur.
Generellt sett är denna begäran från parlamentet definitivt motiverad.
Men parlamentet går också miste om en möjlighet med Garriga Polledo-betänkandet.
Vi skulle kunna bli mer trovärdiga om vi visade var EU kan vara mer effektivt och var pengar kan sparas.
Här ingår definitivt det stora antalet byråer som för en oerhört kostsam självständig tillvaro, och jordbruket, där vissa medlemsstater ännu inte lyckats införa ett mer marknadsanpassat system för schablonmässigt beräknat hektarstöd.
Som föredragande för strukturpolitikens framtid vill jag också säga att även EU:s sammanhållningspolitik bör ingå här.
Många regioner har lyckligtvis kunnat överskrida finansieringströskeln på 75 procent.
Men om fattigdomen minskar i EU:s olika regioner kan den europeiska solidariteten också avta.
Sparade pengar skulle hellre kunna investeras i europeiskt mervärde, exempelvis i en smart koppling mellan strukturfonderna och gränsöverskridande nät i gränsregionerna.
Detta diskuteras för närvarande i utskottet för regional utveckling, tillsammans med ett förslag om en mellankategori på 75-90 procent av BNP, såsom föreslås i Garriga Polledo-betänkandet.
Constanze Angela Krehl kanske drömde om hon trodde att vi redan enats om en kompromiss i utskottet för regional utveckling.
Jag tycker inte att det tillfälliga särskilda utskottet för de politiska utmaningarna och budgetmedlen för en hållbar Europeisk union efter 2013 är det rätta forumet för rekommendationer om en sådan mellankategori.
Vi gör det för enkelt för oss om vi bara säger att även de rikare regionerna behöver särskilt stöd.
Som jag ser det är det är en uppmaning till slöseri med pengar.
Vi lämnar det beprövade in- och utfasningssystemet men erbjuder inte längre något incitament.
Vi garanterar ett permanent stöd till alla regioner upp till en nivå som nästan motsvarar genomsnittlig ekonomisk styrka.
Det kan inte finnas någon framtid för ett system som det här i EU:s regionalpolitik.
Vi måste därför stryka punkt 73 i betänkandet.
Annars kan det inte godtas.
(Talaren godtog att besvara en fråga (blått kort) i enlighet med artikel 149.8 i arbetsordningen.)
(DE) Herr talman, herr Pieper! Det förvånar mig att du, Markus Pieper, påstår att Constanze Angela Krehl drömmer.
En stor majoritet röstade för att införa mellankategorier när omröstningen ägde rum i utskottet för regional utveckling.
Jag anser att vi även här i parlamentet kommer att få stöd av majoriteten eftersom det finns ett majoritetsstöd för solidaritet mellan regionerna.
Därför behöver vi detta mål med mellankategorier.
Det vore intressant att få veta varför du kallar denna majoritet en dröm.
Markus Pieper, kan du förklara varför det är en dröm?
(DE) Herr talman, fru Schroedter! Där här är ditt sätt att uppfatta frågan.
Vi i utskottet för regional utveckling har ett annat förslag än det som ingår i Salvador Garriga Polledos betänkande.
Detta är min första punkt.
Min andra punkt är att det fortfarande finns ett stort grundläggande motstånd mot mellankategorin inom de politiska grupperingarna.
Du är säkert medveten om detta.
Därför är jag förvånad över din fråga.
Jag anser att du drömmer när du helt enkelt påstår att vi har föreslagit kompromisser och att de är entydiga.
I alla händelser är detta ett ärende som utskottet för regional utveckling ska förbereda för att debattera i plenum.
Jag är mycket förvånad över din synnerligen optimistiska uppfattning att vårt arbete är slutfört.
(FR) Herr talman! Debatten om EU:s kommande budgetram ger upphov till frågor om EU-projektet, om dess räckvidd och ambitioner.
Detta betänkande är berömvärt eftersom man strävar efter att mobilisera unionens budgetmedel för att uppfylla målen i Europa 2020-strategin.
Detta gör att betänkandet strider mot de flesta medlemsstaters snäva åsikter.
Under det att medlemsstaterna, när det gäller deras ekonomiska bidrag som de vill inskränka och de ekonomiska intäkterna som de vill ha mer av, betraktar EU utifrån sina finansiella bidrag, förordar man i detta betänkande en stark och integrerad unionspolitik, vare sig det handlar om en sedan länge genomförd politik eller nya befogenheter enligt Lissabonfördraget.
Följaktligen bör detta initiativbetänkande från parlamentet utgöra grunden för framtida diskussioner, även om man, enligt min åsikt, gör fel när det gäller samförstånd och försiktighet.
Visserligen vore en ökning av EU-budgeten på 5 procent bättre än medlemsstaternas budgetramar för 2012.
Men problemet - och antagligen stötestenen - är att komma överens om en siffra som överensstämmer med den politik som beskrivs i betänkandet.
Vi är medvetna om de negativa sidorna av åtstramningspolitiken: Att den påverkar sysselsättningen och att ett växande antal medborgare misströstar.
Vi har ett ansvar för att finansiera en kontracyklisk politik, inte minst genom en stark sammanhållningspolitik genom vilken man främjar offentliga investeringar och sysselsättning i alla EU-regioner.
Jag vill betona betydelsen av att skapa en mellankategori av regioner för att se till att tilldelningen av strukturfonder på ett korrekt sätt återspeglar de ekonomiska och sociala realiteterna i regionerna.
Avslutningsvis vill jag säga att vi måste införa en skatt på finansiella spekulationer, något som skulle öka våra medborgares stöd för ett välfinansierat EU.
(EN) Herr talman! Först och främst vill jag gratulera föredraganden till att ha belyst de många utmaningar som väntar oss.
Jag välkomnar också det mycket tydliga budskapet i betänkandet där man kräver en betydande ökning av forskning och vetenskap, eftersom det är en av de prioriteringar vi behöver.
Jag vill särskilt säga till kommissionen att politik och ledarskap handlar om prioriteringar.
Utan prioriteringar finns det inget ledarskap.
Det finns alltid uppgifter och utmaningar som är viktigare än andra.
Detta är fallet med EU:s budget, och det gäller också medlemsstaterna.
Vi måste öka anslagen till forskning och vetenskap ytterligare, men vi måste också öka anslagen till vetenskap och forskning vid finansieringen av regionerna.
Vi måste ta hänsyn till utvecklingen av jordbruksmarknaderna och minska utgifterna där.
Men vi måste komma ihåg att vi måste prioritera på alla nivåer, både på EU-nivå och i medlemsstaterna.
Jag måste säga att jag ogillar attacker mot EU eller Bryssel, men jag ogillar också attacker mot medlemsstaterna, eftersom man därigenom minskar betydelsen av de utgifter vi har i medlemsstaterna: sjukvård, social trygghet, pensioner och utbildning.
Detta är ingen konflikt mellan EU och medlemsstaterna.
Detta är en pågående kamp om ledarskap och prioriteringar.
Om vi inte uppställer dessa prioriteringar visar vi inte ledarskap.
Jag måste säga att om vi inte förstår den svåra situation som medlemsstaterna befinner sig i i dag förstår vi inte den verklighet EU-medborgarna befinner sig i.
Vi måste fastställa prioriteringar och inte lösa problem bara genom att öka budgetarna.
Därför vill jag be kommissionsledamoten att visa ledarskap och mod och att komma ihåg att forskning och vetenskap, infrastruktur ...
(Talmannen avbröt talaren.)
(IT) Herr talman, mina damer och herrar! Vi ska rösta om ett mycket viktigt strategiskt dokument där man tillhandahåller en fast referens för budgetramen efter 2013.
Det inleds med en begäran om samstämmighet mellan mål och instrument och mellan den nya roll som EU-institutionerna måste spela - mot bakgrund av Lissabonfördraget och den ekonomiska tillbakagången - och de medel som vi tillsammans beslutar att investera.
En sådan samstämmighet inbegriper också ett allvarligt svar på begäran om innovation från allmänheten, från mottagarna av EU-politiken och från EU:s sociala grupper och industrier.
Vi gjorde samma sak när det gällde sammanhållningen, som är en avgörande fråga för att besluta vad vi vill att EU ska vara under de kommande åren.
Erfarenheten visar att sammanhållning nu utgör en livsviktig och central del av EU-projektet och en viktig tillgång som alla måste värna, skydda och förnya.
I detta avseende är den ansträngning man gör för att införa en mellankategori av regioner särskilt viktig, framför allt därför att de år av ekonomisk tillbakagång som vi har kommit ut ur i flera fall har förstärkt de inre skiljaktigheterna, vilket ytterligare har ökat betydelsen av ett effektivt och tillräckligt stöd till de mindre utvecklade regionerna i EU genom att bekämpa slöseri och på allvar fokusera på utvecklingspolitiken.
Jag anser emellertid att vi måste anta utmaningen med mellankategorier och med en skyddsklausul för att inleda en ny fas i EU:s sammanhållningspolitik och för att inom sammanhållningspolitiken förverkliga den mer balanserade och hållbara utveckling som vi vill säkerställa för EU under de kommande åren.
(FR) Herr talman! De 500 miljonerna EU-medborgare utgör för närvarande över 8 procent av världens befolkning.
År 2050 kommer denna siffra att uppgå till 5 eller 6 procent.
År 2100 kommer vi att utgöra 3 procent av denna befolkning.
Denna mängd EU-medborgare fortsätter att, till största delen genom nationella budgetar, underhålla bl.a. 2 000 ambassader, 27 arméer och 50 gemensamma styrkor.
Jag tror att Kina för närvarande har anställt extra vice ministrar bara för att ta emot alla de mäktiga EU-ministrar som kommer för att hos regeringen i Peking anhålla om förmåner och bilaterala överenskommelser.
Allt detta börjar se löjeväckande ut på världsarenan.
Att fördela 8 procent av världens befolkning mellan 30 självständiga nationella budgetar är idiotiskt.
I grunden är denna självständighet fortfarande absolut.
EU förvaltar 2,5 procent eller en fyrtiondel av de totala budgetutgifterna i EU.
Medlemsstaternas bidrag utgör en fyrtiondel av deras nationella utgifter.
Ändå är detta tydligen för mycket.
Låt oss nu, eller kanske någon annan gång, överväga frågan om våra egna medel.
Låt oss sluta gnata om de 2,5 procent offentliga utgifter med vilka vi antas underhålla hela den apparat som krävs för att genomföra Europa 2020-strategin och fullgöra allt det ansvar vi har tilldelats enligt Lissabonfördraget.
Vi har inte utformat strategin och behörigheterna: Det har medlemsstaterna gjort.
Mot bakgrund av denna verklighet är Salvador Garriga Polledos betänkande anspråkslöst.
Ändå finns det de som vill inskränka det ytterligare och som anser att betänkandet är ambitiöst.
Därför bör parlamentet anta detta betänkande.
(FR) Herr talman, herr kommissionsledamot, mina damer och herrar! Detta betänkande är viktigt för EU-projektets framtid, ett projekt som skulle inbegripa solidaritet och ambitiösa mål, framför allt med tanke på den budgetkris som medlemsstaterna för närvarande kämpar med.
Genom att inta en ultraliberal strategi väljer de flesta stats- och regeringschefer i rådet att fortsätta att vilt skära ner budgetarna och är villiga att offra investeringar i sådana viktiga framåtsyftande politikområden som dem som finansieras genom EU-budgeten.
En frysning av budgeten kommer att innebära en försvagning av tillväxten, oavsett vad andra ledamöter kan säga.
En ökning på åtminstone 5 procent, vilket rekommenderas i detta samförståndsbetänkande, är ett minimum om vi vill ta itu med utmaningarna och stå enade.
I den europeiska solidariteten ingår behovet av att finansiera Europa 2020-strategin, inte minst dess sociala målsättningar, som inbegriper bekämpandet av fattigdomen.
Genom betänkandet har jag också blivit övertygad om att den europeiska solidariteten bör stärkas genom skapandet av mellanregioner som en garanti för att man genom sammanhållningspolitiken täcker hela EU på ett rättvist sätt.
Ytterligare ett exempel är slutligen Europeiska fonden för justering för globaliseringseffekter genom vilken man erbjuder verklig solidaritet för arbetstagarna i EU.
I betänkandet erkänner man den stora betydelsen av denna fond.
Ökningen av den fleråriga budgetramen är nödvändig.
Detta bör inte betraktas som en börda för medlemsstaterna eftersom man genom EU-budgeten får ett mervärde och eftersom den i framtiden kommer att inbegripa en skatt på finansiella transaktioner.
(EL) Genom Lissabonfördraget skapades nya behörighetsområden och EU-politiken förstärktes, vilket framgår av den nya fleråriga budgetramen för perioden 2013-2020.
Jag gratulerar föredraganden, Salvador Garriga Polledo, till detta integrerade betänkande där man fastställer de politiska prioriteringarna för ett EU som skiljer sig från det EU vi känner.
På grund av de stora inre utmaningar som unionen och EU-medborgarna står inför och med tanke på den ökade internationella karaktären av dessa utmaningar inser vi att det viktigaste målet för EU-politiken måste vara att minska de befintliga sociala, ekonomiska och territoriella ojämlikheterna.
En planerad och framgångsrik sammanhållningspolitik utgör i sig ett EU-mervärde och kommer säkert att bli till fördel för alla medlemsstater i unionen.
Det nya programmet och den nya sjuåriga budgetramen är grundade på åtgärder inom Europa 2020-strategin och är avsedda att hjälpa EU att återhämta sig från krisen genom att främja en smart, hållbar och övergripande tillväxt.
De fastställda politiska prioriteringarna och målsättningarna är avsedda att främja sysselsättningen, stärka innovation, forskning och tillväxt, ta itu med klimatförändringarna, förbättra utbildningsnivåerna och bekämpa fattigdomen jämsides med invandringspolitiken och att garantera medel för att utveckla otillgängliga områden och gränsområden.
EU-budgeten är den viktigaste mekanismen för att skapa solidaritet mellan medlemsstaterna och är ett kraftfullt verktyg för en reform genom vilken man skulle kunna mobilisera ytterligare privata och offentliga medel för att stödja investeringar som kommer att verka som en katalysator för den exponentiella effekten av EU-utbetalningarna.
EU-budgeten måste ökas och baseras på egna medel om vi vill ha ett starkt EU för medborgarna och mot resten av världen.
EU-budgeten är ett verktyg för global och integrerad utveckling vid en tid då medlemsstaterna inte ensamma kan ...
(Talmannen avbröt talaren.)
(FR) Herr talman, mina damer och herrar! Man säger ofta att krigets nerv är pengar.
Vi måste komma ihåg att pengar också är ryggraden i ett fredsprojekt som EU.
Om EU verkligen har för avsikt att genomföra en politik som står inskriven i fördragen, däribland den nya politik som ingår i Lissabonfördraget, behöver unionen finansiella medel för att förverkliga dessa mål.
Därför röstar jag för att vi inför egna medel och en skatt på finansiella transaktioner.
Den nödvändiga ökningen av EU-budgeten måste åtföljas av betydande besparingar genom att vi optimerar våra utgifter.
Låt oss t.ex. skapa en verklig gemensam utrikes- och säkerhetspolitik för att ge EU mer inflytande på världsarenan, men också för att använda de allmänna medlen på bästa sätt.
Salvador Garriga Polledos betänkande är viktigt, nästan en fullständig omarbetning: Där förordas en mycket stark politisk och finansiell ram för EU.
Dessutom får två mycket väsentliga europeiska politikområden sin vederbörliga plats.
När det gäller den gemensamma jordbrukspolitiken (GJP), som är avgörande för livsmedelssäkerheten och självförsörjningen, rekommenderar man i betänkandet att budgeten för detta område förnyas.
När det gäller sammanhållningspolitiken, det finansiella instrument som används för att skapa regional solidaritet och uppmuntra regional ekonomisk utveckling, föreslår man i betänkandet att stärka målsättningarna genom att införa en mellankategori av regioner så att regioner på samma utvecklingsnivå kan dra fördel ...
(Talmannen avbröt talaren.)
(EN) Herr talman! Jag vill säga några ord om behovet av att röra sig i riktning mot en reform med egna medel.
Jag anser att den dominerade rollen av BNI-baserade inkomster gör att ett beslut om EU-budgeten blir överpolitiserat och mindre effektivitetsorienterat.
Därigenom underlättas kraven på att frysa eller minska EU-utgifterna.
Det leder till den logik som kom till uttryck under förhandlingarna om 2011 års budget, dvs. att om vi skär ner våra nationella budgetar på grund av krisen bör vi tillämpa samma strategi för EU-budgeten.
Det är emellertid inte självklart att vi, med ytterligare egna medel som minskar beroendet av BNI, kan förvänta oss en revolution av EU:s förmåga att finansiera tillväxt och strukturförändringar.
Det finns alltid en risk att samma koalition som antar budgetbeslutet i rådet också kan anta samma beslut i Europaparlamentet.
Om vi värnar om EU bör vi avhålla oss från att reagera på finansministrarnas förväntningar och i stället närma oss medborgarnas förväntningar.
Framgången för en nationell politiker som återvänder hem från förhandlingar i Bryssel bör inte baseras på budskapet att regeringen kommer att betala mindre till EU-budgeten, utan t.ex. på budskapet att EU kommer att hjälpa småföretag att finansiera nyskapande projekt.
Det är uppenbart att sättet att finansiera EU-kostnader ska vara helt öppet.
Detta kunde vara lättare att uppnå med bara en skatt, men det är också möjligt att basera inkomsterna på en grupp av skatter som motsvarar kriterierna för öppenhet, rättvisa, synlighet, effektivitet och tillräcklig harmonisering.
(PT) Herr talman, herr kommissionsledamot! Jag vill börja med att gratulera föredraganden till hans utmärkta arbete.
Jag välkomnar att de prioriteringar som har lagts fram i detta betänkande är i linje med Europa 2020-strategin och att tillväxten därigenom får en central plats i EU-politiken.
Vi behöver mer EU och ett bättre.
Därför bör vi främja de områden som mest bidrar till konkurrenskraft, t.ex. forskning, innovation och energi.
Vi behöver därför i stor utsträckning öka finansieringen av vetenskap och innovation för att främja vetenskaplig expertis i hela EU.
Det är också viktigt att stärka det europeiska systemet för finansiering av forskning för att förverkliga målet att investera 3 procent av BNP.
Den nya budgeten bör också främja ökad energieffektivitet och stödja uppbyggnaden av framtida infrastruktur, framför allt energiinfrastruktur, och därigenom skapa de nödvändiga villkoren för att den europeiska industrin ska bli effektiv.
Vi måste öka industrins roll, framför allt den som bedrivs av små och medelstora företag, och därigenom bidra till att stärka EU:s ledande ställning i en globaliserad värld.
(IT) Herr talman! Jag vill gratulera föredraganden Salvador Garriga Polledo till hans utmärkta årslånga arbete som har fått ett brett politiskt stöd.
Jag välkomnar det budskap som man har lyckats framföra i detta betänkande: Lösningen på krisen är att hävda EU:s ställning som global aktör.
Den framtida budgetramen återspeglar de mål som har fastställts i Europa 2020-strategin och är fast förankrad i Lissabonfördraget.
Lämplig finansiering krävs emellertid för att EU-prioriteringarna ska bli trovärdiga.
För utveckling av infrastruktur för transport och industri, investeringar i forskning och utveckling, utbildning och ungdomspolitik måste man skapa ny stimulans genom EU:s framtida budgetar, samtidigt som de grundläggande pelare som utgörs av sammanhållnings- och jordbrukspolitiken bör fortsätta att ta emot nuvarande finansieringsbelopp.
EU och dess stora projekt är i konflikt med budgetåtstramningarna på nationell nivå, vilket innebär att större engagemang från den privata sektorn genom projektförbindelser eller offentliga-privata partnerskap är det bästa sättet att öka konkurrenskraften och tillväxten.
I likhet med den övriga italienska delegationen är jag oroad över förslagen att även föra över dessa så kallade ”mellankategorier” till regionalpolitiken, eftersom man därigenom riskerar att skada de svagaste regionerna i EU.
Avslutningsvis försäkrar jag att det enda sättet att garantera EU:s framtid och utveckling är att finansiera unionen helt genom ett system som baseras på egna medel.
(DE) Herr talman, herr kommissionsledamot, mina damer och herrar! Reformen av tjänsteföreskrifterna kommer att läggas fram tillsammans med paketet för den fleråriga budgetramen.
Frågan om hur EU i själva verket förvaltas behandlas mycket kortfattat i punkterna 125 och 126 i Garriga Polledos betänkande.
Janusz Lewandowski, jag ber dig vara ambitiös när du lägger fram tjänsteföreskrifterna.
När allt kommer omkring är frågan om vad vi gör, som här har diskuterats i detalj, minst lika viktig som frågan om hur vi arbetar.
Frågan är vilken roll kommissionen kommer att spela i framtiden när den genomför alla punkterna i det program för 2020 som vi har lagt fram i dag.
Jag skulle vilja se att kommissionen väljer en starkare roll för sig själv i stället för att delegera alla uppgifter till andra.
Därför är det, i samband med reformen av tjänsteföreskrifterna, viktigt att det skapas lediga tjänster för dessa nya uppgifter så att också kommissionen själv kan engageras.
Vi har ett mycket stort antal lediga dagar.
Kommissionens tjänstemän har upp till 13 veckors betald ledighet.
Janusz Lewandowski, jag föreslår att du tar några av dessa lediga dagar och omfördelar dem till genomförandet av budgeten så att vi verkligen kan uppnå de politiska mål vi har föresatt oss.
Jag ber att vi också förses med en Europa 2020-strategi för förvaltningen av EU.
Detta skulle kräva åtgärder inte bara av dig utan också av hela kollegiet och av kommissionens ordförande.
(PL) Herr talman! Jag vill gratulera Salvador Garriga Polledo till att ha utarbetat ett utmärkt betänkande om den fleråriga budgetramen.
Betänkandet fick ett mycket starkt stöd i det särskilda utskottet för de politiska utmaningarna och budgetmedlen för en hållbar Europeisk union efter 2013.
Jag hoppas att betänkandet kommer att tjäna som en viktig grund för de förhandlingar om den nya fleråriga EU-budgeten som kommer att inledas inom kort.
Det gläder mig mycket att parlamentsledamöterna har beslutat stödja det ändringsförslag jag lade fram om att stärka ungdomspolitiken.
Vid en tid då unga EU-medborgare är bland de största offren för den ekonomiska krisen bör vi stödja alla initiativ som syftar till att förbättra situationen för ungdomar och framför allt dem som syftar till att förbättra tillgången på utbildning och ungdomarnas yrkessituation.
Program som ”Aktiv ungdom” och ”Livslångt lärande”, som kostar mycket lite per förmånstagare och är mycket effektiva, bör därför behållas som en separat del av framtida fleråriga budgetramar. Dessa program förtjänar också betydligt mer finansiering.
Samtidigt rekommenderar jag förslaget att behålla en hög finansieringsnivå för sammanhållningspolitiken.
Sammanhållningspolitiken spelar inte bara en viktig roll för att uppnå målen i Europa 2020-strategin. Dess huvuduppgift är att stärka den europeiska integrationen och solidariteten genom att minska de sociala, ekonomiska och territoriella skillnader som tyvärr fortfarande finns inom EU.
(RO) Herr talman! Föredraganden inledde sin presentation med ett mycket viktigt påpekande genom att säga att vi måste förena den traditionella EU-politiken med våra nya prioriteringar.
Ingendera kan verka utan den andra.
I detta sammanhang välkomnar jag den syn på den gemensamma jordbrukspolitiken som framgår av betänkandet.
Låt mig påminna er om några viktiga idéer, av vilka den viktigaste är att behålla nivån för budgeten för den gemensamma jordbrukspolitiken under den kommande budgetperioden.
Det europeiska jordbrukets traditionella roll, tillsammans de nya målsättningar vi har satt upp, gör att det är helt berättigat att behålla nivån för denna budget.
För det andra är behovet att behålla ett system för den gemensamma jordbrukspolitiken (GJP) baserat på två pelare, samtidigt som vi främjar landsbygdsområdena som en del av den andra pelaren, ett behov som är nära knutet till målen med Europa 2020-strategin.
Den sista punkten gäller behovet av en framtida reformerad gemensam jordbrukspolitik, där man syftar till att använda budgeten på ett effektivare sätt, baserat på en rättvis fördelning av utbetalningarna som ett av alternativen för att uppnå denna politik.
(LT) Herr talman! Först av allt vill jag tacka alla föredragandena för det enastående arbete de har utfört.
I dag har vi en tydlig ståndpunkt i parlamentet om vad vi och våra medborgare väntar oss av den kommande budgetperioden.
Vi förstår alla att vi kommer att bli tvungna att i grunden ändra inriktningen av den nuvarande politiken, och detta avspeglas tydligt i Europa 2020-strategin.
Vi måste utveckla en säker gemensam europeisk energimarknad, se till att hela EU är sammankopplat genom transportnät och utrota de återstående skillnaderna mellan de olika EU-regionerna.
Vi måste göra en fullständig översyn av den gemensamma jordbrukspolitiken som gör att man kan garantera ett enhetligt system med direktutbetalningar, utan vilket vi inte kommer att kunna skapa ett konkurrenskraftligt och starkt EU.
Detta kommer naturligtvis att kräva stora investeringar, framför allt inom forskningen.
Därför är det nödvändigt att söka efter nya finansiella instrument, t.ex. att införa en skatt på finansiella transaktioner.
Jag anser att ...
(Talmannen avbröt talaren.)
(NL) Herr talman! En av de viktigaste frågorna som har kommit upp under den här debatten är följande: ”Vad är egentligen europeiskt mervärde?”
Jag hoppas att kommissionen, när den i slutet av denna månad lägger fram sina förslag, kommer att ge en tydlig förklaring till varför vissa budgetrubriker har ett klart mervärde.
Enligt min uppfattning är det exakt detta vi behöver få veta, eftersom vi då kommer att kunna motivera vad vi röstar om.
För det andra kommer debatten också att i hög grad påverkas av debatterna om EU:s egna medel.
En av de frågor som har förgiftat debatten är beslutet om den brittiska rabatten som fattades 1984.
Hur har detta kunnat fortsätta så här länge?
Jag anser att den brittiska regeringen antingen inte bör vara berättigad till någon rabatt över huvud taget eller att andra länder, som befinner sig i samma situation som Storbritannien 1984, bör behandlas lika.
Jag hoppas att kommissionen kommer att lägga fram ett förslag i denna riktning.
(ES) Herr talman! Denna ständiga fokusering på den mängd nedskärningar som ska göras och inte på hur eller vad man ska skära ned, och ännu mindre på hur man ska öka inkomsterna, ger redan anledning till oro.
Först och främst betyder mer EU ett bättre EU, eftersom detta innebär mindre ekonomisk makt till medlemsstaterna.
För det andra måste vi naturligtvis också se över utgifterna.
Men vi måste vara noga med var vi ska göra detta: Ett förslag vore att minska de militära utgifterna.
Vi anser att detta är de viktigaste förslagen.
För det tredje blev jag mycket bekymrad över att se Janusz Lewandowski le på ett för mig oroande sätt när frågan om skatten på finansiella transaktioner nämndes.
Det oroade mig, och jag vill fråga honom hur det kunde vara så fel, så skadligt att be dem som har blivit rika genom att spekulera att betala för krisen, i stället för att be dem som bär den minsta skulden för denna situation att betala, och inte som du gjorde i går be Spanien att minska de sociala utgifterna genom att skära ned utgifterna för ...
(Talmannen avbröt talaren.)
Jag vill påminna mina kolleger om en sak. När vi godkänner budgeten måste vi komma ihåg att det bland EU-medborgarna finns en växande misstro mot vad vi gör här i parlamentet.
I detta hänseende anser jag att budgeten inte är tillräckligt samordnad med de ambitiösa målen i Europa 2020-programmet.
Jag har också en fråga: Du, kommissionsledamot Lewandowski, lovade de lettiska jordbrukarna att direktbetalningarna skulle jämnas ut med denna budget.
Men om budgeten godkänns i sin nuvarande form blir det svårt för dig att hålla ditt löfte.
Jag vill att allt vi talar om och allt vi diskuterar också ska motsvara våra väljares intressen.
(EN) Herr talman! Jag trodde inte att EU kunde bli värre förrän jag såg det här betänkandet.
Det börjar med en kraftig portion självbedrägeri: ”EU-medborgarna har aldrig förr ställt så höga krav på EU.”
Nåväl, ett ökande antal av det brittiska folket kräver att vi går ur unionen.
Detta är kanske vad de menar.
I betänkandet avfärdas helt tanken på att frysa budgeten efter 2013, och man insisterar på att till och med en ökning på 5 procent bara skulle möjliggöra ett begränsat bidrag till EU-målen.
Ja, vi måste vara tacksamma för små nådegåvor.
Undangömd i mitten av punkt 166 finns ett krav på att rabatterna ska upphöra.
Genom denna anordning betalar Storbritannien bara ett oacceptabelt nettobidrag i stället för ett skandalöst nettobidrag.
Att insistera på att Storbritannien ska betala ut sina surt förvärvade pengar är illa nog, men i punkt 169 föreslår man att EU ska ha makt att ta ut sina egna skatter utan vårt samtycke och utan vår kontroll.
Detta är helt enkelt oacceptabelt.
(PL) Herr talman! Vi har nått ett viktigt samförstånd.
Det betänkande som har lagts fram är en nödvändig fortsättning på det som har skett tidigare, samtidigt som man också föreslår de väntade ändringarna.
Stabilitet är ett karakteristiskt drag i EU-politiken, vilket förklarar förslaget att behålla den nuvarande budgeten för sammanhållningspolitiken och den gemensamma jordbrukspolitiken.
Genom att skapa lika villkor för utveckling bidrar man på ett betydande sätt till att stärka den gemensamma marknaden, vilket får positiva resultat för alla EU-medlemsstater.
Den gemensamma jordbrukspolitiken är till gagn för alla konsumenter i EU.
Det är värt att komma ihåg att jordbrukarna har mycket låga inkomster, trots det stöd de tar emot från EU-budgeten.
De nya uppgifter som jordbruket nu står inför när det gäller miljön, klimatet, djurens välbefinnande och orealistiska WTO-förhandlingar innebär ytterligare kostnader för jordbrukarna.
Vem ska betala?
De förändringar vi väntar oss inbegriper en ökning av finansieringen av en hållbar och intelligent utveckling och en tonvikt på innovation, forskning och utbildning.
(Talmannen avbröt talaren.)
(EL) Herr talman, herr kommissionsledamot! Parlamentet sänder i dag ut ett tydligt budskap, både till kommissionen och till EU:s premiärministrar, om en budget fram till 2020 som motsvarar unionens ansvar och allmänhetens förväntningar.
När det gäller sammanhållningspolitiken är budskapet tydligt. ”Ja” till en sammanhållningspolitik med tillräcklig finansiering för att lämna ett avgörande bidrag till utveckling, nya arbetstillfällen och innovation. ”Ja” till en oberoende sammanhållningspolitik. ”Ja” till samordning på alla nivåer av politiken, från strategisk planering till genomförande. ”Ja” till inrättandet av en mellankategori för stöd till regionerna. ”Ja” till särskilda åtgärder för öar och bergsområden i EU.
Det finns emellertid också två tydliga och viktiga ”nej”. ”Nej” till all uppsplittring av denna politik i olika sektorer, ”nej” till införandet av sanktioner i samband med stabilitets- och tillväxtpakten.
Härmed avslutas ögonkontaktsförfarandet, och jag ber de 11 eller 12 ledamöter som fanns på listan och inte har fått tala om ursäkt, men det finns uppenbarligen ingen tid för deras anföranden.
Jag har redan använt min talartid, och därför ska jag bara komma med två påpekanden.
För det första kan man inte, på grund av den nuvarande internationella krisen, klandra EU-budgeten, som inte har något underskott, för bristande förvaltning av de nationella finanserna.
EU-budgeten kan emellertid bidra till att skapa arbetstillfällen och tillväxt, eftersom den handlar om investeringar.
I detta avseende skiljer den sig från de nationella budgetarna, som huvudsakligen handlar om sociala transfereringar.
För det andra är successiv konvergens realistiskt när det gäller löftena till jordbrukarna i EU.
En enhetstaxa är inte genomförbar för tillfället, och jag anser att det kommer att fortsätta på detta sätt under de kommande åren.
På kommissionens vägnar väntar jag mig slutligen att man under den förestående omröstningen visar den breda enighet i parlamentet som kommer att göra Europaparlamentets röst stark och inflytelserik.
Vi kommer att avsluta denna debatt med ett anförande av föredraganden Salvador Garriga Polledo, som jag helhjärtat gratulerar till ett utmärkt arbete med denna fråga.
föredragande. - (ES) Herr talman! Jag vill först tacka de nationella delegationerna, som enligt vad jag förstår har stått emot påtryckningarna i sina medlemsstater och kommer att rösta för detta betänkande.
Jag anser att detta inte är en debatt om budgetvolym utan snarare om unionsmetodens överlägsenhet, och jag anser att de som har inriktat denna debatt på ansträngningar att minska EU-budgeten har gjort ett misstag.
De vill ha nya prioriteringar och en minskad budget. Jag säger till dem att denna väg leder till att de får en minskad budget och färre prioriteringar.
Jag förstår verkligen inte hur de kan sitta i denna plenisal och försvara en mellanstatlig strategi.
Låt rådet ta detta steg. Ni bör försvara EU med dess politik, dess prioriteringar, dess ansvar och en lämplig budget.
Vi vill inte ha någon ökning på 5 procent av de offentliga EU-utgifterna. I stället strävar vi efter att lindra de nationella budgetbördorna och samla vissa transnationella investeringar i EU-budgeten där de kan användas på ett effektivare sätt.
Detta är det europeiska mervärde som alla grupper i parlamentet i år accepterade i det särskilda utskottet för politiska utmaningar (SURE).
Jag anser att detta är ett mycket långtgående förslag. Det är ett ambitiöst förslag som innebär att man måste fatta viktiga beslut i medlemsstaterna, och vi vill be dem att möta den utmaning detta innebär.
Jag vill ge mitt erkännande till det konstruktiva i förslagen och i debatten, som enligt min mening har varit tillräckligt livlig, och där man till fullo har uttryckt de skilda åsikter som förenar Europaparlamentet.
Jag anser att vi i varje fall avslutar denna debatt med en mycket starkare ställning som parlament och med en mycket förbättrad politisk profil.
Debatten är härmed avslutad.
Omröstningen kommer att äga rum i dag kl. 12.00.
(Sammanträdet avbröts en stund.)
Skriftliga förklaringar (artikel 149 i arbetsordningen)
skriftlig. - (RO) På grund av den nuvarande krisen och de drastiska offentliga utgiftsrestriktionerna finner medlemsstaterna att det är allt svårare att notera någon ekonomisk tillväxt.
Jag måste betona att EU måste reagera på de demografiska utmaningarna.
Den minskade andelen av den arbetande befolkningen i kombination med det ökade antalet pensionerade kommer att innebära en påfrestning för de sociala trygghetssystemen.
Jag stöder tanken på att den finansiering som tillhandahålls av EU ska bidra till att förbättra det allmänna tillståndet för miljön i EU.
Därför bör de positiva och negativa inverkningarna på klimatet och miljön och användningen av EU-medlen analyseras på varje nivå.
Genom investeringar på EU-nivå kan man uppnå avsevärt större besparingar på nationell nivå, framför allt inom områden där EU otvivelaktigt ger större mervärde än de nationella budgetarna.
skriftlig. - (FR) I Salvador Garriga Polledos betänkande definieras Europaparlamentets politiska prioriteringar för den fleråriga budgetramen för perioden efter 2013, både när det gäller lagstiftning och budget.
Jag har särskilt noterat två saker: Först och främst att sammanhållning för tillväxt och sysselsättning är en politisk prioritering.
Jag stöder helt att man skapar en mellankategori av regioner.
Detta skulle gälla alla regioner där BNP per invånare ligger mellan 75 och 90 procent av BNP i EU.
Därigenom skulle man kunna skapa en bättre balans mellan regionerna.
Förslaget innebär ett genomförande av principen om territoriell sammanhållning enligt artikel 174 i fördraget om Europeiska unionens funktionssätt.
Vad gäller frågan om budgetramen är jag för en beskattning av finansiella transaktioner för att skapa egna medel för EU.
Jag vill fästa uppmärksamheten på förslaget om en EU-skatt på finansiella transaktioner i detta betänkande.
Genom en skatt på finansiella transaktioner skulle man samtidigt kunna hantera två problem - hur man finansierar de ständigt växande kraven på att genomföra ny EU-politik och hur man får finanssektorn att bidra till att lösa den ekonomiska kris som den har bidragit till.
Genom skatteintäkterna skulle man kunna minska de inbetalningar som EU-medlemsstaterna för närvarande gör till EU-budgeten.
Samtidigt möjliggör man därigenom en smidig utveckling av politiken för att trygga EU:s ekonomiska framtid.
Vi skulle få medel för investeringar i forskning och utveckling, för att bekämpa klimatförändringarna och för att skapa solidaritet mellan regionerna i EU.
EU bör vara världsledande genom att uppbära denna skatt inom sina gränser och genom att förespråka att den införs i resten av världen.
Jag uppmanar kommissionen att agera snabbt på detta betänkande och att uppfylla kraven från detta demokratiskt valda parlament att genomföra lämpliga åtgärder.
Under ekonomiskt svåra tider förväntar man sig mer än annars att EU ska komma med konkreta resultat.
Vi behöver bättre, enklare lagstiftning som tjänar EU-medborgarnas intressen.
Förordningarna bör skäras ned.
Vi ska inte skapa EU-lagar som inte är alldeles nödvändiga.
EU:s framtida budget bör svara mer effektivt på de vardagsproblem som vanligt folk står inför.
Budgeten bör stödja tillväxt och nya arbetstillfällen, men framför allt bör den tillföra europeiskt mervärde.
I slutet av den här månaden ska kommissionen offentliggöra förslaget till EU-budget efter 2014.
Genom den ekonomiska krisen har EU:s medlemsstater tvingats att fatta svåra beslut när det gäller de egna budgetarna.
I kristider borde EU-budgeten inte heller öka.
Tvärtom, den borde skäras ned.
Jag hoppas att vi äntligen ska lyckas avskaffa några av de rena dumheter som är förknippade med EU.
Parlamentets förflyttning mellan Bryssel och Strasbourg varje månad kostar EU:s skattebetalare drygt 200 miljoner euro varje år.
De pengarna kan användas bättre.
Rabatter som beviljats Storbritannien, Sverige, Österrike, Nederländerna och Tyskland borde avskaffas.
Bara Storbritannien kommer i år att få en rabatt på ca 3 miljarder euro tack vare en bidragsrabatt som förhandlades fram 1984.
Det är dags att reformera EU och dess budget.
De pengar som EU:s skattebetalare betalar måste användas mer effektivt och tillföra europeiskt mervärde till medlemsstaterna.
Att öka administrationen, byråkratin och onödig EU-lagstiftning ger inte något sådant mervärde.
Föredraganden skriver att EU-bidrag är nödvändiga för att medlemsstaterna ska kunna möta kommande utmaningar.
I Europa 2020-strategin pekar man ut områden dit bidragen bör riktas genom att sammanfatta prioriteringar och ge en vision av ett starkt, stabilt och modernt Europa, som har lärt sig läxan efter den senaste tidens ekonomiska problem och som kommer att garantera arbetstillfällen, en tryggad energiförsörjning och sunda livsmedel för medborgarna.
I budgetplanerna bör man ta hänsyn till de viktigaste målen för hållbar utveckling, samtidigt som budgetplanerna ska vara flexibla och inriktade på konkreta åtgärder.
Jag behöver bara nämna att pengar måste spenderas på ett sätt som medger insyn och på starka grunder.
Allmänhetens acceptans och förståelse är numera en oskiljaktig del av EU:s politik och är grunden för EU:s funktioner.
EU:s fattigaste regioner utvecklas just nu snabbt, och en av orsakerna är EU-finansiering.
Även om många vägar har byggts eller reparerats och internetanslutningar har installerats finns det fortfarande många behov att fylla, eftersom gapet är mycket stort mellan de mycket fattiga och de mycket högutvecklade regionerna.
När vi kom med i EU fick vi höra farhågor om att Polen och de nya medlemsstaterna inte skulle kunna utnyttja de möjligheter som de tilldelades genom medlemskapet, och att man skulle göra slut på EU-medlen utan tillräcklig eftertanke.
Vi fick också höra farhågor om korruption, eftersom tillfället gör tjuven - och här fanns det ju pengar.
Med tiden har analyser visat att EU-medlen har använts på ett mycket klokt sätt i Polen, utan kopplingar till ohederlig verksamhet.
Med tanke på de skillnader som vi försöker överbrygga och med tanke på EU:s målsättningar, kan vi inte minska varken EU-budgeten eller medlen för att genomföra sammanhållningspolitiken.
Men om Europaparlamentet röstar igenom en ökning av EU-budgeten, vilket jag hoppas inte blir fallet, blir det viktigt att övertyga de enskilda medlemsstaterna om att parlamentets politiska ståndpunkt är värd att stödja.
Jag vill uppriktigt gratulera Salvador Garriga Polledo till ett mycket innehållsrikt betänkande och för det imponerande arbete som han lagt ner på att utarbeta kompromissändringsförslag.
Jag instämmer med föredraganden om att sammanhållningspolitiken, som har visat sig vara effektiv, bör få en plats i den nya fleråriga budgetramen, som står i rimligt förhållande till dess betydelse.
Men beträffande enskilda fonder måste vi sträva efter bättre samordning och komplementaritet och efter förenklade förfaranden.
Förändringar i systemen för övervakning och hantering av medel, för att öka insatsernas effektivitet, bör baseras på en grundlig analys av hur de fungerar för närvarande.
Jag stöder också synpunkten att outnyttjade medel bör stå kvar i den budget som öronmärkts för sammanhållning och inte gå tillbaka till medlemsstaterna, och jag anser att vi behöver en grundlig analys av de eventuella konsekvenserna av att ta in Europeiska utvecklingsfonden i EU:s budget, särskilt med tanke på EU:s åtaganden gentemot tredjeländer.
Europa går igenom en kris.
Förlorade skatteintäkter från självstyrande regioner utgör mer än 20 procent av budgeten, jämfört med perioden före krisen.
Detta är ohållbart. Kommunernas inkomstunderskott ser ut på ungefär samma sätt: De kan inte finansiera sina kärnkompetenser, de friställer personal och de sätter sig i skuld.
I den situationen vore det inte särskilt förvånande om de inte kan förstå varför Europaparlamentet ber om ännu mer penningmedel.
Men om medlemsstaterna skulle samordna sin politik och sin finansiering inom prioritetsområden skulle de nå bättre resultat och spara mer pengar än den summa som vi vill få för att öka den gemensamma EU-budgeten.
Det finns alltså inget bättre alternativ än det som vi diskuterar just nu.
Vi måste diskutera och debattera det här ännu mer, inte bara i Europaparlamentet utan i synnerhet med ministrar i rådet, med medlemmar av nationella parlament och dessutom i regionerna, så att man inser att en gemensam lösning inte bara kommer att ge bäst resultat för medborgarna utan också kommer att leda till besparingar i de nationella budgetarna.
Parlamentet tagit ett viktigt steg framåt genom att anta Salvador Garriga Polledos betänkande: det är en tydlig, pragmatisk och realistisk redogörelse för Europaparlamentets budgetambitioner efter 2013, först och främst beträffande sammanhållningspolitiken, som är nyckeln till den regionala utvecklingen.
Jag anser att vi måste behålla budgeten för sammanhållningspolitiken och skapa en skälig biståndsmodell för alla regioner på mellaninkomstnivå så att framtida EU-investeringar i regionerna ska bli öppna och rättvisa.
Den 5-procentiga budgetökningen är rimlig.
Den är inte, som euroskeptikerna hävdar, ett exempel på EU-slöseri, utan ett modigt erkännande av att om vi inte tilldelar oss de här medlen för att tillsammans bygga Europa kommer vi att förbli isolerade och maktlösa.
För att kunna finansiera de åtgärder som hör samman med EU:s nya behörigheter under Lissabonfördraget stöder jag följaktligen begäran om att frågan om egna medel ska undersökas, och om nya former för gemenskapsinkomster, för att lätta trycket på de nationella budgetarna och för att göra slut på tron på en ”rättvis avkastning”, vilket är ekonomiskt felaktigt och politiskt ohållbart.
Europaparlamentet har för första gången framlagt sin vision om EU:s prioriteringar för perioden 2014-2020, för kommissionen och rådet.
Nu är det kommissionens tur att ta in parlamentets yttrande i sitt lagförslag.
Jag vill särskilt understryka att utveckling av en konkurrenskraftig jordbrukssektor samt ekonomisk och social sammanhållning bör förbli en prioritering för den kommande perioden.
Kollegerna har också uppmärksammat EU:s forskningsinsatser.
Europaparlaments hela vision är fast förankrad i Europa 2020-strategin.
När vi beslutar om ramen för nästa budget är min första fråga om vi vill ha ett svagare eller ett starkare Europa.
Enligt min mening har parlamentet redan tagit ställning i den frågan.
Vi har redan fastställt att vi behöver ett starkare Europa genom att godkänna de ambitiösa målen i Europa 2020-strategin.
Nu måste vi förklara högt och tydligt att målen bara kan uppnås om vi tilldelar dem tillräckliga resurser.
Under en period när många medlemsstater lider av ”medelhavsproblemet”, med länder som behöver finanspolitisk expansion för att stimulera tillväxt, men där detta inte är möjligt eftersom den oundvikliga följden skulle bli aldrig sinande åtstramningsåtgärder på grund av skuldsättning, kan vi inte reagera genom att minska eller godkänna den nu gällande EU-budgeten, vars grundläggande mål är utveckling.
Det går inte, eftersom det skulle betyda att eftersatta regioner berövas sin enda chans att leda in sina ekonomier på rätt spår mot tillväxt.
Att skapa ”genomsnittsregioner” såsom föreslås i betänkandet betyder att relativt rika områden i fattiga medlemsstater fortfarande skulle få stöd, och att de gradvis kan förbereda sig för den tidpunkt då de helt förlorar den här extra finansieringen.
Möjligheten att skapa en sådan grupp av regioner är utan tvekan en välkommen utveckling för sammanhållningspolitikens största stödmottagare, som måste planera på lång sikt.
Om parlamentet antar det här förslaget i dag skulle det skicka ut ett viktigt meddelande till debatten om sammanhållningspolitikens framtida utformning.
(DE) Herr talman! Jag ville bara säga att mikrofonen vid min pulpet, nummer 759, inte fungerar.
Jag bad redan i går om att få den att lagad.
Jag skulle behöva hjälp av en tekniker.
Tack.
Kolleger! Som ni vet blev omröstningen och röstförklaringarna uppskjutna i går på grund av brandövningen, så vi tar det i dag, som del av omröstningen.
De har lagts in i den ordning som finns på era omröstningslistor.
Bortfallna skriftliga förklaringar: se protokollet
14.
Tillämpningen av förfarandet vid alltför stora underskott (
Inkomna dokument: se protokollet
3.
Situationen i Syrien (
Undertecknande av rättsakter som antagits i enlighet med det ordinarie lagstiftningsförfarandet: se protokollet
Kommissionens åtgärder till följd av parlamentets åtgärder och resolutioner: se protokollet
Föredragningslista för nästa sammanträde: se protokollet
8.
Övervakningen av de offentliga finanserna samt övervakningen och samordningen av den ekonomiska politiken (
Muntliga frågor och skriftliga förklaringar (ingivande): se protokollet
5.
Alternativ tvistlösning i civil-, handels- och familjerättsliga ärenden (
Situationen i Egypten och Syrien, särskilt för kristna (ingivna resolutionsförslag): se protokollet
Inkomna dokument: se protokollet
9.
Demografiska förändringar och konsekvenserna av dessa för EU:s framtida sammanhållningspolitik (
Rättelser/avsiktsförklaringar till avgivna röster: se protokollet
(Posiedzenie zostało otwarte o godz.
15.00)
