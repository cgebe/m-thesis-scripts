SAMARBETSAVTAL mellan Rådet för arabisk ekonomisk enhet (CAEU) och Europeiska gemenskaperna (82/726/EKSG, EEG, Euratom)
RÅDET FÖR ARABISK EKONOMISK ENHET,
(nedan kallat Rådet), företrätt av dess generalsekreterare,
och
EUROPEISKA GEMENSKAPERNA,
företrädda av kommissionens ordförande,
SOM ÄR MEDVETNA OM att det finns ett behov av ett effektivt och positivt deltagande i utvecklingen och utbyggnaden av förbindelserna mellan organisationer som har kompetens på området för ekonomisk utveckling,
SOM ÖNSKAR göra sitt yttersta för att samordna sina åtgärder till gagn för båda parternas gemensamma intressen,
HAR ENATS OM FÖLJANDE.
Artikel I
Rådets generalsekretariat och Europeiska gemenskapernas kommission skall ställa undersökningar, dokument och information som är tillgängliga för spridning till varandras förfogande inom ramen för deras samarbete om frågor av gemensamt intresse.
Artikel II
Rådets generalsekretariat och Europeiska gemenskapernas kommission skall med lämpliga mellanrum sända experter som ställer sin sakkunskap och erfarenhet till förfogande och som deltar i seminarier av gemensamt intresse så att parterna kan dra ömsesidig nytta av sin respektive erfarenhet på praktiska områden.
Artikel III
Rådets generalsekreterare och Europeiska gemenskapernas kommission skall inbjuda varandra att delta i sammanträden som kan vara av särskilt intresse.
Artikel IV
Rådets generalsekretariat och Europeiska gemenskapernas kommission skall hålla varandra underrättade om pågående eller planerade program i frågor av gemensamt intresse.
Artikel V
Detta avtal är giltigt för en tid av fem år från och med dagen för undertecknandet och förnyas automatiskt för en motsvarande tid såvida inte en av parterna skriftligt uttrycker en önskan om att säga upp avtalet sex månader före dess utlöpande.
Artikel VI
Bestämmelserna i detta avtal får ändras eller revideras helt eller delvis efter gemensam överenskommelse mellan parterna.
Artikel VII
Detta avtal träder i kraft den dag det undertecknas av generalsekreteraren för Rådet för arabisk ekonomisk enhet och av ordföranden för Europeiska gemenskapernas kommission.
Artikel VIII
Detta avtal upprättas i två original på arabiska och engelska, vilka båda är lika giltiga.
SKRIFTVÄXLING mellan Europarådet och Europeiska gemenskapen om befästande och utvidgning av samarbetet (87/476/EEG)
A. Brev från Europarådet
Strasbourg den 16 juni 1987
Ministerkommittén har i sin resolution (85) 5 om samarbete mellan Europarådet och Europeiska gemenskapen, som antogs den 25 april 1985 på dess sammanträde, förklarat att den är övertygad om att den europeiska solidariteten kommer att stärkas genom befästande och utvidgning av samarbetet mellan Europarådet och Europeiska gemenskapen, vilka är det europeiska samfundets väsentligaste organisationer. Den uttryckte sin fasta vilja att med hänsyn till organisationernas särprägel och skilda förfaranden främja ett närmare samarbete mellan dem för att således verka för bredast möjliga samarbete på europeiskt plan.
I denna anda har ministerkommittén uppdragit åt mig att inleda kontakter med europeiska gemenskapens behöriga organ för att med dessa utarbeta konkreta förslag för att stärka samarbetet mellan våra organisationer.
Ministerkommittén har genom min rapport underrättats om resultatet av dessa kontakter och har utan att den inbördes fördelningen av behörighet mellan gemenskapen och dess medlemsstater åsidosätts kommit överens om följande:
a) Europeiska gemenskapen skall företrädd av kommissionen inbjudas att delta i arbete av ömsesidigt intresse i de kommittéer som inrättats av ministerkommittén och som består av personer som utnämnts av medlemsstaternas regeringar, däribland kommittéer av denna art som upprättats inom ramen för delöverenskommelser.
I de fall där gemenskapen har deltagit i utarbetandet av ett förslag till en europeisk konvention eller ett europeiskt avtal skall gemenskapen företrädd av kommissionen inbjudas att låta sig företrädas på de möten som ministrarnas ställföreträdare håller och där ett sådant förslag diskuteras.
b) Beträffande varje nytt förslag till konvention eller europeiskt avtal skall bedömas om det är lämpligt att infoga en klausul som tillåter Europeiska gemenskapen att bli part till konventionen eller avtalet. Infogandet av en sådan klausul föregriper inte på något sätt det beslut som gemenskapens behöriga organ kan fatta i fråga om gemenskapens ingående av konventionen eller avtalet.
c) Europeiska gemenskapen företrädd av kommissionen skall inbjudas att delta i arbete av ömsesidigt intresse vid fackministerkonferenser med vilka Europarådet har upprättat särskilda arbetsförbindelser, utan att detta påverkar de beslut som dessa konferensers behöriga organ kan komma att fatta.
Mot bakgrund av resultaten av våra kontakter och för att gå pragmatiskt tillväga utan att inrätta nya byråkratiska strukturer har ministerkommittén godkänt följande ordning, vilken utan att föregripa ett senare ingående av ett helhetsavtal med Europeiska gemenskapen kan accepteras av båda parter och vilken med beaktande av vad som anges ovan kan ersätta den ordning av den 18 augusti 1959 som kom till stånd genom skriftväxling mellan generalsekreteraren för Europarådet och ordförandena för Europeiska ekonomiska gemenskapen och Europeiska atomenergigemenskapen.
A. Vad beträffar förbindelserna mellan ministerkommittén och Europeiska gemenskapernas kommission:
1. Kommissionen skall till ministerkommittén vidarebefordra den årliga allmänna rapport som anges i artikel 18 i Fördraget om upprättandet av ett gemensamt råd och en gemensam kommission för Europeiska gemenskaperna. I gengäld mottar kommissionen ministerkommittén stadgeenliga rapporter och de rapporter som Europarådets generalsekreterare lägger fram för ministerkommittén om utvecklingen av det europeiska samarbetet.
2. Ministerkommittén får inbjuda kommissionen att delta i dess diskussioner om utvecklingen av det europeiska samarbetet samt om andra frågor av ömsesidigt intresse.
3. Kommissionen får inbjudas att låta sig företrädas och delta i sammanträden för ministrarnas ställföreträdare om frågor av ömsesidigt intresse.
4. Ministerkommittén får till kommissionen rikta de anmärkningar den kan ha rörande de rapporter som kommissionen lämnar och om alla andra frågor av ömsesidigt intresse.
5. Kommissionens generalsekreterare skall som regel en gång om året delta i ett utbyte av synpunkter med ministrarnas ställföreträdare för att överblicka läget för samarbetet mellan Europarådet och gemenskapen.
B. Vad beträffar förbindelserna mellan Europarådets generalsekreterare och Europeiska gemenskapernas kommission:
1. Generalsekreteraren och kommissionen skall vid behov samråda i frågor av ömsesidigt intresse. Detta samråd skall så långt som möjligt syfta till samordning och samförstånd samt gemensam verksamhet och bredast möjliga tillämpning av innehållet i de handlingar och andra dokument som båda parterna har antagit.
2. Möten på hög nivå skall vid behov äga rum mellan tjänstemän från Europarådets sekretariat och kommissionen i syfte att undersöka frågor av ömsesidigt intresse inom bestämda områden, underrätta sig om den andra partens program, överblicka läget för samarbetet och eventuellt bestämma om projekt som kan genomföras gemensamt jämte en tidsplan och en finansieringsplan för deras genomförande. Sådana möten skall regelmässigt anordnas särskilt angående rättsliga och sociala frågor, hälsovård, utbildning och kultur samt det europeiska gemensamma arvet och miljöfrågor utan att detta påverkar möjligheten att kalla till sådana möten inom andra områden av gemensamt intresse.
3. Kommissionen skall när det är lämpligt inbjuda företrädare för Europarådets sekretariat att delta som observatörer i arbetet i dess expertkommittéer och rådgivande grupper för att överlägga om frågor av gemensamt intresse.
4. Europarådets generalsekreterare och kommissionen skall vidta de åtgärder som krävs för att säkerställa nära förbindelser och samarbete mellan tjänstemän i de två organisationerna inom områden av ömsesidigt intresse. En hög tjänsteman skall av båda parterna utnämnas för att följa utvecklingen av samarbetet mellan de två organisationerna och tjäna som kontaktperson i detta syfte.
Jag skulle vara tacksam om Ni ville meddela mig huruvida kommissionen finner ovan nämnda regler acceptabla.
Högaktningsfullt
Marcelino OREJA
Generalsekreterare för Europarådet
B. Brev från Europeiska gemenskapernas kommission
Bryssel den 16 juni 1987
Jag har äran att bekräfta mottagandet av Ert brev av dagens datum om samarbetet mellan Europarådet och Europeiska gemenskapen.
Europeiska gemenskapernas kommission delar ministerkommitténs övertygelse att den europeiska solidariteten kommer att stärkas genom befästande och utvidgning av samarbetet mellan Europarådet och Europeiska gemenskapen, vilka är det europeiska samfundets väsentligaste organisationer. Kommissionen har uttryckt sin fasta vilja att med hänsyn till de två organisationernas särprägel och skilda förfaranden främja ett närmare samarbete mellan dem för att således verka för bredast möjliga samarbete på europeiskt plan.
Kommissionen är ytterst tillfredställd med de bestämmelser som ministerkommittén har beslutat anta enligt den rapport som Ni har bifogat i syfte att underlätta gemenskapens deltagande i Europarådets arbete, och den beaktar rapportens innehåll.
Dessutom har jag mot bakgrund av resultaten av våra kontakter och för att gå pragmatiskt tillväga utan att inrätta nya byråkratiska strukturer glädjen att på Europeiska gemenskapernas kommissions vägnar kunna underrätta Er om att jag godtar de regler i Ert brev som anges nedan och som utan att föregripa ett senare ingående av ett helhetsavtal med Europeiska gemenskapen träder ersätter den ordning som kom till stånd den 18 augusti 1959 genom en skriftväxling mellan generalsekreteraren för Europarådet och ordförandena för Europeiska ekonomiska gemenskapen och Europeiska atomenergigemenskapen.
A. Förbindelserna mellan ministerkommittén och Europeiska gemenskapernas kommission:
1. Kommissionen skall till ministerkommittén vidarebefordra den årliga allmänna rapport som anges i artikel 18 i Fördraget om upprättandet av ett gemensamt råd och en gemensam kommission för Europeiska gemenskaperna. I gengäld mottar kommissionen ministerkommitténs stadgeenliga rapporter och de rapporter som Europarådets generalsekreterare lägger fram för ministerkommittén om utvecklingen av det europeiska samarbetet.
2. Ministerkommittén får inbjuda kommissionen att delta i dess diskussioner om utvecklingen av det europeiska samarbetet samt om andra frågor av ömsesidigt intresse.
3. Kommissionen får inbjudas att låta sig företrädas och delta i sammanträden för ministrarnas ställföreträdare om frågor av ömsesidigt intresse.
4. Ministerkommittén får till kommissionen rikta de anmärkningar den kan ha rörande de rapporter som kommissionen lämnar och om alla andra frågor av ömsesidigt intresse.
5. Kommissionens generalsekreterare skall som regel en gång om året delta i ett utbyte av synpunkter med ministrarnas ställföreträdare för att överblicka läget för samarbetet mellan Europarådet och gemenskapen.
B. Förbindelserna mellan Europarådets generalsekreterare och Europeiska gemenskapernas kommission:
1. Generalsekreteraren och kommissionen skall vidr behov samråda i frågor av ömsesidigt intresse. Detta samråd skall så långt som möjligt syfta till samordning och samförstånd samt gemensam verksamhet och bredast möjliga tillämpning av innehållet i de handlingar och andra dokument som båda parterna har antagit.
2. Möten på hög nivå skall vid behov äga rum mellan tjänstemän från Europarådets sekretariat och kommissionen i syfte att undersöka frågor av ömsesidigt intresse inom bestämda områden, underrätta sig om den andra partens program, överblicka läget för samarbetet och eventuellt bestämma om projekt som kan genomföras gemensamt jämte en tidsplan och en finansieringsplan för deras genomförande. Sådana möten skall regelmässigt anordnas särskilt angående rättsliga och sociala frågor, hälsovård, utbildning och kultur samt det europeiska gemensamma arvet och miljöfrågor utan att detta påverkar möjligheten att kalla till sådana möten inom andra områden av gemensamt intresse.
3. Kommissionen skall när det är lämpligt inbjuda företrädare för Europarådets sekretariat att delta som observatörer i arbetet i dess expertkommittéer och rådgivande grupper för att överlägga om frågor av gemensamt intresse.
4. Europarådets generalsekreterare och kommissionen skall vidta de åtgärder som krävs för att säkerställa nära förbindelser och samarbete mellan tjänstemän i de två organisationerna inom områden av ömsesidigt intresse. En hög tjänsteman skall av båda parterna utnämnas för att följa utvecklingen av samarbetet mellan de två organisationerna och tjäna som kontaktperson i detta syfte. Högaktningsfullt
Jacques DELORS
Ordförande för Europeiska gemenskapernas kommission
WIPO:s fördrag om upphovsrätt
(WCT)
Genève (1996)
Innehåll
%gt%Plats för tabell%gt%
INLEDNING
DE FÖRDRAGSSLUTANDE PARTERNA,
HAR EN STRÄVAN ATT så effektivt och enhetligt som möjligt utveckla och upprätthålla skyddet av upphovsmännens rättigheter till deras litterära och konstnärliga verk,
ÄR MEDVETNA OM behovet av att införa nya internationella bestämmelser och av att förtydliga tolkningen av vissa redan befintliga bestämmelser i syfte att erbjuda ändamålsenliga lösningar till de frågor som den senaste ekonomiska, sociala, kulturella och teknologiska utvecklingen gett upphov till,
ÄR MEDVETNA OM den djupgående inverkan som utvecklingen och samverkan av informations- och kommunikationsteknik har på skapandet och användningen av litterära och konstnärliga verk,
UNDERSTRYKER DEN stora betydelse det upphovsrättsliga skyddet har som drivfjäder för litterärt och konstnärligt skapande,
ÄR MEDVETNA OM behovet att behålla en balans mellan upphovsmännens rättigheter och allmänhetens intresse, särskilt beträffande utbildning, forskning och tillgång till information, såsom det avspeglas i Bernkonventionen, och har
KOMMIT ÖVERENS OM FÖLJANDE.
Artikel 1
Sambandet med Bernkonventionen
1. Detta fördrag är en sådan särskild överenskommelse som avses i artikel 20 i Bernkonventionen för skydd av litterära och konstnärliga verk, med avseende på de fördragsslutande parter som ingår i den union som upprättats genom Bernkonventionen. Detta fördrag är inte förbundet med något annat fördrag än Bernkonventionen, och det inskränker inte rättigheter och skyldigheter enligt andra fördrag.
2. Bestämmelserna i detta fördrag inskränker inte de skyldigheter de fördragsslutande parterna har gentemot varandra enligt Bernkonventionen för skydd av litterära och konstnärliga verk.
3. I det följande avses med Bernkonventionen Bernkonventionen för skydd av litterära och konstnärliga verk, Paris den 24 juli 1971.
4. De fördragsslutande parterna skall iaktta artiklarna 1-21 i och bihanget till Bernkonventionen.
Artikel 2
Det upphovsrättsliga skyddets räckvidd
Det upphovsrättsliga skyddet omfattar uttryck men inte idéer, förfaranden, tillvägagångssätt eller matematiska begrepp som sådana.
Artikel 3
Tillämpning av artiklarna 2-6 i Bernkonventionen
Avseende det skydd som anges i fördraget skall de fördragsslutande parterna med vederbörliga ändringar tillämpa bestämmelserna i artiklarna 2-6 i Bernkonventionen.
Artikel 4
Datorprogram
Datorprogram skyddas som sådant litterärt verk som avses i artikel 2 i Bernkonventionen. Detta skydd gäller datorprogram oavsett på vilket sätt och i vilken form de kommer till uttryck.
Artikel 5
Sammanställning av data (databaser)
Sammanställningar av data eller annat material, oavsett form, som genom urvalet eller dispositionen av innehållet utgör intellektuella skapelser skyddas som sådana. Skyddet gäller inte denna data eller materialet som sådant och påverkar inte eventuell existerande upphovsrätt till den data eller det material som ingår i sammanställningen.
Artikel 6
Spridningsrätten
1. Upphovsmän till litterära och konstnärliga verk äger uteslutande rätt att låta göra originalet och exemplar av verket tillgängligt för allmänheten genom försäljning eller annan överlåtelse.
2. Detta fördrag påverkar inte möjligheten för de fördragsslutande parterna att bestämma under vilka omständigheter rätten enligt första stycket skall upphöra efter en första försäljning eller annan överlåtelse av originalet eller exemplar av verket som företagits med upphovsmannens medgivande.
Artikel 7
Uthyrningsrätten
1. Upphovsmän till
i) datorprogram,
ii) filmverk, och
iii) verk i form av fonogram, så som definieras i de fördragsslutande parternas nationella rätt,
äger uteslutande rätt att i vinstsyfte låta hyra ut originalet eller exemplar av sitt verk till allmänheten.
2. Första punkten gäller inte
i) datorprogram, när programmet som sådant inte är det huvudsakliga föremålet för uthyrningen; och
ii) filmverk, utom när sådan uthyrning i vinstsyfte har lett till utbredd kopiering av sådana verk och detta i väsentlig grad skadar den uteslutande rätten till mångfaldigande.
3. Utan hinder av bestämmelserna i första punkten kan en fördragsslutande part, som den 15 april 1994 upprätthöll och alltjämt upprätthåller en gällande ordning för skälig ersättning till upphovsmän för uthyrning av exemplar av deras verk i form av fonogram, vidmakthålla denna ordning under förutsättning att sådan uthyrning i vinstsyfte inte i väsentlig grad skadar upphovsmannens uteslutande rätt till mångfaldigande.
Artikel 8
Överföringsrätten
Utan att det påverkar tillämpningen av artikel 11.1.1, artikel 11a.1.1 och artikel 11a.1.2, artikel 11b.1.1, artikel 14.1.1 och artikel 14a.1 i Bernkonventionen, äger upphovsmän till litterära och konstnärliga verk uteslutande rätt att låta överföra verken till allmänheten, med tråd- eller trådlös överföring, inbegripet att göra verken tillgängliga för allmänheten på ett sådant sätt att personer ur allmänheten kan få tillgång till verken på platser och vid tidpunkter som var och en själv väljer.
Artikel 9
Skyddstiden för fotografiska verk
Med avseende på fotografiska verk skall de fördragsslutande parterna inte tillämpa bestämmelserna i artikel 7.4 i Bernkonventionen.
Artikel 10
Begränsningar och undantag
1. De fördragsslutande parterna kan i den nationella lagstiftningen föreskriva begränsningar av eller undantag från de rättigheter som enligt detta fördrag tillkommer upphovsmän till litterära och konstnärliga verk i vissa särskilda fall som inte gör intrång i det normala utnyttjandet av verket och inte heller på ett oskäligt sätt inkräktar på upphovsmannens rätt.
2. De fördragsslutande parterna skall vid tillämpningen av Bernkonventionen inskränka begränsningar av eller undantag från de rättigheter som anges i konventionen till vissa särskilda fall som inte gör intrång i det normala utnyttjandet av verket och inte heller på ett oskäligt sätt inkräktar på upphovsmannens rätt.
Artikel 11
Skyldigheter angående tekniska åtgärder
De fördragsslutande parterna skall vidta alla erforderliga åtgärder för att bereda ett tillräckligt rättsligt skydd och möjlighet att påkalla rättsliga åtgärder mot kringgåendet av verksamma tekniska åtgärder som upphovsmän använder i samband med att de utövar sina rättigheter enligt detta fördrag eller Bernkonventionen och som, med avseende på deras verk, begränsar handlingar som inte har medgivits av upphovsmännen i fråga och ej heller är tillåtna enligt lag.
Artikel 12
Skyldigheter angående information för förvaltning av rättigheter
1. De fördragsslutande parterna skall vidta alla erforderliga åtgärder för att bereda ett tillräckligt rättsligt skydd och möjlighet att påkalla rättsliga åtgärder mot personer som avsiktligen utfört någon av följande handlingar och som insåg eller såvitt avser civilrättsliga åtgärder borde ha insett att det medför, möjliggör, underlättar eller döljer ett intrång i en rättighet som följer av detta fördrag eller Bernkonventionen:
i) Att olovligen avlägsna eller ändra elektronisk information för förvaltning av rättigheter.
ii) Att olovligen sprida, importera i spridningssyfte, sända i radio eller överföra till allmänheten verk eller exemplar av verk med vetskap om att elektronisk information för förvaltning av rättigheter olovligen har avlägsnats eller ändrats.
2. Med information för förvaltning av rättigheter avses i denna artikel information som identifierar verket, verkets upphovsman, innehavare av rättighet till verket, eller information om villkoren för användning av verket, och siffror eller koder som betecknar sådan information, när sådan information bifogas ett exemplar av verket eller förekommer i samband med överföring av verket till allmänheten.
Artikel 13
Tillämpning i tidshänseende
De fördragsslutande parterna skall tillämpa bestämmelserna i artikel 18 i Bernkonventionen på allt skydd som omfattas av detta fördrag.
Artikel 14
Bestämmelser om upprätthållande av rättigheter
1. De fördragsslutande parterna åtar sig att i enlighet med sina rättssystem vidta erforderliga åtgärder för att säkerställa tillämpningen av detta fördrag.
2. De fördragsslutande parterna skall säkerställa att det i den nationella lagstiftningen finns föreskrifter om förfarande för upprätthållande så att verksamma åtgärder kan vidtas mot intrång i de rättigheter som omfattas av detta fördrag, inbegripet skyndsamma åtgärder för att förhindra intrång samt preventiva åtgärder.
Artikel 15
Församlingen
1. a) De fördragsslutande parterna skall ha en församling.
b) Varje fördragsslutande part skall företrädas av ett ombud som kan bistås av biträdande ombud, rådgivare och sakkunniga.
c) Kostnaderna för varje delegation skall bäras av den fördragsslutande part som utsett delegationen. Församlingen kan be Världsorganisationen för den intellektuella äganderätten (nedan kallad WIPO) att bevilja finansiellt stöd för att underlätta deltagandet för delegationer från fördragsslutande parter som anses som utvecklingsländer enligt den definition som fastställts av Förenta nationernas generalförsamling eller som är länder under övergång till marknadsekonomi.
2. a) Församlingen skall behandla frågor som rör upprätthållandet och utvecklingen av detta fördrag och dess tilllämpning och funktion.
b) Församlingen skall utföra sina åligganden enligt artikel 17.2 vad gäller upptagning av vissa mellanstatliga organisationer som parter till detta fördrag.
c) Församlingen skall besluta om sammankallande av diplomatkonferens för revidering av detta fördrag och ge WIPO:s generaldirektör alla erforderliga instruktioner för förberedandet av en sådan diplomatkonferens.
3. a) Varje fördragsslutande part som utgör en stat skall ha en röst och skall enbart rösta i sitt eget namn.
b) Fördragsslutande part som utgör en mellanstatlig organisation får delta i omröstning i sina medlemsstaters ställe, med ett antal röster som är lika med det antal av dess medlemsstater som är fördragsslutande parter. Sådan mellanstatlig organisation får inte delta i omröstning om en av dess medlemsstater utövar sin rösträtt och vice versa.
4. Församlingen skall sammanträda till ordinarie möte en gång vartannat år på kallelse av WIPO:s generaldirektör.
5. Församlingen antar själv sin arbetsordning, inbegripet sammankallande av extra ordinarie möte, bestämmelser om beslutsmässighet och, med förbehåll för bestämmelserna i detta fördrag, den majoritet som krävs för olika typer av beslut.
Artikel 16
Internationella byrån
WIPO:s internationella byrå skall utföra förvaltningsuppgifterna angående fördraget.
Artikel 17
Krav för att tillträda fördraget
1. Stater som är medlemmar i WIPO får tillträda fördraget.
2. Församlingen får besluta att låta en mellanstatlig organisation tillträda fördraget, om organisationen förklarar sig behörig i ärenden som omfattas av detta fördrag och har egen för medlemsstaterna bindande lagstiftning för sådana ärenden och den i vederbörlig ordning fått befogenhet att tillträda fördraget.
3. Europeiska gemenskapen, som avgivit en sådan förklaring som anges i föregående stycke under den diplomatkonferens som antagit detta fördrag, får tillträda fördraget.
Artikel 18
Rättigheter och skyldigheter enligt fördraget
Om inte annat särskilt föreskrivs i detta fördrag har varje fördragsslutande part utan inskränkningar de rättigheter och skyldigheter som följer av fördraget.
Artikel 19
Undertecknande av fördraget
Detta fördrag skall stå öppet för undertecknande till och med den 31 december 1997 för de stater som är medlemmar i WIPO och för Europeiska gemenskapen.
Artikel 20
Fördragets ikraftträdande
Detta fördrag träder i kraft tre månader efter det att trettio stater deponerat sina ratifikations- eller anslutningsinstrument hos WIPO:s generaldirektör.
Artikel 21
Faktiskt datum för tillträdet till fördraget
Detta fördrag är bindande för
i) de trettio stater som anges i artikel 20, från och med den dag då fördraget träder i kraft,
ii) övriga stater, tre månader från och med den dag då staten deponerade sitt instrument hos WIPO:s generaldirektör,
iii) Europeiska gemenskapen, tre månader efter det att den deponerat sitt ratifikations- eller anslutningsinstrument om sådant instrument deponerats efter detta fördrags ikraftträdande enligt artikel 20, eller, tre månader efter detta fördrags ikraftträdande om instrumentet deponerats före fördragets ikraftträdande,
iv) annan mellanstatlig organisation som får tillträda fördraget, tre månader efter det att den deponerat sitt anslutningsinstrument.
Artikel 22
Förbehåll mot fördraget
FörbehåIl mot detta fördrag är inte tillåtna.
Artikel 23
Uppsägning av fördraget
Fördragsslutande part kan säga upp fördraget genom meddelande till WIPO:s generaldirektör. Uppsägningen blir gällande ett år från och med den dag då WIPO:s generaldirektör mottagit meddelandet.
Artikel 24
Fördragets språk
1. Detta fördrag är undertecknat i ett original på engelska, arabiska, kinesiska, franska, ryska och spanska, och samtliga dessa versioner skall äga lika vitsord.
2. Officiella texter på andra språk än de som nämns i första stycket skall, på begäran av berörd part, efter samråd med alla berörda parter upprättas av WIPO:s generaldirektör. Med berörd part avses i detta stycke stat som är medlem i WIPO och vars officiella språk, eller något av dess officiella språk, berörs, och Europeiska gemenskapen och annan mellanstatlig organisation som får tillträda fördraget om något av dess officiella språk berörs.
Artikel 25
Depositarie
WIPO:s generaldirektör är depositarie för detta fördrag.
Eniga uttalanden
Beträffande artikel 1.4
Mångfaldiganderätten som fastställs i artikel 9 i Bernkonventionen och de undantag som tillåts enligt denna artikel gäller i sin helhet i den digitala miljön, framför allt för användningen av verk i digital form. Lagring av ett skyddat verk i digital form i ett elektroniskt medium utgör mångfaldigande enligt artikel 9 i Bernkonventionen.
Beträffande artikel 3
Vid tillämpning av artikel 3 i detta fördrag, skall uttrycket unionsland i artiklarna 2-6 i Bernkonventionen förstås som att det syftar på en fördragsslutande part till detta fördrag, när dessa artiklar i Bernkonventionen tillämpas avseende skydd som omfattas av detta fördrag. Uttrycket land utanför unionen i dessa artiklar i Bernkonventionen skall under samma omständigheter förstås som om det syftar på ett land som inte är fördragsslutande part till detta fördrag, och denna konvention i artikel 2.8, artikel 2a.2 och artiklarna 3, 4 samt 5 i Bernkonventionen skall förstås som att det syftar på Bernkonventionen och detta fördrag. Slutligen är hänsyftningen i artiklarna 3-6 i Bernkonventionen på upphovsmän som tillhör ett unionsland, vid de tillfällen då dessa artiklar tillämpas på detta fördrag och avseende mellanstatlig organisation som är fördragsslutande part, att förstå som medborgare i ett land som är medlem i denna organisation.
Beträffande artikel 4
Räckvidden för skyddet för datorprogram enligt artikel 4 i detta fördrag, jämfört med artikel 2, är förenlig med artikel 2 i Bernkonventionen och jämställd med vederbörliga bestämmelser i Trips-avtalet.
Beträffande artikel 5
Räckvidden för skyddet för insamling av data (databaser) enligt artikel 5 i detta fördrag, jämfört med artikel 2, är förenlig med artikel 2 i Bernkonventionen och jämställd med vederbörliga bestämmelser i Trips-avtalet.
Beträffande artiklarna 6 och 7
I dessa artiklar avses med uttrycken exemplar och originalet och exemplar, som föremål för spridnings- och uthyrningsrätten enligt dessa artiklar, endast fasta exemplar som kan sättas i omlopp som föremål.
Beträffande artikel 7
Förpliktelsen i artikel 7.1 innebär inte att en fördragsslutande part måste förbehålla upphovsmän uteslutande rätt till uthyrning i vinstsyfte, när dessa enligt den fördragsslutande partens lagstiftning inte har rättigheter beträffande fonogram. Denna förpliktelse är förenlig med artikel 14.4 i Trips-avtalet.
Beträffande artikel 8
Enbart tillhandahållandet av materiella hjälpmedel för att möjliggöra eller göra en överföring innebär i sig inte sådan överföring som avses i detta fördrag eller Bernkonventionen. Bestämmelserna i artikel 8 hindrar inte fördragsslutande part att tillämpa artikel 11a.2.
Beträffande artikel 10
Bestämmelserna i artikel 10 gör det möjligt för fördragsslutande parter att in i den digitala miljön föra vidare och vederbörligen utsträcka de begränsningar och undantag i sin nationella lagstiftning som har ansetts förenliga med Bernkonventionen. På samma sätt möjliggör dessa bestämmelser för de fördragsslutande parterna att skapa nya undantag och begränsningar som är lämpade för den digitala nätverksmiljön.
Artikel 10.2 varken begränsar eller utvidgar tillämpbarheten av begränsningar och undantag som är förenliga med Bernkonventionen.
Beträffande artikel 12
Uttrycket intrång i en rättighet som följer av detta fördrag eller Bernkonventionen innefattar både uteslutande rätt och rätt till ersättning.
Fördragsslutande parter kan inte med stöd av denna artikel skapa eller genomföra regleringar för förvaltning av rättigheter som skulle medföra formkrav som inte är tillåtna enligt Bernkonventionen eller detta fördrag och som förbjuder den fria rörligheten för varor eller hindrar åtnjutande av rättigheter som följer av detta fördrag.
Gemensamma EES-kommitténs beslut
nr 9/2005
av den 8 februari 2005
om ändring av bilaga II (Tekniska föreskrifter, standarder, provning och certifiering) till EES-avtalet
GEMENSAMMA EES-KOMMITTÉN HAR BESLUTAT FÖLJANDE
med beaktande av avtalet om Europeiska ekonomiska samarbetsområdet, ändrat genom protokollet med justeringar av avtalet om Europeiska ekonomiska samarbetsområdet, nedan kallat "avtalet", särskilt artikel 98 i detta, och
av följande skäl:
(1) Bilaga II till avtalet ändrades genom avtalet om Republiken Tjeckiens, Republiken Estlands, Republiken Cyperns, Republiken Lettlands, Republiken Litauens, Republiken Ungerns, Republiken Maltas, Republiken Polens, Republiken Sloveniens och Republiken Slovakiens deltagande i Europeiska ekonomiska samarbetsområdet, undertecknat i Luxemburg den 14 oktober 2003 [1]..
(2) Europaparlamentets och rådets direktiv 2003/17/EG av den 3 mars 2003 om ändring av direktiv 98/70/EG om kvaliteten på bensin och dieselbränslen [2] bör införlivas med avtalet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Följande skall läggas till i punkt 6a (Europaparlamentets och rådets direktiv 98/70/EG) i kapitel XVII i bilaga II till avtalet:
"— 32003 L 0017: Europaparlamentets och rådets direktiv 2003/17/EG av den 3 mars 2003 (EUT L 76, 22.3.2003, s. 10).
Bestämmelserna i direktivet skall, inom ramen för detta avtal, tillämpas med följande anpassningar:
a) I artikel 2.4 (yttersta randområden) skall "för Islands del hela dess territorium," införas efter "territorierna,".
b) I artikel 6.1 skall "artikel 95.10 i fördraget" ersättas med en hänvisning till "artikel 75 i avtalet"."
Artikel 2
Texterna till direktiv 2003/17/EG på isländska och norska, som skall offentliggöras i EES-supplementet till Europeiska unionens officiella tidning, skall vara giltiga.
Artikel 3
Detta beslut träder i kraft den 9 februari 2005 under förutsättning att alla anmälningar enligt artikel 103.1 i avtalet har gjorts till Gemensamma EES-kommittén [3].
Artikel 4
Detta beslut skall offentliggöras i EES-delen av och EES-supplementet till Europeiska unionens officiella tidning.
Gemensamma EES-kommitténs beslut
nr 19/2005
av den 8 februari 2005
om ändring av bilaga XXI (Statistik) till EES-avtalet
GEMENSAMMA EES-KOMMITTÉN HAR BESLUTAT FÖLJANDE
med beaktande av avtalet om Europeiska ekonomiska samarbetsområdet, anpassat genom protokollet med justeringar av avtalet om Europeiska ekonomiska samarbetsområdet, nedan kallat "avtalet", särskilt artikel 98 i detta, och
av följande skäl:
(1) Bilaga XXI till avtalet ändrades genom gemensamma EES‐kommitténs beslut nr 175/2004 av den 3 december 2004 [1].
(2) Europaparlamentets och rådets förordning (EG) nr 1267/2003 av den 16 juni 2003 om ändring av rådets förordning (EG) nr 2223/96 med avseende på tidsfrister för sändningen av huvudaggregaten i nationalräkenskaperna, undantag när det gäller sändningen av huvudaggregaten i nationalräkenskaperna och sändning av uppgifter om sysselsättning angivna i arbetade timmar [2] bör införlivas med avtalet.
(3) Rådets förordning (EG, Euratom) nr 1287/2003 av den 15 juli 2003 om harmonisering av bruttonationalinkomsten till marknadspris ("BNI‐förordning") [3] bör införlivas med avtalet.
(4) Europaparlamentets och rådets beslut nr 1608/2003/EG av den 22 juli 2003 om produktion och utveckling av gemenskapsstatistik om vetenskap och teknik [4] bör införlivas med avtalet.
(5) Detta beslut bör inte gälla Liechtenstein.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga XXI till avtalet skall ändras på följande sätt:
1. Följande strecksats skall läggas till i punkt 19d (rådets förordning (EG) nr 2223/96):
"— 32003 R 1267: Europaparlamentets och rådets förordning (EG) nr 1267/2003 av den 16 juni 2003 (EUT L 180, 18.7.2003, s. 1).
Bestämmelserna i förordningen skall, inom ramen för detta avtal, tillämpas med följande anpassning:
Denna förordning skall inte gälla Liechtenstein."
2. Följande punkt skall införas efter punkt 19o (Europaparlamentets och rådets förordning (EG) nr 501/2004):
"19p. 32003 R 1287: Rådets förordning (EG, Euratom) nr 1287/2003 av den 15 juli 2003 om harmonisering av bruttonationalinkomsten till marknadspris ("BNI‐förordning") (EUT L 181, 19.7.2003, s. 1).
Bestämmelserna i förordningen skall, inom ramen för detta avtal, tillämpas med följande anpassning:
Denna förordning skall inte gälla Liechtenstein"
3. Följande skall införas efter punkt 28 (Europaparlamentets och rådets förordning (EG) nr 808/2004):
"STATISTIK OM VETENSKAP OCH TEKNIK
29. 32003 D 1608: Europaparlamentets och rådets beslut nr 1608/2003/EG av den 22 juli 2003 om produktion och utveckling av gemenskapsstatistik om vetenskap och teknik (EUT L 230, 16.9.2003, s. 1).
Bestämmelserna i beslutet skall, inom ramen för detta avtal, tillämpas med följande anpassning:
Detta beslut skall inte gälla Liechtenstein."
Artikel 2
Texterna till förordning (EG) nr 1267/2003, förordning (EG, Euratom) nr 1287/2003 och beslut nr 1608/2003/EG på isländska och norska, som skall offentliggöras i EES‐supplementet till Europeiska unionens officiella tidning, skall vara giltiga.
Artikel 3
Detta beslut träder i kraft den 9 februari 2005 under förutsättning att alla anmälningar enligt artikel 103.1 i avtalet har gjorts till gemensamma EES‐kommittén [5].
Artikel 4
Detta beslut skall offentliggöras i EES‐delen av och EES‐supplementet till Europeiska unionens officiella tidning.
Information om ikraftträdandet av protokollet till Europa–Medelhavsavtalet mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Arabrepubliken Egypten, å andra sidan, med anledning av Republiken Tjeckiens, Republiken Estlands, Republiken Cyperns, Republiken Lettlands, Republiken Litauens, Republiken Ungerns, Republiken Maltas, Republiken Polens, Republiken Sloveniens och Republiken Slovakiens anslutning till Europeiska unionen [1] Den 22 september 2005 utväxlades instrumenten för anmälan om avslutandet av de förfaranden som krävs för ikraftträdandet av protokollet, undertecknat i Bryssel den 20 december 2004, till Europa–Medelhavsavtalet mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Arabrepubliken Egypten, å andra sidan, med anledning a
Sedan förhandlingar inletts mellan Europeiska gemenskapen (EG) och Konungariket Thailand i enlighet med artikel XXIV.6 och artikel XXVIII i GATT 1994 om ändring av medgivanden i Republiken Tjeckiens, Republiken Estlands, Republiken Cyperns, Republiken Lettlands, Republiken Litauens, Republiken Ungerns, Republiken Maltas, Republiken Polens, Republiken Sloveniens och Republiken Slovakiens bindningslistor inom ramen för deras anslutning till Europeiska unionen, avtalas följande mellan EG och Konungariket Thailand i syfte att avsluta dessa förhandlingar, som inleddes som en följd av EG:s anmälan till WTO av den 19 januari 2004 enligt artikel XXIV.6 i GATT 1994. EG samtycker till att i sin bindningslista för tullområdet för EG med 25 medlemsstater införliva de medgivanden som ingick i den tidigare bindningslistan för EG med 15 medlemsstater.
EG samtycker till att i sin bindningslista för EG med 25 medlemsstater införliva de medgivanden som är uppförda i bilagan till detta avtal. Konungariket Thailand godtar de grundläggande delarna av EG:s tillvägagångssätt när det gäller att anpassa de skyldigheter inom ramen för GATT som gäller för EG med 15 medlemsstater och de som gäller för Republiken Tjeckien, Republiken Estland, Republiken Cypern, Republiken Lettland, Republiken Litauen, Republiken Ungern, Republiken Malta, Republiken Polen, Republiken Slovenien och Republiken Slovakien efter EG:s senaste utvidgning, nämligen tillämpning av nettometoden när det gäller exportåtaganden, tillämpning av nettometoden när det gäller tullkvoter och sammanslagning av åtaganden beträffande inhemskt stöd.
Med utmärkt högaktning För Europeiska gemenskapen
Avtal
mellan Republiken Albaniens ministerråd och Europeiska gemenskapen om vissa luftfartsaspekter
REPUBLIKEN ALBANIENS MINISTERRÅD,
å ena sidan, och
EUROPEISKA GEMENSKAPEN,
å andra sidan,
nedan kallade "parterna", som
KONSTATERAR att bilaterala luftfartsavtal har slutits mellan flera medlemsstater i Europeiska gemenskapen och Republiken Albanien med bestämmelser som strider mot EG-rätten,
KONSTATERAR att endast Europeiska gemenskapen är behörig i fråga om många av de aspekter som kan omfattas av bilaterala luftfartsavtal mellan medlemsstater i Europeiska gemenskapen och tredjeländer,
KONSTATERAR att enligt EG-rätten har lufttrafikföretag från gemenskapen som är etablerade i en medlemsstat rätt till icke diskriminerande tillgång till flygrutter mellan medlemsstaterna i Europeiska gemenskapen och tredjeländer,
BEAKTAR de avtal mellan Europeiska gemenskapen och vissa tredjeländer som innebär att medborgare i dessa tredjeländer får förvärva äganderätt i lufttrafikföretag som har tillstånd utfärdade i enlighet med EG rätten,
INSER att bestämmelser i de bilaterala luftfartsavtalen mellan medlemsstaterna i EG och Republiken Albanien som står i strid med EG-rätten måste ändras så att de blir förenliga med denna för att en sund rättslig grund skall kunna skapas för flygtrafiken mellan Europeiska gemenskapen och Republiken Albanien och för att kontinuiteten i denna flygtrafik skall kunna upprätthållas,
KONSTATERAR att Europeiska gemenskapen inte har som mål att som ett led i dessa förhandlingar öka totalvolymen för flygtrafik mellan Europeiska gemenskapen och Republiken Albanien, påverka balansen mellan lufttrafikföretag från gemenskapen och lufttrafikföretag från Albanien eller förhandla fram ändringar i de befintliga bilaterala luftfartsavtalen när det gäller trafikrättigheter,
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Allmänna bestämmelser
1. I detta avtal avses med "medlemsstat" en medlemsstat i Europeiska gemenskapen.
2. Hänvisningar i något av de avtal som ingår i förteckningen i bilaga I till medborgare i en medlemsstat som är part i det avtalet skall innebära hänvisningar till medborgare i Europeiska gemenskapens medlemsstater.
3. Hänvisningar i något av de avtal som ingår i förteckningen i bilaga I till lufttrafikföretag i en medlemsstat som är part i det avtalet skall innebära hänvisningar till lufttrafikföretag som har utsetts av den medlemsstaten.
Artikel 2
Lufttrafikföretag utsedda av en medlemsstat
1. Bestämmelserna i punkterna 2 och 3 i den här artikeln skall äga företräde framför motsvarande bestämmelser i de artiklar som förtecknas i bilaga II a respektive b, när det gäller den berörda medlemsstatens utseende av ett lufttrafikföretag, godkännanden och tillstånd som Republiken Albanien beviljat för det företaget samt vägran, återkallande, tillfälligt upphävande eller begränsning av godkännanden eller tillstånd för lufttrafikföretaget.
2. När Republiken Albanien har underrättats om att ett lufttrafikföretag har utsetts av en medlemsstat, skall Republiken Albanien utfärda de tillämpliga godkännandena och tillstånden med så kort handläggningstid som möjligt, under förutsättning att i) lufttrafikföretaget i enlighet med fördraget om upprättandet av Europeiska gemenskapen är etablerat i den medlemsstat där det har utsetts och har en giltig operativ licens i enlighet med EG-rätten,
ii) att den medlemsstat som utfärdar drifttillstånd (AOC) utövar faktisk tillsyn över lufttrafikföretaget och att dess luftfartsmyndighet finns tydligt angiven i den handling där lufttrafikföretaget utses, och
iii) lufttrafikföretaget ägs och skall fortsätta att ägas direkt eller genom majoritetsägande av medlemsstater och/eller medborgare i medlemsstater och/eller av andra stater som är förtecknade i bilaga III och/eller av medborgare i sådana andra stater och att det alltid står under faktisk kontroll av dessa stater och/eller dessa medborgare.
3. Republiken Albanien får vägra, återkalla, tillfälligt upphäva eller begränsa godkännanden och tillstånd för ett lufttrafikföretag som har utsetts av en medlemsstat om
i) lufttrafikföretaget i enlighet med fördraget om upprättandet av Europeiska gemenskapen inte är etablerat i den medlemsstat där det har utsetts eller inte har en giltig operativ licens i enlighet med EG-rätten,
ii) den medlemsstat som utfärdar AOC (Air Operator Certificate) inte utövar faktisk tillsyn över lufttrafikföretaget eller om dess luftfartsmyndighet inte är tydligt angiven i den handling där lufttrafikföretaget utses, eller
iii) lufttrafikföretaget inte ägs eller står under kontroll direkt eller genom majoritetsägande av medlemsstater och/eller medborgare i medlemsstater och/eller av andra stater som är förtecknade i bilaga III och/eller av medborgare i sådana andra stater.
Vid utövandet av sina rättigheter enligt denna punkt får Republiken Albanien inte diskriminera EU lufttrafikföretag på grundval av nationalitet.
Artikel 3
Rättigheter i fråga om tillsyn
1. Bestämmelserna i punkt 2 i den här artikeln skall komplettera de artiklar som förtecknas i bilaga II c.
2. Om en medlemsstat har utsett ett lufttrafikföretag för vilket tillsynen utövas av en annan medlemsstat, skall Republiken Albaniens rättigheter enligt säkerhetsbestämmelserna i avtalet mellan den medlemsstat som har utsett lufttrafikföretaget och Republiken Albanien tillämpas på samma sätt när det gäller säkerhetsnormer som antas och tillämpas av den andra medlemsstaten samt när det gäller tillståndet för nämnda lufttrafikföretags trafik.
Artikel 4
Beskattning av flygbränsle
1. Bestämmelserna i punkt 2 i den här artikeln skall komplettera de artiklar som förtecknas i bilaga II d.
2. Utan hinder av eventuella andra bestämmelser med annat innehåll skall ingenting i de avtal som förtecknas i bilaga II d hindra en medlemsstat från att beskatta eller tull- eller avgiftsbelägga flygbränsle som tillhandahålls på dess territorium och som är avsett för luftfartyg som tillhör ett lufttrafikföretag som har utsetts av Republiken Albanien och som går i trafik mellan en ort i den medlemsstaten och en annan ort i den medlemsstaten eller i en annan medlemsstat.
Artikel 5
Priser för transporter inom Europeiska gemenskapen
1. Bestämmelserna i punkt 2 i den här artikeln skall komplettera de artiklar som förtecknas i bilaga II e.
2. De priser som tas ut av lufttrafikföretag som utses av Republiken Albanien enligt ett avtal i förteckningen i bilaga I med en bestämmelse som finns förtecknad i bilaga II e för transport helt och hållet inom Europeiska gemenskapen skall vara förenliga med EG-rätten.
Artikel 6
Bilagor till avtalet
Bilagorna till detta avtal utgör en integrerad del av detta.
Artikel 7
Översyn och ändring
Parterna får när som helst genom överenskommelse se över eller ändra detta avtal.
Artikel 8
Ikraftträdande och provisorisk tillämpning
1. Detta avtal skall träda i kraft när parterna skriftligen har underrättat varandra om att de respektive interna förfaranden som krävs för ikraftträdandet har slutförts.
2. Utan hinder av vad som sägs i punkt 1 skall parterna vara överens om att provisoriskt tillämpa detta avtal från och med den första dagen i den månad som följer på den dag då parterna har underrättat varandra om att de förfaranden som är nödvändiga för detta ändamål har slutförts.
3. Avtal och andra överenskommelser mellan medlemsstaterna och Republiken Albanien som ännu inte har trätt i kraft när det här avtalet undertecknas och som inte preliminärt tillämpas förtecknas i bilaga I b. Det här avtalet skall tillämpas på alla sådana avtal och överenskommelser när de har trätt i kraft eller tillämpas provisoriskt.
Artikel 9
Upphörande
1. Om ett avtal som förtecknas i bilaga I upphör att gälla, skall alla bestämmelser i det här avtalet som avser det avtal som förtecknas i bilaga I upphöra att gälla vid samma tidpunkt.
2. Om alla de avtal som förtecknas i bilaga I upphör att gälla, skall det här avtalet upphöra att gälla vid samma tidpunkt.
Gemensamma EES-kommitténs beslut
nr 2/2006
av den 27 januari 2006
om ändring av bilaga II (Tekniska föreskrifter, standarder, provning och certifiering) till EES-avtalet
GEMENSAMMA EES-KOMMITTÉN HAR BESLUTAT FÖLJANDE
med beaktande av avtalet om Europeiska ekonomiska samarbetsområdet, ändrat genom protokollet med justeringar av avtalet om Europeiska ekonomiska samarbetsområdet, nedan kallat %quot%avtalet%quot%, särskilt artikel 98, och
av följande skäl:
(1) Bilaga II till avtalet ändrades genom gemensamma EES-kommitténs beslut nr 112/2005 av den 30 september 2005 [1].
(2) Kommissionens direktiv 2005/30/EG av den 22 april 2005 om ändring, för att anpassa dem till den tekniska utvecklingen, av Europarlamentets och rådets direktiv 97/24/EG och 2002/24/EG avseende typgodkännande av två- och trehjuliga motorfordon [2] bör införlivas med avtalet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Kapitel I i bilaga II till avtalet skall ändras på följande sätt:
1) Följande strecksats skall läggas till i punkterna 45x (Europaparlamentets och rådets direktiv 97/24/EG) och 45za (Europaparlamentets och rådets direktiv 2002/24/EG):
- %quot%— 32005 L 0030: Kommissionens direktiv 2005/30/EG av den 22 april 2005 (EUT L 106, 27.4.2005, s. 17)%quot%.
2) Följande punkt skall införas efter punkt 45zf (kommissionens direktiv 2004/104/EG):
%quot%45zg. 32005 L 0030: Kommissionens direktiv 2005/30/EG av den 22 april 2005 om ändring, för att anpassa dem till den tekniska utvecklingen, a
Gemensamma EES-kommitténs beslut
nr 96/2006
av den 7 juli 2006
om ändring av bilaga XXI (Statistik) till EES-avtalet
GEMENSAMMA EES-KOMMITTÉN HAR BESLUTAT FÖLJANDE
med beaktande av avtalet om Europeiska ekonomiska samarbetsområdet, ändrat genom protokollet med justeringar av avtalet om Europeiska ekonomiska samarbetsområdet, nedan kallat "avtalet", särskilt artikel 98, och
av följande skäl:
(1) Bilaga XXI till avtalet ändrades genom gemensamma EES-kommitténs beslut nr 71/2006 av den 2 juni 2006 [1].
(2) Kommissionens förordning (EG) nr 341/2006 av den 24 februari 2006 om antagande av specifikationer för 2007 års ad hoc-modul om olycksfall i arbetet och arbetsrelaterade hälsoproblem i enlighet med rådets förordning (EG) nr 577/98 och om ändring av förordning (EG) nr 384/2005 [2] bör införlivas med avtalet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga XXI till avtalet skall ändras på följande sätt:
1. Följande punkt skall införas efter punkt 18ai (kommissionens förordning (EG) nr 430/2005):
"18aj. 32006 R 0341: Kommissionens förordning (EG) nr 341/2006 av den 24 februari 2006 om antagande av specifikationer för 2007 års ad hoc-modul om olycksfall i arbetet och arbetsrelaterade hälsoproblem i enlighet med rådets förordning (EG) nr 577/98 och om ändring av förordning (EG) nr 384/2005 (EUT L 55, 25.2.2006, s. 9)".
2. Följande skall läggas till i punkt 18ag (kommissionens förordning (EG) nr 384/2005):
", ändrad genom
- 32006 R 0341: Kommissionens förordning (EG) nr 341/2006 av den 24 februari 2006 (EUT L 55, 25.2.2006, s. 9)".
Artikel 2
Texten till förordning (EG) nr 341/2006 på isländska och norska, som skall offentliggöras i EES-supplementet till Europeiska unionens officiella tidning, skall vara giltig.
Artikel 3
Detta beslut träder i kraft den 8 juli 2006 under förutsättning att alla anmälningar enligt artikel 103.1 i avtalet har gjorts till gemensamma EES-kommittén [3].
Artikel 4
Detta beslut skall offentliggöras i EES-delen av och EES-supplementet till Europeiska unionens officiella tidning.
Beslut nr 3/2006 av AVS–EG-ambassadörskommittén
av den 27 september 2006
om budgetförordning för Teknikcentrum för jordbruks- och landsbygdssamarbete
(2006/877/EG)
AVS–EG-AMBASSADÖRSKOMMITTÉN HAR BESLUTAT FÖLJANDE
med beaktande av partnerskapsavtalet mellan medlemmarna i gruppen av stater i Afrika, Västindien och Stillahavsområdet, å ena sidan, och Europeiska gemenskapen och dess medlemsstater, å andra sidan, undertecknat i Cotonou den 23 juni 2000 [1] (nedan kallat "avtalet"), särskilt artikel 3.4 b och d i bilaga III,
med beaktande av det interna avtalet av den 18 september 2000 mellan företrädarna för medlemsstaternas regeringar, församlade i rådet, om finansiering och förvaltning av gemenskapens bistånd inom ramen för finansprotokollet till partnerskapsavtalet mellan staterna i Afrika, Västindien och Stillahavsområdet, å ena sidan, och Europeiska gemenskapen och dess medlemsstater, å andra sidan, undertecknat i Cotonou (Benin) den 23 juni 2000, och om tilldelning av ekonomiskt stöd till de utomeuropeiska länder och territorier på vilka den fjärde delen av EG-fördraget är tillämplig [2],
med beaktande av budgetförordningen av den 27 mars 2003 för den nionde Europeiska utvecklingsfonden [3],
med beaktande av kommissionens förslag, som utarbetats i samarbete med Teknikcentrum för jordbruks- och landsbygdssamarbete, och
av följande skäl:
(1) Enligt artikel 3.4 b i bilaga III till avtalet skall ambassadörskommittén, efter avtalets undertecknande, fastställa budgetförordningen för Teknikcentrum för jordbruks- och landsbygdssamarbete (nedan kallat "centrumet").
(2) Enligt artikel 3.4 d i bilaga III till avtalet skall ambassadörskommittén fastställa förfaranden för antagande av centrumets budget. HÄRIGENOM FÖRESKRIVS FÖLJANDE.
KAPITEL I
ALLMÄNNA PRINCIPER
AVSNITT 1
Principer om enhet, riktighet och jämvikt i budgeten och en enda beräkningsenhet
Artikel 1
1. Alla centrumets inkomster och utgifter skall beräknas på grundval av ett kostnadsberäknat årligt arbetsprogram, som skall upprättas för varje budgetår och tas upp i budgeten.
2. Budgetens inkomster och utgifter skall balansera varandra.
Artikel 2
Budgeten skall upprättas och genomföras i euro och räkenskaperna skall redovisas i euro. För behov som avser förvaltning får centrumet dock genomföra transaktioner i medlemsstaternas och AVS-staternas nationella valutor.
Artikel 3
1. Inkomsterna skall bestå av bidragen från Europeiska utvecklingsfonden (nedan kallad "EUF") det belopp som tas ut i form av skatter på löner och annan ersättning från centrumet samt andra intäkter.
2. Inkomsterna kan också bestå av bidrag från andra givare till centrumets budget.
3. Centrumet får även på tredje parts vägnar förvalta medel avsedda för samfinansiering av de verksamheter som fastställs i bilaga III till avtalet. De finansiella reglerna för förvaltningen av dessa medel fastställs i artikel 34 i det här beslutet.
Artikel 4
Utgiftsberäkningen skall omfatta administrations- och driftskostnader. Det skall göras en klar åtskillnad mellan dem i budgeten.
Artikel 5
1. Budgetåret skall inledas den 1 januari och avslutas den 31 december.
2. De anslag som tas upp i budgeten skall beviljas för ett budgetår.
Anslag för vilka åtaganden gjorts i vederbörlig ordning under ett budgetår, men som inte betalats ut per den 31 december det året, skall dock automatiskt överföras till det närmast följande budgetåret. Anslag som överförts på detta sätt skall klart framgå av räkenskaperna för det löpande budgetåret.
De anslag som dras tillbaka vid utgången av ett budgetår skall återföras till den femåriga finansram som fastställts för centrumet i avtalet.
3. Vid utgången av varje finansprotokoll till avtalet skall anslag för vilka åtaganden gjorts, men som inte utbetalats, automatiskt överföras till nästa finansprotokoll till avtalet. Anslag för vilka åtaganden gjorts, men som inte utbetalats när avtalet löper ut, skall överföras endast under övergångsperioden mellan avtalet och nästa avtal eller, vid behov, under avräkningsperioden på tolv månader.
4. Om beslut om den slutgiltiga budgeten ännu inte föreligger vid budgetårets början får direktören, i syfte att sörja för kontinuitet i centrumets verksamhet, godkänna månatliga utgifter på upp till en tolftedel av de motsvarande anslag för artikeln i fråga som beviljats i budgeten för det föregående året.
När det gäller driftskostnader som skall betalas i förväg för varje kvartal och godkänts i budgeten för det föregående budgetåret, får åtaganden göras per artikel för upp till en fjärdedel av det totala anslag som beviljats för artikeln i fråga för det föregående budgetåret.
AVSNITT 2
Principer om en sund ekonomisk förvaltning
Artikel 6
1. Budgetanslagen skall användas i enlighet med principen om en sund ekonomisk förvaltning, dvs. enligt principerna om sparsamhet, effektivitet och ändamålsenlighet.
2. Principen om sparsamhet innebär att medlen skall göras tillgängliga i rätt tid till lägsta möjliga kostnad samt vara av den kvantitet och kvalitet som behövs.
Principen om effektivitet åsyftar bästa möjliga förhållande mellan de resurser som används och de resultat som uppnås.
Principen om ändamålsenlighet avser hur väl specifika mål med en åtgärd och förväntade resultat uppnås.
3. Tydliga mål skall fastställas och genomförandet av dem skall övervakas med hjälp av mätbara indikatorer. Vid behov skall de projekt som skall finansieras med medel från EUF bygga på bedömningar i förväg. Resultatet av dessa bedömningar skall införas i de handlingar som läggs fram för kommissionen till stöd för det årliga bidrag från EUF som begärs av centrumet.
KAPITEL II
UPPRÄTTANDE AV BUDGETEN
Artikel 7
1. Inom ramen för det övergripande strategidokumentet och den samlade budget som avsatts för centrumet genom finansprotokollet skall direktören upprätta ett utkast till ett årligt arbetsprogram och ett budgetförslag. Utkastet och förslaget skall godkännas av styrelsen senast den 1 juli året före arbetsprogrammets och budgetens genomförande och överlämnas till ambassadörskommittén för antagande.
2. Centrumet skall överlämna ett exemplar av utkastet till årligt arbetsprogram och budgetförslaget till kommissionen, som skall inleda de förfaranden som krävs för deras godkännande.
3. Åtaganden skall kunna göras från budgeten från och med den dag då gemenskapsmyndigheten antar beslutet om finansiering av det begärda bidraget från EUF. Centrumet skall underrättas om detta beslut.
Artikel 8
1. Villkoren för utbetalning av bidrag från EUF skall fastställas i en överenskommelse om bidrag, som skall undertecknas av centrumet och kommissionen.
2. Centrumet skall till EUF återbetala de bidrag för föregående budgetår som motsvarar anslag vilka förfallit enligt reviderade årsbokslut.
3. Budgeten skall delas in i avdelningar (budgetrubriker), kapitel, artiklar och punkter allt efter inkomstens eller utgiftens slag eller ändamål.
Artikel 9
Direktören får vid behov lägga fram ett förslag till tilläggs- eller ändringsbudget, som skall upprättas på samma sätt och underkastas samma förfaranden som den budget som innehöll de ursprungliga beräkningarna.
KAPITEL III
GENOMFÖRANDE AV BUDGETEN
Artikel 10
1. Direktören skall genomföra budgeten under eget ansvar och inom ramarna för beviljade anslag. Direktören skall rapportera till styrelsen om förvaltningen av budgeten.
2. Direktören skall använda budgetanslagen i enlighet med de principer om en sund ekonomisk förvaltning som avses i artikel 6.
Artikel 11
1. Alla inkomster och utgifter skall medföra att en artikel i budgeten krediteras eller debiteras.
Åtagande om eller godkännande av utgifter utöver beviljade anslag för det berörda budgetåret eller utöver de anslag som överförts från det föregående budgetåret får inte göras.
2. Alla inkomster och utgifter skall tas upp som bruttobelopp i räkenskaperna utan att avräknas mot varandra.
Trots denna bestämmelse får följande avdrag göras från beviljade belopp:
a) Böter som förelagts en part i ett avtal.
b) Justering av ett felaktigt betalat belopp, vilket kan göras genom avdrag när en senare utgiftskontroll görs under samma kapitel, artikel och budgetår som den felaktiga betalningen.
c) Värdet av fordon, utrustning och anläggningar som använts som dellikvid vid köp av ny utrustning av samma slag; nettoinköpspriset skall i räkenskaperna tas upp som anskaffningskostnad med tanke på inventarieförteckningen.
d) Rabatter och andra avdrag som räknats av i fakturor och räkningar.
Likaledes trots denna bestämmelse får följande belopp återanvändas inom samma budgetrubrik som den ursprungliga utgiften:
a) Inkomster från återbetalning av belopp som utbetalats felaktigt.
b) Mottagna försäkringsersättningar.
c) Förtjänster från försäljning av fordon, utrustning och anläggningar som avyttrats när de bytts ut.
d) Intäkter från försäljning av publikationer och filmer.
e) De valutakursförändringar som inträffat under genomförandet av budgeten får kompenseras. Den slutliga vinsten eller förlusten skall tas upp i bokslutet.
Artikel 12
Överföringar från en avdelning till en annan skall godkännas av styrelsen. Beslut om överföringar från ett kapitel till ett annat och från en artikel till en annan inom ett kapitel skall fattas av direktören, som skall underrätta styrelsen.
Artikel 13
Centrumets inkomster skall sättas in på ett eller flera konton som öppnats i centrumets namn.
KAPITEL IV
FINANSIELL KONTROLL
Artikel 14
1. En styrekonom som utses av styrelsen skall vara ansvarig för förhandsgodkännandet av åtagandet och godkännandet när det gäller alla utgifter, inkomster och förskott.
2. Styrekonomen skall bevisligen ha erfarenhet av budgetregler för internationella organisationer och av revision.
3. Styrekonomen skall uppfylla anställningsvillkoren för centrumets personal. Han skall för administrativa ändamål rapportera till centrumets direktör. Alla beslut som rör disciplinära åtgärder, avstängning, upphörande av tjänstgöringen eller rättsliga förfaranden skall dock antas av styrelsen på grundval av ett motiverat förslag från direktören.
4. De kontroller som utförs av styrekonomen skall leda fram till att ett godkännande ges eller förvägras. Syftet med godkännandet skall vara att se till att
a) utgifterna eller inkomsterna är förenliga med budgeten och förordningarna,
b) de principer om sund ekonomisk förvaltning som avses i artikel 6 har tillämpats.
Kontrollerna skall utföras i enlighet med de regler för det interna förfarandet som direktören har lagt fram för styrelsen och som godkänts av denna.
5. Om godkännande förvägras skall en skriftlig motivering lämnas till direktören. Om inte skälet är att det saknas tillräckliga anslag, får direktören genom ett motiverat beslut och på eget ansvar bortse från styrekonomens vägran att lämna sitt godkännande. Direktören skall skriftligen underrätta styrelsen om varje sådant beslut vid nästa möte.
6. Styrekonomen skall ha tillgång till alla styrkande handlingar och alla andra handlingar som rör utgifter eller inkomster som skall kontrolleras. Styrekonomen får utföra kontroller på plats.
7. Styrekonomen skall vara fullständigt oberoende i sitt arbete. Styrekonomen får inte ta emot instruktioner och får inte åläggas några restriktioner i sitt arbete.
8. Direktören får inhämta styrekonomens åsikter om frågor som rör analys, organisation och förbättring av centrumets interna förfaranden. Direktören får även uppmana styrekonomen att granska handlingar för att förvissa sig om huruvida verksamhet som finansierats genom budgeten har utförts på ett korrekt sätt.
9. I slutet av varje budgetår och senast den 30 april det påföljande året skall styrekonomen utarbeta en årlig rapport där han uttalar sig om den finansiella administrationen och genomförandet av budgeten. Styrekonomen skall överlämna rapporten till direktören som vid nästa möte skall överlämna den till styrelsen med sina egna kommentarer.
KAPITEL V
FÖRVALTNING AV BUDGETEN
Artikel 15
1. Centrumets budget skall förvaltas i enlighet med principen om åtskillnad mellan utanordnarens och räkenskapsförarens uppgifter. Anslagen skall förvaltas av utanordnaren, som ensam har befogenhet att göra utgiftsåtaganden, fastställa fordringar samt utfärda betalningskrav och betalningsorder.
2. Räkenskapsföraren skall svara för mottagande av inkomster och betalning av utgifter.
3. Utanordnaren får inte utföra räkenskapsförarens uppgifter.
Artikel 16
1. Alla åtgärder som kan ge upphov till en utgift som skall betalas av centrumet skall föregås av ett förslag till åtagande, vilket tillsammans med styrkande handlingar i original skall överlämnas till styrekonomen för förhandskontroll.
2. För återkommande utgifter får ett preliminärt åtagande göras.
3. Åtaganden och betalningsorder skall bokföras. Det skall finnas bokföringsuppgifter om åtaganden och godkännanden.
Artikel 17
1. Syftet med utanordnarens kontroll av utgifter skall vara att
a) kontrollera att borgenärens anspråk existerar,
b) fastställa eller kontrollera att fordran existerar och vilket belopp den uppgår till,
c) kontrollera fordrans förfallovillkor.
2. Varje betalning av utgifter skall grundas på styrkande handlingar som bekräftar borgenärens anspråk på betalning för tjänster som tillhandahållits, varor som levererats eller entreprenader som utförts, eller andra styrkande handlingar som berättigar till betalning.
Alla beslut om betalningar skall godkännas av den behörige utanordnaren.
Artikel 18
1. Godkännandet är den handling genom vilken utanordnaren, genom utfärdande av en betalningsorder, beordrar räkenskapsföraren att betala en utgift som utanordnaren har kontrollerat.
2. Betalningsordern skall åtföljas av samtliga styrkande handlingar i original, som skall innehålla eller åtföljas av ett intyg från utanordnaren om att de belopp som skall betalas är korrekta, att varorna har mottagits och att tjänsterna har utförts.
3. Kopior av de styrkande handlingarna, vilkas överensstämmelse med originalet har bestyrkts av utanordnaren, får i vissa fall godtas i stället för original.
4. Betalningsorder skall överlämnas till räkenskapsföraren för betalning.
5. I förekommande fall skall den betalningsorder som överlämnas till räkenskapsföraren åtföljas av ett intyg om att de berörda tillgångarna har förts upp i inventarieförteckningen.
Artikel 19
1. Betalningen är den slutliga handling genom vilken centrumet befrias från förpliktelserna gentemot sina borgenärer.
2. Betalning skall utföras av räkenskapsföraren inom ramen för de disponibla medlen.
3. Räkenskapsföraren skall hålla inne betalningen om sakfel föreligger, om befrielsen från förpliktelser gentemot borgenären ifrågasätts eller om de formaliteter som föreskrivs i denna budgetförordning inte iakttas. Räkenskapsföraren skall i så fall omedelbart underrätta utanordnaren och styrekonomen om att betalningen hålls inne och ange skälen till detta.
Om betalningen hålls inne får direktören på eget ansvar skriftligen begära att betalningen verkställs. Direktören skall i så fall vid nästa möte skriftligen underrätta styrelsen.
Artikel 20
1. Betalningar skall i princip verkställas via bank- eller postgirokonto, helst genom banköverföring eller, om det är motiverat, med check. Transaktionerna skall ske i euro, utom i välgrundade undantagsfall som godkänts av centrumet.
2. Checkar och bank- eller postgireringar skall undertecknas av två personer: räkenskapsföraren och utanordnaren eller ett ombud.
3. I välgrundade fall får direktören godkänna kontanta betalningar. För sådana betalningar skall ett kvitto erhållas.
4. Om inkomster och utgifter hanteras via dator, får undertecknandet ske på elektronisk väg.
5. Om uppgifter om faktiska valutakurser saknas, skall omräkningskursen för beräkningen i euro av de betalningar som skall göras eller de inkomster som skall mottas i lokal valuta i en AVS-stat vara den som gällde den första arbetsdagen i den månad under vilken den faktiska transaktionsdagen inföll, enligt vad som noterats av centrumets bank- eller postkontor.
Artikel 21
1. För betalning av vissa kategorier av utgifter, som fastställts genom tillämpningsföreskrifter för arbetsordningen, får förskottskonton inrättas i enlighet med de villkor som fastställs av centrumet.
2. Alla beslut om inrättande av ett förskottskonto skall fattas av direktören på grundval av ett förslag om åtagande från den handläggare som ansvarar för ärendet. Innan förslaget läggs fram för direktören skall det godkännas av räkenskapsföraren och styrekonomen.
3. I varje beslut om inrättande av ett förskottskonto skall följande anges:
a) Förskottsförvaltarens namn.
b) Den angivna förvaltarens ansvarsområde.
c) Det maximala belopp som får beviljas som förskott.
d) Slag och maximalt belopp för varje utgift som skall betalas.
e) Det sätt på vilket styrkande handlingar skall lämnas och tidsfristen för detta.
4. Utanordnaren och räkenskapsföraren skall vidta nödvändiga åtgärder för att beviljade förskott inom fastställda tidsfrister skall utfärdas för de exakta belopp det gäller.
Artikel 22
1. Direktören skall vara utanordnare för de anslag som tas upp i centrumets budget.
2. Direktören får delegera en del av sina uppgifter till underställd personal. I varje beslut om delegering av befogenheter skall det anges hur länge och hur omfattande uppdraget skall vara.
Artikel 23
1. Direktören skall utse en räkenskapsförare som skall ansvara för att
a) betalningar verkställs korrekt samt att inkomster uppbärs och fordringar betalas in,
b) sammanställa och redovisa räkenskaper i enlighet med artikel 25,
c) föra räkenskaper i enlighet med artikel 25,
d) genomföra regler och metoder för hur räkenskaperna skall föras samt genomföra kontoplanen på grundval av regler som utformats av kommissionens räkenskapsförare,
e) utforma och godkänna redovisningssystemen och, i förekommande fall, godkänna de system som fastställs av utanordnaren med syftet att leverera eller styrka bokföringsuppgifter,
f) förvalta likvida medel i samförstånd med direktören.
2. Räkenskapsföraren skall från utanordnaren få alla de uppgifter som krävs för att sammanställa räkenskaper som ger en rättvisande bild av centrumets tillgångar och skulder och budgetgenomförande, varvid utanordnaren skall ansvara för de lämnade uppgifternas tillförlitlighet.
3. I enlighet med punkt 1 och artikel 21 skall endast räkenskapsföraren ha befogenhet att förvalta finansiella medel och andra tillgångar. Räkenskapsföraren skall ansvara för förvaringen av medlen och tillgångarna.
4. Vid utförandet av sina arbetsuppgifter och med direktörens samtycke får räkenskapsföraren delegera vissa uppgifter till tjänstemän vid centrumet som är direkt underställda räkenskapsföraren. I den handling genom vilken delegeringen sker skall de uppgifter anges som överlåts på dessa personer liksom deras rättigheter och skyldigheter.
Artikel 24
1. För inkassering av en fordran till centrumet skall ett betalningskrav utfärdas av utanordnaren. Betalningskrav skall godkännas av styrekonomen.
2. Räkenskapsföraren skall ansvara för betalningskrav som utanordnaren överlämnat till honom.
3. För alla kontanta betalningar till räkenskapsföraren eller förskottsförvaltaren skall ett kvitto utfärdas.
KAPITEL VI
RÄKENSKAPER, UPPRÄTTANDE OCH KONTROLL AV BOKSLUT, REVISION, REVISIONSRÄTTEN, OLAF
Artikel 25
1. Räkenskaperna skall föras i euro enligt metoden för dubbel bokföring och på grundval av kalenderåret. De skall visa samtliga inkomster och utgifter från och med den 1 januari till och med den 31 december varje år och inbegripa styrkande handlingar i original.
Räkenskaperna skall avslutas vid utgången av budgetåret för att centrumets årsbokslut skall kunna upprättas.
2. Bokföringsposter skall registreras på grundval av ett redovisningssystem som omfattar en kontoplan, i vilken en klar åtskillnad görs mellan de konton som skall användas för upprättandet av balansräkningen och de konton som skall användas för upprättandet av inkomst- och utgiftsredovisningen. Dessa poster skall införas i böcker eller på kort med hjälp av vilka en samlad månatlig balansställning kan uppställas. Alla förskottsbetalningar skall bokföras på ett bevakningskonto och regleras senast vid utgången av det följande budgetåret, utom när det gäller stående förskott.
3. Centrumet skall senast den 30 april år N+1 upprätta en balansräkning och en inkomst- och utgiftsredovisning.
Balansräkningen skall visa centrumets tillgångar och skulder per den 31 december det senast utlöpta budgetåret.
Inkomst- och utgiftsredovisningen skall omfatta följande:
a) En tabell över "inkomster" som omfattar:
- Beräknade inkomster under kalenderåret.
- Ändringar när det gäller beräknade inkomster.
- Fordringar som uppkommer under kalenderåret.
- Belopp som skall betalas in i slutet av kalenderåret.
- Ytterligare inkomster.
b) En tabell över "utgifter" som omfattar:
- En sammanfattande tabell över anslag som avsatts för åtaganden, anslag som överförts från år N och förfallna anslag.
- En sammanfattande tabell över anslag som överförts från år N-1 och förfallna anslag.
- En tabell med en samlad översikt över åtaganden och godkännanden för år N.
- En tabell med en samlad översikt över åtaganden och godkännanden för anslag som överförts från år N-1.
c) Anmärkningar till bokslutet som omfattar:
- Tillämpade redovisningsprinciper.
- Noggranna anmärkningar och beräkningar som förklarar de enskilda posterna i bokslutet.
- Förklaringar som krävs för att säkerställa öppenhet och insyn i räkenskaperna.
4. Varje kvartal skall det utarbetas och översändas till ambassadörskommittén en redovisning som visar situationen när det gäller genomförandet av den löpande budgeten och användningen av överförda anslag; denna redovisning skall godkännas av styrekonomen och överlämnas till styrelsen.
Artikel 26
1. På rekommendation av centrumets direktör och på grundval av ett anbudsförfarande skall styrelsen utse en internationellt ansedd revisionsbyrå för en period av högst tre år.
2. Revisorerna skall granska centrumets böcker och kassaförvaltning, kontrollera att inventarieförteckningar och balansräkningar har upprättats på ett korrekt sätt och i god tro samt förvissa sig om att uppgifterna om centrumets räkenskaper är korrekta.
3. Syftet med revisionen, som skall bygga på bokföringsmaterial och vid behov ske på platsen, skall vara att fastställa att alla inkomster har uppburits och alla utgifter uppkommit på ett lagligt och korrekt sätt och att den ekonomiska förvaltningen har varit sund.
4. Revisorerna skall intyga att bokslutet är uppställt korrekt och i enlighet med internationella redovisningsstandarder och att det ger en sann och rättvisande översikt av centrumets finansiella ställning.
5. Revisorerna skall utarbeta en rapport senast den 30 juni efter varje budgetårs slut. Rapporten skall överlämnas till direktören, som skall vidarebefordra den med sina eventuella kommentarer till styrelsen, som skall lägga fram den för ambassadörskommittén med sina rekommendationer.
På grundval av denna rapport och bokslutet skall ambassadörskommittén bevilja direktören ansvarsfrihet när det gäller genomförandet av budgeten.
6. Revisorerna skall ge råd till centrumet när det gäller riskhanteringen genom att lämna oberoende omdömen om förvaltningens och kontrollsystemens kvalitet och genom att utfärda rekommendationer för förbättring av villkoren för genomförandet av transaktioner och främjande av en sund ekonomisk förvaltning.
Revisorerna skall vara ansvariga för
a) bedömningen av de interna förvaltningssystemens lämplighet och effektivitet samt av centrumets arbete när det genomför program och vidtar de åtgärder som krävs, mot bakgrund av de därmed förbundna riskerna,
och
b) bedömningen av lämplighet och kvalitet när det gäller de interna kontrollsystemen för budgetens genomförande.
7. Revisorerna skall granska all verksamhet som utförs av centrumet samt alla dess enheter. De skall ha fullt och obegränsat tillträde till all information som behövs för att de skall kunna utföra sina uppgifter.
Artikel 27
I enlighet med budgetförordningen för nionde EUF får kommissionen (på gemenskapens vägnar), revisionsrätten och Europeiska byrån för bedrägeribekämpning (Olaf) kontrollera användningen av de medel som centrumet mottagit från EUF.
Revisionsrätten får kontrollera att inkomsterna och utgifterna är lagliga och formellt korrekta och att bestämmelserna i avtalet och i budgetförordningen för nionde EUF har följts.
KAPITEL VII
UTANORDNARES, RÄKENSKAPSFÖRARES OCH FÖRSKOTTSFÖRVALTARES ANSVAR
Artikel 28
Disciplinära åtgärder och vid behov krav på ekonomisk kompensation kan riktas mot utanordnare som fastställer fordringar, utfärdar betalningskrav, gör utgiftsåtaganden eller undertecknar betalningsorder utan att följa denna budgetförordning. Detsamma gäller om utanordnare försummar att upprätta ett dokument som fastställer en skuld eller om de utan giltig orsak försummar att utfärda ett betalningskrav eller utfärdar dessa dokument för sent.
Ett sådant ansvar får endast åberopas gentemot utanordnaren om uppsåt eller allvarlig försumlighet från dennes sida har orsakat detta fel.
Artikel 29
1. Disciplinära åtgärder och vid behov krav på ekonomisk kompensation kan riktas mot en räkenskapsförare som gör betalningar i strid med artikel 19.
Disciplinära åtgärder och krav på ekonomisk kompensation kan riktas mot räkenskapsföraren på grund av förlust eller skada i fråga om de medel, tillgångar och dokument som han ansvarar för, om uppsåt eller allvarlig försumlighet från hans sida har orsakat denna förlust eller skada.
Räkenskapsföraren skall på samma villkor vara ansvarig för att de order han får beträffande användning och förvaltning av bankkonton blir korrekt utförda, särskilt i följande fall:
a) Om inbetalda belopp eller gjorda utbetalningar inte överensstämmer med beloppen på motsvarande betalningskrav eller betalningsorder.
b) Om de betalar till en annan person än den berättigade betalningsmottagaren.
2. Disciplinära åtgärder och vid behov krav på ekonomisk kompensation skall riktas mot förskottsförvaltare i följande fall:
a) Om de inte med formellt korrekta dokument kan styrka betalningar de gjort.
b) Om de betalar till en annan person än den berättigade betalningsmottagaren.
Disciplinära åtgärder och krav på ekonomisk kompensation skall riktas mot förskottsförvaltare på grund av förlust eller skada i fråga om de medel, tillgångar och dokument som de ansvarar för, om denna förlust eller skada har orsakats av uppsåt eller allvarlig försumlighet från deras sida.
Artikel 30
1. Räkenskapsförare och förskottsförvaltare skall vara försäkrade mot de risker som avses i artikel 29.
Centrumet skall täcka de försäkringskostnader som därigenom uppstår. Det skall ange vilka tjänstemän som fungerar som räkenskapsförare och förskottsförvaltare och de villkor på vilka det kommer att täcka denna personals kostnader för att försäkra sig mot de risker som är förenade med deras uppgifter.
2. Särskilda bidrag skall beviljas räkenskapsförare och förskottsförvaltare. Nivån på dessa bidrag skall fastställas i bestämmelser som utarbetas av centrumet och godkänns av styrelsen. Ett belopp motsvarande detta bidrag skall varje månad tillföras ett konto som öppnas av centrumet för var och en av dessa tjänstemäns räkning i syfte att skapa en garantifond som skall täcka eventuella brister i kassa eller bank som den berörda personen skulle kunna göras ansvarig för, i den mån sådana brister inte täcks genom ersättning från försäkringsbolag.
Tillgodohavandet på dessa garantikonton skall betalas ut till de berörda personerna när deras uppdrag som räkenskapsförare eller förskottsförvaltare upphör och efter det att de har beviljats slutgiltig ansvarsfrihet för sin förvaltning.
3. Direktören skall på grundval av de externa revisorernas rapport bevilja räkenskapsföraren och förskottsförvaltaren ansvarsfrihet inom två år efter framläggandet av årsbokslutet för ambassadörskommittén.
Artikel 31
De krav på ekonomisk kompensation och de disciplinära åtgärder som kan riktas mot utanordnare, räkenskapsförare och förskottsförvaltare skall fastställas i enlighet med centrumets tjänsteföreskrifter.
Artikel 32
Tjänstemän får när det gäller budgetens genomförande inte vidta några åtgärder i de fall deras egna intressen skulle kunna strida mot centrumets intressen. Om en sådan situation uppstår skall den berörda tjänstemannen avstå från alla handlingar och vända sig till sin överordnade.
En intressekonflikt skall anses föreligga om en tjänsteman i samband med budgetens genomförande av familjeskäl eller på grund av personliga förhållanden, på grund av nationell eller politisk koppling eller av ekonomiskt intresse eller varje annat gemensamt intresse med mottagaren, inte kan utföra sina arbetsuppgifter på ett opartiskt och objektivt sätt.
KAPITEL VIII
ALLMÄNNA BESTÄMMELSER OCH SLUTBESTÄMMELSER
Artikel 33
Tilldelning av kontrakt skall ske i enlighet med de allmänna bestämmelser för upphandling av varor, tjänster och byggentreprenader som fastställts genom AVS-EG-ministerrådets beslut nr 2/2002 av den 7 oktober 2002 om genomförande av artiklarna 28, 29 och 30 i bilaga IV till Cotonouavtalet [4].
På vilket sätt de ovannämnda allmänna bestämmelserna skall genomföras skall fastställas i interna föreskrifter som skall godkännas av styrelsen efter yttrande av kommissionen.
Artikel 34
1. Centrumet får också förvalta medel på tredje parts vägnar, i enlighet med sitt uppdrag. Förteckningen över dessa medel skall tas upp i en bilaga till centrumets budget.
2. Dessa medel skall förvaltas i enlighet med denna budgetförordning.
3. Separata räkenskaper skall föras över förvaltningen av dessa medel på tredje parts vägnar.
4. Årsboksluten för var och en av de fonder som förvaltas av centrumet på tredje parts vägnar skall omfatta en balansräkning och en inkomst- och utgiftsredovisning, i vilka situationen per den 31 december det berörda budgetåret anges. De skall attesteras i enlighet med bestämmelserna i det avtal som ingåtts mellan centrumet och den tredje parten.
Om det inte finns några sådana bestämmelser skall attesteringen göras av centrumets externa revisorer.
5. Dessa årsbokslut skall utgöra en bilaga till centrumets årsbokslut.
Artikel 35
1. En löpande inventarieförteckning skall föras över all lös och fast egendom som tillhör centrumet. Endast lös egendom till ett värde av minst 350 EUR skall införas i förteckningen. Löpnumret i förteckningen skall anges på varje faktura innan denna betalas.
2. All försäljning av lös egendom och utrustning vars anskaffningsvärde per enhet översteg 350 EUR skall offentliggöras på lämpligt sätt.
3. En rapport som undertecknats av både direktören och den person som ansvarar för utrustningen skall upprättas närhelst en artikel i inventarieförteckningen avyttras, skrotas eller konstateras saknad på grund av förlust eller stöld eller annat skäl.
4. Den fysiska och den bokföringsmässiga inventarieförteckningen skall avstämmas i slutet av varje budgetår. Avstämningen skall godkännas av de externa revisorerna.
Artikel 36
AVS-staterna, medlemsstaterna och gemenskapen skall, var och en i den mån parten berörs, vidta de åtgärder som krävs för att genomföra detta beslut.
Artikel 37
Den budgetförordning för centrumet som godkänns i AVS–EG-ambassadörskommitténs beslut nr 2/91 av den 19 april 1991 skall upphöra att gälla.
Artikel 38
Detta beslut träder i kraft samma dag som det antas.
RÅDETS DIREKTIV av den 4 juni 1974 om att uppnå etableringsfrihet och frihet att tillhandahålla tjänster som egenföretagare och agent inom handel med och distribution av giftiga ämnen (74/557/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 54.2, 54.3, 63.2 och 63.3 i detta,
med beaktande av Allmänna handlingsprogrammet för upphävande av begränsningar av etableringsfriheten (1), särskilt avdelning IV A och C i detta,
med beaktande av Allmänna handlingsprogrammet för upphävande av begränsningar av friheten att tillhandahålla tjänster (2), särskilt avdelning V C i detta,
med beaktande av rådets direktiv 64/223/EEG (3) av den 25 februari 1964 om att uppnå etableringsfrihet och frihet att tillhandahålla tjänster inom partihandel,
med beaktande av rådets direktiv 64/224/EEG (4) av den 25 februari 1964 om att uppnå etableringsfrihet och frihet att tillhandahålla tjänster som agent inom handel, industri och hantverk,
med beaktande av rådets direktiv 68/363/EEG (5) av den 15 oktober 1968 om att uppnå etableringsfrihet och frihet att tillhandahålla tjänster som egenföretagare inom detaljhandel, med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande (6),
med beaktande av Ekonomiska och sociala kommitténs yttrande (7), och
med beaktande av följande:
I de allmänna handlingsprogrammen påpekas att all särbehandling som grundar sig på nationalitet skall upphävas i fråga om etablering och erbjudande av tjänster - vad gäller partihandel eller agenturverksamhet inom handel, industri och hantverk före utgången av andra året av andra etappen,
- vad gäller detaljhandel efter utgången av andra året av övergångsperiodens andra etapp och före utgången av andra etappen.
Direktiven 64/223/EEG, 64/224/EEG och 68/363/EEG tillämpas inte på området giftiga ämnen som på grund av de särskilda problem som uppstår på grund av skyddet av den allmänna hälsan regleras genom bestämmelser i medlemsstaternas lagar och andra författningar.
De ovannämnda direktiven 64/223/EEG och 68/363/EEG tillämpas inte heller på former av verksamhet inom partihandel, agenturverksamhet och detaljhandel med sjukdomsalstrande ämnen. Bortsett från de sjukdomsalstrande ämnen som är klassificerade som medicinska preparat för användning på människor och djur i den bemärkelse som avses i rådets direktiv 65/65/EEG (8) av den 26 januari 1965 om tillnärmning av bestämmelserna i lagar och andra författningar rörande medicinska produkter med ändringar i direktiv 66/454/EEG (9) omfattas emellertid endast de sjukdomsalstrande ämnen som betecknas som %quot%biologiska bekämpningsmedel för användning inom jordbruket%quot% av de nämnda verksamhetsformerna. I fråga om sjukdomsalstrande ämnen kan därför upphävandet av begränsningar av friheten att erbjuda tjänster och friheten att etablera sig begränsas till att omfatta handel med och distribution av de nämnda bekämpningsmedlen.
Det förefaller vara både önskvärt och lämpligt att vidta åtgärder för att på gemenskapsnivå reglera de områden som avses i ovanstående stycken med avseende på den farliga inverkan som giftiga ämnen kan ha på människors, djurs och växters hälsa antingen direkt eller indirekt genom den omgivande miljön. Agenturverksamhet inom handel, industri och hantverk omfattas av direktiven 64/224/EEG och 68/363/EEG. Agenturverksamhet vad gäller giftiga ämnen och sjukdomsalstrande ämnen är undantagna från dessa direktivs räckvidd. Syftet med det här direktivet är att även liberalisera dessa former av agenturverksamhet; följaktligen omfattar begreppen %quot%handel och distribution%quot% i det här direktivet även agenturverksamhet på dessa områden.
I Allmänna handlingsprogrammet för upphävande av begränsningar av etableringsfriheten föreskrivs att begränsningar av rätten att ansluta sig till yrkes- eller handelsorganisationer skall upphävas i de fall då vederbörandes yrkesverksamhet oundvikligen medför att denna rätt utövas.
Den ställning som tillkommer anställda, vilka medföljer den som erbjuder tjänster eller utför arbete för dennes räkning, kommer att regleras genom bestämmelser som fastställts i enlighet med artikel 48 och 49 i fördraget.
Särskilda direktiv har antagits eller kommer att antas, som är tillämpliga på alla former av verksamhet som egenföretagare, med bestämmelser om förmånstagarnas fria rörlighet och vistelse och, där så krävs, ett direktiv om samordning av de garantier som i medlemsstaterna avkrävs bolag och enskilda firmor till skydd för medlemsstaternas och tredje mans intressen.
I vissa medlemsstater regleras handel, distribution och yrkesmässig användning av giftiga ämnen genom bestämmelser om rätten att påbörja den hanteringen medan andra stater där så är nödvändigt kommer att tillämpa sådana regler. Därför behandlas vissa speciella övergångsåtgärder, vars syfte är att underlätta för medborgare i andra medlemsstater att påbörja och utöva verksamhet inom handel med giftiga ämnen, i ett särskilt direktiv.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Medlemsstaterna skall i fråga om de fysiska personer och bolag eller enskilda firmor (här nedan kallade förmånstagarna) som nämns i avdelning I i de allmänna handlingsprogrammen för upphävande av begränsningar av etableringsfriheten och friheten att tillhandahålla tjänster upphäva de begränsningar som avses i avdelning III i dessa handlingsprogram, vilka påverkar rätten att påbörja och utöva den verksamhet som närmare anges i artikel 2 i detta direktiv.
Artikel 2
1. Detta direktiv skall tillämpas på verksamhet som egenföretagare inom handel med och distribution av giftiga ämnen (substanser och preparat) och biologiska bekämpningsmedel för användning inom jordbruket som har undantagits från tillämpningen av direktiv 64/223/EEG genom artikel 2.1 i detta, av direktiv 64/224/EEG, genom artikel 4.1 femte strecksatsen i detta och av direktiv 68/363/EEG genom artikel 2.1 i detta.
2. De varor som avses i punkt 1 är på grund av den farliga inverkan de kan ha på människors, djurs och växters hälsa allt efter medlemsstaternas lagstiftningar underkastade särskilda direktiv (varorna i fråga finns uppräknade i bilagan). De ändringar i denna förteckning som en medlemsstat gör skall anmälas till kommissionen som kommer att underrätta medlemsstaterna om detta.
3. Detta direktiv skall inte tillämpas på handel med och distribution av de medicinska varor som finns definierade i direktiv 65/65/EEG eller på handelsresande, gatuförsäljare eller gårdfarihandlare.
Artikel 3
1. Begränsningarna i fråga om de former av verksamhet som anges i artikel 2 skall upphävas oavsett den benämning som används på personer som utövar någon av dessa verksamhetsformer.
2. De vanliga benämningar som för närvarande används i medlemsstaterna för att definiera personer som utövar någon form av verksamhet som agent inom handel är de som finns uppräknade i artikel 3 i rådets direktiv 64/224/EEG.
Artikel 4
1. Medlemsstaterna skall i synnerhet upphäva de begränsningar som a) hindrar förmånstagarna från att etablera sig eller erbjuda tjänster i värdlandet på samma villkor och med samma rättigheter som medborgarna i den staten,
b) härrör från en förvaltningspraxis som innebär att förmånstagarna utsätts för särbehandling jämfört med medborgarna i staten i fråga.
2. Till de begränsningar som skall upphävas hör i synnerhet de som härrör från åtgärder som hindrar eller begränsar förmånstagarnas möjligheter att etablera sig eller erbjuda tjänster på följande sätt: a) I Belgien:
- skyldigheten att inneha ett carte professionnelle (artikel 1, lagen av den 19 februari 1965). b) I Frankrike:
- skyldigheten att inneha ett carte d'identité d'étranger commerçant (décret-loi av den 12 november 1938, décret av den 2 februari 1939, lagen av den 8 oktober 1940, lagen av den 10 april 1954, décret nr 59-852 av den 9 juli 1959),
- uteslutning från rätten att förnya arrendeavtal (artikel 38 i décret av den 30 september 1953).
c) I Luxemburg:
- den begränsade giltighetstiden för tillstånd som beviljas utländska medborgare (artikel 21 i lagen av den 2 juni 1962).
Artikel 5
1. Medlemsstaterna skall se till att förmånstagarna har rätt att ansluta sig till yrkes- eller handelsorganisationer på samma villkor och med samma rättigheter och skyldigheter som de egna medborgarna.
2. Vid etablering skall rätten att ansluta sig till yrkes- eller handelsorganisationer medföra möjlighet att inneha uppdrag inom sådana organisationer. Dessa uppdrag kan dock förbehållas de egna medborgarna, då organisationen i fråga har myndighetsutövande uppgifter i enlighet med en lag eller en förordning.
3. I Luxemburg skall medlemskap i Chambre de commerce eller Chambre des métiers inte medföra rätt för de förmånstagare som omfattas av detta direktiv att delta i valet av förvaltningsorgan inom dessa handelskammare.
Artikel 6
Medlemsstaterna får inte ge de egna medborgare som beger sig till en annan medlemsstat i syfte att där utöva sådan verksamhet enligt artikel 2, något stöd som kan snedvrida etableringsvillkoren.
Artikel 7
1. I de fall då ett värdland av de egna medborgare, som vill påbörja någon form av verksamhet enligt i artikel 2, kräver skötsamhetsbevis och bevis att de inte har varit försatta i konkurs eller ettdera av dessa bevis, skall den staten i fråga om medborgare i andra medlemsstater som tillräckligt bevis på detta godta utdrag ur kriminalregistret eller, om något sådant intyg inte kan uppvisas, motsvarande handling utfärdad av behörig rättsinstans eller förvaltningsmyndighet i utlänningens ursprungsland eller senaste hemvistland, av vilken framgår att dessa villkor är uppfyllda.
2. I de fall då det i ett värdland på de egna medborgarna ställs särskilda krav på god vandel för att kunna utöva någon form av verksamhet enligt artikel 2 och bevis på att dessa krav är uppfyllda inte kan erhållas genom den handling som avses i punkt 1 skall den staten vad gäller medborgare i andra medlemsstater som tillräckligt bevis på detta godta intyg utfärdat av behörig rättsinstans eller förvaltningsmyndighet i utlänningens ursprungsland eller senaste hemvistland, av vilken framgår att dessa villkor är uppfyllda. Ett sådant intyg skall hänföra sig till vissa bestämda fakta som av värdlandet betraktas som relevanta.
3. I de fall då det i utlänningens ursprungsland eller senaste hemvistland inte utfärdas någon sådan handling som avses i punkt 1 eller det intyg som avses i punkt 2 om god vandel eller om att denne inte har varit försatt i konkurs, kan ett sådant bevis ersättas av en försäkran under ed eller, i de stater där detta inte förekommer, av en förklaring på heder och samvete som avgivits inför behörig rättsinstans eller förvaltningsmyndighet eller, där så är lämpligt, inför notarius publicus i utlänningens ursprungsland eller senaste hemvistland; sådan myndighet eller notarius publicus utfärdar ett intyg som styrker äktheten av försäkran under ed eller förklaringen på heder och samvete. En förklaring om att vederbörande inte varit försatt i konkurs kan även avges inför behörig yrkes- eller handelsorganisation i samma land.
4. Handlingar som utfärdats i överensstämmelse med punkt 1 och 2 får inte vara äldre än tre månader.
5. Medlemsstaterna skall inom den tid som anges i artikel 8 utse de myndigheter och organ som är behöriga att utfärda de handlingar som avses i punkt 1 och 2 och genast underrätta övriga medlemsstater och kommissionen om detta.
6. I de fall då bevis om den ekonomiska ställningen krävs i värdlandet skall den staten betrakta intyg som utfärdats av banker i utlänningens ursprungsland eller senaste hemvistland som likvärdiga med intyg som utfärdats inom dess eget territorium.
Artikel 8
Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att följa detta direktiv inom sex månader efter dagen för anmälan och skall genast underrätta kommissionen om detta.
Artikel 9
Detta direktiv riktar sig till medlemsstaterna.
KOMMISSIONENS FÖRORDNING (EEG) nr 2182/77 av den 30 september 1977 om närmare bestämmelser för försäljning av fryst nötkött från interventionslager avsett för bearbetning inom gemenskapen och om ändring av förordning (EEG) nr 1687/76
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 805/68 av den 27 juni 1968 om gemensam organisation av marknaden för nötkött(1), senast ändrad genom förordning (EEG) nr 425/77(2), särskilt artikel 7.3 i denna, och
med beaktande av följande: I rådets förordning (EEG) nr 98/69 av den 16 januari 1969 om allmänna bestämmelser för interventionsorgans avyttring av fryst nötkött(3), senast ändrad genom förordning (EEG) nr 429/77(4), fastställs att sådant kött får säljas om det är avsett för särskild användning. Närmare bestämmelser för avyttring till gemenskapens förädlingsindustri bör fastställas.
I kommissionens förordning (EEG) nr 597/77 av den 18 mars 1977 om tillämpningsföreskrifter för särskilda importordningar för vissa typer av fryst nötkött avsett för bearbetning(5), senast ändrad genom förordning (EEG) nr 1384/77(6), anges de produkter som får framställas genom sådan bearbetning. För att underlätta kontrollen av denna bearbetning bör det fastställas att de produkter som säljs enligt den här förordningen skall bearbetas till de produkter som anges i förordning (EEG) nr 597/77, eller till produkter som omfattas av undernummer 02.06 C 1 a 2 i Gemensamma tulltaxan.
I förordning (EEG) nr 597/77 fastställs dessutom en gynnsammare ordning för kött som skall bearbetas till konserver, för att förbättra sådana konservers konkurrenskraft på marknaden. Det bör fastställas att det kött som avyttras enligt den här förordningen skall säljas till priser som varierar beroende på slutanvändningen.
Försäljning enligt den här förordningen till förutfastställda priser bör regleras av bestämmelserna i kommissionens förordning (EEG) nr 216/69 av den 4 februari 1969 om närmare bestämmelser för avyttring av fryst nötkött som köpts upp av interventionsorgan(7), med vissa särskilda undantag med hänsyn till den specifika användning som dessa produkter är avsedda för.
Förutom den säkerhet som fastställs i artikel 4 i förordning (EEG) nr 216/69 bör det fastställas att en säkerhet skall ställas som garanti för användningen av de produkter som säljs enligt denna förordning. Denna säkerhet bör variera beroende på hur köttet används.
I kommissionens förordning (EEG) nr 1687/76 av den 30 juni 1976(8), senast ändrad genom förordning (EEG) nr 1723/77(9), fastställs närmare bestämmelser för kontroll av interventionsprodukternas användning eller bestämmelseort. Vissa av dessa bestämmelser bör anpassas till försäljning enligt denna förordning.
Enligt artikel 4.2 i rådets förordning (EEG) nr 1134/68 av den 30 juli 1968 om tillämpningsföreskrifter för förordning (EEG) nr 653/68 om villkoren för ändring av värdet på den beräkningsenhet som används inom den gemensamma jordbrukspolitiken(10) skall de belopp, uttryckta i nationell valuta och motsvarande belopp fastställda i beräkningsenheter, som en medlemsstat eller en behörig myndighet är skyldig för transaktioner som genomförs i enlighet med gemenskapens jordbrukspolitik, betalas med utgångspunkt i det förhållande mellan beräkningsenheten och den nationella valutan som gällde då transaktionen eller en del av transaktionen genomfördes.
Med den tidpunkt då transaktionen genomförs avses enligt artikel 6 i förordningen ovan den dag då den händelse inträffar, som leder till att transaktionsbeloppet förfaller till betalning, i enlighet med definitionen i gemenskapens regler, eller i avvaktan på sådana regler, enligt den berörda medlemsstatens regler. Den händelse som leder till att produkternas säkerhet och försäljningspris förfaller till betalning inträffar den dag då köpeavtalet ingås.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för nötkött.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Kött som säljs enligt denna förordning skall användas till tillverkning inom gemenskapen enligt köparens val av antingen a) konserver enligt definitionen i artikel 1.5 i förordning (EEG) nr 597/77, eller
b) andra produkter enligt definitionen i artikel 1.6 i samma förordning eller produkter som omfattas av undernummer 02.06 C I a 2 i Gemensamma tulltaxan.
2. För fryst kött som bearbetas till de produkter som anges i punkt 1 a skall bevis på bearbetning endast godtas om kvantiteten konserver som tillverkats av sådant kött minst motsvarar den inköpta kvantiteten.
Koefficienterna för fastställande av kvantiteten urbenat fryst kött som en viss kvantitet konserverat kött innehåller fastställs i bilagan till denna förordning.
3. Vid tillämpningen av denna förordning anses 100 kg kött med ben motsvara 77 kg urbenat kött.
Vad gäller framkvartsparter anses dock 100 kg framkvartsparter med ben motsvara 70 kg urbenat kött.
Artikel 2
Olika försäljningspriser får fastställas för kött som säljs enligt denna förordning, beroende på om köttet är avsett för tillverkning av sådan konserver som avses i artikel 1.1 a eller för tillverkning av sådana andra produkter som avses i artikel 1.1 b.
Artikel 3
1. Ansökningar om köp eller anbud måste innehålla en skriftlig försäkran från köparen att köttet är avsett för tillverkning av produkterna i artikel 1.1 a eller 1.1 b, och måste ange den eller de medlemsstater där tillverkningen skall äga rum.
2. Innan köpeavtalet ingås måste köparen lämna en skriftlig försäkran till den berörda myndigheten i den medlemsstat där bearbetningen skall äga rum, att han inom 30 dagar efter det att avtalet ingås skall ange den eller de anläggningar där det inköpta köttet skall bearbetas.
3. När artikel 13.3 i förordning (EEG) nr 1687/76 tillämpas skall det interventionsorgan som innehar produkterna utan dröjsmål informera den berörda myndigheten i den medlemsstat där bearbetningen skall äga rum om det datum då avtalet ingicks.
Artikel 4
1. Innan köpeavtalet ingås skall en säkerhet för att garantera att produkterna bearbetas ställas till den berörda myndigheten i den medlemsstat där bearbetningen skall äga rum. Den skall ställas i den medlemsstatens nationella valuta.
Säkerhetsbeloppet får variera med hänsyn till de produkter som utbjuds till försäljning och deras användning.
2. När artikel 13.3 i förordning (EEG) nr 1687/76 tillämpas får avtal inte ingås förrän det interventionsorgan som innehar produkterna har mottagit det intyg som avses i det stycket.
Artikel 5
1. Bearbetningen av kött som köpts enligt denna förordning måste genomföras inom fyra månader från den dag då avtalet ingicks.
2. Det bevis som avses i artikel 12 i förordning (EEG) nr 1687/76 måste lämnas in inom fem månader från den dag då avtalet ingicks.
3. För att säkerheten skall frisläppas enligt artikel 4.1 krävs att det bevis som avses i stycke 2 framläggs och att övriga villkor i denna förordning är uppfyllda.
4. Den säkerhet som avses i artikel 4.1 skall frisläppas omedelbart om ansökan om köp avslås, i proportion till de kvantiteter för vilka avtal inte ingås.
Artikel 6
1. Genom undantag från artikel 5.1 i förordning (EEG) nr 216/69 skall priset betalas efterhand som varorna tas ut från lagret, i proportion till de kvantiteter som tas ut och senast dagen före den dag då varorna tas ut.
2. Priset skall betalas i den nationella valutan i den medlemsstat där interventionsorganet som innehar produkterna är beläget.
3. Genom undantag från artikel 2.2 i förordning (EEG) nr 216/69 skall den minsta tillåtna försäljningskvantiteten uppgå till 10 ton.
Artikel 7
Om köparen på grund av force majeure inte kan iaktta den tidsfrist som fastställts för övertagandet, skall interventionsorganet vidta de åtgärder som det finner nödvändigt med hänsyn till omständigheterna.
Interventionsorganet skall meddela kommissionen varje fall av force majeure och de åtgärder som vidtas på grund av detta.
Artikel 8
Den avgörande händelse som avses i artikel 6 i förordning (EEG) nr 1134/68, då den säkerhet som avses i artikel 4.1 och försäljningspriset förfaller till betalning, skall anses inträffa den dag då köpeavtalet ingås.
Artikel 9
I bilagan till förordning (EEG) nr 1687/76 skall följande punkt 17 med tillhörande fotnot läggas till efter punkt 16 under rubriken %quot%II Produkter avsedda för annan användning eller bestämmelseort än de som avses i I%quot%:
%quot%17. Kommissionens förordning (EEG) nr 2182/77 av den 30 september 1977 om närmare bestämmelser för försäljning av fryst nötkött från interventionslager avsett för bearbetning inom gemenskapen och om ändring av förordning (EEG) nr 1687/76(8): a) kött avsett för tillverkning av konserver:
- ruta 104: %quot%Meat intended for the manufacture of preserved food.
System (a) (Regulation (EEC) No 2182/77)%quot%.
%quot%Kød bestemt til femstilling af konserves.
Ordning (a) (Forordning (EØF) nr. 2182/77)%quot%.
%quot%Fleisch zur Herstellung von Konserven bestimmt.
Regelung (a) (Verordnung (EWG) Nr. 2182/77)%quot%.
%quot%Viandes destinées à la fabrication de conserves.
Régime (a) (Règlement (CEE) n° 2182/77)%quot%.
%quot%Carni destinate alle fabbricazione di conserve.
Regime (a) (Regolamento (CEE) n. 2182/77)%quot%.
%quot%Vlees bestemd voor de vervaardiging van conserve.
Regeling (a) (Verordening (EEG) nr. 2182/77)%quot%.
- ruta 106:
Dagen då avtalet ingås.
b) kött avsett för tillverkning av andra produkter: - ruta 104:
%quot%Meat intended for processing.
System (b) (Regulation (EEC) No 2182/77)%quot%.
%quot%Kød bestemt till forarbejdning.
Ordning (b) (Forordning (EØF) nr. 2182/77)%quot%.
%quot%Zur Verarbeitung bestimmtes Fleisch.
Regelung (b) (Verordnung (EWG) Nr. 2182/77)%quot%.
%quot%Viandes destinées à la transformation.
Régime (b) (Règlement (CEE) n° 2182/77)%quot%.
%quot%Carni destinate alle trasformazione.
Regime (b) (Regolamento (CEE) n. 2182/77)%quot%.
%quot%Vlees bestemd voor de verwerking.
Regeling (b) (Verordening (EEG) nr. 2182/77)%quot%.
- ruta 106:
Dagen då avatalet ingås.
(8) EGT nr L 251, 1.10.1977, s. 60.%quot%
Artikel 10
Denna förordning träder i kraft den 10 oktober 1977.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS FÖRORDNING (EEG) nr 3026/77 av den 28 november 1977 om upprättandet av ett tilläggsprotokoll till avtalet om association mellan Europeiska ekonomiska gemenskapen och Turkiet till följd av nya medlemsstaters anslutning till gemenskapen
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 238 i detta,
med beaktande av avtalet om anslutning av nya medlemsstater till Europeiska ekonomiska gemenskapen och till Europeiska atomenergigemenskapen undertecknat den 22 januari 1972, särskilt artikel 108 i härtill bifogad akt, med beaktande av kommissionens rekommendation,
med beaktande av Europaparlamentets yttrande(1), och
med beaktande av följande:
Det är lämpligt att upprätta ett tilläggsprotokoll som fastställer vissa villkor rörande avtalet om association mellan Europeiska ekonomiska gemenskapen och Turkiet till följd av nya medlemsstaters anslutning till Europeiska ekonomiska gemenskapen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Tilläggsprotokollet till avtalet om association mellan Europeiska ekonomiska gemenskapen och Turkiet till följd av nya medlemsstaters anslutning till gemenskapen samt de förklaringar som bifogats slutakten upprättas härmed och godkänns på gemenskapens vägnar. Texten till protokollet och slutakten bifogas denna förordning.
Artikel 2
Rådets ordförande skall underrätta den andra avtalsparten om att de förfaranden som behövs för att protokollet skall träda i kraft har fullföljts för gemenskapens del(2).
Artikel 3
Denna förordning träder i kraft tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EEG) nr 2077/80 av den 1 augusti 1980 om ändring av förordning (EEG) nr 2973/79 om fastställande av tillämpningsföreskrifter för beviljande av bistånd vid export av nötköttsprodukter som kan komma i fråga för förmånsbehandling vid import till tredje land
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 805/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för nötkött(), senast ändrad genom förordning (EEG) nr 2916/79(), särskilt artikel 15.2 i denna,
med beaktande av rådets förordning (EEG) nr 2931/79 av den 20 december 1979 om beviljande av bistånd vid export av jordbruksprodukter som kan komma i fråga för förmånsbehandling vid import till tredje land(), särskilt artikel 1.2 i denna, och
med beaktande av följande: I kommissionens förordning (EEG) nr 2973/79() fastställs närmare föreskrifter för genomförandet av en årlig export till USA på 5 000 ton nötkött som kan komma i fråga för förmånsbehandling.
I artikel 1.2 i förordningen anges att köttet måste komma från djur som slaktats högst en månad före tullklareringen för export. Denna tid har visat sig vara för kort med tanke på de logistiska förutsättningarna och det är därför lämpligt att förlänga den till två månader.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för nötkött.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 1.2 i förordning (EEG) nr 2973/79 ersätts med följande:
%quot%Det kött som avses i punkt 1 måste uppfylla hälsoskyddskraven i det importerande tredje landet och komma från djur som slaktats högst två månader före tullklareringen för export.%quot%
Artikel 2
Denna förordning träder i kraft den 4 augusti 1980.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS DIREKTIV av den 25 maj 1983 om ändring av direktiv 82/400/EEG om ändring av direktiv 77/391/EEG och om införande av en kompletterande gemenskapsåtgärd för bekämpning av brucellos, tuberkulos och leukos hos nötkreatur (83/253/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 43 i detta,
med beaktande av kommissionens förslag (),
med beaktande av Europaparlamentets yttrande (),
med beaktande av Ekonomiska och sociala kommitténs yttrande (), och
med beaktande av följande: Genom rådets direktiv 82/400/EEG () infördes särskilt en kompletterande gemenskapsåtgärd för bekämpning av brucellos, tuberkulos och leukos hos nötkreatur.
För att skapa en bättre överblick över hur anslagen används är det nödvändigt att under det kapitel som rör utgifter inom jordbrukssektorn samla alla utgifter för gemenskapens olika åtgärder inom det veterinära området.
För att relevanta finansiella och monetära regler och förfaranden skall kunna tillämpas vid genomförandet av ovannämnda åtgärd, bör respektive artiklar i rådets förordning (EEG) nr 729/70 av den 21 april 1970 om finansiering av den gemensamma jordbrukspolitiken (), senast ändrad genom förordning (EEG) nr 3509/80 (), och rådets förordning (EEG) nr 129/78 av den 24 januari 1978 om de valutakurser som skall användas i den gemensamma jordbrukspolitiken (), tillämpas på motsvarande sätt inom detta område.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Följande artikel skall införas i direktiv 82/400/EEG:
%quot%Artikel 7a
Förordning (EEG) nr 129/78 och artiklarna 8 och 9 i förordning (EEG) nr 729/70 skall tillämpas på motsvarande sätt.%quot%
Artikel 2
Detta direktiv riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 3 juli 1984 om fastställande av utformningen av den särskilda märkning av färskt kött som avses i artikel 5 a i direktiv 64/433/EEG (84/371/EEG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, och
med beaktande av rådets direktiv 64/433/EEG av den 26 juni 1964 om hygienproblem som påverkar handeln med färskt kött inom gemenskapen(), senast ändrat genom direktiv 83/90/EEG(), särskilt artikel 5 a i detta, och
med beaktande av följande: Artikel 5 a i direktiv 64/433/EEG föreskriver att vissa slag av kött får sändas från en medlemsstats territorium till en annan medlemsstats territorium endast om köttet är avsett att genomgå en av de behandlingar som avses i rådets direktiv 77/99/EEG(), och om det har en speciell märkning.
Det är nödvändigt att fastställa ett märke som är lätt att känna igen och som ger de garantier som behövs för att särskilja köttet.
De åtgärder som avses i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM BESLUTAS FÖLJANDE.
Artikel 1
Det märke som avses i artikel 5 a i direktiv 64/433/EEG skall vara utformat på det sätt som framgår av bilagan.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT av den 5 juli 1984 om ändring av beslut 83/471/EEG om Gemenskapens kontrollkommitté för tillämpningen av klassificeringsskalan för slaktkroppar av vuxna nötkreatur (84/375/EEG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1208/81 av den 28 april 1981 om fastställande av en gemenskapsskala för klassificering av slaktkroppar av fullvuxna nötkreatur(), särskilt artikel 5.4 i denna, och
med beaktande av följande: Genom kommissionens beslut 83/471/EEG() fastställs närmare bestämmelser för genomförandet av kontroll på plats av den kontrollkommitté från gemenskapen som avses i artikel 5 i förordning (EEG) nr 1208/81.
Genom förordning (EEG) nr 869/84(), beslöt rådet att under en försöksperiod på tre år skall interventionsåtgärder genomföras på grundval av gemenskapens klassificeringsskala som fastställs i förordning (EEG) nr 1208/81. Räckvidden av de kontroller som genomförs av kontrollkommittén bör utökas så att de också täcker klassificering, identifiering och märkning av produkter som omfattas av interventionsåtgärder. Beslut 83/471/EEG bör därför ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Beslut 83/471 ändras på följande sätt:
1. Artikel 1 skall ersättas med följande:
%quot%Artikel 1
Den kontrollkommitté från gemenskapen som föreskrivs i artikel 5 i förordning (EEG) nr 1208/81, i det följande kallad 'kommittén', skall ansvara för genomförandet av kontroll på plats i fråga om
a) tillämpningen av de bestämmelser som rör gemenskapens klassificeringsskala för slaktkroppar av vuxna nötkreatur,
b) registreringen av marknadspriser i enlighet med klassificeringsskalan,
c) klassificeringen, identifieringen och märkningen av produkter som omfattas av de interventionsåtgärder som föreskrivs i artikel 5 i förordning (EEG) nr 805/68.%quot%2. Artikel 3.1 skall ersättas med följande:
%quot%1. Kontroll på plats skall ske vid slakterier, köttmarknader, interventionsorter, prisnoteringsorter och regionala och centrala organ som ansvarar för genomförandet av de bestämmelser som avses i artikel 1.%quot%
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
RÅDETS BESLUT av den 15 september 1986 om slutande av ett tilläggsprotokoll till avtalet mellan Europeiska ekonomiska gemenskapen och Island till följd av Spaniens och Portugals anslutning till gemenskapen (86/543/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 113 i detta, med beaktande av kommissionens rekommendation, och
med beaktande av följande:
Det är nödvändigt att godkänna tilläggsprotokollet till avtalet mellan Europeiska ekonomiska gemenskapen och Island(1), som undertecknades i Bryssel den 22 juli 1972, för att ta hänsyn till Spaniens och Portugals anslutning till gemenskapen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Tilläggsprotokollet till avtalet mellan Europeiska ekonomiska gemenskapen och Island med anledning a
KOMMISSIONENS FÖRORDNING (EEG) nr 1032/86 av den 9 april 1986 om ändring av förordning (EEG) nr 2388/84 om särskilda tillämpningsföreskrifter för exportbidrag för vissa konserverade nötköttsprodukter
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 805/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för nötkött(), senast ändrad genom förordning (EEG) nr 3768/85(), särskilt artikel 18.5 i denna, och med beaktande av följande:
I kommissionens förordning (EEG) nr 2388/84() fastställs att vissa konserver som uppfyller villkoren i den förordningen och som exporteras till tredje land skall komma i fråga för ett särskilt bidrag om de tillverkas i enlighet med bestämmelserna i artikel 4 i rådets förordning (EEG) nr 565/80(). Med tanke på de avsättningsmöjligheter som finns på marknaderna i tredje land bör dessa villkor anpassas på följande sätt.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för nötkött.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I artikel 2 första stycket andra strecksatsen i förordning (EEG) nr 2388/84 skall %quot%80 %%quot% ersättas med %quot%60 %%quot%.
Artikel 2
Denna förordning träder i kraft den 10 april 1986.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EEG) nr 3940/87 av den 21 december 1987 om ändring av rådets förordningar (EEG) nr 103/76, (EEG) nr 104/76, (EEG) nr 105/76, (EEG) nr 2203/82, (EEG) nr 3117/85 och kommissionens förordningar (EEG) nr 3321/82, (EEG) nr 3510/82, (EEG) nr 3598/83, (EEG) nr 3611/84, (EEG) nr 254/86 och (EEG) nr 314/86
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistikklassifikation och om gemensam tulltaxa(), särskilt artikel 15 i denna, och
med beaktande av följande: Med hänsyn till införandet av den kombinerade varunomenklaturen baserad på det harmoniserade systemet har den tullnomenklatur som ingår i rådets förordning (EEG) nr 3796/81() ändrats i överensstämmelse med den nämnda nomenklaturen med verkan från den 1 januari 1988 genom rådets förordning (EEG) nr 3759/87().
Därför är det nödvändigt att ändra vissa förordningar om tillämpning av förordning (EEG) nr 3796/81.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De förordningar som anges i rubriken skall ändras i enlighet med bilagan.
Artikel 2
Denna förordning träder i kraft den 1 januari 1988.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS DIREKTIV av den 3 december 1987 om ändring i direktiv 70/220/EEG om tillnärmning av medlemsstaternas lagstiftning om åtgärder mot luftföroreningar genom avgaser från motorfordon (88/76/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av kommissionens förslag(1),
i samarbete med Europaparlamentet(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
med beaktande av följande: Det är viktigt att vidta åtgärder i syfte att successivt upprätta den inre marknaden under tiden fram till den 31 december 1992. Den inre marknaden skall utgöra ett område utan inre gränser inom vilket ett fritt utbyte av varor, personer, tjänster och kapital är säkerställt.
Enligt de Europeiska gemenskapernas första aktionsprogram om skyddet för miljön, som antogs av rådet den 22 november 1973, skall de senaste vetenskapliga framstegen beaktas när det gäller att bekämpa luftförorening i form av avgaser som släpps ut från motordrivna fordon och tidigare antagna direktiv ändras i enlighet med detta. Enligt det tredje aktionsprogrammet bör ytterligare ansträngningar göras för att avsevärt minska utsläppen av luftföroreningar från motordrivna fordon.
I direktiv 70/220/EEG(4) fastslås gränsvärden för utsläpp av kolmonoxid och oförbrända kolväten från sådana motorer. Dessa gränsvärden sänktes först genom direktiv 74/290/EEG(5) och kompletterades, genom direktiv 77/102/EEG(6), med gränsvärden för utsläpp av kväveoxider. Gränsvärdena för dessa tre föroreningar sänktes ytterligare genom direktiven 78/665/EEG(7) och 83/351/EEG(8).
Kommissionens arbete, som utförts i en strävan att til lämpa en övergripande syn vid utvecklingen av regler för motorfordonsindustrin, har visat att den europeiska industrin redan har tillgång till eller håller på att förfina en motorteknologi som kommer att göra det möjligt att ytterligare sänka gränsvärdena. Under den tidrymd som är aktuell kommer en sådan sänkning inte att äventyra gemenskapens målsättningar inom andra områden, särskilt vad gäller ett effektivt energiutnyttjande. Det är nödvändigt att främja nytänkande och industriell konkurrens på såväl den inre marknaden som på utländska marknader. Det är nödvändigt att gemenskapen vidtar åtgärder mot fordonsutsläpp, vilka innebär en hög ambitionsnivå för miljöskyddet och samtidigt är anpassade till europeiska förhållanden, så att den slutliga effekten på miljön motsvarar den som uppnås med de normer som gäller för utsläpp från fordon i Amerikas Förenta Stater. För att nå detta mål är det lämpligt att tillämpa varierande lösningar för olika motorstorlekar, för att så långt möjligt uppnå att gemenskapens krav kan tillgodoses till rimliga kostnader och med olika tekniska lösningar. De gränsvärden som fastslagits för fordon med en slagvolym mindre än 1,4 liter återspeglar nuvarande tekniska och ekonomiska förhållanden hos de europeiska tillverkarna inom denna sektor av marknaden. De gränsvärden som skall gälla år 1992/93 bör fastställas år 1987.
Gränsvärdena i detta direktiv grundar sig på den provmetod som fastslagits i direktiv 70/220/EEG. Förfarandet måste dock anpassas så att det är representativt inte bara för tätortsområden med hög trafikbelastning utan också utanför sådana områden. Ett beslut om en sådan anpassning bör fattas senast år 1987.
Enligt artikel 5 i direktiv 70/220/EEG är det möjligt att anpassa bestämmelserna i bilagorna med hänsyn till tekniska framsteg.
Bensinmotorer i sådana fordon som omfattas av detta direktiv bör vara konstruerade för att drivas med blyfri bensin, så att användningen av blybaserade tillsatser i bränslen kan upphöra, vilket i hög grad skulle bidra till att minska föroreningen av miljön med detta ämne.
Det är nödvändigt att säkerställa att bestämmelserna om motorer med kompressionständning (dieselmotorer) i fordon som omfattas av detta direktiv fortsättningsvis, med hänsyn till de speciella egenskaperna hos de föroreningar som avges från sådana motorer, överensstämmer med kommande ändringar i de bestämmelser som rör andra föroreningar från sådana motorer, vilka behandlas i direktiv 72/306/EEG(9).
Under tiden från det att de europeiska normerna antas till det att den modifierade europeiska körcykeln införs, är det önskvärt att fordon som erhåller typgodkännande enligt motsvarande normer på gemenskapens exportmarknader också skall anses uppfylla kraven för EEG-typgodkännande.
De medlemsstater som så önskar får, med beaktande av fördragets bestämmelser, i förtid tillämpa de nya värden som fastställs genom detta direktiv. De får dock inte hindra att fordon, av inhemsk tillverkning eller importerade, används eller sprids på marknaden om de uppfyller gemenskapens krav.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga 1-3, 6 och 7 till direktiv 70/220/EEG ändras enligt bilagan till detta direktiv. En ny bilaga 3 A införs.
Artikel 2
1. Från och med den 1 juli 1988 får ingen medlemsstat av skäl som hänför sig till luftförorening genom gaser från en motor eller kvalitetskrav på motorbränsle: - vägra att bevilja EEG-typgodkännande eller att utfärda det dokument som avses i andra strecksatsen i artikel 10.1 i direktiv 70/156/EEG(10), senast ändrat genom direktiv 87/403/EEG(11), eller att bevilja nationellt typgodkännande för en motorfordonstyp, eller
- förbjuda att sådana fordon tas i bruk,
om utsläppen av gasformiga föroreningar från fordonstypen eller från fordonen liksom kraven på motorbränslets kvalitet är sådana att bestämmelserna i direktiv 70/220/EEG i dess lydelse enligt detta direktiv är uppfyllda.
2. Medlemsstaterna får: från och med den 1 oktober 1988 i fråga om fordonstyper med motorer med större slagvolym än 2 000 cm³,
från och med den 1 oktober 1990 i fråga om fordonstyper med motorer med mindre slagvolym än 1 400 cm³,
från och med den 1 oktober 1991 i fråga om fordonstyper med motorer med en slagvolym som uppgår till 1 400 cm³ men inte överstiger 2 000 cm³, samt från och med den 1 oktober 1994 i fråga om fordonstyper med direktinsprutade dieselmotorer med samma slagvolym,
- inte längre utfärda det dokument som avses i sista strecksatsen i artikel 10.1 i direktiv 70/156/EEG för en motorfordonstyp, och
- vägra att bevilja nationellt typgodkännande för en motorfordonstyp,
som släpper ut gasformiga föroreningar i sådana mängder att kraven i bilagorna till direktiv 70/220/EEG, i deras lydelse enligt detta direktiv, inte är uppfyllda.
3. Från och med den 1 oktober 1989 i fråga om fordonstyper med motorer med större slagvolym än 2 000 cm³,
från och med den 1 oktober 1991 i fråga om fordonstyper med motorer med mindre slagvolym än 1 400 cm³,
från och med den 1 oktober 1993 i fråga om fordonstyper med motorer med en slagvolym som uppgår till 1 400 cm³ men inte överstiger 2 000 cm³, samt från och med den 1 oktober 1996 i fråga om fordonstyper med direktinsprutade dieselmotorer med samma slagvolym,
får medlemsstaterna förbjuda att fordon tas i bruk, om utsläppen av gasformiga föreningar från fordonen eller kraven på motorbränslets kvalitet är sådana att bestämmelserna i bilagorna till direktiv 70/220/EEG, i deras lydelse enligt detta direktiv, inte är uppfyllda.
Artikel 3
1. Medlemsstaterna får vägra att utfärda nationellt typgodkännande, EEG-typgodkännande eller det dokument som avses i andra strecksatsen i artikel 10.1 i direktiv 70/156/EEG för en fordonstyp med förbränningsmotor med styrd tändning som behöver ett bränsle som inte överensstämmer med bestämmelserna i bilagorna till direktiv 70/220/EEG i deras lydelse enligt detta direktiv: - från och med den 1 oktober 1988 i fråga om fordonstyper med en motor med större slagvolym än 2 000 cm³, med de undantag som anges i avsnitt 8.1,
- från och med den 1 oktober 1989 i fråga om andra fordonstyper.
2. Från och med den 1 oktober 1990 får medlemsstaterna förbjuda att fordon tas i bruk som är utrustade med förbränningsmotorer med styrd tändning som behöver ett bränsle som inte överensstämmer med bestämmelserna i bilagorna till direktiv 70/220/EEG i deras lydelse enligt detta direktiv, om inte tillverkaren lämnar ett skriftligt intyg som godtas av det tekniska organ som beviljade det första typgodkännandet avseende utsläpp. Av intyget skall framgå att en anpassning av fordonen till de nya kraven på bränsle innebär omfattande konstruktions ändringar i form av andra material i inloppseller avgasventilsätena eller en minskning av kompressionsförhållandet, eller en ökning av motorns storlek för att kompensera för effektförluster. I detta fall kan ett sådant förbud endast tillämpas från de tidpunkter som anges i artikel 2.3.
Artikel 4
Senast den 31 december 1987 skall rådet på förslag från kommissionen: - besluta om en ytterligare sänkning av de gränsvärden som gäller för fordon med en motorstorlek mindre än 1 400 cm³, att tillämpas senast år 1992 i fråga om utfärdande av nya nationella typgodkännanden och år 1993 i fråga om att ta fordon i bruk,
- ändra den provmetod som anges i bilaga 3 till direktiv 70/220/EEG för att anpassa metoden till aktuella förhållanden, främst genom att lägga till körcykler för landsvägskörning,
- besluta om ordningen för ikraftträdandet av den ändrade provmetoden i bilaga 3 och om de villkor som skall gälla vid upphävandet av de nuvarande bilagorna 3 och 3 A till direktiv 70/220/EEG i deras lydelse enligt detta direktiv, inbegripet övergångsperioden.
Artikel 5
Medlemsstaterna skall sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv senast den 1 juli 1988 och genast underrätta kommissionen om detta.
Artikel 6
Detta direktiv riktar sig till medlemsstaterna.
KOMMISSIONENS DIREKTIV av den 22 juni 1988 om anpassning till den tekniska utvecklingen av rådets direktiv 79/622/EEG om tillnärmning av medlemsstaternas lagstiftning om skyddsbågar på jordbruks- eller skogsbrukstraktorer med hjul (statisk provning) (88/413/EEG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets direktiv 74/150/EEG av den 4 mars 1974 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av jordbruks- eller skogsbrukstraktorer med hjul(1), senast ändrat genom direktiv 88/279/EEG(2), särskilt artikel 11 i detta,
och med beaktande av följande: Med hänsyn till de erfarenheter som har vunnits är det nu möjligt att precisera och komplettera vissa bestämmelser i rådets direktiv 79/622/EEG(3), senast ändrat genom direktiv 87/354/EEG(4).
De åtgärder som har införts genom detta direktiv har tillstyrkts av kommittén för anpassning till den tekniska utvecklingen av direktiven om att avskaffa tekniska handelshinder inom sektorn för jordbruks- och skogsbrukstraktorer.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagorna 3 och 4 till direktiv 79/622/EEG skall ändras enligt bilagan till detta direktiv.
Artikel 2
1. Från den 1 oktober 1988 får ingen medlemsstat
- vägra, vad avser en typ av traktor, att bevilja EEG-typgodkännande, att utfärda det dokument som nämns i artikel 10.1, den sista strecksatsen i direktiv 74/150/EEG, eller att bevilja nationellt typgodkännande, eller
- förbjuda att traktorer tas ibruk,
om överrullningsskyddet för denna typ av traktor eller traktorer överensstämmer med bestämmelserna i detta direktiv.
2. Från den 1 oktober 1989 kan medlemsstaterna
- inte längre utfärda det dokument som nämns i artikel 10.1, sista strecksatsen i direktiv 74/150/EEG, med avseende på en typ av traktor vars överrullningsskydd inte överensstämmer med bestämmelserna i detta direktiv,
- vägra att bevilja nationellt typgodkännande med avseende på en traktortyp, vars överrullningsskydd inte överensstämmer med bestämmelserna i detta direktiv.
Artikel 3
Medlemsstaterna skall sätta i kraft de bestämmelser som är nödvändiga för att följa detta direktiv senast den 30 september 1988. De skall genast underrätta kommissionen om detta.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS DIREKTIV av den 18 juni 1991 om ändring för tionde gången av direktiv 76/769/EEG om tillnärmning av medlemsstaternas lagar och andra författningar om begränsning av användning och utsläppande på marknaden av vissa farliga ämnen och preparat (beredningar) (91/338/EEG)
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 100a i detta,
med beaktande av kommissionens förslag(1),
i samarbete med Europaparlamentet(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
med beaktande av följande: Åtgärder bör vidtas för att successivt upprätta den inre marknaden under tiden fram till den 31 december 1992. Den inre marknaden skall vara ett område utan inre gränser inom vilket ett fritt utbyte av varor, personer, tjänster och kapital är säkerställt.
I rådets resolution av den 25 januari 1988(4) uppmanas kommissionen att utan dröjsmål utreda vilka särskilda åtgärder som bör ingå i ett gemenskapsprogram för att bekämpa miljöförorening genom kadmium. Människors hälsa måste också skyddas. En övergripande strategi bör tillämpas, som särskilt syftar till att begränsa användningen av kadmium och stimulera forskningen om ersättningsämnen.
Kunskapen om och metoderna för framställning av ersättningsämnen förbättras. Det är därför lämpligt att systematiskt se över situationen mot bakgrund av de vetenskapliga och tekniska studier som skall utföras enligt den nyss nämnda resolutionen.
Polyvinylklorid (PVC) får inte färgas med kadmiumbaserade pigment. För vissa tillämpningar har dock tekniken ännu inte utvecklats så långt att det är möjligt att använda en icke-kadmiumbaserad stabilisator.
Vissa medlemsstater har redan infört begränsningar i fråga om användning eller saluförande av de ovan nämnda ämnena eller beredningar i vilka de ingår. Sådana begränsningar inverkar direkt på den inre marknadens upprättande och funktion. En tillnärmning av medlemsstaternas lagstiftning på detta område är således nödvändig. Bilaga 1 till direktiv 76/769/EEG(5) senast ändrat genom direktiv 89/678/EEG(6) bör därför ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga 1 till direktiv 76/769/EEG ändras på det sätt som anges i bilagan till det här direktivet. De nya bestämmelserna skall dock inte gälla för kadmiumhaltiga produkter som redan omfattas av annan gemenskapslagstiftning.
Artikel 2
Kommissionen skall mot bakgrund av utvecklingen i fråga om kunskaper och metoder som avser mindre farliga ersättningsämnen för kadmium och dess föreningar och i samråd med medlemsstaterna utvärdera situationen, första gången senast tre år efter den dag som anges i artikel 3.1 och därefter med jämna mellanrum. Förfarandet enligt artikel 2a i direktiv 76/769/EEG skall tillämpas.
Artikel 3
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 31 december 1992. De skall genast underrätta kommissionen om detta.
2. När en medlemsstat antar bestämmelser till följd av punkt 1 skall dessa innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
KOMMISSIONENS FÖRORDNING (EEG) nr 1180/91 av den 6 maj 1991 om ändring av förordning (EEG) nr 1014/90 om närmare tillämpningsföreskrifter för definition, beskrivning och presentation av spritdrycker
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1576/89 av den 29 maj 1989 om allmänna bestämmelser för definition, beskrivning och presentation av spritdrycker(1), särskilt artikel 6.3 i denna, och
med beaktande av följande: Tillämpningsföreskrifter om definition, beskrivning och presentation av spritdrycker finns i kommissionens förordning EEG nr 1014/90 av den 24 april 1990(2). För att vissa termer, som kompletterar försäljningsbeteckningen för ett antal spritdrycker som tillverkas enligt traditionella metoder, skall skyddas mot illojal konkurrens, bör termerna förbehållas de spritdrycker som definieras i bilagan till denna förordning.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för genomförande av regler om spritdrycker. HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1 Följande artikel 7a skall införas i förordning (EEG) nr 1014/90:
%quot%Artikel 7a De tillägg till försäljningsbeteckningen som anges i bilagan till denna förordning skall reserveras för de produkter som definieras där.
Spritdrycker som inte uppfyller kraven för produkterna i bilagan, får inte bära de beteckningar som anges där.%quot% Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS FÖRORDNING (EEG) nr 2155/91 av den 20 juni 1991 om särskilda tillämpningsföreskrifter för artiklarna 37, 39 och 40 i avtalet mellan Europeiska ekonomiska gemenskapen och Schweiz om annan direkt försäkring än livförsäkring
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 57.2 sista meningen och artikel 235 i detta,
med beaktande av kommissionens förslag (1),
i samarbete med Europaparlamentet (2),
med beaktande av Ekonomiska och sociala kommitténs yttrande (3), och
med beaktande av följande: Ett avtal mellan Europeiska ekonomiska gemenskapen och Schweiz om annan direkt försäkring än livförsäkring undertecknades i Luxemburg den 10 oktober 1989.
Enligt avtalet skall en gemensam kommitté inrättas som skall administrera avtalet, säkerställa att det genomförs på ett riktigt sätt samt fatta beslut i de fall som avtalet föreskriver. Gemenskapens företrädare i den gemensamma kommittén måste utses och särskilda bestämmelser måste antas för fastställandet av gemenskapens ståndpunkter i kommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I den gemensamma kommitté som anges i artikel 37 i avtalet skall gemenskapen företrädas av kommissionen som skall biträdas av företrädare för medlemsstaterna.
Artikel 2
Gemenskapens ståndpunkt i den gemensamma kommittén skall beslutas av rådet med kvalificerad majoritet på förslag från kommissionen.
Rådet skall med kvalificerad majoritet på förslag från kommissionen besluta om antagande av de beslut som den gemensamma kommittén fattar i enlighet med artiklarna 37, 39 och 40 i avtalet.
Artikel 3
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS FÖRORDNING (EEG) nr 3578/92 av den 7 december 1992 om ändring av förordning (EEG) nr 1107/70 om stöd till transporter på järnväg, väg och inre vattenvägar
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, särskilt artikel 75 i detta,
med beaktande av kommissionens förslag (),
med beaktande av Europaparlamentets yttrande (),
med beaktande av Ekonomiska och sociala kommitténs yttrande (), och
med beaktande av följande: I förordning (EEG) nr 1107/70 () fastställs att medlemsstaterna får främja utvecklingen av kombinerad transport genom att bevilja stöd till investeringar i infrastruktur och i stationära och rörliga anläggningar som krävs för omlastning, eller till driftskostnader för kombinerad transittrafik inom gemenskapen som passerar genom tredje lands territorium.
Utvecklingen av den kombinerade transporten visar att för gemenskapen som helhet är igångsättningsfasen för denna teknik ännu inte över, och stödordningen måste följaktligen upprätthållas under ytterligare en tid.
Möjligheterna att bevilja stöd för driftskostnader för kombinerad transittrafik som passerar genom tredje land är endast berättigad beträffande Österrike, Schweiz och staterna i det forna Jugoslavien.
Behovet av att snabbt uppnå ekonomisk och social samhörighet inom gemenskapen innebär att tonvikten måste ligga på investeringar i järnvägs- och väganläggningar som är särskilt utformade med hänsyn till kombinerade transporter, i synnerhet om dessa utgör ett alternativ till sådana förbättringar i infrastrukturen som inte kan genomföras på kort sikt.
Beviljande av stöd till väganläggningar för kombinerade transporter kan dessutom vara ett effektivt sätt att få små och medelstora företag att använda kombinerade transporter.
Stöd till utrustning som är särskilt utformat med hänsyn till kombinerade transporter kan främja utvecklingen av ny bimodalteknik och ny omlastningsteknik.
Under en begränsad igångsättningsfas bör möjligheten att bevilja stöd utsträckas till investeringar i transportanläggningar som särskilt är utformade med hänsyn till kombinerade transporter förutsatt att stödet endast går till detta ändamål.
Den nuvarande stödordningen bör upprätthållas till och med den 31 december 1995, och rådet bör i enlighet med villkoren i fördraget besluta vilken ordning som skall tillämpas därefter eller, om nödvändigt, villkoren för avveckling av stödet.
Förordning (EEG) nr 1107/70 bör därför ändras i enlighet med detta.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 3.1 e i förordning (EEG) nr 1107/70 skall ersättas med följande:
%quot%e) när stöd beviljas som en tillfällig åtgärd och i avsikt att underlätta utvecklingen av kombinerade transporter, gäller till och med den 31 december 1995 att sådant stöd skall avse
- investeringar i infrastruktur, eller
- stationära och rörliga anläggningar som krävs för omlastning, eller
- investeringar i transportutrustning som är särskilt utformad med hänsyn till kombinerad transport och används enbart för kombinerad transport, eller
- driftskostnader för kombinerade transporter som passerar genom Österrike, Schweiz eller genom staterna i forna Jugoslavien.
Vartannat år skall kommissionen till rådet överlämna en lägesrapport om tillämpningen av ovannämnda åtgärder och särskilt uppgifter om bl.a. hur stödet används, storleken på stödet och dess betydelse för kombinerade transporter. Medlemsstaterna skall förse kommissionen med de uppgifter som behövs för sammanställning av lägesrapporten.
Senast den 31 december 1995 skall rådet på kommissionens förslag och i enlighet med villkoren i fördraget besluta vilken stödordning som skall tillämpas därefter eller, om nödvändigt, villkoren för avveckling av stödet.%quot%
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Den skall tillämpas från och med den 1 januari 1993. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS BESLUT av den 21 december 1992 om inrättande av en vetenskaplig kommitté för ursprungsbeteckningar, geografiska beteckningar och särartsskydd (93/53/EEG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen, och
med beaktande av följande: För gemenskapens skydd av ursprungsbeteckningar och geografiska beteckningar kan det krävas en granskning dels av en benämnings generiska natur och de faktorer som skall beaktas när ursprungsbeteckning och geografisk beteckning för jordbruksprodukter och livsmedel skall definieras, dels av tillämpningen av kriterierna för sund konkurrens i affärstransaktioner och av faran av att konsumenterna vilseleds i den mening som avses i artiklarna 13 och 14 i rådets förordning (EEG) nr 2081/92(1) i de fall då det råder motsättning mellan ursprungsbeteckning eller geografisk beteckning och varumärke, homonymer eller befintliga produkter som saluförs enligt gällande lagstiftning.
För gemenskapens särartsskydd kan det vid registreringen uppstå behov av en granskning av frågor som gäller bedömningen av jordbruksprodukters och livsmedels traditionella natur.
För att sådana frågor skall kunna avgöras krävs biträde av experter med hög kompetens inom juridik eller jordbruk och i synnerhet inom immaterialrätt.
Det är därför lämpligt att inrätta en vetenskaplig kommitté som skall biträda kommissionen i dess arbete.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
En vetenskaplig kommitté, nedan kallad kommittén, inrättas härmed för att biträda kommissionen i dess arbete.
Artikel 2
Kommitténs uppgift skall vara att, på kommissionens uppdrag, granska alla tekniska frågor som sammanhänger med tillämpningen av förordning (EEG) nr 2081/92 och rådets förordning (EEG) nr 2082/92(2), då det gäller registrering av benämningar på jordbruksprodukter och livsmedel samt motsättningar mellan medlemsstaterna, särskilt i följande frågor:
1. Vilka faktorer som skall beaktas vid definitionen av geografisk beteckning och ursprungsbeteckning samt undantag till sådana, särskilt i fråga om extraordinärt rykte och anseende.
2. Generisk natur.
3. Bedömning av traditionell natur.
4. Bedömning av kriterier för sund konkurrens i affärstransaktioner och av risken att konsumenterna vilseleds i de fall då det råder motsättning mellan ursprungsbeteckning eller geografisk beteckning och varumärke, homonymer eller befintliga produkter som saluförs enligt gällande lagstiftning.
Artikel 3
1. Medlemmarna i kommittén skall utses av kommissionen bland experter med hög kompetens inom de områden som avses i artikel 2.
2. Kommittén skall bestå av sju ordinarie medlemmar och sju suppleanter med rätt att delta i sammanträdena.
Artikel 4
1. Kommittén skall bland sina medlemmar utse en ordförande och en vice ordförande.
Dessa skall väljas med enkel majoritet.
2. Kommissionen skall tillhandahålla sekretariattjänster till kommittén.
Artikel 5
Kommittén är beslutför endast då samtliga medlemmar är närvarande. Kommittén skall tillstyrka förslag, när antalet röster för förslaget överstiger antalet röster mot. Vid lika röstetal skall nedläggning av röst räknas som röst för förslaget.
Artikel 6
1. Medlemmarna skall utses för en period på fem år, och deras mandat får förnyas. Ordföranden och vice ordföranden skall dock utses på två år. De får inte återväljas omedelbart efter två efterföljande mandatperioder på vardera två år. Medlemmarna skall inte ersättas för sina tjänster.
2. Efter utgången av femårs- eller tvåårsperioderna skall medlemmarna, ordföranden och vice ordföranden sitta kvar tills de ersätts eller deras mandat förnyas.
3. Om en medlem, ordföranden eller vice ordföranden är förhindrad att fullgöra sina uppgifter eller avgår, skall en ersättare utses för återstoden av mandattiden enligt det förfarande som föreskrivs i artikel 3 eller artikel 4.
Artikel 7
1. Kommittén skall sammanträda på begäran av en företrädare för kommissionen.
2. Kommissionens företrädare samt berörda tjänstemän och andra anställda vid kommissionen skall närvara vid kommitténs sammanträden.
3. Kommissionens företrädare får inbjuda framstående experter med särskilt hög kompetens i de frågor som behandlas att delta i sammanträdena.
Artikel 8
1. Kommittén skall behandla ärenden där kommissionen har begärt ett yttrande.
Kommissionen får bestämma en tidsfrist för yttrandet.
2. När det råder enighet i kommittén om det yttrande som skall avges skall kommittén utarbeta ett gemensamt yttrande. Om enighet inte uppnås, skall de olika synpunkter som uttryckts under arbetet tas med i en rapport som skall utarbetas under ansvar av kommitténs sekretariat.
Artikel 9
Kommitténs medlemmar är skyldiga att inte avslöja uppgifter som kommit till deras kännedom genom arbete i kommittén, om kommissionens företrädare underrättar dem om att det yttrande som begärts gäller ett ärende av konfidentiell natur.
KOMMISSIONENS FÖRORDNING (EEG) nr 1718/93 av den 30 juni 1993 om den avgörande faktorn för jordbruksomräkningskurserna för utsäde
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska ekonomiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 3813/92 av den 28 december 1992 om den beräkningsenhet och de omräkningskurser som skall tillämpas avseende den gemensamma jordbrukspolitiken(1), särskilt artikel 6.2 i denna, och
med beaktande av följande: I enlighet med artikel 3 i rådets förordning (EEG) nr 2358/71 av den 26 oktober 1971 om den gemensamma organisationen av marknaden för utsäde(2), senast ändrad genom förordning (EEG) nr 3695/92(3), kan stöd beviljas för de produkter som anges i bilagan till den förordningen.
I kommissionens förordning (EEG) nr 1546/75 av den 18 juni 1975 om fastställande av den faktor som ligger till grund för rätten till stöd för utsäde(4), senast ändrad genom förordning (EEG) nr 2811/86(5), anges den avgörande faktorn för jordbruksomräkningskursen på grundval av rättsliga kriterier och bestämmelser som har ändrats väsentligt i samband med den nya agromonetära ordning som infördes genom förordning (EEG) nr 3813/92. Enligt de nya bestämmelserna infaller den tidpunkt då verksamhetens mål uppnås under skördetiden och kan därför anses vara den 1 augusti varje regleringsår. Denna dag anses därför som den avgörande faktorn för jordbruksomräkningskursen i fråga om stöd till producenter av utsäde.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för utsäde.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Den kurs som skall tillämpas i samband med det stöd som fastställs i artikel 3 i förordning (EEG) nr 2358/71 skall vara den jordbruksomräkningskurs som gäller den 1 augusti det regleringsår för vilket stödet gäller.
Artikel 2
Förordning (EEG) nr 1546/75 skall upphöra att gälla.
Artikel 3
Denna förordning träder i kraft den 1 juli 1993.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS BESLUT av den 19 april 1994 om en av rådet enligt artikel J 3 i Fördraget om den Europeiska unionen beslutad gemensam åtgärd till stöd för fredsprocessen i Mellanöstern (94/276/GUSP)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om Europeiska unionen, särskilt artiklarna J 3 och J 11 i detta,
med beaktande av de allmänna riktlinjer som utfärdades av Europeiska rådet den 29 oktober 1993,
med beaktande av ramen för den gemensamma åtgärd som Europeiska rådet enades om den 10 och 11 december 1993, och
med beaktande av artikel C i Fördraget om Europeiska unionen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
a) I syfte att verka för att en heltäckande fred i Mellanöstern sluts på grundval av FN:s säkerhetsråds resolutioner skall Europeiska unionen
- delta i de internationella arrangemang som parterna kommer överens om för att säkerställa fred inom ramen för den process som startades i Madrid,
- använda sitt inflytande för att uppmuntra alla parter att ovillkorligt stödja fredsprocessen på grundval av inbjudningar till Madrid-konferensen och arbeta för att stärka demokratin och respekten för de mänskliga rättigheterna,
- bidra till utformningen av de framtida förbindelserna mellan regionens parter i arbetsgruppen för vapenkontroll och regional säkerhet.
b) Europeiska unionen skall
- utveckla sin roll i den särskilda sambandskommitté som ansvarar för samordningen av internationellt stöd till de ockuperade områdena,
- bevara sin ledande roll i arbetsgruppen för regional ekonomisk utveckling (REDWG) och utveckla sitt deltagande i andra multinationella grupper,
- överväga andra sätt att bidra till regionens utveckling.
c) Europeiska unionen skall
- fortsätta att driva frågan om de förtroendeskapande åtgärder som den har förelagt parterna,
- fortsätta att rikta demarscher till de arabiska staterna i syfte att få till stånd ett slut på bojkotten mot Israel,
- följa utvecklingen vad avser israeliska bosättningar inom samtliga ockuperade områden och fortsätta att rikta demarscher till Israel i denna fråga.
Artikel 2
Rådet skall i enlighet med relevanta gemenskapsförfaranden behandla de förslag som kommissionen lägger fram om
- ett snabbt genomförande av biståndsprogrammen för utveckling av de ockuperade områdena och en palestinsk driftsbudget, i nära samråd med palestinierna och en lika nära samverkan med andra biståndsgivare,
- lämnande av stöd enligt befintliga riktlinjer till de andra parterna i de bilateral förhandlingarna, allteftersom dessa gör betydande framsteg mot fred.
Artikel 3
För att aktivt och snabbt bidra till att en palestinsk polisstyrka upprättas skall
a) Europeiska unionen lämna bistånd,
b) presidiet i nära samverkan med kommissionen underlätta samordningen genom utbyte av information mellan medlemsstaterna om deras bilaterala bistånd,
c) ett belopp på högst 10 miljoner ecu från gemenskapens budget som en brådskande åtgärd ställas till förfogande som bistånd till upprättandet av en palestinsk polisstyrka.
Artikel 4
Europeiska unionen skall på begäran av parterna medverka till att det palestinska folket skyddas genom tillfällig internationell närvaro på de ockuperade områdena i överensstämmelse med säkerhetsrådets resolution 904 (1994).
De praktiska arrangemangen och den finansiering som följer av denna artikel skall behandlas i ett särskilt, separat beslut.
Artikel 5
På begäran av parterna skall Europeiska unionen genomföra ett samordnat program för bistånd till förberedelse och övervakning av de val på de ockuperade områdena som påbjöds i principdeklarationen av den 13 september 1993. De exakta praktiska arrangemangen och finansieringen skall fastställas i ett särskilt rådsbeslut när Israel och PLO har enats om hur valet skall arrangeras. Europaparlamentet kommer att inbjudas att delta i dessa arrangemang.
Artikel 6
Europeiska unionen bekräftar att den är villig att fatta ytterligare praktiska beslut inom ramen för denna gemensamma åtgärd allteftersom fredsprocessen utvecklas.
Artikel 7
Detta beslut skall ha verkan från och med denna dag.
Artikel 8
Detta beslut skall offentliggöras i Europeiska gemenskapernas officiella tidning.
RÅDETS BESLUT av den 17 juni 1994 om bemyndigande för Europeiska gemenskapen och Europeiska atomenergigemenskapen att underteckna och sluta konventionen med stadga för Europaskolorna (94/557/EG, Euratom)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 235 i detta,
med beaktande av Fördraget om upprättandet av Europeiska kol- och stålgemenskapen, särskilt artikel 203 i detta,
med beaktande av kommissionens förslag (),
med beaktande av Europaparlamentets yttrande (), och
med beaktande av följande:
För europeiska gemenskaperna är det angeläget att tillhandahålla gemensam utbildning för sin personals barn i Europaskolor för att säkerställa att gemenskapens institutioner fungerar tillfredsställande och för att underlätta för personalen att fullgöra sina uppgifter. I detta syfte undertecknade de ursprungliga medlemsstaterna den 12 april 1957 konventionen angående stadgan för Europaskolorna.
Den 31 maj 1990 efterlyste rådet och utbildningsministrarna, församlade i rådet, en ny konvention om Europaskolorna som skulle utarbetas för att effektivisera skolornas verksamhet och i högre grad erkänna gemenskapens roll i skolorna.
Gemenskapernas deltagande i genomförandet av konventionen är nödvändig för att säkerställa att Europeiska gemenskapens och Europeiska atomenergigemenskapens mål uppnås.
Europeiska gemenskapen och Europeiska atomenergigemenskapen kommer att delta i genomförandet av konventionen genom att utöva de befogenheter som följer av de bestämmelser som fastställs genom konventionen och av sådana framtida rättsakter som de kan anta i enlighet med konventionens villkor.
Det är följaktligen nödvändigt för Europeiska gemenskaperna att sluta denna konvention. De enda befogenheter som finns för antagandet av detta beslut är de som fastställs i artikel 235 i Fördraget om upprättandet a
KOMMISSIONENS FÖRORDNING (EG) nr 180/94 av den 28 januari 1994 om ändring av förordning (EEG) nr 1756/93 om avgörande händelser för den jordbruksomräkningskurs som tillämpas för mjölk och mjölkprodukter
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 3813/92 av den 28 december 1992 om beräkningsenheten och de omräkningskurser som skall tillämpas inom den gemensamma jordbrukspolitiken(1), särskilt artikel 6.2 i denna, och
med beaktande av följande: Syftet med kommissionens förordning (EEG) nr 1756/93(2), senast ändrad genom förordning (EG) nr 114/94(3), är att fastställa den exakta jordbruksomräkningskurs som skall tilllämpas på belopp som fastställs i ecu inom sektorn för mjölk och mjölkprodukter. Den nämnda förordningen måste därför kompletteras genom fastställande av avgörande händelser för de belopp som avses i artikel 1.3 i kommissionens förordning (EG) nr 3582/93 av den 21 december 1993 om tillämpningsföreskrifter för rådets förordning (EEG) nr 2073/92 om främjande av konsumtionen inom gemenskapen och breddande av marknaderna för mjölk och mjölkprodukter(4).
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från förvaltningskommittén för mjölk och mjölkprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Följande punkt 14 skall läggas till i del D i bilagan till förordning (EEG) nr 1756/93:
%quot%%gt%Plats för tabell%gt% %quot%
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning. Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EG) nr 1026/94 av den 2 maj 1994 om ändring av förordning (EEG) nr 1538/91 om tillämpningsföreskrifter för rådets förordning (EEG) nr 1906/90 om vissa handelsnormer för fjäderfäkött
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1906/90 av den 26 juni 1990 om vissa handelsnormer för fjäderfäkött(1), senast ändrad genom förordning (EG) nr 3204/93(2), särskilt artikel 9 i denna, och
med beaktande av följande: I kommissionens förordning (EEG) nr 1538/91(3), senast ändrad genom förordning (EEG) nr 2891/93(4), anges det referens-laboratorium i gemenskapen som ansvarar för kontrollen av vattenhalten i fryst och djupfryst kyckling och dess befogenheter och uppgifter. Det bör fastställas vilket finansiellt stöd gemenskapen skall ge till referenslaboratoriet så att det kan utföra sina uppgifter.
Gemenskapens finansiella stöd bör inledningsvis fastställas för en period på tre år. Stödet kommer att ses över med syftet att förlängning skall beviljas före utgången av den inledande perioden.
Ett kontrakt bör ingås mellan Europeiska gemenskapen och gemenskapens referenslaboratorium som fastställer villkoren för utbetalning av finansiellt stöd.
Förvaltningskommittén för fjäderfäkött och ägg har inte avgivit något yttrande inom den tid som dess ordförande bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I artikel 14a i förordning (EEG) nr 1538/91 skall följande punkt 14 läggas till:
%quot%14. Gemenskapen skall bevilja gemenskapens referenslaboratorium %quot%Het Spelderholt%quot%, Centre for Poultry Research and Information Services, Beekbergen, Nederländerna, ett finansiellt stöd på högst 75 000 ecu för en period på tre år för fullgörandet av de uppgifter som avses i bilaga 9 punkt 1.
Det finansiella stödet skall betalas till referens-laboratoriet i enlighet med villkoren i ett kontrakt som sluts mellan kommissionen på uppdrag a
KOMMISSIONENS FÖRORDNING (EG) nr 2714/94 av den 8 november 1994 om ändring av förordning (EEG) nr 2054/89 om tillämpningsföreskrifter för systemet med minimipriser vid import av torkade druvor
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av av rådets förordning (EEG) nr 426/86 av den 24 februari 1986 om den gemensamma organisationen av marknaden för bearbetade produkter av frukt och grönsaker(1), senast ändrad genom kommissionens förordning (EG) nr 1490/94(2), särskilt artikel 9.6 i denna, och
med beaktande av följande: I artikel 2.3 i kommissionens förordning (EEG) nr 2054/89(3), senast ändrad genom förordning (EEG) nr 3821/92(4), föreskrivs de villkor på vilka det viktade genomsnittet av återförsäljningspriserna för torkade druvor anses vara importpriset. För att förhindra en artificiell minskning av skyddet bör det föreskrivas att importpålagor motsvarande införselskatt och indirekta skatter som faktiskt betalas vid import skall dras av från de noterade återförsäljningspriserna. I artikel 2.6 i samma förordning definieras %quot%slutanvändare%quot%. De tillverkare som förpackar produkten i detaljhandelsförpackning kan inte omfattas av detta begrepp, för även om sådan förpackning och presentation resulterar i en förändring av KN-numret kan detta inte anses vara bearbetning vid tillämpningen av den här förordningen.
I artikel 6 i förordning (EEG) nr 2054/89 föreskrivs om ett särskilt kontrollförfarande. Erfarenheten visar att när det förfarandet tillämpas bör varornas övergång till fri omsättning endast tillåtas efter ställande av den säkerhet som föreskrivs i artikel 248 i kommissionens förordning (EEG) nr 2454/93 av den 2 juli om tillämpningsföreskrifter för rådets förordning (EEG) nr 2913/92 om inrättandet av en tullkodex för gemen-skapen(5), senast ändrad genom förordning (EEG) 2193/94(6). Den säkerheten bör krävas om tullmyndigheterna hyser några tvivel om att importpriset är korrekt, även före de kontroller som föreskrivs i artikel 248. I fråga om kontroller i efterhand bör det klargöras att mått och steg avses vidtas för att återvinna förfallna tullavgifter i enlighet med artikel 220 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(7). Därutöver bör det klargöras att ränta skall betalas på förfallna tullavgifter enligt samtliga kontrollförfaranden.
I artikel 7.1 i förordning (EEG) nr 2054/89 föreskrivs de villkor enligt vilka det bedöms att minimipriset vid import skall följas. Erfarenheten visar att för undvikande av störningar måste hänsyn tas till de importpålagor som faktiskt betalas och till kostnaden för eventuell behandling som den importerade produkten genomgår efter import och före försäljning till slutkonsumenten.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för bearbetade produkter av frukt och grönsaker.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 2054/89 ändras på följande sätt:
1. Artikel 2 skall ändras enligt följande:
a) Punkt 3 skall ersättas med följande:
%quot%3. Om det upptäcks att priserna vid detaljhandelsförsäljning eller via mellanhänder, efter avdrag för de importpålagor som faktiskt betalats, är lägre än minimipriset i fråga om mer än 15 % av en importerad försändelse, skall det viktade genomsnittet av dessa justerade priser anses vara importpriset.%quot%
b) Punkt 6 skall ersättas med följande:
%quot%6. Vid tillämpningen av denna förordning avses med slutanvändare antingen en tillverkare som använder den berörda produkten för att bearbeta den på annat sätt än genom förpackning till en produkt som omfattas av ett annat KN-nummer än det som anges i försäkran om övergång till fri omsättning, eller en detaljhandlare som säljer endast till konsumenter.%quot%
2. Artikel 6 skall ersättas med följande:
%quot%Artikel 6
1. När tullmyndigheterna hyser välgrundade tvivel om att det pris som anges i försäkran om övergång till fri omsättning avspeglar det faktiska importpriset, skall de tillåta övergång till fri omsättning först efter det att importören har ställt den säkerhet som avses i artikel 248.1 i förordning (EEG) nr 2454/93, plus ränta för den period på sex månader som avses i andra stycket. Den tillämpliga räntesatsen skall vara den dröjsmålsränta som gäller enligt nationell lagstiftning.
Importörer skall ha sex månader på sig att bevisa att produkten har avsatts på villkor som säkerställer att minimipriset vid import följs. Om denna tidsfrist inte iakttas skall detta leda till att säkerheten förverkas, utan att det påverkar tillämpningen av bestämmelserna i punkt 2.
2. Den tidsfrist som fastställs i punkt 1 får av de behöriga myndigheterna förlängas med upp till tre månader efter en välgrundad ansökan från importören, förutsatt att säkerheten justeras i enlighet härmed.%quot%
3. Artikel 7.1 skall ersättas med följande:
%quot%1. Minimipriset vid import skall anses följas om importören företer bevis avseende minst 95 % av den importerade försändelsen om att produkten i alla saluföringsled har sålts till ett pris som lägst motsvarar minimipriset vid import efter avdrag för de faktiskt betalade importpålagorna. Om produkten genomgår behandling efter dess övergång till fri omsättning och innan den säljs till slutkonsumenten, skall kostnaden för den behandlingen avspeglas i försäljningspriset till slutanvändaren.%quot%
4. Artikel 10 skall ersättas med följande:
%quot%Artikel 10
Om den behöriga myndigheten vid en kontroll upptäcker att minimipriset vid import inte har följts skall de driva in de förfallna avgifterna i enlighet med artikel 220 i förordning (EEG) nr 2913/92. Vid fastställandet av det avgiftsbelopp som skall återvinnas eller som återstår att återvinna skall de ta hänsyn till den ränta som uppkommer från och med dagen för varornas övergång till fri omsättning till dagen för återvinning. Den räntesats som skall tillämpas skall vara den dröjsmålsränta som gäller enligt nationell lagstiftning.%quot%
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS FÖRORDNING (EG) nr 2965/94 av den 28 november 1994 om upprättande av ett översättningscentrum för Europeiska unionens organ
EUROPEISKA GEMENSKAPERNAS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 235 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande, och
med beaktande av följande: I samband med antagandet av beslutet av den 29 oktober 1993, som träffades genom ett gemensamt avtal mellan representanterna för medlemsstaternas regeringar, samlade på stats- och regeringschefsnivå, om lokaliseringen av vissa av de europeiska gemenskapernas organ och tjänster samt av Europol (), antog dessa representanter genom ett gemensamt avtal en deklaration om upprättande under kommissionens översättningstjänst i Luxemburg av ett översättningscentrum för unionens organ, som skall utföra det nödvändiga översättningsarbetet för de organ vars lokalisering fastställs genom beslutet av den 29 oktober 1993, med undantag för det Europeiska monetära institutet.
Upprättandet av ett gemensamt centrum är en praktisk lösning på problemet med att tillfredsställa översättningsbehoven för ett stort antal organ som ligger utspridda över hela unionens område.
Reglerna för översättningscentrumet skall göra det möjligt för detta att arbeta åt organ som har status som juridisk person, självständig förvaltning och egen budget, samtidigt som den arbetsmässiga förbindelsen mellan centrumet och kommissionen upprätthålls.
Fördraget anger inte andra befogenheter för antagandet av denna förordning än de som finns i artikel 235.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Ett översättningscentrum för unionens organ (i det följande betecknat %quot%centrumet%quot%) inrättas härmed.
Artikel 2
1. Centrumet skall utföra det nödvändiga översättningsarbetet för följande organ:
- Europeiska miljöbyrån,
- Europeiska yrkesutbildningsstiftelsen,
- Europeiska centrumet för kontroll av narkotika och narkotikamissbruk,
- Europeiska läkemedelsmyndigheten,
- Europeiska arbetsmiljöbyrån,
- Byrån för harmonisering av den inre marknaden (varumärken, mönster och modeller),
- Europol och Europols narkotikaenhet.
Centrumet och vart och ett av de ovannämnda organen skall utarbeta ordningar för det inbördes samarbetet.
2. Andra organ inrättade av rådet, förutom de i punkt 1 nämnda, kan också anlita centrumet på grundval av överenskommelser med centrumet.
Artikel 3
1. Centrumet skall vara en juridisk person.
2. För att centrumet skall kunna utföra de uppgifter som det tilldelas, skall det i varje medlemsstat ha den mest vittgående rättskapacitet som tillerkänns juridiska personer enligt den nationella lagstiftningen.
Artikel 4
1. Centrumet skall ha en styrelse som består av
a) en representant från vart och ett av de organ som nämns i artikel 2.1; var och en av de överenskommelser som avses i artikel 2.2 kan innehålla bestämmelser om att det organ som överenskommelsen gäller för skall vara representerat
b) en representant från var och en av Europeiska unionens medlemsstater, och
c) två representanter från kommissionen.
2. Det skall utses suppleanter för de i punkt 1 nämnda representanterna.
3. En av kommissionens representanter skall besätta ordförandeposten i styrelsen.
Artikel 5
1. Styrelseledamöterna skall utses för tre år.
2. Styrelseledamöterna kan väljas om.
Artikel 6
1. Ordföranden skall sammankalla ett styrelsemöte minst två gånger om året och när minst en tredjedel av de ledamöter som avses i artikel 4.1 a så kräver.
2. Styrelsens beslut skall fattas med två tredjedels majoritet.
3. Varje styrelseledamot skall ha en röst.
4. Ordföranden skall inte delta i omröstningar.
Artikel 7
Styrelsen skall anta sin egen arbetsordning.
Artikel 8
1. Styrelsen skall anta centrumets årliga arbetsprogram på grundval av ett utkast utarbetat av direktören.
2. Programmet kan anpassas under årets lopp i enlighet med förfarandet i punkt 1.
3. Senast den 31 januari varje år skall styrelsen anta en årsberättelse om centrumets verksamhet. Direktören skall skicka denna till de organ som anges i artikel 2 och till Europaparlamentet, rådet, kommissionen och revisionsrätten.
Artikel 9
1. Centrumet skall ledas av en direktör som utnämns av styrelsen på förslag av kommissionen för en femårsperiod, som kan förlängas.
2. Direktören skall vara laglig företrädare för centrumet. Han eller hon skall ansvara för
- utarbetande och genomförande på lämpligt sätt av arbetsprogrammet och av styrelsens beslut,
- den löpande förvaltningen,
- utförandet av de uppgifter som åläggs centrumet,
- genomförandet av budgeten,
- alla personalfrågor,
- förberedelse av styrelsens möten.
3. Direktören skall avlägga rapport till styrelsen om sin verksamhet.
Artikel 10
1. För varje budgetår, vilket motsvarar kalenderåret, skall det utarbetas beräkningar över alla centrumets inkomster och utgifter, vilka uppförs i centrumets budget.
2. a) Det skall råda balans mellan inkomster och utgifter i budgeten.
b) Om inte annat följer av bestämmelserna i c) skall centrumets inkomster bestå av betalning för tjänster från de organ som centrumet betjänar.
c) Under inkörningsperioden, som inte skall överstiga tre budgetår
- bidrar de organ som centrumet betjänar med ett fast belopp som på grundval av så goda faktaupplysningar som möjligt beräknas som en viss procentandel av deras budget, och som kommer att justeras med ledning av det faktiskt utförda arbetet,
- kan det utbetalas ett driftsbidrag till centrumet från Europeiska gemenskapernas allmänna budget.
3. Centrumets utgifter omfattar bl.a. löner till personalen, utgifter för administration och infrastruktur samt driftsutgifter.
Artikel 11
1. Före den översyn som behandlas i artikel 19 kan vart och ett av de i artikel 2.1 nämnda organen som känner av särskilda svårigheter när det gäller centrumets tjänster, vända sig till centrumet för att försöka finna bästa möjliga lösning på dessa svårigheter.
2. Om det visar sig omöjligt att finna en lösning inom tre månader, kan organet sända kommissionen ett meddelande med utförliga motiveringar så att kommissionen kan vidta nödvändiga åtgärder och vid behov under centrumets insyn och med dess bistånd ordna så att tredje man på ett mer systematiskt sätt tas till hjälp vid översättning av dokumenten i fråga.
Artikel 12
Kommissionen skall på grundval av avtal som ingås med centrumet mot återbetalning av kostnaderna förse centrumet med följande bistånd:
1) Stödfunktioner: terminologi, databaser, dokumentation, maskinöversättning, utbildning och listor över frilansöversättare samt utstationering av medarbetare till tjänster vid centrumet.
2) Förvaltning av grundläggande administrativa tjänster: utbetalning av löner, sjukförsäkring, pensionsplaner, social service.
Artikel 13
1. Direktören skall senast den 31 mars varje år utarbeta ett utkast till beräkningar av centrumets inkomster och utgifter för det kommande budgetåret. Utkastet skall överlämnas till styrelsen tillsammans med en tjänsteförteckning.
2. Styrelsen skall anta beräkningarna tillsammans med tjänsteförteckningen och omedelbart överlämna dessa till kommissionen, som på grundval därav skall göra beräkningar, motsvarande stödet till de organ som förtecknas i artikel 2, i det preliminära budgetförslag som skall föreläggas rådet i enlighet med artikel 203 i fördraget.
3. Styrelsen skall anta centrumets budget före budgetårets början, och vid behov anpassa den till utbetalningarna från de organ som nämns i artikel 2.
Artikel 14
1. Direktören skall genomföra budgeten.
2. Kommissionens styrekonom skall övervaka åtaganden och betalningar av alla centrumets utgifter samt att alla centrumets inkomster fastställs och inkasseras.
3. Senast den 31 mars varje år skall direktören överlämna räkenskaperna för centrumets inkomster och utgifter för det föregående året till kommissionen, styrelsen och revisionsrätten. Revisionsrätten skall granska dessa i enlighet med artikel 188c i fördraget.
4. Styrelsen skall bevilja direktören ansvarsfrihet för genomförandet av budgeten.
Artikel 15
Styrelsen skall efter att ha hört kommissionen och revisionsrätten anta interna finansiella bestämmelser, som bl.a. närmare anger hur centrumets budget skall ställas upp och genomföras.
Artikel 16
Protokollet om immunitet och privilegier för Europeiska gemenskaperna skall tillämpas på centrumet.
Artikel 17
1. Centrumets personal skall omfattas av de regler och föreskrifter som gäller för tjänstemän och övriga anställda inom Europeiska gemenskaperna.
2. Centrumet skall gentemot sin personal utöva de befogenheter som tillkommer en anställande myndighet.
3. Styrelsen skall anta lämpliga tillämpningsbestämmelser i samråd med kommissionen, bl.a. för att säkerställa skyddet av vissa uppgifters förtrolighet.
Artikel 18
1. Centrumets ansvar i kontraktsförhållanden skall bestämmas av den lagstiftning som tillämpas på kontraktet i fråga.
Europeiska gemenskapernas domstol skall vara behörig att träffa avgöranden i enlighet med en skiljedomsklausul som ingår i ett kontrakt som centrumet ingått.
2. Vad gäller ansvar utanför kontraktsförhållanden skall centrumet gottgöra alla skador som orsakats av dess anställda under tjänsteutövning, i enlighet med de allmänna principer som är gemensamma för medlemsstaternas lagstiftning.
Europeiska gemenskapernas domstol skall ha behörighet att pröva tvister som rör ersättning för sådana skador.
3. Det personliga ansvaret för centrumets anställda skall regleras av de bestämmelser som gäller för dem.
Artikel 19
Rådet kan på förslag av kommissionen och efter att ha hört Europaparlamentet ta upp denna förordnings regler för centrumets drift och funktion till översyn senast tre år efter utgången av centrumets inkörningsperiod, vilken inte får överstiga tre budgetår.
Artikel 20
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS FÖRORDNING (EG) nr 3383/94 av den 19 december 1994 om vissa förfaranden för tillämpning av Europaavtalet om associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Bulgarien, å andra sidan
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 113 i detta,
med beaktande av kommissionens förslag, och
med beaktande av följande: Ett Europaavtal om associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Bulgarien, å andra sidan, nedan kallat %quot%avtalet%quot%, undertecknades i Bryssel den 8 mars 1993.
I avvaktan på att Europaavtalet skall träda i kraft har dess bestämmelser om handel och handelsfrågor trätt i kraft sedan den 31 december 1993 genom ett interimsavtal om handel och handelsfrågor mellan Europeiska ekonomiska gemenskapen och Europeiska kol- och stålgemenskapen, å ena sidan, och Bulgarien, å andra sidan, som undertecknades i Bryssel den 8 mars 1993(1).
I enlighet med slutsatserna från Europeiska rådets möte i Köpenhamn den 21 och 22 juni 1993 om nya handelsåtaganden för länderna i central- och östeuropa undertecknades ett tilläggsprotokoll den 20 december 1993(2) av Europeiska gemenskaperna och Europeiska kol- och stålgemenskapen, å ena sidan, och Bulgarien, å andra sidan.
Det är nödvändigt att fastställa förfaranden för tillämpning av vissa av avtalets bestämmelser.
I fråga om skyddsåtgärder vid handel är det lämpligt att, i de fall bestämmelserna i Europaavtalet så kräver, fastställa särskilda bestämmelser avseende de allmänna regler som särskilt föreskrivs i rådets förordning (EG) nr 518/94 av den 7 mars 1994 om gemenskapsregler för import(3) och i rådets förordning (EG) nr 521/94 av den 7 mars 1994 om skydd mot dumpad eller subventionerad import från länder som inte är medlemmar i Europeiska ekonomiska gemenskapen(4).
Vid övervägandet av huruvida en skyddsåtgärd bör införas, bör hänsyn tas till de åtaganden som föreskrivs i Europaavtalet.
De förfaranden avseende skyddsklausuler som fastställs i Fördraget om upprättandet av Europeiska gemenskapen är likaledes tillämpliga.
Särskilda bestämmelser om skyddsåtgärder har antagits för textilprodukter som omfattas av protokoll 1 till avtalet.
Vissa särskilda förfaranden bör införas för tillämpningen av skyddsåtgärder på jordbruksområdet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
AVDELNING I Jordbruksprodukter
Artikel 1
För de jordbruksprodukter som omfattas av bilaga II till fördraget och som inom ramen för organisationen av den gemensamma marknaden är belagda med importavgifter, och för de produkter som omfattas av KN-numren 0711 90 50 och 2003 10 10 skall bestämmelser för tillämpning av artikel 21.2 och 21.4 i avtalet antas i enlighet med det förfarande som föreskrivs i artikel 23 i förordning (EG) nr 1766/92(5) eller i motsvarande bestämmelser i andra förordningar om upprättandet av en gemensam organisation av jordbruksmarknaderna. Dessa bestämmelser kan föreskriva införandet av ett system med importlicenser på de områden där den gemensamma organisationen av jordbruksmarknaderna inte föreskriver sådana licenser.
AVDELNING II Skyddsåtgärder
Artikel 2
I enlighet med de förfaranden som föreskrivs i artikel 113 i fördraget får rådet hänskjuta beslut om de åtgärder som fastställs i artiklarna 29 och 118.2 i avtalet till det associationsråd som inrättats genom avtalet. Vid behov skall rådet vidta dessa åtgärder i enlighet med samma förfarande.
Kommissionen kan på eget initiativ eller på begäran av en medlemsstat lägga fram de förslag som är nödvändiga för detta ändamål.
Artikel 3
1. I händelse av ett förfarande som kan berättiga gemenskapen att vidta de åtgärder som föreskrivs i artikel 64 i avtalet, skall kommissionen, efter att ha utrett ärendet, på eget initiativ eller på begäran av en medlemsstat avgöra om ett sådant förfarande är förenligt med avtalet. Vid behov skall den föreslå rådet att vidta skyddsåtgärder, och rådet skall då handla i enlighet med förfarandet i artikel 113 i fördraget, utom i de fall det gäller stöd som omfattas av förordning (EG) nr 521/94, då åtgärder skall vidtas i enlighet med de förfaranden som fastställs i den förordningen. Åtgärder skall endast vidtas på de villkor som fastställs i artikel 64.6 i avtalet.
2. I händelse av ett förfarande som kan medföra att Bulgarien vidtar åtgärder mot gemenskapen på grundval av artikel 64 i avtalet, skall kommissionen efter att ha utrett ärendet avgöra om förfarandet är förenligt med de principer som fastställs i avtalet. Vid behov skall den fatta lämpliga beslut på grundval av de kriterier som följer av tillämpningen av artiklarna 85, 86 och 92 i fördraget.
Artikel 4
I händelse av ett förfarande som kan berättiga gemenskapen att tillämpa de åtgärder som fastställs i artikel 30 i avtalet, skall beslut om införandet av antidumpningsåtgärder fattas i enlighet med bestämmelserna i förordning (EG) nr 521/94 och förfarandena i artikel 34.2 och 34.3 b eller 34.3 d i avtalet.
Artikel 5
1. Om en medlemsstat begär att kommissionen skall vidta skyddsåtgärder i enlighet med artiklarna 31 eller 32 i avtalet, skall den till stöd för sin begäran förse kommissionen med de upplysningar som är nödvändiga för att berättiga detta. Om kommissionen beslutar att inte vidta skyddsåtgärder skall den meddela rådet och medlemsstaterna detta inom fem arbetsdagar efter det att medlemsstatens begäran mottagits.
Varje medlemsstat får hänskjuta ett sådant kommissionsbeslut till rådet senast tio arbetsdagar efter meddelandet om detta beslut.
Om rådet med kvalificerad majoritet tillkännager att det avser att fatta ett annat beslut skall kommissionen omedelbart underrätta Bulgarien om detta och meddela att samråd i associationsrådet skall inledas i enlighet med artikel 34.2 och 34.3 i avtalet.
Rådet kan med kvalificerad majoritet fatta ett annat beslut senast tjugo arbetsdagar efter det att samråden med Bulgarien har avslutats i associationsrådet.
2. Kommissionen skall biträdas av den kommitté som inrättats genom förordning (EG) nr 3491/93(6), nedan kallad %quot%kommittén%quot%.
Kommittén skall sammanträda på kallelse av dess ordförande. Denne skall snarast möjligt förse medlemsstaterna med alla ändamålsenliga upplysningar.
3. Om kommissionen på eget initiativ eller på begäran av en medlemsstat beslutar att de skyddsåtgärder som fastställs i artiklarna 31 eller 32 i avtalet bör vidtas, skall den
- omedelbart underrätta medlemsstaterna om den handlar på eget initiativ eller om den efterkommer en medlemsstats begäran inom fem arbetsdagar efter det att denna begäran mottagits,
- samråda med kommittén,
- samtidigt informera Bulgarien om detta och meddela associationsrådet att samråd inleds i enlighet med artikel 34.2 och 34.3 i avtalet,
- samtidigt förse associationsrådet med samtliga upplysningar som är nödvändiga för dessa samråd.
4. Under alla omständigheter skall samråden inom associationsrådet anses vara avslutade inom 30 dagar efter det meddelande som avses i punkt 1 fjärde stycket och i punkt 3.
När samråden avslutas eller när tidsfristen om 30 dagar löper ut kan kommissionen, om det visar sig att inga andra arrangemang är möjliga, efter samråd med kommittén vidta lämpliga åtgärder för att sätta artiklarna 31 och 32 i avtalet i kraft.
5. Det beslut som avses i punkt 4 skall omedelbart meddelas rådet, medlemsstaterna och Bulgarien. Det skall även meddelas associationsrådet.
Beslutet skall vara direkt tillämpligt.
6. Varje medlemsstat får hänskjuta kommissionens beslut enligt punkt 4 till rådet inom tio dagar efter det att beslutet meddelats.
7. Om kommissionen inte har fattat ett beslut i enlighet med punkt 4 andra stycket inom 10 arbetsdagar efter det att den tidsfrist om 30 dagar som anges i den punkten har löpt ut, kan varje medlemsstat som har hänskjutit ärendet till kommissionen i enlighet med punkt 3 hänskjuta det till rådet.
8. I de fall som avses i punkterna 6 och 7 kan rådet med kvalificerad majoritet fatta ett annat beslut inom två månader.
Artikel 6
1. Vid undantagsfall enligt artikel 34.3 d i avtalet kan kommissionen vidta omedelbara skyddsåtgärder för de fall som anges i artiklarna 31 och 32 i avtalet.
2. Om kommissionen får en begäran av en medlemsstat skall den fatta beslut senast fem arbetsdagar efter det att begäran mottagits.
Kommissionen skall meddela rådet och medlemsstaterna sitt beslut.
3. Varje medlemsstat kan hänskjuta kommissionens beslut till rådet i enlighet med förfarandet i artikel 5.6.
Förfarandet i artikel 5.7 och 5.8 skall tillämpas.
Om kommissionen inte har fattat något beslut inom den tidsfrist som anges i punkt 2, kan varje medlemsstat som hänskjutit ärendet till kommissionen hänskjuta det till rådet i enlighet med de förfaranden som fastställs i första och andra stycket i denna punkt.
Artikel 7
Förfarandena i artiklarna 5 och 6 skall inte tillämpas på de produkter som omfattas av protokoll 1 till avtalet.
Artikel 8
När omständigheterna kräver att åtgärder vidtas för jordbruksprodukter på grundval av artiklarna 22 eller 31 i avtalet eller på grundval av bestämmelserna i de bilagor som omfattar dessa produkter, skall dessa åtgärder, trots artiklarna 5 och 6, vidtas i enlighet med de förfaranden som fastställs i bestämmelserna om upprättandet av den gemensamma organisationen av jordbruksmarknaderna, eller i de särskilda bestämmelser som antagits enligt artikel 235 i fördraget för produkter som framställs genom bearbetning av jordbruksprodukter, under förutsättning att de villkor som fastställs i artiklarna 22 eller 34.2 och 34.3 i avtalet uppfylls.
Artikel 9
Meddelanden till associationsrådet i enlighet med avtalet skall lämnas av kommissionen på gemenskapens vägnar.
Artikel 10
Denna förordning utesluter inte att de skyddsåtgärder som föreskrivs i Fördraget om upprättandet a
RÅDETS DIREKTIV 95/7/EG av den 10 april 1995 om ändring av direktiv 77/388/EEG och om införande av nya förenklingsåtgärder avseende mervärdeskatt - tillämpningsområde för vissa undantag från beskattning och praktiska åtgärder för genomförandet
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 99 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande,
med beaktande av Ekonomiska och sociala kommitténs yttrande, och
med beaktande av följande: Den inre marknadens effektivitet kan förbättras genom att gemensamma regler införs som klargör tillämpningsområdet och de närmare reglerna för genomförandet av några av de undantag från beskattning som behandlas i artiklarna 14.1, 15.2 och 16.1 i rådets sjätte direktiv (77/388/EEG) av den 17 maj 1977 om harmonisering av medlemsstaternas lagstiftning rörande mervärdeskatt: enhetlig beräkningsgrund (1). Fastställandet av sådana gemensamma regler föreskrivs i direktivet, särskilt i artiklarna 14.2 och 16.3.
Enligt artikel 3 i rådets direktiv 92/111/EEG av den 14 december 1992 om ändring av direktiv 77/388/EEG och om vidtagande av åtgärder för att förenkla mervärdeskatten (2), skall särskilda regler för beskattning av kedjetransaktioner mellan skattskyldiga antas. Dessa regler skall garantera såväl att principen om det allmänna mervärdeskattesystemets neutralitet med avseende på varors och tjänsters ursprung respekteras som att de principer som valts för mervärdeskatten och kontrollsystemet under övergångsperioden respekteras.
Alla omkostnader som avser transport av varor till destinationsorten inom gemenskapen, i de fall då orten är känd vid den tidpunkt då importen görs, bör inkluderas i skatteunderlaget avseende import. Dessa tjänster skall därför undantas från beskattning enligt vad som föreskrivs i artikel 14.1 i) i direktiv 77/388/EEG.
I artikel 15.2 i det nämnda direktivet föreskrivs att kommissionen skall lägga fram förslag för rådet att fastställa gemensamma skatteregler som klart anger tillämpningsområdet och de praktiska åtgärderna vid genomförandet av de undantag från beskattning vid export som är tillämpliga på leveranser av varor som medförs med resandes personliga bagage.
Den period som ligger till grund för den beräkning av jämkningen som anges i artikel 20.2 i nämnda direktiv bör av medlemsstaterna kunna förlängas till 20 år när det gäller fasta anläggningstillgångar, med hänsyn till dessas ekonomiska livslängd.
Medlemsstater som den 1 januari 1993 tillämpade den skattesats som gäller för varor som framställs genom beställningsarbete bör få fortsätta att göra det.
Reglerna om leveransort och beskattning på området för tillhandahållande av transporttjänster inom gemenskapen fungerar smidigt och tillfredsställande både för företagarna och myndigheterna i medlemsländerna.
Om transporter av varor inom ett medlemsland, som är direkt anknutna till transporter mellan medlemsländerna jämställs med transporter inom gemenskapen, blir det möjligt att förenkla principerna och reglerna för beskattning inte bara av dessa inre transporttjänster utan också för andra tjänster som är knutna till dessa, liksom för de tjänster som utförs av mellanhänder.
Förfarandet att anse vissa arbeten på lös egendom som beställningsarbeten har givit upphov till vissa svårigheter, varför det bör upphöra.
För att underlätta handeln inom gemenskapen på området för arbete på lösegendom bör beskattningsformerna för dessa arbeten ändras när de utförs för kunder som är registrerade för mervärdeskatt i en annan medlemsstat än den där arbetet faktiskt utförs.
Bestämmelserna i artikel 16.1 punkterna B-E i direktivet jämförda med bestämmelserna i artikel 22.9, som rör viss skattebefrielse, gör det möjligt att lösa de problem som företagare möter när de deltar i kedjetransaktioner som avser egendom som har placerats och lagrats i enlighet med ett upplagsförfarande.
I detta sammanhang är det nödvändigt att säkerställa att den skattemässiga behandling som tillämpas på leveranser av varor och på till vissa varor knutna tillhandahållanden av tjänster, som kan hänföras till ett tullupplagsförfarande, också kan gälla för transaktioner rörande varor som är föremål för annat upplagsförfarande än tullupplagsförfarande.
Eftersom dessa transaktioner framför allt avser råvaror och andra varor som inköpts på de internationella terminsmarknaderna bör det upprättas en förteckning över alla varor som omfattas av dessa bestämmelser.
Förutsatt att samrådsförfarandet med Rådgivande kommittén för mervärdeskatt iakttas, ankommer det på medlemsstaterna att ange vilka dessa andra lagringsförfaranden är. Icke desto mindre är det nödvändigt att utesluta varor, som är avsedda för leverans i detaljhandelsledet, från sådana förfaranden.
Det är nödvändigt att närmare ange vissa beskattningsregler enligt de i artikel 16.1 punkterna B-E i direktivet nämnda förfarandena, särskilt såvitt avser beräkningen av avgiftsbeloppen.
Det är nödvändigt att närmare ange innebörden av bestämmelserna i artikel 17.2 a) i direktivet om vilka åtgärder som kan användas under den i artikel 28 l nämnda övergångsperioden.
Följaktligen bör direktiv 77/388/EEG ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 77/388/EEG ändras på följande sätt:
1) Artikel 5.5 skall ersättas med följande text:
%quot%5. Medlemsstaterna får betrakta överlämnandet av vissa byggnadsarbeten som en leverans i den betydelse som begreppet har enligt punkt 1.%quot%
2) Artikel 11B.3b), tredje stycket, skall ersättas med följande:
%quot%De bikostnader som avses ovan skall också inkluderas i det beskattningsunderlaget på de härrör från transport till en annan bestämmelseort inom gemenskapens territorium om denna är känd när skattskyldigheten inträder.%quot%
3) Artikel 15.2, andra och tredje styckena, skall ersättas med följande tre stycken:
%quot%I fall leveransen avser varor som medförs i resenärers personliga bagage skall detta undantag tillämpas förutsatt att:
- resenären inte är etablerad inom gemenskapen,
- varorna transporteras ut ur gemenskapen före utgången av den tredje månaden efter den månad då leveransen genomförs,
- leveransen sammanlagda värde inklusive mervärdeskatt överstiger motvärdet i nationell valuta av 175 ecu, fastställt i enlighet med artikel 7.2 i direktiv 69/169/EEG (*). Medlemsstaterna får emellertid undanta en leverans vars sammanlagda värde är lägre än detta belopp.
För tillämpningen av andra stycket gäller följande:
- med en resenär som inte är etablerad inom gemenskapen avses en resenär vars hemvist eller stadigvarande vistelseort inte är belägen inom gemenskapen. I denna bestämmelse avses med %quot%hemvist eller stadigvarande vistelseort%quot% den plats som anges som sådan i pass, identitetskort eller någon annan identitetshandling som den medlemsstat, inom vilken leveransen äger rum, godkänner som identitetshandling,
- bevis om utförsel skall framläggas i form av fakturan eller jämförbar handling som skall vara påtecknad av det tullkontor där varorna lämnade gemenskapen.
Varje medlemsstat skall till kommissionen översända prov på de stämplar som den använder för det påtecknande som anges i tredje stycket andra strecksatsen. Kommissionen skall vidarebefordra denna information till skattemyndigheterna i de övriga medlemsstaterna.
(*) EGT nr L 133, 4.6.1969, s. 6, senast ändrat genom direktiv 94/4/EG (EGT nr L 60, 3.3.1994, s. 14).%quot%4) I artikel 20.2 skall det sista stycket ersättas med följande text: %quot%När det gäller fast egendom förvärvad som anläggningstillgångar kan jämkningsperioden förlängas till högst 20 år.%quot%
5) I artikel 28.2h) skall följande led läggas till:
%quot%h) Medlemsstaterna som den 1 januari 1993 använde sig av den i artikel 5.5a) i dess dåvarande lydelse angivna möjligheten får på leveranser enligt avtal om beställningsarbete tillämpa den skattesats som är tillämplig på den vara som frambringas genom beställningsarbetet.
För tillämpningen av denna bestämmelse avses med leveranser enligt ett avtal leverans av beställningsarbete att den som har åtagit sig arbetet till sin kund levererar lös egendom som han har gjort färdigt eller satt samman med hjälp av material eller föremål som kunden i detta syfte har ställt till hans förfogande, oavsett om den som har åtagit sig arbetet har levererat en del av det använda materialet eller inte.%quot%
6) Artikel 28a.5 skall ändras på följande sätt:
- den inledande meningen skall ersättas med följande:
%quot%Följande skall betraktas som leverans av varor mot vederlag:%quot%,
- a) skall utgå,
- fjärde strecksatsen i andra stycket av b) skall utgå,
- femte strecksatsen i andra stycket av b) skall erstättas med följande text:
%quot%- tillhandahållande av en tjänst som utförts åt den skattskyldiga personen och som innebär att arbete på varorna faktiskt har utförts i den medlemsstat dit de skickats eller transporterats förutsatt att varorna sedan arbetet utförts återsänds till den skattskyldige i den medlemsstat från vilken de ursprungligen avsändes eller transporterades%quot%.
7) Artikel 28b skall ändras på följande sätt:
- i den första strecksatsen i C 1 skall följande stycke införas:
%quot%Transport av varor där avgångsorten och ankomstorten är belägna inom landets territorium skall jämställas med transport av varor inom gemenskapen när sådan transport är direkt förbunden med en transport av varor där avgångsorten och ankomstorten är belägna inom två olika medlemsstaters territorier.%quot%
- följande avsnitt skall införas:
%quot%F. Platsen för utförande av tjänster i fråga om värderingar av eller arbete på lösegendom Genom undantag från artikel 9.2c) skall platsen för utförande av tjänster som innefattar värderingar eller arbete på lös egendom som tillhandahålls kunder som är registrerade för mervärdeskatt i en annan medlemsstat än den där dessa tjänster faktiskt utförs vara belägen i den medlemsstat som till kunden utfärdade det registreringsnummer för mervärdeskatt under vilket tjänsterna utfördes för denne.
Detta undantag skall inte tillämpas när varorna inte sänds eller transporteras ut ur den medlemsstat där tjänsterna utfördes.%quot%
8) I artikel 28c.Aa) första punkten skall orden %quot%såsom det definieras i artikel 28a.5a)%quot% utgå.
9) Artikel 28c.E första stycket skall ersättas med följande:
%quot%1) I artikel 16,
- skall punkt 1 ersättas med följande:
'1. Utan att det påverkar tillämpningen av gemenskapens övriga skattebestämmelser får medlemsstaterna efter det samråd som föreskrivs i artikel 29 vidta särskilda åtgärder i syfte att undanta alla eller några av följande transaktioner, om de inte syftar till slutlig användning och/eller konsumtion och att summan av den mervärdeskatt som förfaller till betalning när varorna lämnar de i A och E uppräknade förfarandena eller ordningarna motsvarar det skattebelopp som skulle ha betalats om var och en av dessa transaktioner skulle ha beskattats inom landets territorium:
A. Införsel av varor som är avsedda att placeras i andra lager än tullager,
B. Leveranser av varor som är avsedda att:
a) visas upp för tullen och, i tillämpliga fall, placeras i tillfällig förvaring,
b) placeras i en frizon eller ett frilager,
c) placeras i tullagerförfarande eller aktivt förädlingsförfarande,
d) släppas in i territorialvattnen:
- för att införlivas i borrnings- eller produktionsplattformar i avsikt att konstruera, reparera, underhålla, ändra eller utrusta sådana plattformar, eller för att förbinda sådana borrnings- eller produktionsplattformar med fastlandet,
- för bunkring eller proviantering för borrnings- eller produktionsplattformar,
e) inom landets territorium behandlas enligt annat lagringsförfarande än tull-lagring.
Vid tillämpningen av denna artikel avses med andra lager än tullager:
- för punktskattepliktiga varor, de platser som definieras skatteupplag i artikel 4b) i rådets direktiv 92/12/EEG,
- för andra varor än punktskattepliktiga varor, de platser som av medlemsstaterna definieras som sådana. Medlemsstaterna får emellertid inte föreskriva om något annat lagringsförfarande än tullagring när de ifrågavarande varorna är avsedda att levereras till detaljhandelsledet.
Medlemsstaterna får ändå föreskriva om ett sådant förfarande för varor som är avsedda för:
- skattskyldiga personer med avseende på leveranser som genomförs enligt de villkor som anges i artikel 28k,
- butiker för skattefri försäljning i den betydelse som begreppet har enligt artikel 28k, och som är avsedda för tillhandahållande till resenärer som med flyg eller sjövägen beger sig till ett tredje land, och som är undantagna enligt artikel 15,
- skattskyldiga personer med avseende på leverans av varorna ombord på flygplan eller fartyg under en flygning eller överfart till en ankomstort som är belägen utanför gemenskapen,
- skattskyldiga personer såvitt avser skattefria leveranser som genomförs i enlighet med artikel 15.10.
De platser som avses i a), b), c) och d) skall vara de som definieras i gemenskapens gällande tullbestämmelser.
C. Tillhandahållande av tjänster som hänför sig till de leveranser av varor som avses i B,
D. leveranser av varor och tillhandahållande av tjänster som utförs:
a) på de platser som anges i B a), b), c) och d) som fortfarande omfattas av en av de situationer som anges där,
b) på de platser som anges i B e), inom landets territorium, omfattas av den situation som anges däri.
I den mån som de använder den möjlighet som anges i a) för transaktioner som genomförs i tullager skall medlemsstaterna vidta de nödvändiga åtgärderna för att säkerställa att de har definierat begreppet annat lagringsförfarande än tullagring på ett sätt som gör det möjligt att tillämpa bestämmelserna i b) på samma transaktioner avseende de varor som räknas upp i bilaga J och som genomförs i sådana lager som inte är tullager.
E. leveranser:
- av varor som avses i artikel 7.1a) som även i fortsättningen omfattas av förfaranden för tillfällig införsel med total befrielse från importtull eller av externt transiteringsförfarande,
- av varor som avses i artikel 7.1b) som fortfarande omfattas av gemenskapens interna transiteringsförfarande som anges i artikel 33a,
samt tillhandahållande av tjänster som hänför sig till sådana leveranser.
Genom undantag från artikel 21.1.a), första stycket, skall den person som är betalningsskyldig för den skatt som skall erläggas i enlighet med första stycket vara den person som är ansvarig för att varorna upphör att omfattas av de förfaranden eller situationer som anges i denna punkt.
När det förhållandet att varor upphör att omfattas av de förfaranden eller situationer som avses i denna punkt medför att import enligt artikel 7.3 föreligger, skall importmedlemsstaten vidta de nödvändiga åtgärderna för att undvika dubbelbeskattning inom landets territorium.`
- följande punkt skall tilläggas:
'1a. I den mån som de använder den möjlighet som anges i punkt 1 skall medlemsstaterna vidta de nödvändiga åtgärderna för att säkerställa att gemenskapsinterna förvärv av varor som är avsedda att omfattas av ett av de förfaranden eller en av de situationer som avses i punkt 1 B omfattas av samma bestämmelser som leveranser av varor som genomförs inom landet under motsvarande villkor.`%quot%
10) I artikel 28f.1 skall artikel 17.2 a) ersättas med följande:
%quot%a) mervärdeskatt som förfaller till betalning eller betalats inom landets territorium avseende varor eller tjänster som tillhandahållits, eller kommer att tillhandahållas, till honom av en annan skattskyldig person.%quot%
11) I artikel 28g skall artikel 21.1 b) ersättas med följande text:
%quot%b) personer till vilka tjänster som avses i artikel 9.2 e) tillhandahålls eller personer som är registrerade för mervärdeskatt inom landets territorium till vilka tjänster som avses i artikel 28 b, C, D, E och F tillhandahålls, om tjänsterna utförs av en skattskyldig person som är etablerad utomlands. Medlemsstaterna får emellertid kräva att den som tillhandahåller tjänsten skall vara solidariskt ansvarig för betalningen av skatten.%quot%
12) Artikel 28h skall ändras på följande sätt:
- artikel 22.2 b) skall ersättas med följande:
%quot%b) Varje skattskyldig person skall föra register över de varor som denne har avsänt eller transporterat eller som har avsänts eller transporterats för dennes räkning ut ur det territorium som anges i artikel 3 men inom gemenskapen med avseende på de transaktioner som avses i femte, sjätte och sjunde strecksatserna i artikel 28a.5 b).
Varje skattskyldig person skall föra tillräckligt detaljerade räkenskaper för att göra det möjligt att identifiera varor som avsänts till honom från en annan medlemsstat av en skattskyldig person eller på en skattskyldig persons vägnar, som är registrerad för mervärdeskatt i den andra medlemsstaten, i samband med tillhandahållande av en tjänst som avses i den tredje eller fjärde strecksatsen i artikel 9.2 c).%quot%
- den första strecksatsen i artikel 22.3 b) andra stycket skall ersättas med följande:
%quot%- vad gäller de transaktioner som avses i artikel 28b, C, D, E och F, det nummer under vilket den skattskyldiga personen är registrerad inom landets territorium och det nummer under vilket kunden är registrerad och under vilket tjänsten har överlämnats till denne.%quot%
- artikel 22.6 b) första stycket skall ersättas med följande:
%quot%Varje skattskyldig person som är registrerad för mervärdeskatt skall också överlämna en sammanställning över de köpare som är registrerade för mervärdeskatt till vilka han har levererat varor enligt de villkor som anges i artikel 28c.A a) och d) och över varumottagare som är registrerade för mervärdeskatt för de transaktioner som avses i femte stycket.%quot%
- andra strecksatsen i artikel 22.6 b) tredje stycket skall ersättas med följande:
%quot%- det nummer under vilket varje person som förvärvar varor registreras för mervärdeskatt i en annan medlemsstat och under vilket varorna levererades till honom%quot%,
- femte stycket i artikel 22.6 b) utgår.
13) Bilaga J som finns som bilaga till detta direktiv skall läggas till.
Artikel 2
1. Medlemsstaterna skall sätta i kraft de lagar, förordningar och bestämmelser som är nödvändiga för att följa detta direktiv den 1 januari 1996. De skall genast underrätta kommissionen om dessa.
När medlemsstaterna antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Utan hinder av punkt 1 första stycket får medlemsstater vidta åtgärder genom lagar, förordningar och bestämmelser för att sätta i kraft bestämmelserna i artikel 1.3, 1.4 och 1.9 senast den 1 januari 1996.
Tyskland och Luxemburg är emellertid berättigade att vidta åtgärder genom lagar, förordningar och andra bestämmelser för att tillämpa bestämmelserna i artikel 1.9 senast den 1 januari 1997.
3. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 3
Detta direktiv träder i kraft den tjugonde dagen efter det att det offentliggjorts i Europeiska gemenskapernas officiella tidning.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
KOMMISSIONENS FÖRORDNING (EG) nr 2931/95 av den 19 december 1995 om ändring av förordningarna (EEG) nr 804/68, (EEG) nr 2730/75, (EEG) nr 776/78, (EEG) nr 570/88, (EEG) nr 584/92, (EEG) nr 2219/92, (EG) nr 2883/94, (EG) nr 1466/95, (EG) nr 1598/95, (EG) nr 1600/95 och (EG) nr 1713/95 till följd av ändring av Kombinerade nomenklaturen i fråga om vissa mjölkprodukter
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 234/79 av den 5 februari 1979 om förfarandet vid anpassning av Gemensamma tulltaxenomenklaturen för jordbruksprodukter (1), ändrad genom förordning (EEG) nr 3209/89 (2), särskilt artikel 2.1 i denna,
med beaktande av rådets förordning (EEG) nr 804/68 av den 27 juni 1968 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter (3), senast ändrad genom förordning (EG) nr 1538/95 (4), särskilt artiklarna 13.3, 15.4, 16.1, 16.4 och 17.14 i denna,
med beaktande av rådets förordning (EEG) nr 518/92 av den 27 februari 1992 om vissa förfaranden vid tillämpning av interimsavtalet om handel och handelsfrågor mellan Europeiska ekonomiska gemenskapen och Europeiska kol- och stålgemenskapen å ena sidan och Polen å andra sidan (5), ändrad genom förordning (EEG) nr 2233/93 (6), särskilt artikel 1 i denna,
med beaktande av rådets förordning (EEG) nr 519/92 av den 27 februari 1992 om vissa förfaranden vid tillämpning av interimsavtalet om handel och handelsfrågor mellan Europeiska ekonomiska gemenskapen och Europeiska kol- och stålgemenskapen å ena sidan och Ungern å andra sidan (7), ändrad genom förordning (EEG) nr 2234/93 (8), särskilt artikel 1 i denna,
med beaktande av rådets förordning (EEG) nr 520/92 av den 27 februari 1992 om vissa förfaranden för tillämpningen av interimsavtalet om handel och handelsfrågor mellan Europeiska ekonomiska gemenskapen och Europeiska kol- och stålgemenskapen å ena sidan och Tjeckien och Slovakien å andra sidan (9), ändrad genom förordning (EEG) nr 2235/93 (10), särskilt artikel 1 i denna,
med beaktande av rådets förordning (EEG) nr 1600/92 av den 15 juni 1992 om särskilda bestämmelser för Azorerna och Madeira angående vissa jordbruksprodukter (11), senast ändrad genom kommissionens förordning (EG) nr 2537/95 (12), särskilt artiklarna 10 och 24.6 i denna,
med beaktande av rådets förordning (EEG) nr 1601/92 av den 15 juni 1992 om särskilda åtgärder för Kanarieöarna rörande vissa jordbruksprodukter (13), senast ändrad genom förordning (EG) nr 2537/95, särskilt artikel 3.4 i denna,
med beaktande av rådets förordning (EG) nr 1275/95 av den 29 maj 1995 om vissa förfaranden för tillämpning av avtalet om liberalisering av handeln och inrättandet av kompletterande åtgärder mellan Europeiska gemenskapen, Europeiska atomenergigemenskapen och Europeiska kol- och stålgemenskapen å ena sidan och Estland å andra sidan (14),
med beaktande av rådets förordning (EG) nr 1276/95 av den 29 maj 1995 om vissa förfaranden för tillämpning av avtalet om liberalisering av handeln och inrättandet av kompletterande åtgärder mellan Europeiska gemenskapen, Europeiska atomenergigemenskapen och Europeiska kol- och stålgemenskapen å ena sidan och Lettland å andra sidan (15),
med beaktande av rådets förordning (EG) nr 1277/95 av den 29 maj 1995 om vissa förfaranden för tillämpning av avtalet om liberalisering av handeln och inrättandet av kompletterande åtgärder mellan Europeiska gemenskapen, Europeiska atomenergigemenskapen och Europeiska kol- och stålgemenskapen å ena sidan och Litauen å andra sidan (16), och
med beaktande av följande: I kommissionens förordning (EG) nr 2448/95 om ändring av bilaga I till rådets förordning (EEG) nr 2658/87 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (17) fastställs ändringar i fråga om vissa mjölkprodukter från och med den 1 januari 1996. Även vissa andra KN-nummer för mjölkprodukter har senare ändrats.
Följaktligen bör de förordningar som berörs av ändringar av undernummer till dessa KN-nummer ändras, särskilt följande:
- Rådets förordning (EEG) nr 804/68.
- Rådets förordning (EEG) nr 2730/75 av den 29 oktober 1975 om glukos och laktos (18), ändrad genom kommissionens förordning (EEG) nr 222/88 (19).
- Kommissionens förordning (EEG) nr 776/78 av den 18 april 1978 om tillämpning av det lägsta bidragsbeloppet vid export av mejeriprodukter och om upphävande och ändring av vissa förordningar (20), senast ändrad genom förordning (EG) nr 1586/95 (21).
- Kommissionens förordning (EEG) nr 570/88 av den 16 februari 1988 om försäljningen av smör till sänkta priser och beviljandet av stöd för smör och koncentrerat smör avsett att användas i framställningen av konditorivaror, glass och andra livsmedel (22), senast ändrad genom förordning (EG) nr 1802/95 (23).
- Kommissionens förordning (EEG) nr 584/92 av de 6 mars 1992 om tillämpningsföreskrifter för importordningen i interimsavtalen mellan gemenskapen å ena sidan och Polen, Ungern, Tjeckien och Slovakien (24) å den andra vad avser mjölk och mjölkprodukter, senast ändrad genom förordning (EG) nr 2416/95 (25).
- Kommissionens förordning (EEG) nr 2219/92 av den 30 juli 1992 om tillämpningsföreskrifter för det särskilda försörjningssystemet för Madeira avseende mjölkprodukter och om fastställande av den förhandsberäknade försörjningsbalansen (26), senast ändrad genom förordning (EG) nr 2835/95 (27).
- Kommissionens förordning (EG) nr 2883/94 av den 28 november 1994 om upprättande av en prognostiserad försörjningsbalans för försörjningen av Kanarieöarna med de jordbruksprodukter som omfattas av den särskilda ordning som föreskrivs i artikel 2-5 i rådets förordning (EEG) nr 1601/92 (28), senast ändrad genom förordning (EG) nr 1820/95 (29).
- Kommissionens förordning (EG) nr 1466/95 av den 27 juni 1995 om särskilda tillämpningsföreskrifter för exportbidrag inom sektorn för mjölk och mjölkprodukter (30), ändrad genom förordning (EG) nr 2452/95 (31).
- Kommissionens förordning (EG) nr 1598/95 av den 30 juni 1995 om tillämpningsföreskrifter för systemet med tilläggsavgifter vid import inom sektorn för mjölk och mjölkprodukter (32).
- Kommissionens förordning (EG) nr 1600/95 av den 30 juni 1995 om tillämpningsföreskrifter för importordningen och om öppnande av tullkvoter inom sektorn för mjölk och mjölkprodukter (33), senast ändrad genom förordning (EG) nr 2537/95 (34).
- Kommissionens förordning (EG) nr 1713/95 av den 13 juli 1995 om tillämpningsföreskrifter inom sektorn för mjölk och mjölkprodukter för den ordning som fastställs i avtalen om liberalisering av handelsutbytet mellan gemenskapen och de tre baltiska staterna (35).
För klarhetens skull bör det fastställas att dessa ändringar träder i kraft den 1 januari 1996.
Förvaltningskommittén för mjölk och mjölkprodukter har inte yttrat sig inom den tid som dess ordförande har bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 804/68 ändras på följande sätt:
1. I artikel 1 skall uppgifterna i c, e och g ersättas med följande:
%gt%Plats för tabell%gt%
2) I artikel 17.12 skall KN-nummer %quot%2106 90 99%quot% ersättas med KN-nummer %quot%2106 90 98%quot%.
3) I artikel 26.5 skall KN-nummer %quot%0405 00%quot% ersättas med KN-nummer %quot%0405%quot%.
4) I bilagan skall följande ändringar göras:
- Följande uppgifter skall föras in efter uppgifterna enligt KN-nummer 0403:
%gt%Plats för tabell%gt%
- Uppgifterna enligt KN-nummer 1702 10 skall ersättas med följande:
%gt%Plats för tabell%gt%
- Uppgifterna enligt KN-nummer ex 1901 90 90 skall ersättas med följande:
%gt%Plats för tabell%gt%
- Uppgifterna enligt KN-nummer ex 1904 skall ersättas med följande:
%gt%Plats för tabell%gt%
- Uppgifterna enligt KN-nummer 1905 90 50 skall ersättas med följande:
%gt%Plats för tabell%gt%
- Uppgifterna enligt KN-nummer ex 2008 92 och ex 2008 99 skall utgå.
- Uppgifterna enligt KN-nummer ex 2101 10 och ex 2101 20 skall ersättas med följande:
%gt%Plats för tabell%gt%
- Uppgifterna enligt KN-nummer ex 2106 skall ersättas med följande:
%gt%Plats för tabell%gt%
- Uppgifterna enligt KN-nummer 2208 skall ersättas med följande:
%gt%Plats för tabell%gt%
- Följande uppgifter enligt KN-nummer 3302 skall införas före KN-nummer 3501:
%gt%Plats för tabell%gt%
- Uppgifterna enligt KN-nummer ex 3502 skall ersättas med följande:
%gt%Plats för tabell%gt%
Artikel 2
I artiklarna 2 och 3 i förordning (EEG) nr 2730/75 skall - KN-nummer %quot%1702 10 10%quot% ersättas med KN-nummer %quot%1702 11 00%quot%,
- KN-nummer %quot%1702 10 90%quot% ersättas med KN-nummer %quot%1702 19 00%quot%.
Artikel 3
I bilaga II till förordning (EEG) nr 776/78 skall uppgifterna enligt KN-nummer 0405 ersättas med följande:
%gt%Plats för tabell%gt%
Artikel 4
Förordning (EEG) nr 570/88 ändras på följande sätt:
- I artikel 4.2 b skall KN-nummer %quot%2106 90 99%quot% ersättas med KN-nummer %quot%2106 90 98%quot%.
- I artikel 4.4 skall
- i första strecksatsen KN-nummer %quot%1902 20 90%quot% ersättas med KN-nummer %quot%1902 20 99%quot%,
- i andra strecksatsen KN-nummer %quot%2104 10 00%quot% ersättas med KN-nummer %quot%2104 10%quot%.
Artikel 5
I bilagorna I A (Polen), I B.1 (Tjeckien) och I B.2 (Slovakien) till förordning (EEG) nr 584/92 skall KN-nummer %quot%0405 00 11 och 0405 00 19%quot% ersättas med KN-nummer %quot%0405 10 11 respektive 0405 10 19%quot%.
Artikel 6
I bilaga I till förordning (EEG) nr 2219/92 och i bilaga IV till förordning (EG) nr 2883/94 skall uppgifterna enligt KN-nummer 0405 ersättas med följande:
%gt%Plats för tabell%gt%
Artikel 7
I artikel 8.3 i förordning (EG) nr 1466/95 skall KN-nummer %quot%0405 00 90 och 0405 00 19%quot% ersättas med KN-nummer %quot%0405 10 90, 0405 90 10, 0405 90 90 och 0405 10 19%quot%.
Artikel 8
I bilagan till förordning (EG) nr 1598/95 skall uppgifterna enligt KN-nummer 0403 10, 0404 90 och 0405 ersättas med de uppgifter enligt KN-nummer 0403 10, 0404 90 och 0405 som anges i bilaga I till den här förordningen.
Artikel 9
Förordning (EG) nr 1600/95 ändras på följande sätt:
- I bilaga I, punkt 28, skall KN-nummer %quot%ex 0405 00 11 och ex 0405 00 19%quot% ersättas med KN-nummer %quot%ex 0405 10 11 och ex 0405 10 19%quot%.
- I bilaga IV, punkt 1, skall KN-nummer %quot%ex 0404 90 53 och ex 0404 90 93%quot% ersättas med KN-nummer %quot%0404 90 83%quot%.
- I bilaga VI, led A, skall KN-nummer %quot%ex 0404 90 53 och ex 0404 90 93%quot% ersättas med KN-nummer %quot%0404 90 83%quot%.
- I bilaga VII skall
- i det avsnitt som avser Nya Zeeland KN-nummer %quot%0405 00 11 och 0405 00 19%quot% ersättas med KN-nummer %quot%0405 10 11 respektive 0405 10 19%quot%,
- i det avsnitt som avser Schweiz KN-nummer %quot%ex 0404 90 53 och ex 0404 90 93%quot% ersättas med KN-nummer %quot%0404 90 83%quot%,
- I översiktstabellen skall
- uppgifterna enligt KN-nummer %quot%0403 10-0403 10 36%quot% ersättas ned de uppgifter enligt KN-nummer %quot%0403 10-0403 10 39%quot% som anges i bilaga II till den här förordningen,
- uppgifterna enligt KN-nummer %quot%0404 90-0405 00 90%quot% ersättas med de uppgifter enligt KN-nummer %quot%0404 90-0405 90 90%quot% som anges i bilaga II till den här förordningen,
- uppgifterna enligt KN-nummer %quot%1702 10%quot% ersättas med de uppgifter enligt KN-nummer %quot%1702 11 00-1702 19 00%quot% som anges i bilaga II till den här förordningen.
Artikel 10
I bilaga I led A, B och C i förordning (EG) nr 1713/95 skall KN-nummer %quot%0405 00 11 och 0405 00 19%quot% ersättas med KN-nummer %quot%0405 10 11 respektive 0405 10 19%quot%.
Artikel 11
Denna förordning träder i kraft den 1 januari 1996.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS BESLUT av den 6 februari 1996 om utsläppande på marknaden av en produkt bestående av en genetiskt modifierad organism, en herbicidtolerant hybridsort av raps (Brassica napus L. oleifera Metzg. MS1Bn × RF1Bn) enligt rådets direktiv 90/220/EEG (Text av betydelse för EES) (96/158/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 90/220/EEG av den 23 april 1990 om avsiktlig utsättning av genetiskt modifierade organismer i miljön (1), senast ändrat genom kommissionens direktiv 94/15/EG (2), särskilt artikel 13 i detta, och
med beaktande av följande: I direktiv 90/220/EEG, artikel 10-18, fastställs ett gemenskapsförfarande som bemyndigar en medlemsstats behöriga myndighet att medge utsläppande på marknaden av levande produkter som består av genetiskt modifierade organismer.
En anmälan om utsläppande på marknaden av en sådan produkt (en herbicidtolerant hybridsort av raps saluförd som utsäde) har inlämnats till den behöriga myndigheten i Förenade kungariket för produktion av utsäde men inte för saluföring som livsmedel eller foder.
Förenade kungarikets behöriga myndighet har överlämnat handlingarna i ärendet till kommissionen med tillstyrkan.
Kommissionen har sänt handlingarna till de behöriga myndigheterna i alla medlemsstater. De behöriga myndigheterna i andra medlemsstater har rest invändningar mot handlingarna.
Invändningarna berör
- bedömningen av produktens inverkan på bruket av herbicider och osäkerheten rörande tänkbara långsiktiga miljökonsekvenser,
- bedömningen av toxikologiska hälsoeffekter av produkten om den kommer att användas som livsmedel eller foder, och
- märkningen av produkten.
Enligt artikel 13.3 skall kommissionen därför besluta enligt förfarandet i artikel 21 i direktiv 90/220/EEG.
Tillstånd för användning av herbicider i miljön är underkastade annan gemenskapslagstiftning, särskilt rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande på marknaden av växtskyddsprodukter (3), senast ändrat genom kommissionens direktiv 94/43/EG (4). Tillämpningsområdet för direktiv 90/220/EEG omfattar därför inte frågor rörande tillstånd för herbicider.
I den anmälan som inlämnats enligt direktiv 90/220/EEG gjordes en bedömning av risken för människors hälsa och för miljön av den herbicidtoleranta rapsens överlevnad och spridning samt av ett överförande av den herbicidtoleranta genen eller andra modifierande gener till mottagliga arter. Det konstaterades att risken för etablering var ringa och att spridning eller överförande av den herbicidtoleranta genen kunde kontrolleras genom tillämpning av existerande hanteringsmetoder.
Efter att ha granskat de handlingar som inlämnats enligt direktiv 90/220/EEG och beaktat all den information som överlämnats av medlemsstaterna har kommissionen funnit att den information om miljörisker som finns i handlingarna är tillfyllest för att kommissionen skall kunna fatta ett positivt beslut om utsläppande på marknaden av nämnda produkt som utsäde, förutsatt att föreskrivna villkor för användning och märkning följs.
Artiklarna 11.6 och 16.1 i direktivet 90/220/EEG ger ytterligare stöd om ny kunskap blir tillgänglig om risker förknippade med produkten.
Detta besluts föreskrifter är förenliga med yttrandet från den kommitté som inrättats enligt artikel 21 i direktiv 90/220/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Under de villkor som fastställs i rådets direktiv 69/208/EEG (5) samt de villkor som anges i stycke 2, skall Förenade kungarikets behöriga myndighet lämna medgivande enligt artikel 13 i direktiv 90/220/EEG till utsläppande på marknaden av följande produkt, anmäld av Plant Genetic Systems (ref. C/UK/94/M1/1).
Produkten omfattar levande frön av en hybridsort av raps (Brassica napus L. oleifera Metzg.) med användande av:
a) Avkomman av den hansterila rapslinjen MS1Bn (B91-4) av sorten Drakkar innehållande barnase-genen från Bacillus amyloliquefaciens som kodar för ribonunkleas, bar-genen från Streptomyces hygroscopicus som kodar för fosfinotricinacetyltransferas, neo-genen från Escherichia coli som kodar för neomycinfosfotransferas II, promotorn PSsuAra från Arabidopsis thaliana, promotorn PNos från Agrobacterium tumefaciens, promotorn PTA29 från Nicotiana tabacum, och
b) avkomman av den fertilitetsåterställande rapslinjen RF1Bn (B93-101) av sorten Drakkar innehållande barstar-genen från Bacillus amyloliquefaciens som kodar för ribonukleasinhibitor, bar-genen från Streptomyces hygroscopicus som kodar för fosfinotricinacetyltransferas, neo-genen från Escherichia coli som kodar för neomycinfosfotransferas II, promotorn PSsuAra från Arabidopsis thaliana, promotorn PNos från Agrobacterium tumefaciens, promotorn PTA29 från Nicotiana tabacum.
2. Följande villkor gäller för medgivandet:
a) Medgivandet avser utsäde av alla hybrider mellan icke genetiskt modifierad raps och den genetiskt modifierade raps som beskrivs i punkt 1 men omfattar inte utsäde av hybrider som kan uppkomma genom korsning mellan andra genetiskt modifierade växter än de som beskrivs i punkt 1.
b) Medgivandet avser endast användning av produkten för fröproduktion enligt anmälan och inte användning som livsmedel eller foder, utan att detta påverkar en eventuell framtida bedömning av produkten för sådan användning.
c) Utöver annan märkning skall det anges på etiketten till varje utsädesförpackning att produkten är tolerant mot herbicidenglufosinatammonium och att den endast får användas för produktion av frö och inte som livsmedel eller foder.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
RÅDETS BESLUT av den 4 mars 1996 om ett varnings- och beredskapsförfarande för ansvarsfördelning vid mottagande av och tillfällig vistelse för fördrivna personer (96/198/RIF)
EUROPEISKA UNIONENS RÅD HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om Europeiska unionen, särskilt artikel K.3.2 a i detta,
med beaktande av rådets resolution av den 25 september 1995 om ansvarsfördelning vid mottagande av fördrivna personer och tillfälligt uppehälle för fördrivna personer (1) och
med beaktande av följande: Den ovannämnda resolutionen bör kompletteras för att göra det möjligt att effektivt tillämpa dess principer i krissituationer som kräver snabba åtgärder.
Ett varnings- och beredskapsförfarande bör fastställas i detta syfte.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
1. Igångsättning av förfarandet
På initiativ av ordförandeskapet, en medlemsstat eller kommissionen kan den samordningskommitté som avses i artikel K.4 i fördraget genast sammankallas, sedan dess medlemmar rådgivits av medlemsstaternas asyl- och invandringsansvariga, för att konstatera om situationen är sådan att det krävs ett samordnat handlande från Europeiska unionens för mottagande av och tillfällig vistelse för fördrivna personer.
Ett handlande av sådant slag kan endast planeras om de villkor som anges i punkterna 1 och 2 i rådets resolution av den 25 september 1995 är uppfyllda.
Ordförandeskapet skall regelmässigt och i alla händelser före mötet utarbeta en lägesrapport i samarbete med kommissionen, mot bakgrund av FN:s flyktingkommissaries yttrande och med bistånd av rådets generalsekretariat. Denna rapport skall överlämnas till medlemsstaterna.
2. Dagordning för mötet
Dagordningen för mötet kan omfatta särskilt följande punkter:
- undersökning av situationen och bedömning av folkförflyttningarnas omfattning,
- bedömning av det lämpliga i ett brådskande ingripande på Europeiska unionens nivå,
- undersökning av andra möjligheter, inklusive eventuella åtgärder på plats,
- upprättande av en tidsplan och planläggning i flera steg för det beräknade mottagningsbehovet,
- angivande av varje medlemsstat om hur många personer den kan ta emot och när den kan ta emot dem, på grundval av punkt 4 i rådets resolution av den 25 september 1995,
- samordning med kommissionens åtgärder inom området för humanitär hjälp,
- informationsutbyte med Förenta nationernas flyktingkommissarie och samordning av planen för mottagandet,
- samordning med tredje länder.
3. Beslut om ansvarsfördelning
Ett förslag efter resultatet av arbetet från den ovannämnda samordningskommitténs möte skall utarbetas och förläggas rådet för godkännande.
Om det bedöms som nödvändigt, kan de föreskrifter som anges i rådets arbetsordning för nödsituationer tillämpas, i enlighet med punkt 3 i rådets resolution av den 25 september 1995 och om en månad förflyter utan att samordningskommittén når fram till en överenskommelse.
4. Uppföljning av situationen
Formerna för mottagandet av de fördrivna personerna skall fastställas av varje medlemsstat.
Så länge som krissituationen består, kan den ovannämnda samordningskommittén mötas ofta, med mellanrum som den själv bestämmer och enligt villkoren i punkt 2.
RÅDETS BESLUT av den 11 juni 1996 om tillämpning av artikel 8 i avtalet genom skriftväxling mellan Europeiska ekonomiska gemenskapen och Furstendömet Andorra (96/366/EG)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 113 i detta,
med beaktande av kommissionens förslag, och
med beaktande av följande: I artikel 8.1 a i avtalet genom skriftväxling mellan Europeiska ekonomiska gemenskapen och Furstendömet Andorra (1), som undertecknades i Luxemburg den 28 juni 1990, föreskrivs att Furstendömet Andorra bemyndigar gemenskapen att för Furstendömet Andorras räkning under en tid av fem år, eller därutöver om någon överenskommelse inte går att nå enligt b, låta produkter med ursprung i tredje land och avsedda för Furstendömet Andorra övergå till fri omsättning.
I 1 b i samma artikel föreskrivs att Furstendömet Andorra vid utgången av denna tid och inom ramen för artikel 20 i avtalet, kan förbehålla sig att utöva sin rätt att låta dessa varor övergå till fri omsättning efter det att de avtalsslutande parterna slutit avtal därom.
Furstendömet Andorra har begärt att få utöva denna rätt till övergång till fri omsättning.
Rådet markerade i en förklaring som antogs den 30 oktober 1995 sitt principiella godkännande till att Furstendömet Andorra utöver denna rätt.
Det är lämpligt att rådet som avtalsslutande part formellt fastställer gemenskapens ståndpunkt.
Det är lämpligt att fastställa en frist för att genomförandet av rätten till övergång till fri omsättning skall kunna förberedas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Enda artikel
Från och med den 1 juli 1996 upphör Europeiska gemenskapen att på Furstendömet Andorras vägnar och för dess räkning låta varor med ursprung i tredje land och avsedda för Furstendömet Andorra övergå till fri omsättning.
GEMENSAM ÅTGÄRD av den 4 mars 1996 beslutad av rådet på grundval av artikel K.3 i Fördraget om Europeiska unionen, om ett system för flygplatstransitering (96/197/RIF)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT OM FÖLJANDE GEMENSAMMA ÅTGÄRD
med beaktande av Fördraget om Europeiska unionen, särskilt artikel K.3.2 b,
med beaktande av Frankrikes förslag av den 23 februari 1995, och
med beaktande av följande: Att bestämma villkoren för inresa i och rörlighet inom medlemsstaternas territorium för medborgare i tredje land samt kampen mot olaglig invandring av medborgare från tredje land är en fråga av gemensamt intresse med stöd av artikel K.1.3 a respektive c i fördraget.
Flyget utgör, särskilt när det gäller ansökningar om inresa eller faktisk inresa vid flygplatstransitering, en betydande möjlighet till intrång, särskilt för illegal bosättning inom medlemsstaternas territorium, och det är därför lämpligt att sträva efter att förbättra kontrollen av detta.
I bilaga IX till Chicagokonventionen angående internationell civil luftfart fastläggs principen om fri passage vid transitering via internationella flygplatsområden. Staterna kan trots detta avvika från denna allmänna princip genom att anmäla denna avvikelse till Internationella civila luftfartsorganisationen (ICAO) och genom att kräva innehav av visering för flygplatstransitering. Denna möjlighet bör i görligaste mån begränsas för att undvika att utvecklingen av luftfarten hindras i onödan.
Harmoniseringen av medlemsstaternas politik på detta område svarar mot målen att uppnå säkerhet och kontroll av illegal invandring, samtidigt som den bidrar till att harmonisera konkurrensvillkoren för medlemsstaternas flygbolag och flygplatser.
Denna fråga berör inte de viseringar som krävs vid passage av medlemsstaternas yttre gränser och omfattas således inte av artikel 100c. 1 i Fördraget om upprättandet av Europeiska gemenskapen, men den är trots detta av gemensamt intresse och skulle kunna regleras på ett mer effektivt sätt genom en gemensam åtgärd.
De medlemsstater som inte har några regler för flygplatstransitvisering bör få tillräcklig tid för att införa sådana regler.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I denna gemensamma åtgärd avses med visering för flygplatstransitering ett tillstånd som skall innehas av medborgare i vissa tredje länder, med avvikelse från principen om fri transitering enligt bilaga IX till Chicagokonventionen angående internationell civil luftfart, vid transitering via medlemsstaternas internationella flygplatsområden.
Artikel 2
1. Visering för flygplatstransitering skall utfärdas av medlemsstaternas konsulära myndigheter.
2. Varje medlemsstat bestämmer villkoren för utfärdande av visering för flygplatstransitering, under förutsättning att rådet antar kriterier för handläggning och utfärdande av viseringar.
De konsulära myndigheterna skall i alla händelser kontrollera att det inte finns någon risk för säkerheten eller för illegal invandring. De skall i synnerhet försäkra sig om att ansökningen om visering för flygplatstransitering är berättigad, på grundval av de handlingar som den sökande lämnat in och att dessa handlingar i möjligaste mån garanterar inresa i det slutliga bestämmelselandet, särskilt genom företeende av visering när sådan krävs.
3. Så snart genomförandet av de bestämmelser som anges i rådets förordning (EG) nr 1683/95 av den 29 maj 1995 om en enhetlig utformning av visumhandlingar (1) blivit tillämpliga skall medlemsstaterna utfärda visering för flygplatstransitering med användning av denna enhetliga utformning av viseringshandlingar.
Artikel 3
Varje medlemsstat skall kräva en visering för flygplatstransitering av medborgare i de tredje länder som finns uppräknade i den gemensamma förteckning som bifogas, om de inte redan innehar en inresevisering eller en transitvisering för denna medlemsstat när de passerar via de internationella flygplatsområdena på dess territorium.
Artikel 4
En medlemsstat får föreskriva undantag från skyldigheten att inneha visering för flygplatstransitering när det gäller medborgare i de tredje länder som finns uppräknade i den gemensamma förteckning som bifogas, särskilt för
- besättningsmedlemmar på luftfartyg och fartyg,
- innehavare av diplomatpass: officiella eller tjänstepass,
- innehavare av uppehållstillstånd eller motsvarande handlingar som utfärdats av en medlemsstat,
- innehavare av visering som utfärdats av en medlemsstat eller av en stat som är part i avtalet om Europeiska ekonomiska samarbetsområdet.
Artikel 5
Varje medlemsstat skall själv bestämma om det finns anledning att kräva visering för flygplatstransitering när det gäller medborgare i stater som inte finns nämnda i den gemensamma förteckning som bifogas.
Artikel 6
Varje medlemsstat skall själv bestämma vilket system för flygplatstransitering som skall tillämpas på statslösa och personer med flyktingstatus.
Artikel 7
Inom en tidsfrist av tio arbetsdagar efter den gemensamma åtgärdens ikraftträdande skall varje medlemsstat underrätta övriga medlemsstater och rådets generalsekretariat om de åtgärder som den har vidtagit med tillämpning av artiklarna 4, 5 och 6. Dessa åtgärder skall för kännedom offentliggöras i EGT.
Artikel 8
Varje år skall rådets ordförandeskap utarbeta en lägesrapport om harmoniseringen av systemet för flygplatstransiteringen inom Europeiska unionen.
Rådet skall granska alla förslag till justering av den förteckning över länder som bifogas.
Artikel 9
Denna gemensamma åtgärd skall inte utgöra något hinder för en mer långtgående harmonisering i fråga om flygplatstransitering mellan vissa medlemsstater, en harmonisering med en räckvidd utöver den i den gemensamma förteckning som bifogas.
Artikel 10
Denna gemensamma åtgärd träder i kraft den första dagen i den sjätte månaden efter det att den har offentliggjorts i EGT.
För Danmark, Finland och Sverige träder den emellertid i kraft den första dagen i den artonde månaden efter det att den har offentliggjorts i EGT.
RÅDETS DIREKTIV 96/49/EG av den 23 juli 1996 om tillnärmning av medlemsstaternas lagstiftning om transport av farligt gods på järnväg
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 75 i detta,
med beaktande av kommissionens förslag (1),
med beaktande av Ekonomiska och sociala kommitténs yttrande (2),
i enlighet med det i artikel 189c i fördraget angivna förfarandet (3), och
med beaktande av följande: 1. Omfattningen av transporter av farligt gods på järnväg har under senare år ökat kraftigt och därmed har olycksrisken ökat. Åtgärder bör följaktligen vidtas för att denna typ av transporter skall kunna utföras under sådana betingelser som ger största möjliga säkerhet.
2. Alla medlemsstater är fördragsslutande parter i Fördraget om internationell järnvägstrafik (COTIF), som i sitt bihang B fastställer enhetliga regler för avtalet om internationell järnvägsbefordran av gods (CIM), vars bilaga I utgör reglementet om internationell järnvägsbefordran av farligt gods (RID). Fördragets geografiska tillämpningsområde sträcker sig utanför gemenskapen.
3. Det fördraget omfattar inte nationell transport av farligt gods på järnväg. Följaktligen är det viktigt att säkerställa en enhetlig tillämpning av harmoniserade säkerhetsbestämmelser i hela gemenskapen. Det lämpligaste sättet att nå detta mål är att anpassa medlemsstaternas lagstiftningar till RID.
4. Med iakttagande av subsidiaritetsprincipen bör denna tillnärmning av lagstiftningarna ske för att kunna säkerställa en hög säkerhetsnivå hos nationella och internationella transporter, för att garantera att snedvridna konkurrensförhållanden undanröjs och för att underlätta den fria rörligheten för varor och tjänster i hela gemenskapen, samt för att säkerställa enhetlighet med annan gemenskapslagstiftning.
5. Bestämmelserna i detta direktiv påverkar inte gemenskapen och dess medlemsstaters åtagande att i framtiden i englighet med de mål som anges i kapitel 19 i Agenda 21 från UNCED-konferensen i Rio de Janeiro i juni 1992 harmonisera systemen för klassificering av farliga ämnen.
6. Det finns ännu inte någon särskild gemenskapslagstiftning som reglerar de säkerhetsmässiga förhållandena för transport av biologiska agens och genetiskt modifierade mikroorganismer, som omfattas av rådets direktiv 90/219/EEG (4), 90/220/EEG (5) och 90/679/EEG (6).
7. Bestämmelserna i detta direktiv är tillämpliga utan att de påverkar tillämpningen av andra gemenskapsbestämmelser om arbetstagarnas säkerhet och miljöskydd.
8. Medlemsstaterna måste på sina territorier kunna tillämpa särskilda regler för rörligheten avseende transport av farligt gods på järnväg.
9. Medlemsstaterna bör vad gäller nationella transporter av farligt gods på järnväg behålla rätten att provisoriskt tillämpa regler som överensstämmer med Förenta nationernas multimodala rekommendationer för transport av farligt gods i den utsträckning som RID ännu inte har harmoniserats med dessa regler, vilka bör underlätta intermodal transport av farligt gods.
10. Varje medlemsstat bör, enbart av andra skäl än säkerhetsmässiga, behålla rätten att reglera och förbjuda nationell transport av visst farligt gods på järnväg.
11. Hänsyn bör tas till de strängare säkerhetsåtgärder som tillämpas i tunneln under Engelska kanalen på grund av dennas särskilda egenskaper, framför allt dess sträckning och längd, och medlemsstaterna bör ges möjlighet att införa samma slags åtgärder när liknande situationer uppstår. Vissa medlemsstater bör kunna tillämpa strängare regler för gods som skall transporteras på grund av temperaturen i godsets omgivning.
12. För att kunna beakta vikten av nödvändiga investeringar på detta område bör en övergångsperiod fastställas, så att medlemsstaterna tillfälligt kan upprätthålla vissa särskilda nationella bestämmelser om konstruktions- eller användningskrav för tankar, behållare, förpackningar, eller nödåtgärdskod.
13. Utnyttjandet av den nya tekniska och industriella utvecklingen får inte hämmas och bestämmelser om tillfälliga undantag bör därför införas.
14. RID-bestämmelserna tillåter bestämmelser om avvikelser härifrån och det stora antalet avtal som har ingåtts bilateralt mellan medlemsstaterna hindrar det fria tillhandahållandet av tjänster för transport av farligt gods. Införandet av de nödvändiga bestämmelserna i bilagan till detta direktiv bör göra det möjligt att undvika sådana avvikelser. Det är viktigt att medlemsstaterna under en övergångsperiod kan fortsätta att tillämpa befintliga avtal mellan sig.
15. Järnvägstransporter av farligt gods till eller från tredje land är tillåtna i den mån som de utförs i enlighet med RID-bestämmelserna. Vad gäller transporter från eller till republikerna i det forna Sovjetunionen, som inte är fördragsslutande parter i COTIF, bör medlemsstaterna emellertid införa lämpliga bestämmelser om dessa transporter för att säkerställa att säkerhetsnivån motsvarar den som fastlagts i RID.
16. Detta direktiv bör snabbt kunna anpassas till den tekniska utvecklingen, särskilt genom antagande av de nya bestämmelser om vilka beslut fattas inom ramen för RID. En kommitté bör därför upprättas och ett förfarande införas som innebär ett nära samarbete mellan medlemsstaterna och kommissionen inom denna kommitté.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
KAPITEL I Tillämpningsområde
Artikel 1
1. Detta direktiv skall tillämpas på transport av farligt gods med järnväg inom eller mellan medlemsstaterna. Medlemsstaterna får dock från tillämpningsområdet undanta transport av farligt gods som genomförs med hjälp av transportmedel som tillhör de väpnade styrkorna eller för vilka dessa är ansvariga.
2. Bestämmelserna i detta direktiv skall inte påverka medlemsstaternas rätt att, med iakttagande av gemenskapsrätten, ställa särskilda säkerhetskrav för nationell eller internationell transport av farligt gods på järnväg, i den mån bilagan till det här direktivet inte täcker detta område, särskilt såvitt avser
- tågtrafik,
- utanordning av godsvagnar i tåg i nationell trafik,
- driftsbestämmelser i samband med transportrelaterade operationer som till exempel rangering och parkering,
- personalutbildning och administration av information beträffande farligt gods som transporteras,
- särskilda regler för transport av farligt gods med passagerartåg.
Artikel 2
I detta direktiv avses med
- RID: reglementet om internationell järnvägsbefordran av farligt gods, som finns i bilaga I till bihang B till Fördraget om internationell järnvägstrafik (COTIF), inklusive ändringar,
- CIM: de enhetliga rättsreglerna för avtal om internationell järnvägsbefordran av gods, som finns i bihang B till Fördraget om internationell järnvägstrafik (COTIF), med ändringar,
- farligt gods: de ämnen och föremål som inte får transporteras på järnväg eller som endast får transporteras på särskilda villkor i enlighet med bilagan till detta direktiv,
- transport: sådan järnvägstransport av farligt gods som helt eller delvis utförs inom en medlemsstats territorium, inbegripet såväl lastning och lossning av gods som omlastning till eller från ett annat transportslag samt stopp, som är nödvändiga på grund av betingelserna för transporten, och som omfattas av bilagan till detta direktiv, utan att det påverkar medlemsstaternas bestämmelser om ansvar som är en följd av sådana operationer. Transporter som endast sker inom ett företags område skall inte omfattas av denna definition.
Artikel 3
1. Utan att det påverkar tillämpningen av artikel 6, får farligt gods som är förbjudet att transportera enligt bestämmelserna i bilagan inte transporteras på järnväg.
2. Om inte annat föreskrivs i detta direktiv, och utan att det påverkar tillämpningen av bestämmelserna om järnvägsföretagens tillträde till marknaden eller bestämmelser som på ett allmänt sätt är tillämpliga på transport av gods på järnväg, är transport på järnväg av annat farligt gods tillåtet, om den är förenlig med bestämmelserna i bilagan.
KAPITEL II Avvikelser, begränsningar och undantag
Artikel 4
I fråga om nationella transporter på järnväg, kan en medlemsstat upprätthålla de bestämmelser i sin nationella lagstiftning om transport av farligt gods på järnväg som är förenliga med Förenta nationernas rekommendationer om transport av farligt gods, tills bilagan till detta direktiv har revideras så att den överensstämmer med dessa rekommendationer. I detta fall skall den berörda medlemsstaten underrätta kommissionen om detta.
Artikel 5
1. Utan att det påverkar tillämpningen av andra gemenskapsbestämmelser, skall medlemsstaterna endast av andra skäl än transportsäkerhetsmässiga, som har samband med den nationella säkerheten eller skyddet av miljön, behålla rätten att reglera eller förbjuda transport av visst farligt gods inom sitt territorium.
2. a) Beträffande transport genom tunneln under Engelska kanalen kan Frankrike och Förenade kungariket införa strängare bestämmelser än de som anges i bilagan. Kommissionen skall få meddelande om dessa bestämmelser och meddela de övriga medlemsstaterna om detta.
b) Om en medlemsstat bedömer att dessa strängare bestämmelser bör tillämpas på transport inom dess territorium genom tunnlar med liknande egenskaper som de som avses i punkt 1, skall den underrätta kommissionen om detta. Denna skall i enlighet med förfarandet i artikel 9 besluta om den ifrågavarande tunneln har liknande egenskaper. De bestämmelser som en medlemsstat antar skall meddelas kommissionen, som skall underrätta de övriga medlemsstaterna om detta.
c) De medlemsstater vilkas omgivningstemperatur regelbundet är lägre än -20° C får, tills bestämmelser om lämpliga referenstemperaturer för vissa bestämda klimatzoner införs i bilagan, införa strängare bestämmelser med avseende på ett materials möjlighet att fungera vid vissa temperaturer för användning vid nationell transport av farligt gods.
3. Om en medlemsstat till följd av en olyckshändelse eller en incident finner att säkerhetsbestämmelserna kan förbättras så att de risker som är förbundna med transporten minskas och att åtgärder måste vidtas omedelbart, skall den på planeringsstadiet underrätta kommissionen om de åtgärder den avser att vidta. Kommissionen skall i enlighet med förfarandet i artikel 9 besluta huruvida ett genomförande av dessa åtgärder kan tillåtas och bestämma hur länge de skall tillämpas.
4. Medlemsstaterna kan upprätthålla de nationella bestämmelser som den 31 december 1996 gäller för transport och förpackning av ämnen som innehåller dioxiner eller furaner.
Artikel 6
1. I de fall där transporten innefattar ett sjö- eller luftavsnitt får medlemsstaterna tillåta järnvägstransport på sina territorier av farligt gods som är klassificerat, förpackat och märkt i överensstämmelse med internationella krav för sjö- eller lufttransport.
Om det ingår ett sjöavsnitt i en nationell eller internationell transport, får medlemsstaterna för att ta hänsyn till internationella regler om sjötransport, däribland internationella regler om färjetransport, tillämpa bestämmelser som kompletterar bestämmelserna i bilagan.
2. Bestämmelserna i bilagan om användning av transportdokument och om vilka språk som skall användas vid märkningen eller i transportdokumenten skall inte gälla för transport som är begränsad till en enda medlemsstats territorium. Medlemsstaterna får tillåta att andra dokument och språk än de som anges i bilagan används för transporter som är begränsade till deras eget territorium.
3. En medlemsstat får på sitt territorium tillåta användning av järnvägsvagnar som är tillverkade före den 1 januari 1997 och som inte är i enlighet med detta direktiv men vilkas konstruktion följer de bestämmelser i den nationella lagstiftningen som är i kraft den 31 december 1996, under förutsättning att dessa vagnar uppfyller säkerhetskraven.
4. En medlemsstat får upprätthålla de nationella bestämmelser om tillverkning, användning och transportvillkor för nya tankar och nya behållare som motsvarar klass 2 i bilagan, som är i kraft den 31 december 1996 och som avviker från bestämmelserna i bilagan tills hänvisningar till normer för konstruktion och användning av sådana tankar och behållare införs i bilagan med samma bindande verkan som de bestämmelser den innehåller, dock längst till och med den 31 december 1998. Behållare och tankar som tillverkats före den 1 januari 1999 och som uppfyller säkerhetskraven, får även i fortsättningen användas på de ursprungliga villkoren.
5. En medlemsstat får upprätthålla andra nationella bestämmelser än de som finns i bilagan i fråga om referenstemperaturen vid transport inom sitt territorium av flytande gaser eller av blandningar av flytande gaser, tills bestämmelser om lämpliga referenstemperatur för bestämda klimatzoner har införlivats med europeiska standarder och hänvisning till dessa standarder har gjorts i bilagan.
6. Varje medlemsstat får vid transport inom sitt territorium tillåta användning av förpackningar som är tillverkade före den 1 januari 1997 men som inte är godkända i överensstämmelse med RID, förutsatt att förpackningen är märkt med tillverkningsdagen, kan klara de relevanta provningarna i enlighet med kraven i de nationella bestämmelser som gäller den 31 december 1996, och uppfyller säkerhetskraven (vilket i förekommande fall innebär provningar och kontroller), enligt följande ordning: stora metallbehållare för bulkvaror samt metallfat med en kapacitet på mer än 50 liter får användas under en tidsperiod på högst 15 år från och med tillverkningsdagen. Andra metallförpackningar och alla plastförpackningar får användas under en tidsperiod på högst fem år från och med tillverkningsdagen, dock inte efter den 31 december 1998.
7. En medlemsstat får till och med den 31 december 1998 tillåta transport på sitt territorium av visst farligt gods som förpackats före den 1 januari 1997, förutsatt att godset är klassificerat, förpackat och märkt i enlighet med kraven i de nationella bestämmelser som gällde före den 1 januari 1997.
8. Varje medlemsstat får för nationella transporter på järnväg inom sitt territorium upprätthålla de bestämmelser i sin lagstiftning som gäller den 31 december 1996 för märkning med en nödåtgärdskod i ställe för det faronummer som anges i bilagan.
9. Varje medlemsstat får efter samråd med kommissionen upprätthålla mindre stränga bestämmelser än de i bilagan för transport på järnväg på sitt territorium av små mängder av visst farligt gods, med undantag för ämnen som har en hög eller mellanhög grad av radioaktivitet.
10. En medlemsstat får på sitt territorium tillåta enstaka transporter av farligt gods eller transporter som är förbjudna enligt bestämmelserna i bilagan eller som utförs på andra villkor än de som anges i bilagan.
11. Med iakttagande av gemenskapslagstiftningen påverkar detta direktiv inte medlemsstaternas rätt att, efter samråd med kommissionen och på vederbörligen angivna sträckor inom sina territorier tillåta regelbundna transporter av farligt gods, som utgör en del av en angiven industriell process som antingen kan vara förbjuden enligt bestämmelserna i bilagan eller utföras på andra villkor än de som anges i bilagan, när dessa operationer är av lokal karaktär och är underkastade sträng kontroll på klart angivna villkor.
12. Medlemsstaterna får medge tillfälliga undantag från bilagan för att på sina territorier utföra de provningar som är nödvändiga för ändringar av dessa bestämmelser för att anpassa dem till den tekniska och industriella utvecklingen, förutsatt att säkerheten inte åsidosätts. Kommissionen skall underrättas om detta och skall i sin tur underrätta de andra medlemsstaterna.
Tillfälliga undantag som medlemsstaternas behöriga myndigheter kommer överens om på grundval av bilagan, skall ges formen av ett multilateralt avtal som den myndighet som tar initiativ till avtalet föreslår samtliga medlemsstaters behöriga myndigheter att ingå. Kommissionen skall underrättas om detta.
De undantag som avses i första och andra styckena skall medges utan diskriminering på grund av avsändarens, operatörens eller mottagarens nationalitet eller etableringsort. De skall gälla under en tid av högst fem år och kan inte förlängas.
13. En medlemsstat får längst till och med den 31 december 1998 tillämpa avtal som har ingåtts med andra medlemsstater utan diskriminering på grund av avsändarens, operatörens eller mottagarens nationalitet eller etableringsort. Alla framtida undantag skall vara i överensstämmelse med punkt 12.
14. Med iakttagande av gemenskapslagstiftningen skall detta direktiv inte påverka medlemsstaternas rätt att efter samråd med kommissionen tillåta transporter av farligt gods under mindre stränga villkor än de som anges i bilagan när det gäller lokala transporter på korta sträckor och som är begränsade till hamnområden, flygplatser eller industriområden.
Artikel 7
1. Med förbehåll för nationella bestämmelser eller gemenskapsbestämmelser om tillträde till marknaden, kan järnvägstransport av farligt gods mellan gemenskapens territorium och tredje länders territorium tillåtas i den utsträckning som transporten sker i enlighet med RID bestämmelserna.
2. Det här direktivet påverkar inte medlemsstaternas rätt att på sina territorier och efter underrättelse till kommissionen införa bestämmelser om transport på järnväg av farligt gods, som sker från eller till republiker i det forna Sovjetunionen som inte är fördragsslutande parter till COTIF. Dessa bestämmelser gäller bara transport på järnväg av farligt gods (som kolli, bulklast eller i tankar) med järnvägsvagner som godkänts av en stat som inte är fördragsslutande part i COTIF. Genom lämpliga åtgärder och förpliktelser skall de berörda medlemsstaterna säkerställa att säkerhetsnivån motsvarar den som föreskrivs i RID-bestämmelserna. För vissa medlemsstater gäller bestämmelserna i detta stycke endast cisternvagnar.
KAPITEL III Slutbestämmelser
Artikel 8
De ändringar som är nödvändiga för att anpassa bilagan till den vetenskapliga och tekniska utvecklingen på de områden som omfattas av detta direktiv och som syftar till att anpassa dem till de nya RID-bestämmelserna skall antas enligt det förfarande som anges i artikel 9.
Artikel 9
1. Kommissionen skall biträdas av kommittén för transport av farligt gods, som inrättas genom artikel 9 i direktiv 94/55/EG (7), nedan kallad kommittén, som består av företrädare för medlemsstaterna och har en företrädare för kommissionen som ordförande.
2. Kommissionens företrädare skall förelägga kommittén ett förslag till åtgärder. Kommittén skall yttra sig över förslaget inom den tid som ordföranden bestämmer med hänsyn till hur brådskande frågan är. Yttrandet skall avges med den majoritet som enligt artikel 148.2 i fördraget skall tillämpas vid beslut som rådet skall fatta på förslag av kommissionen. Vid röstning i kommittén skall de röster som avges av medlemsstaterna vägas enligt samma artikel. Ordföranden får inte rösta.
3. a) Kommissionen skall anta de föreslagna åtgärderna när dessa är förenliga med kommitténs yttrande.
b) Om de föreslagna åtgärderna inte är förenliga med kommitténs yttrande eller om inget yttrande avges, skall kommissionen utan dröjsmål föreslå rådet vilka åtgärder som skall vidtas. Rådet skall fatta sitt beslut med kvalificerad majoritet.
Om rådet inte har fattat något beslut inom tre månader från det att förslaget mottagits, skall kommissionen själv besluta att de föreslagna åtgärderna skall vidtas.
Artikel 10
1. Medlemsstaterna skall före den 1 januari 1997 sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser, skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 11
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
Artikel 12
Detta direktiv riktar sig till medlemsstaterna.
KOMMISSIONENS FÖRORDNING (EG) nr 216/96 av den 5 februari 1996 om processordningen för överklagningsnämnderna vid Byrån för harmonisering inom den inre marknaden (varumärken och mönster)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 40/94 av den 20 december 1993 om gemenskapsvarumärken (1), ändrad genom förordning (EG) nr 3288/94 (2), särskilt artikel 140.3 i denna, och
med beaktande av följande: Genom förordning (EG) nr 40/94 (nedan kallas %quot%förordningen%quot%) införs ett nytt varumärkessystem som gör det möjligt att, på grundval av en ansökan till Byrån för harmonisering inom den inre marknaden (varumärken och mönster) (nedan kallad %quot%byrån%quot%), förvärva ett varumärke med rättsverkan inom hela gemenskapen.
I detta syfte innehåller förordningen framförallt de nödvändiga bestämmelserna avseende förfarandet vid registrering av ett gemenskapsvarumärke, administrationen av gemenskapsvarumärken, överklaganden av byråns beslut och förfarandet för att upphäva eller ogiltigförklara ett gemenskapsvarumärke.
Enligt artikel 130 i förordningen ankommer det på överklagningsnämnderna att besluta om överklaganden av beslut av granskarna, invändningsavdelningarna, avdelningen för varumärkesrätt och övriga juridiska frågor och annulleringsavdelningarna.
Avdelning VII i förordningen innehåller grundprinciper för överklaganden av beslut av granskare, invändningsavdelningarna, avdelningen för varumärkesrätt och övriga juridiska frågor och annuleringsavdelningarna.
Avdelning X i kommissionens förordning (EG) nr 2868/95 av den 13 december 1995 om genomförande av rådets förordning (EG) nr 40/94 om gemenskapsvarumärke (3) innehåller genomförandebestämmelser till avdelning VII i förordningen.
Den här förordningen kompletterar de övriga bestämmelserna, framförallt dem som gäller nämndernas organisation och muntliga förhandlingar.
Före varje verksamhetsår bör en plan för fördelning av ärenden mellan överklagningsnämnderna fastställas av ett organ som inrättats i detta syfte. Nämnda organ bör tillämpa objektiva kriterier, såsom varu- och tjänsteklasser eller begynnelsebokstäverna i de sökandes namn.
För att underlätta handläggningen och expedieringen av överklaganden bör för varje ärende en referent utses som skall vara ansvarig bl.a. för att förbereda meddelanden till parterna och utarbeta förslag till beslut.
Parterna inför överklagningsnämnderna har kanske inte förutsättningarna eller viljan att göra överklagningsnämnderna uppmärksamma på frågor av allmänt intresse för ett pågående ärende. Överklagningsnämnderna bör därför ha befogenhet att, på eget initiativ eller på begäran av byråns direktör, ge direktören tillfälle att framföra synpunkter på frågor av allmänt intresse som rör pågående ärenden vid överklagningsnämnderna.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från den kommitté som inrättats enligt artikel 141 i förordningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Fördelning av arbetsuppgifter samt det organ som är behörigt att göra denna fördelning
1. Före varje verksamhetsårs början skall ärendena fördelas mellan överklagningsnämnderna i enlighet med objektiva kriterier och ledamöterna i varje nämnd och deras suppleanter skall utses. Varje ledamot i en överklagningsnämnd kan utses som ledamot eller suppleant i flera överklagningsnämnder. Dessa åtgärder kan i förkommande fall ändras under det ifrågavarande verksamhetsåret.
2. De åtgärder som anges i punkt 1 skall vidtas av ett organ bestående av byråns direktör som ordförande, vice direktören för den byrå som är ansvarig för överklagningsnämnderna, ordförandena för överklagningsnämnderna och tre andra ledamöter av överklagningsnämnderna valda av samtliga ledamöter i dessa nämnder, med undantag för ordförandena, för det ifrågavarande verksamhetsåret. För att organet skall vara beslutfört krävs att minst fem av dess ledamöter är närvarande, inklusive byråns direktör eller vice direktör och två ordförande i överklagningsnämnderna. Organets beslut skall fattas med en majoritet av rösterna. Vid lika röstetal skall ordförandens röst vara utslagsgivande. Organet kan själv fastställa sin arbetsordning.
3. Det organ som avses i punkt 2 skall avgöra tvister som rör fördelningen av arbetsuppgifter mellan olika överklagningsnämnder.
4. Fram till dess att fler än tre överklagningsnämnder har inrättats skall det organ som avses i punkt 2 bestå av byråns direktör, som skall fungera som ordförande, byråns vice direktör, som är ansvarig för överklagningsnämnderna, ordföranden eller ordförandena i den eller de överklagningsnämnder som redan har inrättats, och en annan ledamot av överklagningsnämnderna, vald av samtliga ledamöter i nämnderna, med undantag av ordföranden eller ordförandena, för verksamhetsåret i fråga. För att organet skall vara beslutfört krävs att minst tre av dess ledamöter är närvarande, inklusive byråns direktör eller vice direktör.
Artikel 2
Ersättande av ledamöter
1. En ledamot kan ersättas av en suppleant bl.a. vid ledighet, sjukdom och åtaganden som måste fullgöras samt vid de jävsgrunder som avses i artikel 132 i förordningen.
2. Varje ledamot som begär att ersättas av en suppleant skall genast underrätta ordföranden i den berörda nämnden om sitt förhinder.
Artikel 3
Jäv och jävsanmälan
1. Om en nämnd har kännedom om en möjlig grund för jäv eller jävsanmälan enligt artikel 132.3 i förordningen och denna grund inte har åberopats av ledamoten själv eller av någon av parterna skall förfarandet i artikel 132.4 i förordningen tillämpas.
2. Den berörda ledamoten skall beredas tillfälle att yttra sig om huruvida det finns grund för jäv eller jävsanmälan.
3. Handläggningen skall ställas in till dess att ett beslut om vilka åtgärder som skall vidtas har fattats i enlighet med artikel 132.4 i förordningen.
Artikel 4
Referent
1. Ordföranden i varje nämnd skall för varje överklagande utse en ledamot i sin egen nämnd eller sig själv som referent.
2. Referenten skall genomföra en preliminär undersökning av överklagandet. Han kan avfatta meddelanden till parterna enligt ordförandens instruktioner. Meddelanden skall undertecknas av referenten för nämndens räkning.
3. Referenten skall förbereda nämndens egna sammanträden och de muntliga förhandlingarna.
4. Referenten skall utarbeta förslag till beslut.
Artikel 5
Registratorskontor
1. Registratorskontor skall inrättas för överklagningsnämnderna. Registratorer skall ansvara för alla funktioner på registratorskontoren. En av registratorerna kan utses till förste registrator.
2. Det organ som avses i artikel 1.2 kan anförtro registratorerna uppgifter som inte innefattar några svårigheter av rättslig eller teknisk art i synnerhet vad avser företrädare, inleverering av översättningar, granskning av akter och delgivningar.
3. Registratorn skall till ordföranden i den berörda nämnden för varje nytt överklagande överlämna en redogörelse för huruvida överklagandet kan tas upp till prövning.
4. Protokoll över muntliga förhandlingar och bevisupptagning skall föras av registratorn eller, efter medgivande av byråns direktör, av någon annan av byråns anställda, som har utsetts av överklagningsnämndens ordförande.
Artikel 6
Ändring av en överklagningsnämnds sammansättning
1. Om en nämnds sammansättning ändras efter muntliga förhandlingar, skall parterna underrättas om att, på begäran av någon part, nya muntliga förhandlingar skall hållas inför nämnden i dess nya sammansättning. Nya muntliga förhandlingar skall även hållas om den nya ledamoten begär detta och de övriga ledamöterna i nämnden har samtyckt till detta.
2. Den nya ledamoten skall i samma utsträckning som de övriga ledamöterna vara bunden av ett redan fattat interimistiskt beslut.
3. Om en ledamot, när en nämnd redan har fattat ett slutgiltigt beslut, är förhindrad att delta, skall denne inte ersättas av en suppleant. Om ordföranden är förhindrad att delta skall den ledamot av den berörda nämnden som har tjänstgjort längst i nämnden eller, om ledamöterna har samma tjänstgöringstid, den äldsta ledamoten underteckna beslutet för ordförandens räkning.
Artikel 7
Sammanförande av överklaganden
1. Om flera överklaganden görs av samma beslut, skall dessa överklaganden handläggas gemensamt.
2. Om överklagandena gäller olika beslut och om alla överklaganden skall handläggas av en nämnd bestående av samma ledamöter, kan den nämnden med parternas samtycke behandla dessa överklaganden gemensamt.
Artikel 8
Återförvisning till första instans
Om handläggningen vid den första instansen, vars beslut överklagandet gäller, är behäftad med allvarliga brister, skall nämnden upphäva beslutet och, om det inte föreligger skäl mot detta, återförvisa ärendet till den instansen eller själv fatta beslut i ärendet.
Artikel 9
Muntlig förhandling
1. Om muntlig förhandling skall hållas, skall nämnden sörja för att parterna har lämnat alla relevanta uppgifter och handlingar före förhandlingen.
2. Nämnden kan, tillsammans med kallelsen till muntlig förhandling, underrätta parterna om frågor som kan vara av särskild vikt eller om den omständigheten att vissa frågor inte längre verkar vara tvistiga eller ge andra upplysningar som kan bidra till att den muntliga förhandlingen kan koncentreras på de viktigaste frågorna.
3. Nämnden skall sörja för att beslut i ärendet kan fattas efter det att den muntliga förhandlingen har avslutats, om inte särskilda skäl talar mot detta.
Artikel 10
Meddelanden till parterna
Om en nämnd anser det lämpligt att meddela parterna hur nämnden kan komma att bedöma vissa sakfrågor eller rättsliga frågor skall ett sådant meddelande utformas så att det inte kan tolkas som att nämnden på något sätt är bunden av det.
Artikel 11
Synpunkter på frågor av allmänt intresse
Nämnden kan på eget initiativ eller på en skriftlig motiverad begäran av byråns direktör ge denne tillfälle att skriftligen eller muntligen framföra sina synpunkter på frågor av allmänt intresse som uppkommer i samband med handläggningen av ett ärende i nämnden. Parterna skall ha rätt att yttra sig över direktörens synpunkter.
Artikel 12
Överläggningar inför beslut
Referenten skall överlämna ett förslag till beslut till nämndens övriga ledamöter och ange en rimlig tidsfrist inom vilken invändningar kan göras eller ändringar kan föreslås. Nämnden skall sammanträda för att överlägga om det beslut som skall fattas, om det visar sig att inte alla ledamöter i nämnden har samma uppfattning. Endast nämndens ledamöter skall delta i överläggningarna. Ordföranden i den berörda nämnden kan dock tillåta andra anställda, såsom registratorer eller tolkar att närvara. Överläggningarna skall vara hemliga.
Artikel 13
Omröstningsförfarande
1. Under överläggningarna mellan en nämnds ledamöter skall referenten yttra sig först och ordföranden, såvida han själv inte är referent, sist.
2. Om omröstning är nödvändig skall rösterna avges i samma ordning, men om ordföranden även är referent skall han rösta sist. Det är inte tillåtet att avstå från att rösta.
Artikel 14
Ikraftträdande
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EG) nr 691/96 av den 16 april 1996 om klassificering av vissa varor i Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan (1), senast ändrad genom kommissionens förordning (EG) nr 586/96 (2), särskilt artikel 9 i denna, och med beaktande av följande:
För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som utgör bilaga till ovannämnda förordning är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till den här förordningen.
I förordning (EEG) nr 2658/87 fastställs allmänna bestämmelser för tolkningen av Kombinerade nomenklaturen. Dessa bestämmelser gäller också varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder som rör varuhandeln.
Enligt dessa allmänna bestämmelser måste de varor som beskrivs i kolumn 1 i tabellen i bilagan till den här förordningen klassificeras enligt motsvarande KN-nummer som anges i kolumn 2 med de motiveringar som anges i kolumn 3.
Det är lämpligt att bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter beträffande klassificeringen av varor i Kombinerade nomenklaturen och som inte överensstämmer med de rättigheter som fastställs i denna förordning fortfarande kan åberopas av innehavaren enligt bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen (3) under en period av tre månader.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Tullkodexkommitténs sektion för tulltaxe- och statistiknomenklatur.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 2
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
Artikel 3
Denna förordning träder i kraft den tjugoförsta dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EG) nr 904/96 av den 21 maj 1996 om ändring för andra gången av förordning (EG) nr 1802/95 om anpassning och ändring av de bestämmelser inom sektorn för mjölk och mjölkprodukter som innan den 1 februari 1995 fastställde vissa priser och belopp vars värde i ecu har ändrats till följd av avskaffandet av korrigeringsfaktorn för jordbruksomräkningskurserna
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 804/68 av den 27 juni 1968 om den gemensamma organisation av marknaden för mjölk och mjölkprodukter (1), senast ändrad genom kommissionens förordning (EG) nr 2931/95 (2), särskilt artikel 5c.7 i denna, och
med beaktande av följande: I bilagan till kommissionens förordning (EG) nr 1802/95 (3), ändrad genom förordning (EG) nr 2700/95 (4), har ett fel uppstått som bör rättas till.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för mjölk och mjölkprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I bilagan till förordning (EG) nr 1802/95 skall följande rad införas efter förordning (EEG) nr 1547/87 och före förordning (EEG) nr 570/88:
%gt%Plats för tabell%gt%
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EG) nr 1485/96 av den 26 juli 1996 om närmare bestämmelser för tillämpningen av rådets direktiv 92/109/EEG vad gäller kundförsäkran om särskild användning av vissa ämnen som används vid illegal tillverkning av narkotiska preparat och psykotropa ämnen (Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 92/109/EEG av den 14 december 1992 om tillverkning och utsläppande på marknaden av vissa ämnen som används vid illegal tillverkning av narkotiska preparat och psykotropa ämnen (1), ändrat genom kommissionens direktiv 93/46/EEG (2), särskilt artikel 2.1 b i detta, och med beaktande av följande:
Fastställandet av bestämmelser om kundförsäkran kommer att underlätta säkerställandet av att vid varje transaktion kundens avsedda användning av ett listat ämne, enligt definitionen i artikel 1.2 a i direktiv 92/109/EEG, klart preciseras. En sådan precisering kommer att bidra till att förhindra att listade ämnen avleds till den illegala tillverkningen av narkotiska preparat. Alla transaktioner som leder fram till att listade ämnen släpps ut på marknaden måste dokumenteras på ett tillfredsställande sätt. Dokumentationen måste dessutom innehålla en försäkran från kunden som preciserar hur ämnena skall användas.
För att ta hänsyn till regelbundna transaktioner mellan samma leverantörer och en kund bör det finnas möjlighet för kunden att lämna en enda försäkran som omfattar alla transaktioner som avser ett ämne listat i kategori 2 under en period av högst ett år, på vissa villkor.
Åtgärderna i denna förordning är förenliga med yttrandet från den kommitté som har inrättats enligt artikel 10 i rådets förordning (EEG) nr 3677/90 (3), senast ändrad genom kommissionens förordning (EEG) nr 3769/92 (4).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Försäkran för enskilda transaktioner
1. Fysiska och juridiska personer som är etablerade inom gemenskapen och som tillhandahåller kunder med något av de listade ämnena i kategori 1 eller 2 enligt bilaga I till direktiv 92/109/EEG och som är skyldiga att dokumentera varje enskild transaktion enligt artikel 2 i direktivet skall, om inte annat anges i artikel 2 i denna förordning, från kunden erhålla en försäkran om särskild användning av ämnet. Separata försäkringar skall utfärdas för varje listat ämne.
2. Försäkran skall innehålla de uppgifter som anges i exemplaret i punkt 1 i bilagan till denna förordning. Juridiska personer skall utfärda försäkran på eget brevpapper.
Artikel 2
Försäkran för flera transaktioner med ämnen i kategori 2
1. Fysiska och juridiska personer som är etablerade inom gemenskapen och som regelbundet tillhandahåller kunder med ett ämne listat i kategori 2 enligt bilaga I till direktiv 92/109/EEG och som är skyldiga att dokumentera transaktioner enligt artikel 2 i direktivet får, i stället för försäkran för enskilda transaktioner, acceptera en enda försäkran som omfattar ett antal transaktioner under en period av högst ett år om leverantören är övertygad om att följande villkor är uppfyllda:
- Kunden har erhållit leverans av ämnet vid minst tre tillfällen under de föregående tolv månaderna.
- Det finns ingen anledning att misstänka att ämnet skall användas i illegala syften.
- De beställda kvantiteterna är inte osedvanliga för denna kund.
2. Försäkran skall innehålla de uppgifter som anges i exemplet i punkt 2 i bilagan till denna förordning. Juridiska personer skall utfärda försäkran på eget brevpapper.
Artikel 3
Ikraftträdande
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EG) nr 1503/96 av den 29 juli 1996 om tillämpningsföreskrifter till rådets förordning (EG) nr 3072/95 vad gäller importtullar för ris
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 3072/95 av den 22 december 1995 om den gemensamma organisationen av marknaden för ris (1), särskilt artikel 11.2 och 11.4 i denna, och
med beaktande av följande: I artikel 11.2 tredje stycket i förordning (EG) nr 3072/95 anges metoden för beräkning av den procentsats som skall läggas till det interventionspris som gäller dagen för import, med hänsyn till beräkningen av importtull för helt slipat ris. Vid användning av denna metod skall hänsyn tas till omräkningsfaktorn, förädlingskostnaderna, värdet på biprodukter och beloppet till skydd för industrin. Dag för importen bör fastställas till den dag då deklarationen godkändes av tullmyndigheterna enligt artikel 67 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen (2), senast ändrad genom Anslutningsakten för Österrike, Finland och Sverige.
I artikel 11 i förordning (EG) nr 3072/95 fastställs att tullsatserna i Gemensamma tulltaxan skall gälla vid import av produkter enligt artikel 1 i den förordningen. För produkter enligt punkt 2 i den artikeln är importtullen lika med det interventionspris som gäller för dessa produkter vid tidpunkten för import plus en särskilt procentsats, om det rör sig om råris eller helt ris, indicaris eller japonicaris, minskat med importpriset om denna importtull inte överstiger tullsatsen i Gemensamma tulltaxan.
Det finns speciella svårigheter inom rissektorn gällande kontrollen av de importerade produkternas värde; därför är ett system med fasta värden bäst ägnat att genomföra resultatet av förhandlingarna under Uruguayrundan från och med den 1 september. Å andra sidan pågår det fortfarande tekniska diskussioner mellan de berörda parterna och i väntan på utfallet av dessa diskussioner finns det, för att garantera rättssäkerheten, anledning att behålla det system som tillämpas under 1995/96.
Vid klassificering av importerade partier skall produkterna enligt artikel 11.2 i förordning (EG) nr 3072/95 indelas i flera kvaliteter. Därför är det nödvändigt att ange vilka KN-nummer som motsvarar dessa kvaliteter.
Vid beräkning av importtullen med hjälp av schablonvärdet vid importen bör det föreskrivas att de representativa priserna vid import cif beräknas för var och en av de definierade kvaliteterna. För att detta pris skall kunna fastställas måste prisnoteringarna för de olika riskvaliteterna anges noga. Det är därför lämplig att definiera dessa prisnoteringar.
För tydlighetens och öppenhetens skull utgör prisnoteringarna för de olika ristyperna i USA:s jordbruksdepartements kungörelser en objektiv grundval vid utarbetandet av representativa importpriser cif för ris i bulk. De representativa priserna på USA:s, Thailands och andra ursprungsländers rismarknader får omvandlas till representativa priser för import cif genom tillägg av priserna för sjöfrakt på fraktmarknaden från ursprungshamnarna till en gemenskapshamn. Mot bakgrund av omfattningen av de nordeuropeiska hamnarnas transporter och handel utgör dessa hamnar den gemenskapsdestination för vilken prisnoteringar för sjöfrakt är de mest allmänt kända, mest överskådliga och mest tillgängliga. Därför är de hamnar som kan godtas, de hamnar som ligger i Nordeuropa (ARAG).
I syfte att övervaka utvecklingen av sålunda fastställda representativa importpriser cif är det lämpligt att varje vecka göra en uppföljning av de komponenter som ingår i beräkningen.
Vid fastställande av importtullar på ris enligt artikel 11.2 i förordning (EG) nr 3072/95 beaktas marknadsutvecklingen under en tvåveckors rapporteringsperiod av representativa importpriser cif för ris i bulk utan att osäkra komponenter räknas med. På grundval härav skall importtullarna för produkten fastställas på onsdagar varannan vecka och den sista arbetsdagen i varje månad, med hänsyn till det representativa medelimportpris cif som fastställs under denna period.
Den importtull som beräknas på detta sätt får tillämpas under en tvåveckorsperiod utan att importpriset efter uttagen tull påverkas. Om det för en viss produkt inte finns någon prisnotering tillgänglig under den period som representativa importpriser cif beräknas, eller om dessa representativa importpriser cif till följd av plötsliga förändringar av komponenter som ingår i beräkningen av dem undergår väsentliga fluktuationer under denna period, måste åtgärder vidtas i syfte att upprätthålla representativiteten hos importpriserna cif för den berörda produkten.
Marknadspriset på ris av sorten Basmati med ursprung i Indien och Pakistan ligger vanligtvis högre än det fastställda representativa priset. Under året 1993/94 var skillnaden 250 ecu per ton för basmatiris med ursprung i Indien och 50 ecu per ton för basmatiris med ursprung i Pakistan. Därför bör importtullen för dessa rissorter minskas med de angivna beloppen i syfte att följa principen i artikel 11 i förordning (EG) nr 3072/95 och i syfte att iaktta gemenskapens internationella förpliktelser.
I avsaknad av prisnoteringar är det lämpligt att tills vidare tillämpa den tull som fastställts för föregående period och att, vid stora fluktuationer i prisnoteringarna, sjöfraktskostnaderna eller i den omräkningskurs som tillämpas vid beräkningen av det representativa importpriset cif för produkten i fråga, åter söka göra dessa priser representativa med hjälp av en motsvarande justering av den konstaterade skillnaden i förhållande till gällande fastställda pris för att ta hänsyn till uppkomna förändringar. Även om en sådan ändring kommer till stånd påverkar inte detta tidpunkten för följande prisfastställande.
Förvaltningskommittén för spannmål har inte avgivit något yttrande inom den tidsfrist som dess ordförande bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De importtullar som avses i artikel 11.1 och 11.2 i förordning (EG) nr 3072/95 skall vara de som tillämpas vid den tidpunkt som avses i artikel 67 i förordning (EEG) nr 2913/92.
Artikel 2
Importtullen för helt slipat ris enligt KN-nummer 1006 30 skall motsvara interventionspriset vid tidpunkten för importen ökat med
- 163 % i fråga om indicaris,
- 167 % i fråga om japonicaris
och minskat med importpriset.
I alla händelser får denna importtul inte överstiga tullsatsen enligt Gemensamma tulltaxan.
Artikel 3
1. I denna förordning avses med indicaris ris enligt KN-nummer: 1006 20 17, 1006 20 98, 1006 30 27, 1006 30 48, 1006 30 67, 1006 30 98.
2. Alla andra produkter enligt KN-nummer 1006 20 och 1006 30 skall anses vara japonicaris.
Artikel 4
1. Importtullen för de produkter som avses i artikel 3 skall beräknas varje vecka men fastställas av kommissionen på onsdagen varannan vecka och den sista arbetsdagen i varje månad för tillämpning nästföljande arbetsdag respektive första dagen i nästföljande månad, och för perioden fram till den första torsdagen i juli månad 1995, från och med den 1 juli detta år enligt den metod som avses i artikel 5.
Om det efter fastställandet för följande vecka konstateras att den beräknade importtullen avviker med 10 ecu per ton eller mer från gällande importtull skall dock en motsvarande justering göras av kommissionen.
Det fastställande av importtullen som görs den sista arbetsdagen i varje månad baseras på interventionspriset för följande månad.
Om onsdagen då importtullen skall fastställas inte är en arbetsdag för kommissionen skall fastställandet göras närmast följande arbetsdag.
2. Det gällande världsmarknadspris som skall beaktas vid beräkningen av importtullen skall vara medeltalet av de representativa priserna för import cif i bulk under en vecka, beräknade i enlighet med metoden i artikel 5 och fastställda under de två föregående veckorna.
3. De importtullar som fastställs i enlighet med denna förordning skall tillämpas till dess att ett nytt fastställande träder i kraft.
Om det i fråga om en produkt inte finns någon prisnotering som kan utgöra referenspris i enlighet med artikel 5 under de två veckor som föregår nästa periodiska fastställande, skall den tidigare fastställda importtullen fortsätta att gälla.
Efter varje fastställande eller justering skall kommissionen i Europeiska gemenskapernas officiella tidning offentliggöra importtullarna och de komponenter som ingår i beräkningen av dem.
4. För de basmatiris enligt KN-nummer ex 1006 20 17 och ex 1006 29 98 får en nedsättning av importtullen som fastställs i enlighet med punkt 1 göras med ett belopp på 250 ecu för ris med ursprung i Indien och 50 ecu för ris med ursprung i Pakistan.
Denna nedsättning skall verkställas om en importlicens som utfärdats mot ställande av en säkerhet liksom ett ursprungsintyg för produkten visas upp vid övergången till fri omsättning.
Med undantag från artikel 10 a i kommissionens förordning (EG) nr 1162/95 (3) skall den säkerhet som ställs vara 275 ecu per ton för basmatiris med ursprung i Indien och 75 ecu per ton för basmatiris med ursprung i Pakistan.
Ursprungsintyget skall upprättas enligt förebilden i bilaga II. Det skall utfärdas i enlighet med relevant bestämmelse i kommissionens förordning (EEG) nr 81/92 (4).
De belopp som anges i första stycket i denna punkt får ses över mot bakgrund av marknadsutvecklingen.
Artikel 5
1. I syfte att fastställda det importpris på ris som avses i artikel 11.4 i förordning (EG) nr 3072/95 skall följande komponenter beaktas för olika sorters ris i bulk enligt artikel 3:
a) Priset cif Rotterdam.
b) Det representativa priset på Thailands marknad.
c) Det representativa priset på USA:s marknad.
d) Det representativa priset på övriga marknader.
e) Fraktkostnaderna mellan ursprungshamnen å ena sidan och hamnen i Antwerpen, Rotterdam, Amsterdam eller Gent å andra sidan.
Importpriset skall normalt vara det som anges i a, men i avsaknad av ett sådant pris skall det fastställas på grundval av de komponenter som anges i b, c och e. Det pris som anges i d skall inte användas, utom i avsaknad av priser enligt a, b och c.
I avsaknad av prisnoteringar för sjöfrakt av ris skall de för spannmål användas.
2. Dessa komponenter skall noteras och bekräftas varje vecka på grundval av de källor och den referenskvalitet som återges i bilaga I till denna förordning. Sjöfraktskostnaderna skall noteras på grundval av den offentliga information som finns tillgänglig.
Om det noterade priset anges som c. %amp% f. skall det ökas med 0,75 %.
Artikel 6
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
Förordningen är tillämplig från och med den 1 september 1996.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EG) nr 2400/96 av den 17 december 1996 om upptagandet av vissa namn i %quot%Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar%quot% som föreskrivs i rådets förordning (EEG) nr 2081/92 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel (Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2081/92 av den 14 juli 1992 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel (1), särskilt artikel 6.3 och 6.4 i denna, och med beaktande av följande:
I enlighet med artikel 5 i förordning (EEG) nr 2081/92 har medlemsstaterna till kommissionen lämnat in ansökningar om inregistrering av geografisk eller ursprungsbeteckning för vissa namn.
I enlighet med artikel 6.1 i den förordningen har det konstaterats att dessa är förenliga med den förordningen, särskilt att de innehåller alla de uppgifter som föreskrivs i artikel 4 i den förordningen.
Ingen invändning enligt artikel 7 i den förordningen har framställts till kommissionen efter offentliggörandet av berörda namn i Europeiska gemenskapernas officiella tidning (2).
Följaktligen bör dessa namn tas upp i %quot%Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar%quot% och alltså skyddas på gemenskapsnivå i egenskap av geografisk eller ursprungsbeteckning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De namn som finns upptagna i bilagan skall tas upp i %quot%Register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar%quot% såsom geografiskt skyddad beteckning (PGI) eller skyddad ursprungsbeteckning (PDO) i enlighet med artikel 6.3 i förordning (EEG) nr 2081/92.
Artikel 2
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS BESLUT av den 28 februari 1997 om upprättande av en förteckning över de tredje länder från vilka medlemsstaterna tillåter import av köttprodukter (Text av betydelse för EES) (97/222/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 72/462/EEG av den 12 december 1972 om hälsoproblem och problem som rör veterinärbesiktning vid import från tredje land av nötkreatur, svin och färskt kött (1), senast ändrat genom direktiv 96/91/EG (2), särskilt artiklarna 21a och 22 i detta,
med beaktande av rådets direktiv 92/118/EEG av den 17 december 1992 om djurhälso- och hygienkrav för handel inom gemenskapen med produkter, som inte omfattas av sådana krav i de särskilda gemenskapsbestämmelser som avses i bilaga A.1 till direktiv 89/662/EEG och, i fråga om patogener, i direktiv 90/425/EEG, samt för import till gemenskapen av sådana produkter (3), senast ändrat genom direktiv 96/90/EG (4), särskilt artikel 10 punkt 2 c i detta, och
med beaktande av följande: I rådets beslut 79/542/EEG (5), senast ändrat genom beslut 97/160/EG (6), upprättas en förteckning över de tredje länder från vilka medlemsstaterna tillåter import av bland annat köttprodukter av kött från nötkreatur, svin, hovdjur, får och getter.
I kommissionens beslut 91/449/EG (7), senast ändrat genom beslut 96/92/EG (8), upprättas förteckningar över de tredje länder från vilka medlemsstaterna tillåter import av köttprodukter av nötkreatur, svin, hästdjur, får och getter.
I kommissionens beslut 94/85/EG (9), senast ändrat genom beslut 96/2/EG (10), upprättas en förteckning över de tredje länder från vilka medlemsstaterna tillåter import av färskt fjäderfäkött. Denna förteckning gäller också import av köttprodukter av fjäderfäkött.
I kommissionens beslut 94/86/EG (11), ändrad genom beslut 96/137/EG (12), upprättas en förteckning över de tredje länder från vilka medlemsstaterna tillåter import av viltkött. Denna förteckning gäller import av viltköttsprodukter.
I kommissionens beslut 94/278/EG (13), senast ändrat genom beslut 96/344/EG (14), upprättas en förteckning över de tredje länder från vilka medlemsstaterna tillåter import av bland annat köttprodukter av kaninkött, hägnat fjädervilt och hägnat pälsvilt.
Kommissionens beslut 91/449/EEG upphävs genom kommissionens beslut 97/221/EG (15).
En ändrad förteckning bör upprättas över de godkända tredje länder från vilka import tillåts av köttprodukter som inte enbart framställts av kött från nötkreatur, svin, hästdjur, får och getter utan också av kött från hägnat vilt, tamkaniner och vilt.
Vilka typer av köttprodukter som får importeras från tredje land beror på hälsosituationen i det tredje landet eller delar av tredje land där produkterna framställts. För att få importeras måste vissa köttprodukter ha genomgått en särskild behandling.
I rådets direktiv 77/99/EEG (16), senast ändrat genom rådets direktiv 95/68/EG (17), definieras en köttprodukt genom att lägsta krav för behandlling fastställs. Vissa tredje länder eller delar av tredje land som finns med i ovan nämnda förteckning skall bara godkännas för import av köttprodukter som har genomgått en fullständig värmebehandling.
I beslut 97/221/EG fastställs de djurhälsovillkor och veterinärintyg som skall tillämpas av medlemsstaterna vid import av köttprodukter från tredje land.
Lägsta behandlingskrav bör fastställas för import av dessa produkter från det tredje land där de produceras.
De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Medlemsstaterna skall tillåta import av köttprodukter enligt definition i beslut 97/221/EG från de tredje länder eller delar av tredje land som är upptagna i förteckningarna i delarna I, II och III i bilagan, under förutsättning att de har genomgått en lämplig behandling i enlighet med del IV i bilagan och åtföljs av lämpligt veterinärintyg enligt beslut 97/221/EG.
Artikel 2
Detta beslut skall gälla från och med den 1 mars 1997.
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
RÅDETS FÖRORDNING (EG) nr 1139/98 av den 26 maj 1998 om obligatoriska uppgifter vid märkning av vissa livsmedel som framställs från genetiskt modifierade organismer utöver de uppgifter som föreskrivs i direktiv 79/112/EEG
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 79/112/EEG av den 18 december 1978 om tillnärmning av medlemsstaternas lagstiftning om märkning, presentation och reklam i fråga om livsmedel (1), särskilt artikel 4.2 i detta, med beaktande av kommissionens förslag, och
med beaktande av följande:
(1) Med tillämpning av bestämmelserna i del C i rådets direktiv 90/220/EEG av den 23 april 1990 om avsiktlig utsättning av genetiskt modifierade organismer i miljön (2) har tillstånd för utsläppande på marknaden av vissa genetiskt modifierade organismer beviljats genom kommissionens beslut 96/281/EG av den 3 april 1996 om utsläppande på marknaden av genetiskt modifierade sojabönor (Glycine max L.) med förhöjd tolerans mot bekämpningsmedlet glyfosat enligt rådets direktiv 90/220/EEG (3) och genom kommissionens beslut 97/98/EG av den 23 januari 1997 om utsläppande på marknaden av genetiskt modifierad majs (Zea mays L.) med följande kombinerade modifikation: BT-endotoxin-genens insekticidverkan och ökad tolerans mot herbiciden glufosinatammonium i enlighet med rådets direktiv 90/220/EEG (4).
(2) I enlighet med direktiv 90/220/EEG har det inte funnits några säkerhetsskäl för att vid märkning av genetiskt modifierade sojabönor (Glycine max L.) eller genetiskt modifierad majs (Zea mays L.) nämna att dessa har framställts genom metoder för genetisk modifiering.
(3) Direktiv 90/220/EEG omfattar inte icke-levande produkter som har häletts från genetiskt modifierade organismer (i det följande betecknade %quot%GMO%quot%).
(4) Vissa medlemsstater har vidtagit åtgärder i fråga om märkning av livsmedel och livsmedelsingredienser som har framställts från de berörda produkterna. Skillnaderna mellan dessa åtgärder kan hindra den fria rörligheten för dessa livsmedel och livsmedelsingredienser och därigenom negativt påverka den inre marknadens funktion. Det är därför nödvändigt att anta enhetliga gemenskapsregler om märkning av de berörda produkterna.
(5) I artikel 8 i Europaparlamentets och rådets förordning (EG) nr 258/97 av den 27 januari 1997 om nya livsmedel och nya livsmedelsingredienser (5) meddelas ytterligare särskilda bestämmelser för märkning vilka skall säkerställa att konsumenten erhåller relevant information. Dessa ytterligare särskilda bestämmelser för märkning gäller inte för livsmedel och livsmedelsingredienser som i stor utsträckning användes för konsumtion inom gemenskapen innan förordning (EG) nr 258/97 trädde i kraft och som därför inte betraktas som nya.
(6) För att undvika en snedvridning av konkurrensen bör märkningsregler för livsmedel och livsmedelsingredienser som består av eller har härletts från genetiskt modifierade organismer och som i enlighet med ett enligt direktiv 90/220/EEG beviljat tillstånd släpptes ut på marknaden innan förordning (EG) nr 258/97 trädde i kraft och märkningsregler för livsmedel och livsmedelsingredienser som släpps ut på marknaden efter ikraftträdandet, grundas på samma principer.
(7) Genom kommissionens förordning (EG) nr 1813/97 av den 19 september 1997 om obligatoriska uppgifter vid märkning av vissa livsmedel som framställs av genetiskt modifierade organismer utöver de uppgifter som föreskrivs i direktiv 79/112/EEG (6) har allmänna märkningsregler fastställts för de ovannämnda produkterna.
(8) Det är nu angeläget att snabbt fastställa detaljerade och enhetliga gemenskapsregler för märkning av de livsmedel som omfattas av förordning (EG) nr 1813/97.
(9) Det är nödvändigt att, i enlighet med det tillvägagångssätt som används i artikel 8 i förordning (EG) nr 258/97, se till att den slutliga konsumenten informeras om sådana särdrag och egenskaper hos ett livsmedel eller en livsmedelsingrediens som gör att det inte längre är jämförbart med ett befintligt livsmedel eller en befintlig livsmedelsingrediens, t.ex. dess sammansättning, näringsvärde, näringsmässiga effekter eller avsedda användning. Livsmedel och livsmedelsingredienser som framställs från genetiskt modifierade sojabönor eller från genetiskt modifierad majs och som inte är jämförbara med traditionella motsvarigheter bör därför omfattas av bestämmelser för märkning.
(10) I enlighet med det tillvägagångssätt som används i artikel 8 i förordning (EG) nr 258/97 måste bestämmelserna för märkning grundas på en vetenskaplig bedömning.
(11) Det är nödvändigt att fastställa tydliga märkningsregler för de ovannämnda produkterna som möjliggör en tillförlitlig, enkelt reproducerbar och praktiskt genomförbar offentlig kontroll. Gemensamma, vetenskapligt validerade testmetoder bör därför utvecklas.
(12) Det är också nödvändigt att se till att bestämmelserna för märkning inte blir onödigt betungande men ändå tillräckligt detaljerade för att förse konsumenterna med den information de behöver.
(13) Livsmedlens och livsmedelsingrediensernas innehåll av protein eller DNA som är ett resultat av genetiskt modifiering är idag det kriterium som bäst uppfyller ovannämnda krav. Ett sådant synsätt kan komma att omprövas mot bakgrund av nya vetenskapliga kunskaper.
(14) Oavsiktlig förorening av livsmedel med DNA eller protein som är ett resultat av genetisk modifiering kan inte uteslutas. Märkning till följd av en sådan förorening kan undvikas genom att ett tröskelvärde fastställs för upptäckt av DNA och protein.
(15) Frågan om det är möjligt att bestämma en de-minimiströskel för förekomst av DNA eller protein som ett resultat av genetisk modifiering och, i så fall, på vilken nivå detta kan ske, bör snabbt övervägas mot bakgrund av relevanta vetenskapliga utlåtanden.
(16) Livsmedel och livsmedelsingredienser som framställs från genetiskt modifierade sojabönor (Glycine max L.) eller från genetiskt modifierad majs (Zea mays L.) som innehåller DNA som är ett resultat av genetisk modifiering är inte jämförbara och de bör därför omfattas av bestämmelser för märkning.
(17) Protein eller DNA som är ett resultat av genetiskt modifiering kan ha förstörts genom flera på varandra följande bearbetningssteg. I detta fall bör livsmedlen eller livsmedelsingredienserna betraktas som jämförbara från märkningssynpunkt. De bör därför inte omfattas av bestämmelser för märkning. En förteckning över sådana produkter bör upprättas.
(18) Med vissa bearbetningsmetoder är det emellertid möjligt att eliminera DNA men däremot inte proteiner. Det kan inte uteslutas att sådana metoder kan användas med avseende på livsmedel. Livsmedel och livsmedelsingredienser som inte innehåller DNA som är ett resultat av genetisk modifiering, men däremot proteiner som är ett resultat av sådan modifiering, kan inte betraktas som jämförbara. De bör därför omfattas av bestämmelser för märkning.
(19) De nödvändiga upplysningarna bör framgå av ingrediensförteckningen. Om ingrediensförteckning saknas bör uppgifterna anges tydligt på produktens märkning.
(20) Denna förordning påverkar inte tillverkarens rätt att på produktens etikett göra andra påståenden än dem som föreskrivs i denna förordning (t.ex. påståenden om att produkten inte innehåller livsmedel och livsmedelsingredienser som framställts från genetiskt modifierad soja eller majs, eller uppgifter om att sådana livsmedel och livsmedelsingredienser ingår i produkten, när detta inte kan kontrolleras med vetenskapliga metoder men kan visas på annat sätt), under förutsättning att sådana påståenden görs i enlighet med bestämmelserna i direktiv 79/112/EEG.
(21) Med beaktande av deras räckvidd och effekter är de gemenskapsbestämmelser som införs genom denna förordning inte bara nödvändiga utan också avgörande för att nå de uppställda målen. Dessa mål kan inte nås av medlemsstaterna om de handlar var för sig.
(22) Denna förordning ersätter kommissionens förordning (EG) nr 1813/97 som därför bör upphävas.
(23) I enlighet med det förfarande som anges i artikel 17 i direktiv 79/112/EEG överlämnades denna text till Ständiga livsmedelskommittén, vilken dock inte haft möjlighet att avge något yttrande. Enligt samma förfarande överlämnade kommissionen ett förslag till rådet om de åtgärder som bör vidtas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Denna förordning skall gälla livsmedel och livsmedelsingredienser avsedda att som sådana överlämnas till den slutliga konsumenten (i det följande betecknade %quot%de angivna livsmedlen%quot%) och som helt eller delvis framställts från.
- genetiskt modifierade sojabönor som omfattas av beslut 96/281/EG,
- genetiskt modifierad majs som omfattas av beslut 97/98/EG.
2. Denna förordning skall inte gälla livsmedelstillsatser, aromer för användning i livsmedel eller extraktionsmedel som används vid framställning av livsmedel enligt artikel 2.1 i förordning (EG) nr 258/97.
Artikel 2
1. De angivna livsmedlen skall omfattas av de ytterligare särskilda bestämmelser för märkning som anges i punkt 3.
2. Angivna livsmedel utan förekomst av vare sig protein eller DNA som är ett resultat av genetisk modifiering skall inte omfattas av de ytterligare särskilda bestämmelserna för märkning.
En förteckning över produkter som inte omfattas av de ytterligare särskilda bestämmelserna för märkning skall utarbetas i enlighet med förfarandet i artikel 17 i direktiv 79/112/EEG under beaktande av den tekniska utredningen, yttrandet från Vetenskapliga livsmedelskommittén och relevanta vetenskapliga utlåtanden.
3. De ytterligare särskilda bestämmelserna för märkning skall vara följande:
a) Om livsmedlet består av mer än en ingrediens skall texten %quot%framställd från genetiskt modifierad soja%quot% eller %quot%framställd från genetiskt modifierad majs%quot%, beroende på vilket som är tillämpligt, anges inom parentes omedelbart efter namnet på den berörda ingrediensen i den ingrediensförteckning som avses i artikel 6 i direktiv 79/112/EEG. Alternativt kan denna text placeras i en väl synlig fotnot till ingrediensförteckningen, med en asterisk (*) som hänvisar till ingrediensen i fråga. Om en ingrediens redan återfinns i förteckningen över ingredienser som har framställts från soja eller majs kan texten %quot%framställd från genetiskt modifierad . . .%quot% förkortas till %quot%genetiskt modifierad%quot%. Om den förkortade texten står i en fotnot till ingrediensförteckningen skall asterisken direkt hänvisa till ordet %quot%soja%quot% eller %quot%majs%quot%. Oavsett vilken textvariant som används i fotnoten till ingrediensförteckningen, skall den vara tryckt med ett typsnitt av minst samma storlek som det som finns i ingrediensförteckningen.
b) I fråga om produkter för vilka ingrediensförteckning saknas skall texten %quot%framställd från genetiskt modifierad soja%quot% eller %quot%framställd från genetiskt modifierad majs%quot%, beroende på vilket som är tillämpligt, tydligt anges på livsmedlets märkning.
c) När en ingrediens anges med namnet på en kategori i enlighet med artikel 6.5 b första strecksatsen i direktiv 79/112/EEG skall denna beteckning kompletteras med texten %quot%innehåller . . . (*) framställd(a) från genetiskt modifierad soja/genetiskt modifierad majs
(*) Uppgift om ingrediensen/ingredienserna.%quot%, beroende på vilket som är tillämpligt.
d) Om en beståndsdel av en sammansatt ingrediens har härletts från de angivna livsmedlen, skall den anges på slutproduktens märkning med den tilläggstext som anges i punkt b.
4. Denna artikel skall inte påverka tillämpningen av andra bestämmelser i gemenskapslagstiftningen rörande märkning av livsmedel.
Artikel 3
Kommissionens förordning (EG) nr 1813/97 upphävs.
Artikel 4
1. Bestämmelserna för märkning i denna förordning skall inte gälla produkter som lagligen har tillverkats och märkts i gemenskapen eller som lagligen har importerats till gemenskapen och övergått i fri omsättning innan denna förordning träder i kraft.
2. Tillämpningen av artikel 2 på produkter som släpps ut på marknaden i enlighet med kommissionens förordning (EG) nr 1813/97 med en märkning som anger förekomst av genetiskt modifierat material får uppskjutas till sex månader efter det att denna förordning träder i kraft.
Artikel 5
Denna förordning träder i kraft 90 dagar efter det att den offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EG) nr 1367/98 av den 29 juni 1998 om ändring av förordning (EEG) nr 94/92 om genomförande av den ordning för import från tredje land som föreskrivs i rådets förordning (EEG) nr 2092/91 (Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2092/91 av den 24 juni 1991 om ekologisk produktion av jordbruksprodukter och uppgifter därom på jordbruksprodukter och livsmedel (1), senast ändrad genom kommissionens förordning (EG) nr 1488/97 (2), särskilt artikel 11 i denna, och med beaktande av följande:
I artikel 11.1 i förordning (EEG) nr 2092/91 föreskrivs att produkter som importeras från tredje land endast får marknadsföras om de härrör från ett tredje land som står upptaget i en förteckning som upprättats enligt villkoren i punkt 2 i nämnda artikel. En sådan förteckning har fastställts i bilagan till kommissionens förordning (EEG) nr 94/92 (3), senast ändrad genom förordning (EG) nr 314/97 (4).
Ungern och Schweiz har upptagits i förordning (EG) nr 314/97 i den förteckning som avses i artikel 11.1 i förordning (EEG) nr 2092/91 för en period som löper ut den 30 juni 1998 för att man under denna period noggrant skall granska vissa aspekter gällande genomförandet i dessa länder av regler likvärdiga dem som fastställs i förordning (EEG) nr 2092/91.
Det faktiska genomförandet i Ungern av regler likvärdiga dem som fastställs i förordning (EEG) nr 2092/91 har bekräftats genom en kontroll på plats som utförs av kommissionen.
Schweiz har godkänt ett nytt kontrollorgan som kommer att genomföra de kontroller som krävs enligt schweiziska bestämmelser för ekologiskt jordbruk.
För att systemet skall fungera bör det för varje tredje land fastställas vilka organ som skall utfärda kontrollintyg enligt artikel 11.1 b i förordning (EEG) nr 2092/91.
Australien har meddelat ändringar i sitt kontrollsystem. Kontrollerna av aktörer i Australien görs för närvarande av privata kontrollorgan som övervakas av en offentlig myndighet.
Israel har bekräftat att kontroll och utfärdande av intyg för ekologiska produkter kommer att skötas av jordbruksministeriet.
Genomgången av de uppgifter som har lämnats in av de ovannämnda tredje länderna visar att kraven motsvarar vad som krävs enligt gemenskapsrätten.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från den kommitté som anges i artikel 14 i förordning (EEG) nr 2092/91.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till förordning (EEG) nr 94/92 skall ändras enligt bilagan till denna förordning.
Artikel 2
Denna förordning träder i kraft den 1 juli 1998.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS FÖRORDNING (EG) nr 2767/98 av den 21 december 1998 om ändring av förordning (EG) nr 2300/97 om tillämpningsföreskrifter för rådets förordning (EG) nr 1221/97 om allmänna tillämpningsregler för åtgärder som syftar till att förbättra villkoren för produktion och saluföring av honung
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1221/97 av den 25 juni 1997 om allmänna tillämpningsregler för åtgärder som syftar till att förbättra villkoren för produktion och saluföring av honung (1), ändrad genom rådets förordning (EG) nr 2070/98 (2), särskilt artikel 5 i denna, och
av följande skäl: I kommissionens förordning (EG) nr 2300/97 (3), senast ändrad genom förordning (EG) nr 2633/98 (4), fastställs nödvändiga tillämpningsföreskrifter för åtgärder som syftar till att förbättra villkoren för produktion och saluföring.
För att möjliggöra en viss flexibilitet i genomförandet av programmet får de ekonomiska ramarna för varje åtgärd variera med ett visst procenttal utan att överstiga de totala begränsningarna för det årliga programmet. Om denna flexibilitet utnyttjas inom programmet får finansieringen från gemenskapen inte överstiga 50 % av de kostnader för vilka den berörda medlemsstaten betalar ut ersättning.
De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för fjäderfäkött och ägg.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Följande artikel 4 a skall läggas till i förordning (EG) nr 2300/97:
%quot%Artikel 4 a
De ekonomiska ramarna för varje åtgärd får ökas eller minskas med högst 10 %, utan att vare sig de totala begränsningarna för det årliga programmet överstigs eller gemenskapens finansiering av programmet som avses i artikel 3 överstiger 50 % av de kostnader för vilka den berörda medlemsstaten betalar ut ersättning.%quot%
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS BESLUT av den 22 juni 1998 om ingående av ett avtal om ömsesidigt erkännande mellan Europeiska gemenskapen och Amerikas förenta stater (1999/78/EG)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 113, tillsammans med artikel 228.2 första meningen och 228.3 första stycket, samt artikel 228.4 i detta,
med beaktande av kommissionens förslag, och
av följande skäl: Avtalet om ömsesidigt erkännande mellan Europeiska gemenskapen och Amerikas förenta stater, vilket undertecknades i London den 18 maj 1998, har framförhandlats och bör godkännas.
Vissa genomförandeuppgifter har anförtrotts den gemensamma kommitté som inrättas genom avtalet, särskilt befogenheten att ändra vissa aspekter av de sektoriella bilagorna till detta.
För att säkerställa att avtalet fungerar korrekt bör tillämpliga interna förfaranden fastställas och det är nödvändigt att bemyndiga kommissionen att göra vissa ändringar av teknisk natur i avtalet och att fatta vissa beslut för dess genomförande.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Avtalet om ömsesidigt erkännande mellan Europeiska gemenskapen och Amerikas förenta stater, inbegripet dess bilagor, godkänns härmed på Europeiska gemenskapens vägnar.
Texten till avtalet och bilagorna till det bifogas detta beslut.
Artikel 2
Rådets ordförande skall på gemenskapens vägnar överlämna den skrivelse som avses i artikel 21.1 i avtalet (1).
Artikel 3
1. Gemenskapen skall i den gemensamma kommitté som föreskrivs i artikel 14 i avtalet och i de gemensamma sektoriella kommittéer som inrättas genom de sektoriella bilagorna företrädas av kommissionen, som skall biträdas av den särskilda kommitté som utsetts av rådet. Kommissionen skall efter samråd med denna särskilda kommitté verkställa de utseenden och anmälningar, det informationsutbyte och de framställningar om inspektioner som avses i artiklarna 10 b, 12, 13 och 14.2 i avtalet och i motsvarande bestämmelser i de sektoriella bilagorna.
2. Gemenskapens ståndpunkt vad gäller beslut som skall fattas av den gemensamma kommittén eller i förekommande fall av de gemensamma sektoriella kommittéerna skall, såvitt gäller ändringar i de sektoriella bilagorna (artikel 14.4 b och artiklarna 7 9 i avtalet samt de motsvarande bestämmelserna i de sektoriella bilagorna) samt kontroll enligt artikel 7 d i avtalet av att gällande krav är uppfyllda, fastställas av kommissionen efter samråd med den särskilda kommitté som avses i punkt 1 i den här artikeln.
3. I samtliga övriga fall skall gemenskapens ståndpunkt i den gemensamma kommittén eller i de gemensamma sektoriella kommittéerna fastställas av rådet som skall fatta sina beslut med kvalificerad majoritet på förslag av kommissionen. Samma förfarande skall gälla för beslut som fattas av gemenskapen inom ramen för artiklarna 16 och 21 i avtalet.
KOMMISSIONENS BESLUT av den 17 mars 1999 om ändring av rådets beslut 79/542/EEG och beslut 92/160/EEG och 93/197/EEG när det gäller djurhälsovillkor för import till gemenskapen av registrerade hästar från vissa delar av Kirgizistan [delgivet med nr K(1999) 609] (Text av betydelse för EES) (1999/236/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 90/426/EEG av den 26 juni 1990 om djurhälsovillkor vid förflyttning och import av hästdjur från tredje land (1), senast ändrat genom Anslutningsakten för Österrike, Finland och Sverige, särskilt artiklarna 12, 13, 15 och 16 samt artikel 19 ii i detta, och
av följande skäl: (1) Genom rådets beslut 79/542/EEG (2), senast ändrat genom beslut 1999/227/EG (3), upprättas en förteckning över tredje länder från vilka medlemsstaterna tillåter import av nötkreatur, svin, hästdjur, får och getter samt färskt kött och köttprodukter.
(2) Genom kommissionens beslut 92/160/EEG (4), senast ändrat genom beslut 1999/228/EG regionaliseras vissa tredje länder när det gäller import av hästdjur.
(3) Krav avseende djurhälsa och veterinärintyg vid import av registrerade hästar fastställs i kommissionens beslut 93/197/EEG (5), senast ändrat genom beslut 1999/227/EG.
(4) Efter att representanter för kommissionen gjort en veterinärinspektion i Kirgizistan gjordes bedömningen att de veterinära myndigheterna i detta land har en tillfredsställande kontroll över hälsosituationen för hästdjur.
(5) De veterinära myndigheterna i Kirgizistan har gjort ett skriftligt åtagande att inom 24 timmar meddela kommissionen och medlemsstaterna via fax, telegram eller telex om någon av de smittsamma sjukdomar hos hästdjur som finns upptagna i förteckningen över anmälningspliktiga sjukdomar i bilaga A till direktiv 90/426/EEG har kunnat konstateras i landet i fråga. Åtagandet innebär också att de veterinära myndigheterna inom rimlig tid och på det sätt som anges ovan skall underrätta kommissionen och medlemsstaterna om alla förändringar som görs av vaccinations- eller importbestämmelserna beträffande hästdjur. (6) Hästar i Kirgizistan testas varje år för rots, och under åtminstone sex månader har inga nya fynd gjorts. Vidare har afrikansk hästpest, Venezuelan equine encephalomyelitis och vesikulär stomatit aldrig förekommit i Kirgizistan.
(7) Kontrollen av virusarterit hos häst har just påbörjats, så landets status när det gäller denna sjukdom kan ännu inte fastställas. Okastrerade hingstar som är äldre än 180 dagar och som är avsedda för import till gemenskapen bör därför bli föremål för laboratorietester avseende denna sjukdom.
(8) Beskällarsjuka (dourine) har rapporterats från vissa delar av Kirgizistan. Regionen Issyk-Kul har dock varit fri från beskällarsjuka under minst sex månader, och officiella garantier har lämnats för att transporter och förflyttningar av hästdjur till denna region från resten av landet är föremål för officiella veterinärkontroller.
(9) Med tanke på hälsosituationen för hästdjur i vissa delar av Kirgizistan verkar det lämpligt att regionalisera landet i fråga, så att gemenskapen kan tillåta import till medlemsstaternas territorier av registrerade hästar från de delar av Kirgizistans territorium som är fria från sjukdom.
(10) Kraven avseende djurhälsa och veterinärintyg måste anpassas efter djurhälsosituationen i det berörda tredje landet. Föreliggande beslut avser bara registrerade hästar.
(11) Beslut 79/542/EEG samt beslut 92/160/EEG och 93/197/EEG bör ändras i enlighet med detta.
(12) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I den särskilda kolumnen för registrerade hästar i del 2 i bilagan till beslut 79/542/EEG skall följande rad läggas till, i enlighet med ISO-kodens korrekta alfabetiska placering:
%gt%Plats för tabell%gt%
Artikel 2
Bilagan till beslut 92/160/EEG skall ändras på följande sätt:
1) Följande ord skall läggas till:
%quot%Kirgizistan (4)
Regionen Issyk-Kul.%quot% 2) Följande fotnot skall läggas till:
%quot%(4) Endast permanent import till gemenskapen av registrerade hästar godkänns.%quot%
Artikel 3
Kommissionens beslut 93/197/EEG ändras på följande sätt:
1. I den förteckning över tredje länder tillhörande grupp B som återfinns i bilaga I skall %quot%Kirgizistan (1) (2) (KG)%quot% läggas till, i enlighet med ISO-kodens korrekta alfabetiska placering.
2. I bilaga II skall titeln på hälsointyget för tredje länder som tillhör grupp B ersättas med följande:
%quot%B - HÄLSOINTYG
för import till gemenskapens territorium av registrerade hästar från Kirgizistan (1) och för import av registrerade hästdjur respektive hästdjur för avel och produktion från Australien, Bosnien och Hercegovina, Bulgarien, Vitryssland, Cypern, Tjeckiska republiken, Estland, Kroatien, Ungern, Litauen, Lettland, f.d. jugoslaviska republiken Makedonien, Nya Zeeland, Polen, Rumänien, Ryssland (1), Slovakiska republiken, Slovenien, Ukraina och Förbundsrepubliken Jugoslavien.%quot%
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS BESLUT
av den 31 maj 1999
om ändring av beslut 94/448/EG om särskilda villkor för import av fiskeri- och vattenbruksprodukter med ursprung i Nya Zeeland
[delgivet med nr K(1999) 1404]
(Text av betydelse för EES)
(1999/402/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/493/EEG av den 22 juli 1991 om fastställande av hygienkrav för produktionen och marknadsföringen av fiskprodukter(1), senast ändrat genom direktiv 97/79/EG(2), särskilt artikel 11.1 i detta, och
av följande skäl: (1) I artikel 1 i kommissionens beslut 94/448/EG av den 20 juni 1994 om särskilda villkor för import av fiskeri- och vattenbruksprodukter med ursprung i Nya Zeeland, senast ändrat genom beslut 96/254/EG(3), anges att Ministry of Agriculture and Fisheries (MAF) skall vara den behöriga myndighet i Nya Zeeland som ansvarar för kontrollen av att fiskeri- och vattenbruksprodukterna uppfyller kraven enligt direktiv 91/493/EEG.
(2) Efter omstruktureringen av regeringen i Nya Zeeland har behörigheten att utfärda hälsointyg övergått från Ministry of Agriculture and Fisheries till Ministry of Agriculture and Forestry. Denna nya myndighet har möjlighet att effektivt kontrollera hur gällande lagstiftning tillämpas. Därför är det nödvändigt att ändra utnämningen av den behöriga myndighet som anges i beslut 94/448/EG.
(3) Det är lämpligt att harmonisera ordalydelsen i kommissionens beslut 94/448/EG med lydelsen i kommissionsbeslut av senare datum genom att fastställa särskilda villkor för import av fiskeri- och vattenbruksprodukter med ursprung i vissa tredje länder.
(4) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Kommissionens beslut 94/448/EG ändras på följande sätt:
1) Artikel 1 skall ersättas med följande: %quot%Artikel 1
'The Ministry of Agriculture and Forestry (MAF)' skall vara den behöriga myndighet i Nya Zeeland som ansvarar för att kontrollera och intyga att fiskeri- och vattenbruksprodukterna uppfyller kraven enligt direktiv 91/493/EEG.%quot%
2) Artikel 2 skall ersättas med följande: %quot%Artikel 2
Fiskeri- och vattenbruksprodukter med ursprung i Nya Zeeland skall uppfylla följande villkor:
1) Varje sändning skall åtföljas av ett numrerat hygienintyg i original, vederbörligen ifyllt, undertecknat och daterat, bestående av ett enda blad, enligt förlagan i bilaga A till detta beslut.
2) Produkterna skall komma från godkända anläggningar, fabriksfartyg, kyl- eller fryshus, eller frysfartyg enligt förteckningen i bilaga B till detta beslut.
3) Varje förpackning skall, med undantag för frysta fiskeriprodukter i bulk avsedda för tillverkning av livsmedelskonserver, i outplånlig skrift vara märkt med ordet 'NYA ZEELAND' och med godkännandenumret för den anläggning, det fabriksfartyg, kyl- eller fryshus, eller frysfartyg där produkterna har sitt ursprung.%quot%
3) Bilaga A skall ersättas med bilagan till detta beslut.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
KOMMISSIONENS DIREKTIV 1999/58/EG
av den 7 juni 1999
om anpassning till den tekniska utvecklingen av rådets direktiv 79/533/EEG om kopplingsanordningen och backväxeln på jordbruks- eller skogsbrukstraktorer med hjul
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 74/150/EEG av den 4 mars 1974 om tillnärmning av medlemsstaternas lagstiftning om typgodkännande av jordbruks- eller skogsbrukstraktorer med hjul(1), senast ändrat genom Europaparlamentets och rådets direktiv 97/54/EG(2), särskilt artikel 11 i detta,
med beaktande av rådets direktiv 79/533/EEG av den 17 maj 1979 om tillnärmning av medlemsstaternas lagstiftning om kopplingsanordningen och backväxeln på jordbruks- eller skogsbrukstraktorer med hjul(3), senast ändrat genom Europaparlamentets och rådets direktiv 97/54/EG, särskilt artikel 4 i detta, och
av följande skäl: (1) För att öka säkerheten förefaller det nödvändigt att närmare fastställa kraven rörande kopplingsanordningarna.
(2) De bestämmelser som föreskrivs i detta direktiv är förenliga med yttrandet från Kommittén för anpassning till teknisk utveckling, inrättad genom artikel 12 i direktiv 74/150/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Punkt 3 i bilaga I till direktiv 79/533/EEG skall ändras på följande sätt:
1. Första stycket skall ersättas med följande text: %quot%Anordningen skall vara utformad som en gaffel. Öppningen i låstappens centrum skall vara 60 mm + 0,5/- 1,5 mm och gaffelns djup från tappens centrum skall vara 62 +- 0,5 mm.%quot%
2. Figuren skall utgå.
Artikel 2
1. Från och med den 1 juli år 2000 får medlemsstaterna inte
- vägra att bevilja EG-typgodkännande eller nationellt typgodkännande, eller vägra att utfärda det dokument som avses i artikel 10.1 tredje strecksatsen i direktiv 74/150/EEG för en viss traktortyp,
- förbjuda att traktorer tas i bruk,
om dessa traktorer uppfyller kraven i direktiv 79/533/EEG, i dess lydelse efter att ha ändrats genom det här direktivet.
2. Från och med den 1 januari 2001 får medlemsstaterna
- inte längre utfärda det dokument som avses i artikel 10.1 tredje strecksatsen i direktiv 74/150/EEG för en traktortyp som inte uppfyller kraven i direktiv 79/533/EEG, i dess lydelse efter att ha ändrats genom det här direktivet.
- vägra bevilja nationellt typgodkännande av en traktortyp som inte uppfyller kraven i direktiv 79/533/EEG, i dess lydelse efter att ha ändrats genom det här direktivet.
Artikel 3
1. Medlemsstaterna skall senast den 30 juni år 2000 sätta i kraft de lagar och andra författningar som behövs för att uppfylla detta direktiv. De skall genast underrätta kommissionen om detta.
När medlemsstaterna antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 4
Detta direktiv träder i kraft den tjugonde dagen efter det att det har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Artikel 5
Detta direktiv riktar sig till medlemsstaterna.
RÅDETS FÖRORDNING (EG) nr 2166/1999
av den 8 oktober 1999
om tillämpningsföreskrifter för förordning (EG) nr 2494/95 i fråga om minimistandarder för hur produkter inom sektorerna hälsa, utbildning och social trygghet skall behandlas i det harmoniserade konsumentprisindexet
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 2494/95 av den 23 oktober 1995 om harmoniserade konsumentprisindex(1), särskilt artikel 4 och artikel 5.3 i denna,
med beaktande av kommissionens förslag,
efter samråd med Europeiska centralbanken(2), och
av följande skäl:
1. Enligt artikel 5.1 b i förordning (EG) nr 2494/95 skall varje medlemsstat sammanställa ett harmoniserat konsumentprisindex (HIKP) från och med indexet för januari 1997.
2. I kommissionens förordning (EG) nr 1749/96(3), definieras HIKP:s omfattning som de varor och tjänster som ingår i hushållens slutliga monetära konsumtionsutgifter. Varor och tjänster från sektorerna hälsa, utbildning och social trygghet ingår i HIKP:s omfattning. De utgifter som de personer har som bor på institutioner ingår i hushållens slutliga monetära konsumtionsutgifter och bör grupperas enligt de COICOP/HIKP-kategorier som fastställs i kommissionens förordning (EG) nr 2214/96(4).
3. Enligt kommissionens förordning (EG) nr 1749/96, särskilt artikel 3 och bilaga Ia i denna, bör en utvidgning av omfattningen inom sektorerna hälsa, utbildning och social trygghet genomföras i december 1999 och bli gällande i och med indexet för januari 2000, varvid metodföreskrifterna för införande bör specificeras i enlighet med förfarandet i artikel 14 inom ramen för förordning (EG) nr 2494/95. Tidsplanen för att införa sjukhusvård och de tjänster inom social trygghet som utförs i hemmet samt i ålderdomshem och handikappboende bör specificeras enligt samma förfarande.
4. Det finns stort utrymme för olikheter i förfarandena för hur varor och tjänster inom sektorerna hälsa, utbildning och social trygghet behandlas i HIKP. En harmoniserad metod för dessa varor och tjänster är nödvändig för att garantera att beräknade HIKP uppfyller de krav på jämförbarhet som föreskrivs i artikel 4 i förordning (EG) nr 2494/95.
5. Behandlingen av varor och tjänster inom sektorerna hälsa, utbildning och social trygghet överensstämmer med definitionerna i Europeiska nationalräkenskapssystemet (ENS) 1995 fastställd genom rådets förordning (EG) nr 2223/96(5).
6. Kommittén för det statistiska programmet har inte yttrat sig inom den tid som dess ordförande fastställt. Enligt förfarandet i artikel 14.2 i förordning (EG) nr 2494/95 skall kommissionen därför utan dröjsmål förelägga rådet ett förslag om vilka åtgärder som skall vidtas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Syfte
Syftet med denna förordning är att fastställa minimistandarder för hur varor och tjänster inom sektorerna hälsa, utbildning och social trygghet skall behandlas i de harmoniserade konsumentprisindexen, nedan kallade HIKP, för att garantera att de är tillförlitliga och relevanta samt uppfyller de krav på jämförbarhet som föreskrivs i artikel 4 i förordning (EG) nr 2494/95.
Artikel 2
Defnition
1. Med återbetalningar avses de betalningar som offentliga organ, socialförsäkringssystem eller hushållens ideella organisationer gör till hushållen som direkt följd av inköp av individuella specificerade varor och tjänster som hushållen ursprungligen betalt för själva.
2. Försäkringsföretags betalningar av ersättningar till hushållen skall inte omfattas av begreppet återbetalningar.
3. Andra betalningar och rabatter till hushållen från offentliga organ, socialförsäkringssystem eller hushållens ideella organisationer i form av bidrag för att minska hushållens utgifter, t.ex. bostadsbidrag till hyresgäster eller betalningar i samband med sjukdom, funktionshinder, vård av äldre släktingar eller studiebidrag till studerande, skall anses vara sociala förmåner i form av kontantersättningar. De skall behandlas som överföringar till hushållen och skall inte utgöra en återbetalning.
Artikel 3
Omfattning
1. De varor och tjänster inom sektorerna hälsa, utbildning och social trygghet som räknas till hushållens slutliga monetära konsumtionsutgifter skall omfattas av HIKP och grupperas enligt de COICOP/HIKP-kategorier som föreskrivs i kommissionens förordning (EG) nr 2214/96.
2. Alla leverantörer av varor och tjänster inom sektorerna hälsa, utbildning och social trygghet, såsom statliga och privata institutioner, hushållens ideella organisationer eller egenföretagare, skall omfattas av HIKP oberoende av deras ställning. Detta utesluter enskilda eller grupper av enskilda som producerar varor och icke-finansiella tjänster uteslutande för egen slutlig förbrukning.
3. I enlighet med COICOP/HIKP omfattar utbildning (huvudgrupp 10) endast utbildningstjänster. Om ett totalpris debiteras för utbildningstjänster i vilket ingår läromedel eller stödtjänster till utbildning, skall de olika komponenterna delas upp och föras upp i de berörda undergrupperna i COICOP/HIKP. Om ett totalpris inte kan delas upp i fråga om priserna på de berörda komponenterna, skall totalpriset föras upp under huvudgrupp 10 i COICOP/HIKP.
4. Gränsfall mellan förskoleutbildning och barnomsorg, såsom barnskötare, daghem och lekskolor, skall föras upp i huvudgrupp 10 i COICOP/HIKP, om barnet då det inskolas är över tre år och om verksamheten består i organiserad undervisning i en skolliknande miljö och där syftet är att överbrygga steget mellan hemmet och skolan. Om huvudsyftet däremot inte är av pedagogisk art, utan att tillhandahålla barnomsorg skall den berörda tjänsten föras upp i undergrupp 12.4.0 i COICOP/HIKP.
5. Om det vid sjukhusvård tillhandahålls andra varor och tjänster för intagna patienter än de bastjänster som definieras i COICOP/HIKP 06.3 och dessa debiteras separat, skall de inte föras upp i undergrupp 06.3.0, utan i de berörda undergrupperna i COICOP/HIKP.
Artikel 4
Priser
1. De av HIKP:s delindex som berörs skall beräknas med hjälp av en formel som överensstämmer med den formel av Laspeyres-typ som används för andra delindex. De skall spegla prisförändringen på grundval av hur utgifterna ändras vid ett oförändrat konsumtionsmönster för hushållen och en oförändrad sammansättning av konsumentpopulationen under bas- eller referensperioden.
2. a) De anskaffningspriser på varor och tjänster inom sektorerna hälsa, utbildning och social trygghet som skall användas för HIKP skall vara de belopp som konsumenterna betalar med avdrag för återbetalningar.
b) De förändringar i anskaffningspriserna som speglar förändringar i de regler som fastställer dem, skall framgå som prisförändringar i HIKP.
c) Om anskaffningspriserna är knutna till ett index skall ändringar som följer av förändringar i indexet framgå som prisförändringar i HIKP.
d) Förändringar i anskaffningspriser som följer av förändringar i konsumenternas inkomster skall framgå som prisförändringar i HIKP.
3. Om det rör sig om kvalitetsförändringar, skall priserna behandlas enligt de regler som tillämpas i samband med ändringar i specifikationen, särskilt de som gäller kvalitetsjusteringar i enlighet med artikel 5 i kommissionens förordning (EG) nr 1749/96.
4. Om konsumenterna kostnadsfritt har erhållit en vara eller tjänst inom sektorerna hälsa, utbildning och social trygghet och man därefter tar ut ett faktiskt pris, skall förändringen från nollpris till det faktiska priset, och omvänt, framgå i HIKP.
5. Om varor och tjänster inom sektorerna hälsa, utbildning och social trygghet har tillhandahållits konsumenterna utan kostnad tillsammans med andra varor och tjänster och man därefter tar ut ett pris för dessa separat, skall denna förändring framgå i HIKP.
6. Om det är relevant skall förfarandet i artikel 5 i kommissionens förordning (EG) nr 2646/98(6) avseende tariffer tillämpas i tillämpliga delar.
Artikel 5
Grundläggande uppgifter
De grundläggande uppgifterna skall utgöras av alla anskaffningspriser på varor och tjänster inom sektorerna hälsa, utbildning och social trygghet och deras komponenter, tillsammans med korrigeringskoefficienter som speglar nivå, tidpunkt och struktur på konsumtionen av sådana varor och tjänster, enligt de socioekonomiska karakteristika som är prisbestämmande.
Artikel 6
Uppgiftskällor
1. Medlemsstaterna skall beräkna berörda HIKP-delindex utifrån de grundläggande uppgifterna såsom de definieras i artikel 5.
2. De statistiska enheter, t.ex. statliga organ, socialförsäkringssystem eller hushållens ideella organisationer, som av medlemsstaterna uppmanas att samarbeta vid insamlingen eller tillhandahållandet av de grundläggande uppgifterna skall lämna sann och fullständig information vid den tidpunkt då den begärs, och de organisationer och institutioner som ansvarar för att sammanställa officiell statistik skall på begäran erhålla uppgifter på den detaljnivå som krävs för att utvärdera efterlevnaden av jämförbarhetskraven och kvaliteten på HIKP:s delindex.
Artikel 7
Jämförbarhet
HIKP som konstrueras enligt förfarandena i artiklarna 4 och 5 i denna förordning eller enligt andra förfaranden, som inte leder till ett index som systematiskt avviker med mer än i genomsnitt en tiondels procentenhet för ett år i förhållande till föregående års index som sammanställdes enligt samma förfarande skall anses vara jämförbara.
Artikel 8
Kvalitetskontrol
1. Medlemsstaterna skall innan sådana förfaranden tillämpas förse kommissionen (Eurostat) med de uppgifter om de förfaranden som utarbetats för behandling av varor och tjänster inom sektorerna hälsa, utbildning och social trygghet, om dessa förfaranden avviker från dem som anges i artiklarna 4 och 5 i denna förordning.
2. Medlemsstaterna skall på begäran förse kommissionen (Eurostat) med de uppgifter som är nödvändiga för att bedöma hur de förfaranden som fastställs i artiklarna 4 och 5 i denna förordning fungerar. Resultatet av denna bedömning skall ingå i de rapporter som kommissionen skall överlämna till rådet i enlighet med artikel 2 i rådets förordning (EG) nr 1687/98 och med artikel 2 i rådets förordning (EG) nr 1688/98.
Artikel 9
Genomförande
Medlemsstaterna skall genomföra bestämmelserna i denna förordning i december 1999 och de skall bli gällande i och med indexet för januari 2000, med undantag för följande som skall genomföras i december 2000 och bli gällande i och med indexet för januari 2001:
a) Sjukhusvård (COICOP/HIKP 06.3). b) Tjänster inom social trygghet som tillhandahålls i hemmet, t.ex. städning, måltider, transporter av funktionshindrade (ingår i COICOP/HIKP 12.4.0).
c) Ålderdomshem och handikappboende (ingår i COICOP/HIKP 12.4.0).
Artikel 10
Ikraftträdande
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
RÅDETS FÖRORDNING (EG) nr 2791/1999
av den 16 december 1999
om att upprätta vissa kontrollåtgärder som skall tillämpas i det område som avses i konventionen om framtida multilateralt samarbete om fisket i Nordostatlanten
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 37 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(1), och
av följande skäl:
1. Konventionen om framtida multilateralt samarbete om fisket i Nordostatlanten, nedan kallad %quot%NEAFC-konventionen%quot% godkändes genom beslut 81/608/EEG av den 13 juli 1981(2) och trädde i kraft den 17 mars 1982.
2. Genom NEAFC-konventionen upprättas den ram som behövs för ett multilateralt samarbete på området för ett rationellt bevarande och en rationell förvaltning av fiskeresurserna i det område som definieras i konventionen.
3. Vid sitt 17:e årsmöte den 17-20 november 1998 antog den nordostatlantiska fiskerikommissionen två rekommendationer, i den ena upprättas en tvångs- och kontrollplan för de fiskefartyg som bedriver fiske i områdena utanför gränserna för den nationella jurisdiktionen för avtalsslutande parterna i konventionsområdet (nedan kallat planen), och i den andra upprättas ett program (nedan kallat programmet) med syftet att få icke avtalsslutande parters fartyg att följa dessa rekommendationer för att se till att NEAFC:s bevarande- och förvaltningsåtgärder till fullo iakttas.
4. I planen föreskrivs kontrollåtgärder för fartyg som för en avtalsslutande parts flagg och som bedriver fiske i NEAFC-området samt en plan för inspektion till havs med förfaranden för inspektion och övervakning samt överträdelseförfaranden som skall genomföras av avtalsslutande parterna.
5. I programmet föreskrivs att det är obligatoriskt att inspektera icke-avtalsslutande parters fartyg om dessa fartyg frivilligt lägger till i en hamn som tillhör en avtalsslutande part; landning och omlastning skall förbjudas om det under en sådan inspektion visar sig att fångst har gjorts i strid med de bevarandeåtgärder som NEAFC har antagit.
6. I enlighet med artiklarna 12 och 15 i NEAFC-konventionen träder dessa rekommendationer i kraft den 1 juli 1999 och blir obligatoriska för avtalsslutande parterna. Gemenskapen bör tillämpa dem.
7. För att göra det möjligt att övervaka gemenskapens fiske i det område som NEAFC råder över, samtidigt som de kontrollbestämmelser iakttas som föreskrivs i förordning (EEG) nr 2847/93 av den 12 oktober 1993 om införande av ett kontrollsystem för den gemensamma fiskeripolitiken(3), bör vissa särskilda kontrollåtgärder fastställas för bedrivandet av fiske, för märkning och dokumentation av fartyg och fiskeredskap, för registrering och meddelande om fångst samt för omlastning.
8. I artikel 2.3 i förordning (EEG) nr 2847/93 föreskrivs att medlemsstaterna, utanför gemenskapens fiskeområde, skall se till att deras fartyg är föremål för lämplig övervakning och, om det finns åligganden från gemenskapen i detta avseende, inspektioner och övervakning på ett sätt som garanterar att den gemenskapslagstiftning som gäller för dessa vatten följs. Det bör därför föreskrivas att de medlemsstater vars fiskefartyg har tillåtelse att fiska i NEAFC-området skall utse inspektörer som skall utföra kontroll och övervakning enligt planen, samt tillhandahålla den utrustning som behövs för inspektionen.
9. För att se till att fiskeaktiviteterna i NEAFC-området övervakas, måste medlemsstaterna samarbeta med varandra och med kommissionen vid tillämpningen av planen.
10. Medlemsstaterna har ansvar för att se till att deras inspektörer följer de inspektionsförfaranden som har upprättats av NEAFC.
11. Befälhavarna på gemenskapens fartyg bör samarbeta med inspektören när deras fartyg inspekteras enligt de förfaranden som fastställs i denna förordning.
12. Det bör fastställas förfaranden som skall följas vid misstanke om överträdelser och i synnerhet allvarliga överträdelser. För detta ändamål bör det upprättas en förteckning över vad som skall anses som allvarliga överträdelser.
13. Det bör fastställas tillämpningsföreskrifter för programmet i gemenskapen.
14. I kraft av fördraget bör inre farvatten och hamnar kontrolleras av medlemsstaterna. När det gäller tillträde till hamnanläggningar i gemenskapen för icke avtalsslutande parter som har påträffats verksamma i NEAFC-området, bör enhetliga tilläggsåtgärder vidtas på gemenskapsnivå för att skapa bestämmelser för sådana fartygs verksamhet i gemenskapens hamnar på så sätt att NEAFC:s åtgärder förblir effektiva.
15. Det bör fastställas ett förfarande för att anta tillämpningsföreskrifter för planen.
16. De åtgärder som krävs för att genomföra den här förordningen bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(4).
17. I syfte att uppnå erfarenhet inför den slutgiltiga fördelning av uppgifterna som skall genomföras är det lämpligt att vissa bestämmelser om inspektion och kontroll som skall genomföras i samarbete mellan medlemsstaterna och kommissionen tillämpas under en begränsad period i väntan på ett beslut om den slutgiltiga ordningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Syfte
I denna förordning fastställs allmänna principer och villkor för gemenskapens tillämpning av
a) kontroll- och genomdrivandeplanen för fartyg som bedriver fiske i områden utanför nationell jurisdiktion i NEAFC-området,
b) programmet som främjar att icke avtalsslutande parters fartyg följer mot NEAFC:s rekommendationer.
Artikel 2
Definitioner
I denna förordning skall följande definitioner gälla:
1. kontrollområde: de vatten inom konventionens område som definieras i artikel 1.1 i NEAFC-konventionen och som ligger utanför vattnen under NEAFC-parternas jurisdiktion.
2. fisktillgångar: de fisktillgångar som anges i artikel 1.2 i NEAFC-konventionen.
3. reglerade tillgångar: de fisketillgångar som är föremål för rekommendationer enligt konventionen och som förtecknas i bilagan. Bilagan får ändras enligt förfarandet i artikel 29.2.
4. fiskeverksamhet: fiske, bearbetning av fisk, omlastning av fisk eller fiskeprodukter och all annan verksamhet som syftar till fiske eller har anknytning till fiske i kontrollområdet.
5. NEAFC-inspektör: en inspektör som utsetts för planen av en avtalsslutande part till NEAFC.
6. bordning: NEAFC-inspektörer går ombord på ett fiskefartyg för att genomföra en inspektion.
7. överträdelse: ett fiskefartygs alla handlingar eller underlåtenhet som ger starka skäl att misstänka att ett brott har begåtts mot bestämmelserna i denna förordning eller varje annan förordning som genomför NEAFC-rekommendationerna, och som noterats i en inspektionsrapport enligt planen.
8. allvarlig överträdelse innebär:
a) att fiska utan giltigt tillstånd från flaggstaten,
b) att fiska utan tilldelad kvot eller efter det att kvoten har uttömts,
c) att använda förbjudna fiskeredskap,
d) att göra en grovt felaktig anteckning om fångst,
e) att vid upprepade tillfällen underlåta att lämna uppgifter om förflyttning och fångst,
f) att hindra en inspektör ifrån att fullgöra sina uppgifter,
g) att genomföra riktat fiske mot ett bestånd som omfattas av ett moratorium eller ett fiskeförbud,
h) att förfalska eller dölja ett fiskefartygs märkning, identitet eller registrering,
i) att dölja, förändra eller göra sig av med bevis som behövs vid en undersökning, eller
j) att genom flera överträdelser visa allvarling brist på respekt för bevarande- och förvaltningsåtgärder.
9. vederbörligen godkänd inspektör: en NEAFC-inspektör som vederbörligen godkänts av den medlemsstat vars flagg det fartyg för som misstänks ha begått en allvarlig överträdelse.
10. icke avtalsslutande parts fartyg: ett fartyg som har setts och meddelats vara sysselsatt med fiskeverksamhet i NEAFC-området och
i) som för en flagg som tillhör en stat som inte är avtalsslutande part till NEAFC-konventionen, eller
ii) det finns rimliga skäl att misstänka att det saknar nationalitet.
AVDELNING I
GENOMFÖRANDE AV NEAFC:s KONTROLLPLAN
Artikel 3
Tillämpningsområde
1. Denna avdelning är tillämplig på alla gemenskapens fiskefartyg som används eller avses användas i avsikt att bedriva kommersiell fiskeverksamhet inriktad på fisktillgångarna i kontrollområdet.
2. De gemenskapsfartyg som bedriver fiske i kontrollområdet och som bevarar fisk ombord från detta område skall göra detta i enlighet med målen och principerna i NEAFC-konventionen.
KAPITEL 1
KONTROLLÅTGÄRDER
Artikel 4
Gemenskapens deltagande
1. Endast de av gemenskapsfiskefartygen som innehar ett särskilt fisketillstånd som utfärdats av den medlemsstat vars flagg de för har tillåtelse att, på de villkor som anges i tillståndet, fiska, bevara ombord, lasta om och landa fisktillgångar från kontrollområdet.
2. Medlemsstaterna skall på elektronisk väg till kommissionen översända en förteckning över alla fartyg som för deras flagg och är registrerade i gemenskapen och som har tillåtelse att fiska i kontrollområdet, särskilt de fartyg som har tillåtelse att fiska direkt efter en eller flera arter för vilka särskilda bestämmelser gäller samt eventuella ändringar i förteckningen. Detta skall ske senast den 15 december varje år eller minst 5 dagar innan fartyget ankommer till kontrollområdet. Kommissionen skall utan dröjsmål översända dessa uppgifter till NEAFC:s sekretariat.
3. Beslut om hur den förteckning som avses i punkt 2 samt specifikationerna skall översändas skall fattas i enlighet med förfarandet i artikel 29.2.
Artikel 5
Registrering av fångster och fiskeansträngning
1. Utöver de uppgifter som anges i artikel 6 i förordning (EEG) nr 2847/93 skall befälhavarna på gemenskapens fiskefartyg i sin loggbok skriva in när de ankommer till och lämnar kontrollområdet.
2. Befälhavarna på gemenskapens fiskefartyg skall, för fångst av de reglerade arter som anges i bilagan, bearbetade eller frysta, föra
a) en bearbetningsjournal som anger, per art och bearbetad produkt, den samlade produktionen, eller
b) en lagringsplan per art över bearbetade produkter, med uppgifter om lagringsplats för bearbetade produkter och för produkter i lastrummet.
3. Tillämpningsföreskrifter för denna artikel skall antas i enlighet med förfarandet i artikel 29.2.
Artikel 6
Fångstrapport för reglerade resurser
1. Befälhavarna för gemenskapens fiskefartyg skall till de behöriga myndigheterna i deras flaggmedlemsstat översända en rapport med namnet %quot%fångstrapport%quot% inom den tid som anges i andra stycket.
En fångstrapport för reglerade resurser skall omfatta följande:
a) De kvantiteter som bevaras ombord när befälhavarna på gemenskapens fiskefartyg ankommer till kontrollområdet. Rapporten skall sändas inom 12 timmar och minst 6 timmar före ankomsten till kontrollområdet.
b) Veckofångsten. En sådan rapport måste första gången översändas senast i slutet av den sjunde dagen efter ankomsten till kontrollområdet eller, om fångstresan varar längre än sju dagar, senast på måndagen, för de fångster som gjorts i kontrollområdet under föregående vecka fram till midnatt på söndagen.
c) De kvantiteter som finns ombord när fartyget lämnar kontrollområdet. Rapporten skall sändas tidigast 8 timmar och senast 6 timmar i förväg varje gång kontrollområdet lämnas. Den skall om det är lämpligt innehålla uppgifter om antal fiskedagar och fångster i kontrollområdet.
d) De kvantiteter som lastats och lossats vid varje omlastning av fisk under den period som fartyget stannar i kontrollområdet. Meddelandet skall sändas inom 24 timmar efter omlastningen.
2. Varje medlemsstat skall omedelbart när den har mottagit fångstrapporterna elektroniskt översända dessa till NEAFC:s sekretariat.
3. Fångstrapporterna skall översändas till medlemsstaternas behöriga myndigheter för vidarebefordran till NEAFC:s sekretariat(5).
4. Medlemsstaterna i den databas som anges i artikel 19.2 i förordning (EEG) nr 2847/93 skall registrera uppgifterna i fångstrapporterna.
5. Närmare bestämmelser för tillämpningen av denna artikel, särskilt om den form och de specifikationer för överföringen som avses i punkt 3, skall fastställas enligt förfarandet i artikel 29.2.
Artikel 7
Global rapportering om fångst och fiskeansträngning
1. Medlemsstaterna skall före den 15 varje månad elektroniskt översända uppgifter till kommissionen om de resursmängder som avses i punkt 3 och som har fångats i kontrollområdet och landats eller omlastats under föregående månad.
2. Utan hinder av artikel 3.2 skall denna artikel även tillämpas på reglerade resurser som har fångats i den del av konventionsområdet som står under medlemsstaternas jurisdiktion utan att det påverkar tillämpningen av artikel 15 i förordning (EEG) nr 2847/93.
3. Beslut om den förteckning över resurser som avses i punkt 1 samt formen för översändandet av uppgifter skall antas i enlighet med förfarandet i artikel 29.2.
Artikel 8 (6)
Det satellitbaserade kontrollsystemet
Medlemsstaterna skall se till att de uppgifter som erhålls via det satellitbaserade kontrollsystemet (VMS) om fartyg som för deras flagg och som fiskar i kontrollområdet översänds elektroniskt till NEAFC:s sekretariat i realtid, i den form och med de specifikationer som anges enligt förfarandet i artikel 29.2.
Artikel 9
Omlastning
Gemenskapens fiskefartyg får endast lasta om i kontrollområdet om de har satt tillåtelse i förväg av de behöriga myndigheterna i den medlemsstat vars flagg de för och där de är registrerade.
KAPITEL 2
INSPEKTIONSFÖRFARANDEN
Artikel 10 (7)
Allmänna bestämmelser för inspektion och kontroll
1. De medlemsstater vars fiskefartyg har tillåtelse att fiska i kontrollområdet skall utse inspektörer för genomförande av kontroll och inspektion i enlighet med planen.
2. Varje medlemsstat skall vidta de åtgärder som krävs för att NEAFC:s inspektörer skall kunna genomföra sina inspektioner ombord på de fartyg som för dess flagg.
3. Varje medlemsstat skall se till att de inspektioner som dess inspektörer genomför, görs på ett icke-diskriminerande sätt och i enlighet med planen. Antalet inspektioner skall vara baserat på hur stor del av de avtalsslutande parternas flotta som befinner sig i kontrollområdet och med hänsyn till hur lång tid som dessa fartyg funnits där.
4. Kommissionen får utse gemenskapsinspektörer för planen.
Artikel 11 (8)
Inspektionsutrustning
1. Medlemsstaterna, eller kommissionen i enlighet med artikel 10.4, skall ställa den utrustning som behövs till förfogande för sina inspektörer, så att övervaknings- och inspektionsuppdraget kan genomföras. För detta ändamål skall de tilldela inspektionsfartyg och luftfartyg till planen.
2. Kommissionen skall samordna gemenskapens övervaknings- och inspektionsverksamhet. I detta syfte får kommissionen, i samförstånd med de berörda medlemsstaterna, upprätta gemensamma operationella övervaknings- och inspektionsprogram som gör det möjligt för gemenskapen att fullgöra sina skyldigheter enligt planen. De medlemsstater vars fartyg bedriver fiske med reglerade tillgångar skall vidta nödvändiga åtgärder för att underlätta genomförandet av dessa program, särskilt när det gäller nödvändiga mänskliga och materiella resurser samt de perioder och områden där dessa skall tas i bruk.
3. Medlemsstaterna skall senast den 1 januari 2000 meddela kommissionen namn på de inspektörer och inspektionsfartyg samt de luftfartyg som de avser skall knytas till planen under följande år. På grundval av dessa uppgifter skall kommissionen i samarbete med medlemsstaterna upprätta en verksamhetsplan för gemenskapens deltagande i planen under kalenderåret i fråga och kommissionen skall sedan skicka denna till NEAFC-sekretariatet och till medlemsstaterna.
4. När mer än tio av gemenskapens fiskefartyg samtidigt bedriver fiske riktat mot reglerade tillgångar i kontrollområdet skall kommissionen, vid framtagandet av operationella övervaknings- och inspektionsprogram, se till att en medlemsstats inspektionsfartyg finns i området eller att ett avtal har slutits med en annan avtalsslutande part om att ett inspektionsfartyg skall finnas på plats.
5. Medlemsstaterna skall se till att alla fartyg som omfattas av planen och som har inspektörer ombord samt eventuella hjälpfartyg hissar en särskild flagga eller vimpel för att visa att inspektören genomför en inspektion inom ramen för planen. Luftfartyg som omfattas av planen skall ha den internationella radioanropssignalen tydligt målad och väl synlig. Den särskilda flaggan eller vimpeln skall utformas enligt förfarandet i artikel 29.2.
6. Medlemsstaterna skall underrätta kommissionen elektroniskt och i enlighet med förfarandet i artikel 29.2 om de datum och tider då inspektionsfartygens och luftfartygens verksamhet börjar och slutar.
Artikel 12
NEAFC-inspektörer
1. Medlemsstaterna eller, i enlighet med artikel 10.4, kommissionen skall utfärda ett särskilt identitetskort för varje inspektör. Varje inspektör skall medföra detta när han går ombord på ett fiskefartyg. Det särskilda identitetskortets form skall fastställas enligt förfarandet i artikel 29.2.
2. Medlemsstaterna och kommissionen skall se till att inspektörerna uppfyller sitt uppdrag enligt bestämmelserna i planen. Inspektörerna fortsätter att lyda under sina behöriga myndigheter och ansvarar inför dem.
Artikel 13
Övervakningsförfarande
1. NEAFC-inspektörerna skall från ett fartyg eller ett luftfartyg som omfattas av planen genomföra kontroller baserade på samtliga observationer av fiskefartygen. De skall notera sina observationer i en rapport vars form skall beslutas i enlighet med förfarandet i artikel 29.2 och som skall översändas till den behöriga myndigheten.
2. Medlemsstaterna skall utan dröjsmål på elektronisk väg översända observationsrapporten till den flaggstat som fartyget i fråga hör till eller till de myndigheter som denna stat utsett och anmält till NEAFC-sekretariatet, till NEAFC-sekretariatet och till kommissionen. Medlemsstaterna skall också på begäran skicka originalet till varje observationsrapport och fotografier till den flaggstat som fartyget i fråga tillhör.
Artikel 14
Inspektionsförfarande
1. Medlemsstaterna och kommissionen skall se till att NEAFC-inspektörerna:
a) inte bordar ett fartyg utan föregående anmälan via radio till fartyget eller utan att fartyget fått lämplig signal enligt det internationella signalsystemet med uppgift om inspektionsgruppens identitet,
b) inte beordrar det fartyg som bordas att stanna eller göra manövrar under pågående fiskeverksamhet, eller när fiskeredskap sätts ut eller tas upp. Inspektörerna får dock beordra fartyget att avbryta eller vänta med att sätta ut redskapen till dess att fartyget har bordats, men detta får under inga omständigheter ske senare än 30 minuter efter det att signalen har mottagits,
c) ser till att inspektionen inte pågår längre tid än fyra timmar eller efter det att gamen och fångsten har tagits upp och inspekterats om detta tar längre tid. Om en överträdelse upptäcks får inspektörerna stanna ombord under den tid som krävs för att genomföra uppgifterna enligt artikel 16.1.b. Under särskilda omständigheter, med hänsyn till fartygets storlek och kvantiteterna ombord, får dock inspektionen pågå längre än vad som anges ovan. I detta fall skall inspektörerna inte stanna längre ombord än den tid det tar att genomföra inspektionen. Orsaken till att en inspektion tagit längre tid än normalt skall anges i inspektionsrapporten,
d) under bordningen och inspektionen inte hindrar befälhavaren från att kommunicera med myndigheterna i flaggstaten,
e) manövrerar på ett säkert avstånd från fiskefartyget i enlighet med gott sjömanskap,
f) undviker våld utom om det är absolut nödvändigt för att garantera inspektörernas säkerhet. Inspektörerna får inte medföra skjutvapen ombord på fiskefartyget under inspektion,
g) genomför inspektionen med så liten störning som möjligt för fartyg, fiskeverksamheten och fångsten,
h) upprättar en inspektionsrapport i enlighet med de bestämmelser som antagits enligt förfarandet i artikel 29.2 och skickar den till deras myndigheter.
2. Inspektörerna skall ha befogenhet att undersöka alla relevanta områden, fiskefartygets däck och utrymmen, fångster (bearbetade eller obearbetade), nät och andra redskap, utrustning samt alla relevanta dokument som behövs för att kontrollera att NEAFC:s bevarandeåtgärder har iakttagits samt att förhöra befälhavaren eller en person som har utsetts av befälhavaren.
3. Vid inspektionen har inspektörerna rätt att begära hjälp från befälhavaren. Befälhavaren har rätt att kommentera inspektionsrapporten som skall undertecknas av inspektörerna i slutet av inspektionen. Befälhavaren på fiskefartyget skall få en kopia av inspektionsrapporten.
4. Medlemsstaterna skall se till att inspektionsgruppen skall bestå av högst två NEAFC-inspektörer.
Artikel 15
Befälhavarnas skyldigheter vid inspektion
Befälhavaren på ett av gemenskapens fiskefartyg som blir föremål för bordning och inspektion skall
a) bidra till att bordningen sker effektivt och säkert,
b) samarbeta och ge stöd vid en inspektion av ett fiskefartyg som genomförs i enlighet med förfarandena i denna förordning och får inte hindra inspektörerna att fullgöra sitt uppdrag, hota eller störa dem i arbetet, utan se till att deras säkerhet är garanterad,
c) göra det möjligt för inspektörerna att kommunicera med myndigheterna i flaggstaten och i den stat som genomför inspektionen,
d) ge tillträde till relevanta områden, däck, utrymmen, fångster (bearbetade eller obearbetade), nät och andra redskap, utrustning och alla relevanta dokument,
e) erbjuda inspektörerna rimliga arbetsförhållanden, vid behov även kost och logi om de förblir ombord på fartyget i enlighet med artikel 18.3,
f) göra det möjligt för inspektören att lämna fartyget under säkra förhållanden.
Artikel 16
Förfarande vid överträdelse
1. Om NEAFC-inspektörer har starka skäl att tro att ett fiskefartyg bedriver fiske i strid med de bevarandeåtgärder som NEAFC har antagit skall
a) en anteckning om överträdelse införas i inspektionsrapporten,
b) alla nödvändiga åtgärder vidtas för att säkra och bevara bevisningen. Ett identifieringsmärke skall noga fästas på varje del av de fiskeredskap som vid inspektion misstänks ha använts i strid med bestämmelserna,
c) kontakt omedelbart tas med en inspektör eller den utsedda myndigheten i den stat vars flagg det inspekterade fartyget för,
d) inspektionsrapporten utan dröjsmål skickas till deras myndigheter.
2. Den medlemsstat som genomför inspektionen eller, i förekommande fall, kommissionen skall under den arbetsdag som följer efter den dag då inspektionen påbörjades om möjligt meddela det inspekterade fartygets flaggstat och kommissionen uppgifter om den överträdelse som det inspekterade fartyget har begått.
3. Den medlemsstat som genomför inspektionen skall översända inspektionsrapporten i original med alla underlag till kommissionen som skall vidarebefordra den till behöriga myndigheter i den stat vars flagg det inspekterade fartyget för samt en kopia till NEAFC-sekretariatet.
Artikel 17
Uppföljning av överträdelser
1. Om en medlemsstat får en anmälan från en annan avtalsslutande part eller från en annan medlemsstat om en överträdelse som begåtts av ett fartyg som för den medlemsstatens flagg, skall medlemsstaten snabbt vidta åtgärder i enlighet med nationell rätt för att kunna ta emot och undersöka bevisen samt genomföra de undersökningar som behövs för de åtgärder som skall vidtas till följd av överträdelser samt, om möjligt, inspektera fartyget.
2. Medlemsstaterna skall utse de myndigheter som skall ta emot bevis på överträdelse och meddela kommissionen denna myndighets adress.
Artikel 18
Särskilt förfarande vid allvarliga överträdelse
1. Om en NEAFC-inspektör anser sig ha starka skäl att tro att ett fiskefartyg har begått en allvarlig överträdelse skall han utan dröjsmål underrätta flaggstaten, de egna myndigheterna och NEAFC-sekretariatet.
2. Inspektören skall vidta alla nödvändiga åtgärder för att se till att bevisningen säkras och bevaras utan att fiskeverksamheten störs mer än absolut nödvändigt.
3. Inspektören får stanna ombord på fartyget så länge som behövs för att ge den behörige inspektören upplysningar om överträdelsen eller fram till det att flaggstaten begär att inspektören skall lämna fiskefartyget.
4. Den medlemsstat som genomför inspektionen skall med samtycke av den stat som fartyget tillhör besluta om inspektören skall stanna ombord under fartygets omdirigering. Den medlemsstat som genomför inspektionen skall också besluta om en NEAFC-inspektör skall närvara vid en grundligare inspektion av fartyget i hamn. Medlemsstaten skall utan dröjsmål underrätta kommissionen om de beslut som fattats i enlighet med denna punkt.
Artikel 19
Uppföljning av allvarliga överträdelser
1. Om de behöriga myndigheterna i en flaggmedlemsstat får information av en NEAFC-inspektör om misstanke om att en allvarlig överträdelse har begåtts av ett fiskefartyg som för medlemsstatens flagg eller om kommissionen får sådan information, skall de behöriga myndigheterna och kommissionen utan dröjsmål underrätta varandra om detta.
2. Efter att ha mottagit den information som anges i punkt 1 skall flaggmedlemsstaten se till att fartyget inspekteras inom 72 timmar av en godkänd inspektör.
3. Den godkända inspektören skall gå ombord på fiskefartyget i fråga och granska bevisen på den misstänkta allvarliga överträdelsen som konstaterats av NEAFC-inspektören, och snarast möjligt översända resultaten av granskningen till den behöriga myndigheten i flaggmedlemsstaten och till kommissionen.
4. Efter anmälan av resultaten och om överträdelsen i fråga visat sig vara allvarlig skall den behöriga myndigheten i det inspekterade fartygets flaggmedlemsstat, inom 24 timmar beordra eller utse en godkänd inspektör för att beordra fartyget att gå mot en utsedd hamn, om situationen motiverar detta.
Vid omdirigering skall den godkände inspektören vidta alla åtgärder som behövs för att säkra och bevara bevisningen.
5. Vid ankomsten till den hamn dit fartyget har omdirigerats skall det inspekteras grundligt av flaggmedlemsstatens myndigheter, i närvaro av en NEAFC-inspektör från någon annan avtalsslutande part som vill delta i inspektionen.
Flaggmedlemsstaten skall utan dröjsmål underrätta kommissionen om resultaten av den grundliga inspektionen och om de åtgärder som den har vidtagit till följd av överträdelsen.
6. Om flaggmedlemsstatens behöriga myndighet inte omdirigerar fartyget till en hamn, skall orsakerna till detta utan dröjsmål meddelas kommissionen. Kommissionen skall så snart som möjligt underrätta NEAFC-sekretariatet om beslutet och dess orsaker.
7. Tillämpningsföreskrifter till denna artikel skall fastställas enligt förfarandet i artikel 29.2.
Artikel 20
Behandling av inspektionsrapporterna
1. Medlemsstaterna skall lägga samma vikt vid rapporter som sammanställts av NEAFC-inspektörer från andra avtalsslutande parter och andra medlemsstater som vid de egna inspektörernas rapporter.
2. Medlemsstaterna skall samarbeta med de berörda avtalsslutande parterna för att underlätta rättsliga eller andra förfaranden i enlighet med deras nationella rätt till följd av en rapport från en inspektor i enlighet med planen.
Artikel 21
Rapport om överträdelser
1. Samtliga medlemsstater skall före den 15 september varje år skicka en rapport till kommissionen för det föregående kalenderåret med information om utvecklingen i de ärenden som hänför sig till anmälda överträdelser av NEAFC:s bevarandeåtgärder. Dessa överträdelser skall förtecknas årligen fram tills dess att ett slutgiltigt beslut har fattats i enlighet med relevanta bestämmelser i nationell rätt.
2. Rapporten skall innehålla detaljer av de framsteg som görs i förfarandena (vilande ärende, åtal väckt, under utredning, osv.), påföljder eller böter beskrivna i särskilda termer (dvs. bötesbelopp, värdet på beslagtagen fisk och/eller redskap, skriftlig varning, osv.) och innefatta en förklaring i de fall ingen åtgärd har vidtagits.
Artikel 22
Rapport om inspektionsverksamheten
Medlemsstaterna skall senast den 15 september varje år, angående det föregående kalenderåret, underrätta kommissionen om följande:
a) Antal genomförda inspektioner inom ramen för planen med angivande av antal inspektioner på varje avtalsslutande parts fartyg samt, vid överträdelse, datum och position för inspektionsfartyget i fråga och uppgift om arten av den överträdelse som misstänks.
b) Antal timmar med flygövervakning, antal observationer och antal övervakningsrapporter som har utarbetats och uppföljningen av dessa rapporter.
AVDELNING II
GENOMFÖRANDE AV PROGRAMMET FÖR ATT FRÄMJA EFTERLEVNAD AV FARTYG FRÅN ICKE AVTALSSLUTANDE PARTER
Artikel 23
Översändande av observationsrapport
1. När en medlemsstat har mottagit en observationsrapport från en av sina NEAFC-inspektörer om en icke avtalsslutande parts fartyg, skall medlemsstaten utan dröjsmål översända denna information till NEAFC-sekretariatet och till kommissionen samt, om möjligt, till fartyget med information om att uppgifterna skall översändas till fartygets flaggstat.
2. Kommissionen skall utan dröjsmål underrätta alla medlemsstater om varje observationsrapport som har mottagits genom anmälan till NEAFC-sekretariatet eller till en annan avtalsslutande part.
Artikel 24
Omlastning
Det är förbjudet för gemenskapens fiskefartyg att ta emot omlastningar av fisk från en icke avtalsslutande parts fartyg.
Artikel 25
Kontroll av fiskeverksamheten på fartyg som för icke avtalsslutande parts flagg
1. Medlemsstaterna skall se till att alla icke avtalsslutande parters fartyg som anlöper en hamn som utsetts i enlighet med artikel 28e.2 i förordning (EEG) nr 2847/93 inspekteras av deras behöriga myndigheter. Så länge som inspektionen pågår är det förbjudet att landa eller omlasta fartygets fångst.
2. Om de behöriga myndigheterna i slutet av en sådan inspektion finner att det ombord på en icke avtalsslutande parts fartyg finns tillgångar som omfattas av en NEAFC-rekommendation som överförts till gemenskapslagstiftningen skall medlemsstaten i fråga förbjuda landning och omlastning.
3. Detta förbud gäller dock inte om det inspekterade fartygets befälhavare eller dennes representant på ett tillfredsställande sätt för den berörda medlemsstatens behöriga myndigheter kan påvisa att:
a) den fångst som finns ombord har fångats utanför kontrollområdet, eller
b) den fångst som finns ombord har fångats i enlighet med gemenskapens bevarandeåtgärder.
Artikel 26
Uppföljning av inspektioner
1. Medlemsstaterna skall utan dröjsmål underrätta kommissionen om resultaten av varje inspektion och om eventuella förbud mot landning eller omlastning till följd av inspektionen.
2. Kommissionen skall utan dröjsmål översända denna information till NEAFC-sekretariatet och snarast möjligt till det inspekterade fartygets flaggstat.
AVDELNING III
SLUTBESTÄMMMELSER
Artikel 27
Konfidentialitet
Utöver skyldigheterna som anges i artikel 37 i förordning (EEG) nr 2847/93 skall medlemsstaterna och kommissionen följa bestämmelserna om konfidentialitet som antas enligt förfarandet i artikel 29.2.
Artikel 28
De bestämmelser som krävs för att genomföra denna förordning när det gäller artiklarna 2.3, 4.3, 5.3, 6.5, 7.3, 8, 11.5, 11.6, 12.1, 13.1, 14.1 h, 19.7 och 27 skall antas i enlighet med det förvaltningsförfarande som fastställs i artikel 29.2.
Artikel 29
1. Kommissionen skall biträdas av en förvaltningskommitté för fiske och vattenbruk (nedan kallad kommittén).
2. När det hänvisas till denna punkt, skall i artiklarna 4 och 7 i beslut 1999/468/EG tillämpas. Den tid som avses i artikel 4.3 i beslut 1999/468/EG skall vara en månad.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 30
Ikraftträdande
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas offciella tidning.
De bestämmelser som avses i artiklarna 6.2, 6.3, 8, 10 och 11 skall förbli i kraft på ad hoc-basis till och med den 31 december 2000. Senast den 30 september 2000 skall kommissionen lägga fram eventuella lämpliga förslag för en slutgiltig ordning. Rådet skall i enlighet med förfarandet i artikel 37 i EG-fördraget anta de nödvändiga åtgärderna senast den 31 december 2000.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
KOMMISSIONENS BESLUT
av den 16 december 1999
om fastställande av ekologiska kriterier för tilldelning av gemenskapens miljömärke till kylskåp
[delgivet med nr K(1999) 4522]
(Text av betydelse för EES)
(2000/40/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 880/92 av den 23 mars 1992 om ett gemenskapsprogram för tilldelning av miljömärke(1), särskilt artikel 5.1 andra stycket i denna, och
av följande skäl: 1. I artikel 5.1 i förordning (EEG) nr 880/92 föreskrivs att villkoren för tilldelning av gemenskapens miljömärke skall fastställas för varje produktgrupp för sig.
2. Enligt artikel 10.2 i förordning (EEG) nr 880/92 skall en produkts påverkan på miljön bedömas i enlighet med de särskilda kriterierna för produktgrupper.
3. Det är lämpligt att fastställa kriterier för testmetoder och klassificering för energiförbrukning i enlighet med kommissionens direktiv 94/2/EG av den 21 januari 1994 om genomförande av rådets direktiv 92/75/EEG om märkning som anger energiförbrukning hos elektriska kylskåp och frysar (även i kombination) för hushållsbruk(2) och att dessutom anpassa kraven på energiförbrukning till de tekniska innovationerna och utvecklingen på marknaden.
4. I beslut 96/703/EG(3), fastställde kommissionen ekologiska kriterier för tilldelning av gemenskapens miljömärke till kylskåp, vilka enligt artikel 3 i beslutet gällde till och med den 27 november 1999.
5. Det är lämpligt att fatta ett nytt beslut om fastställande av ekologiska kriterier för denna produktgrupp, så att tillverkare och importörer av kylskåp kan delta i gemenskapens miljömärkningsprogram.
6. I enlighet med artikel 6 i förordning (EEG) nr 880/92 har kommissionen rådgjort med de närmast berörda intressegrupperna i ett samrådsforum.
7. De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från den kommitté som inrättats enligt artikel 7 i förordning (EEG) nr 880/92.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Med produktgruppen kylskåp (nedan kallad produktgruppen) avses
Elektriska nätanslutna kylskåp, frysboxar och frysar (även i kombination) för hushållsbruk.
Apparater som även kan utnyttja andra energikällor, t.ex. batterier, omfattas inte av direktivet.
Artikel 2
Produktgruppens miljöpåverkan och användbarhet skall bedömas mot bakgrund av de kriterier som anges i bilagan.
Artikel 3
Definitionen av och kriterierna för produktgruppen skall gälla från och med dagen för anmälan av detta beslut till den 1 december 2002. Om ett nytt beslut om en definition av och kriterier för denna produktgrupp fortfarande inte antagits den 1 december 2002 skall giltighetsperioden förlängas fram till den 1 december 2003 eller till dess att ett nytt beslut antagits, om detta skulle ske tidigare.
Artikel 4
För administrativa ändamål skall denna produktgrupp tilldelas kodnummer %quot%012%quot%.
Artikel 5
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 3 maj 2000
om ersättning av beslut 94/3/EG om en förteckning över avfall i enlighet med artikel 1 a i rådets direktiv 75/442/EEG om avfall, och rådets beslut 94/904/EG om upprättande av en förteckning över farligt avfall i enlighet med artikel 1.4 i rådets direktiv 91/689/EEG om farligt avfall
[delgivet med nr K(2000) 1147]
(Text av betydelse för EES)
(2000/532/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 75/442/EEG av den 15 juli 1975 om avfall(1), senast ändrat genom direktiv 91/156/EEG(2), särskilt artikel 1 a i detta,
med beaktande av rådets direktiv 91/689/EEG av den 12 december 1991 om farligt avfall(3), särskilt artikel 1.4 andra strecksatsen i detta, och
av följande skäl:
(1) Flera medlemsstater har anmält ett antal avfallskategorier som de anser uppvisar en eller flera av de egenskaper som anges i bilaga III till direktiv 91/689/EEG.
(2) Enligt artikel 1.4 i direktiv 91/689/EEG skall kommissionen granska anmälningar från medlemsstaterna och vid behov revidera den förteckning över farligt avfall som upprättats i enlighet med rådets beslut 94/904/EG(4).
(3) Avfall som ingår i förteckningen över farligt avfall måste också införas i Europeiska avfallskatalogen som upprättats i enlighet med kommissionens beslut 94/3/EG(5). För att systemet skall bli mer överskådligt och för att förenkla gällande bestämmelser är det lämpligt att upprätta en gemenskapsförteckning som integrerar den avfallsförteckning som upprättats genom beslut 94/3/EG och den förteckning över farligt avfall som upprättats genom beslut 94/904/EG.
(4) Kommissionen skall i detta arbete bistås av den kommitté som inrättats genom artikel 18 i direktiv 75/442/EEG.
(5) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från ovannämnda kommitté.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Härmed antas förteckningen i bilagan till detta beslut.
Artikel 2
Avfall som klassificeras som farligt anses uppvisa en eller flera av de egenskaper som avses i bilaga III till direktiv 91/689/EEG och, vad beträffar H3 till H8, H10(6) och H11 i denna bilaga, en eller flera av följande egenskaper:
- flampunkt %amp%lt;= 55 °C,
- ett eller flera ämnen som klassificeras(7) som mycket giftiga vid en total koncentration %amp%gt;= 0,1 %,
- ett eller flera ämnen som klassificeras som mycket giftiga vid en total koncentration %amp%gt;= 3 %,
- ett eller flera ämnen som klassificeras som hälsoskadliga vid en total koncentration %amp%gt;= 25 %,
- ett eller flera frätande ämnen som klassificeras som R35 vid en total koncentration %amp%gt;= 1 %,
- ett eller flera frätande ämnen som klassificeras som R34 vid en total koncentration %amp%gt;= 5 %,
- ett eller flera irriterande ämnen som klassificeras som R41 vid en total koncentration %amp%gt;= 10 %,
- ett eller flera irriterande ämnen som klassificeras som R36, R37 eller R38 vid en total koncentration %amp%gt;= 20 %,
- ett eller flera ämnen som är kända för att vara cancerframkallande (kategori 1 eller 2) vid en total koncentration %amp%gt;= 0,1 %,
- ett eller flera ämnen som är skadliga för fortplantningen (kategori 1 eller 2) vilka klassificeras som R60 eller R61 vid en total koncentration %amp%gt;= 0,5 %,
- ett eller flera ämnen som är skadliga för fortplantningen (kategori 3) vilka klassificeras som R62 eller R63 vid en total koncentration %amp%gt;= 5 %,
- ett eller flera mutagena ämnen i kategori 1 eller 2 vilka klassificeras som R46 vid en total koncentration %amp%gt;= 0,1 %,
- ett eller flera mutagena ämnen i kategori 3 vilka klassificeras som R40 vid en total koncentration %amp%gt;= 1 %.
Artikel 3
Medlemsstaterna får i undantagsfall, på grundval av skriftlig bevisning som på lämpligt sätt tillhandahålls av innehavaren, besluta att en viss typ av avfall som enligt förteckningen är farligt inte uppvisar någon av de egenskaper som anges i bilaga III till direktiv 91/689/EEG. Utan att det påverkar tillämpningen av artikel 1.4 andra strecksatsen i direktiv 91/689/EEG får medlemsstaterna likaså i undantagsfall besluta att avfall som enligt förteckningen inte är farligt uppvisar en eller flera av de egenskaper som anges i bilaga III till direktiv 91/689/EEG. Kommissionen skall en gång per år underrättas om alla sådana beslut som fattas av medlemsstaterna. Kommissionen skall göra en sammanställning av dessa beslut och undersöka huruvida det finns anledning att ändra gemenskapens förteckning över avfall och farligt avfall mot bakgrund av sådana beslut.
Artikel 4
Medlemsstaterna skall vidta de åtgärder som är nödvändiga för att följa detta beslut senast den 1 januari 2002.
Artikel 5
Beslut 94/3/EG och beslut 94/904/EG skall upphöra att gälla från och med den 1 januari 2002.
Artikel 6
Detta beslut riktar sig till medlemsstaterna.
Rådets beslut
av den 28 september 2000
om ingående av ett avtal mellan Europeiska gemenskapen och Konungariket Norge om Norges deltagande i arbetet vid Europeiskt centrum för kontroll av narkotika och narkotikamissbruk
(2000/602/EG)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av europeiska gemenskapen, särskilt artikel 308 tillsammans med artikel 300.2 första stycket andra meningen i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2), och
av följande skäl:
(1) I artikel 13 i rådets förordning (EEG) nr 302/93 av den 8 februari 1993 om upprättande av ett europeiskt centrum för kontroll av narkotika och narkotikamissbruk(3), anges att tredje land som delar gemenskapens och medlemsstaternas intressen och målsättningar med uppgifterna och arbetet inom centrumet skall få möjlighet att delta i centrumets arbete.
(2) Det av kommissionen framförhandlade avtalet mellan gemenskapen och Konungariket Norge om Norges deltagande i arbetet vid Europeiskt centrum för kontroll av narkotika och narkotikamissbruk bör godkännas på gemenskapens vägnar.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Avtalet mellan Europeiska gemenskapen och Konungariket Norge om Norges deltagande i arbetet vid Europeiskt centrum för kontroll av narkotika och narkotikamissbruk godkänns härmed på gemenskapens vägnar.
Texten till avtalet bifogas detta beslut.
Artikel 2
Rådets ordförande bemyndigas härmed att utse den person som skall ha rätt att med för gemenskapen bindande verkan underteckna avtalet och att lämna den diplomatiska not som avses i artikel 12 i avtalet(4).
KOMMISSIONENS FÖRORDNING (EG) nr 452/2000
av den 28 februari 2000
om genomförande av rådets förordning (EG) nr 530/1999 om strukturstatistik över löner och arbetskraftskostnader vid kvalitetsbedömning av arbetskraftskostnadsstatistik
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 530/1999 av den 9 mars 1999 om strukturstatistik över löner och arbetskraftskostnader(1), särskilt artikel 11 i denna, och
av följande skäl:
(1) I enlighet med artikel 11 i förordning (EG) nr 530/1999 är det nödvändigt med tillämpningsåtgärder i fråga om utvärderingskriterier för kvaliteten på statistiken och den rapport där tillämpningen av förordningen beskrivs.
(2) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för det statistiska programmet som upprättades genom rådets beslut 89/382/EEG, Euratom(2).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Utvärderingskriterier för kvalitetsbedömning och anvisningar för innehållet i rapporten om kvalitet
Utvärderingskriterierna för kvalitetsbedömning och anvisningar för innehållet i den rapport om kvalitet som avses i artikel 10 i förordning (EG) nr 530/1999 återfinns i bilagan till denna förordning.
Artikel 2
Ikraftträdande
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 635/2000
av den 24 mars 2000
om ändring av förordning (EG) nr 2571/97 om försäljningen av smör till sänkta priser och om beviljande av stöd för grädde, smör och koncentrerat smör avsett att användas i framställningen av konditorivaror, glass och andra livsmedel
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1255/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter(1), särskilt artiklarna 10 och 15 i denna, och
av följande skäl:
(1) I kommissionens förordning (EG) nr 2571/97(2), senast ändrad genom förordning (EG) nr 494/1999(3) föreskrivs i artikel 3 a att de spårämnen kan användas som anges i bilaga II till den förordningen. Anledningen är att man skall kunna kontrollera att den slutliga användningen av produkterna följer föreskrifterna. Då vissa spårämnen sedan en tid inte längre används inom ramen för förordningen och det i bilaga II till förordningen även anges alternativa spårämnen, bör de berörda spårämnena avskaffas så att kontrollerna kan förenklas genom en minskning av antalet spårämnen. Samma spårämnen granskas också med hänsyn till de senaste forskningsrönen på området.
(2) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för mjölk och mjölkprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I bilaga II förordning (EG) nr 2571/97 skall punkt V utgå.
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Rådets förordning (EG) nr 1673/2000
av den 27 juli 2000
om den gemensamma organisationen av marknaderna för lin och hampa som odlas för fiberproduktion
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artiklarna 36 och 37 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3),
med beaktande av Regionkommitténs yttrande(4), och
av följande skäl:
(1) För att den gemensamma marknaden för jordbruksprodukter skall kunna fungera och utvecklas måste den åtföljas av införandet av en gemensam jordbrukspolitik. Denna politik bör framförallt innefatta gemensam organisation av marknaderna för jordbruksprodukter vilken kan utformas på olika sätt beroende på vilken produkt det är fråga om.
(2) Syftet med den gemensamma jordbrukspolitiken är att nå de mål som anges i fördraget. När det gäller lin och hampa som odlas för fiberproduktion bör det, utöver bestämmelserna om arealersättning i rådets förordning (EG) nr 1251/1999 av den 17 maj 1999 om upprättande av ett stödsystem för producenter av vissa jordbruksgrödor(5), föreskrivas åtgärder med hänsyn till den inre marknaden som omfattar stöd till förste beredare av lin- och hampstrån eller till jordbrukare som låter bereda stråna för egen räkning.
(3) För att säkerställa att lin- och hampstrån verkligen bereds bör stödet endast beviljas på vissa villkor, däribland att den förste beredaren skall vara godkänd och att beredarna åtar sig att ingå avtal om att köpa stråna. För att motverka eventuellt missbruk skall stödet till beredning likaså inte beviljas annat än i förhållande till beredningen av stråna eller användningen av fibrerna på marknaden, om jordbrukaren låter bereda stråna för egen räkning.
(4) För att gemenskapens medel inte skall missbrukas bör det inte beviljas stöd till en förste beredare eller jordbrukare om det kan konstateras att denne på ett konstlat sätt har uppfyllt de villkor som krävs för att få stödet och därmed får en förmån som inte är förenlig med målet för stödsystemet för stråberedning.
(5) Med hänsyn till de särskilda karaktärsdragen för dels marknaden för långa linfibrer, dels för marknaden för korta linfibrer och hampfibrer bör det fastställas olika stödbelopp för de två fiberkategorierna. För att säkerställa att det totalt beviljas ett stöd som gör det möjligt att behålla den traditionella produktionen av långa linfibrer på villkor som liknar dem som föreskrivs i rådets förordning (EEG) nr 1308/70 av den 4 juli 1970 om den gemensamma organisationen av marknaden för lin och hampa(6) bör stödbeloppet gradvis öka i takt med att det hektarstöd som producenter beviljas enligt förordning (EG) nr 1251/1999 gradvis minskar och stödet till korta linfibrer bör på sikt upphöra. För korta linfibrer och hampfibrer bör det beviljas ett stödbelopp som tillåter nya fiberprodukter och de potentiella avsättningsmarknaderna att anpassa sig till varandra under en viss tid. För att stimulera produktionen av korta linfibrer och hampfibrer av god kvalitet bör det föreskrivas en högsta procentandel orenheter och ved samt övergångsbestämmelser för att göra det möjligt för beredningsindustrin att anpassa sig till detta krav.
(6) Med tanke på den särskilda situationen i den traditionella linodlingen inom vissa områden i Nederländerna, Belgien och Frankrike är det nödvändigt att för berörda arealer bevilja ett kompletterande övergångsstöd till de första stråberedarna.
(7) För att undvika bedrägeri i form av ökning av de stödberättigande kvantiteterna bör medlemsstaterna införa en gräns för dessa i förhållande till de arealer för vilka det finns avtal eller åtagande att bereda stråna.
(8) För att begränsa de utgifter som uppstår genom tillämpningen av denna förordning bör det införas en stabiliseringsmekanism för varje typ av fiber, dvs. både för långa linfibrer och för korta linfibrer eller hampfibrer. För att bidra till att det produceras rimliga mängder i varje medlemsstat bör det för varje fibertyp fastställas en garanterad maximikvantitet som fördelas mellan medlemsstaterna i form av garanterade nationella kvantiteter. De garanterade nationella kvantiteterna för korta linfibrer och hampfibrer bör dock vara begränsade till den period som krävs för att nya produkter av dessa skall kunna anpassa sig till marknaden. De garanterade nationella kvantiteterna skall tillämpas för stödet till beredningen och berör inte den ordning som föreskrivs i förordning (EG) nr 1251/1999. De garanterade nationella kvantiteterna bör fastställas särskilt med hänsyn till de senaste genomsnittsarealerna för spånadslin och hampa, som i förekommande fall anpassas till de faktiska produktionsarealerna multiplicerat med den genomsnittliga fiberavkastningen. För de medlemsstater som för närvarande har liten produktion bör det fastställas en gemensam kvantitet som skall fördelas varje regleringsår så att den kan anpassas till deras produktionsutveckling.
(9) Det bör fastställas villkor för överföring mellan de garanterade nationella kvantiteter som tilldelats varje medlemsstat för de båda fiberkvaliteterna så att varje medlemsstat kan justera kvantiteterna i förhållande till skörden. Kvantiteterna överförs enligt en koefficient som säkerställer en oförändrad budgetsituation.
(10) Producentmedlemsstaterna skall vidta de åtgärder som är nödvändiga för att säkerställa att stödsystemet fungerar på ett smidigt sätt. Med hänsyn till den tid som krävs för att bereda all den stråhalm som producerats under regleringsåret bör det dessutom, som en kontrollåtgärd, införas ett system med utbetalning av förskott på stödet.
(11) Åtgärderna i systemet för handel med tredje land bör sammantaget göra det möjligt att avstå från kvantitativa restriktioner och från uttag av avgifter vid gemenskapens yttre gränser. Dessa åtgärder kan emellertid i undantagsfall visa sig otillräckliga. I sådana fall bör gemenskapen, i syfte att skydda marknaden mot störningar som kan uppstå till följd av detta, omedelbart ges möjligheten att vidta alla nödvändiga åtgärder. Dessa åtgärder skall vara förenliga med de åtaganden som följer av Världshandelsorganisationens avtal om jordbruk(7).
(12) För att illegal odling av hampa inte skall störa den gemensamma organisationen av marknaden för hampa som odlas för fiberproduktion, bör det föreskrivas kontroll av import av hampa och hamputsäde för att säkerställa att produkterna i fråga ger vissa garantier i fråga om tetrahydrocannabinolhalt. Import av andra hampfrön än sådana som är avsedda för utsäde bör underkastas kontroll genom att man upprättar ett ackrediteringssystem för de berörda importörerna.
(13) Allteftersom marknaderna för lin och hampa som odlas för fiberproduktion utvecklas skall medlemsstaterna och kommissionen skicka varandra de uppgifter som krävs för tillämpningen av denna förordning.
(14) De åtgärder som krävs för att genomföra denna förordning bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(8).
(15) De utgifter som medlemsstaterna ådrar sig till följd av de åtaganden som uppstår till följd av denna förordning bör finansieras av gemenskapen i enlighet med rådets förordning (EG) nr 1258/1999 av den 17 maj 1999 om finansiering av den gemensamma jordbrukspolitiken(9).
(16) Den gemensamma organisationen av marknaderna för lin och hampa, som fastställs i förordning (EEG) nr 1308/70, har vid ett flertal tillfällen ändrats men överensstämmer inte längre med de genomgripande förändringar som sektorn har genomgått. Förordning (EEG) nr 1308/70 och rådets förordning (EEG) nr 619/71 av den 22 mars 1971 om allmänna bestämmelser för beviljande av stöd för lin och hampa(10) bör därför upphöra att gälla. Rådets förordning (EEG) nr 620/71 av den 22 mars 1971 om rambestämmelser för försäljningsavtal för linstrå och hampstrå(11), rådets förordning (EEG) nr 1172/71 av den 3 juni 1971 om allmänna bestämmelser om stöd för privat lagring av lin- och hampfibrer(12), rådets förordning (EEG) nr 1430/82 av den 18 maj 1982 om importrestriktioner för hampa och hampfrö och om ändring av förordning (EEG) nr 1308/70 vad avser hampa(13), rådets förordning (EEG) nr 2059/84 av den 16 juli 1984 om allmänna bestämmelser för importrestriktioner för hampa och hampfrö och om ändring av förordning (EEG) nr 619/71 med avseende på hampa(14) som grundar sig på förordning (EEG) nr 1308/70 och förordning (EEG) nr 619/71 bör upphöra att gälla och ersättas med de nya bestämmelserna i den här förordningen.
(17) Övergången från systemet i förordning (EEG) nr 1308/70 till det som återges i den här förordningen kan orsaka problem som inte tas upp i den här förordningen. För att sådana problem skall kunna hanteras bör kommissionen anta nödvändiga övergångsåtgärder. Den bör dessutom bemyndigas att lösa specifika praktiska problem.
(18) Med hänsyn till den tidpunkt då denna förordning träder i kraft är det nödvändigt att föreskriva särskilda åtgärder för regleringsåret 2000/2001. Därför bör den ordning som gäller under regleringsåret 1999/2000 fortsätta att tillämpas till och med den 30 juni 2001. Stödbeloppen skall dock fastställas av kommissionen i förhållande till de tillgängliga budgetmedlen så snart de berörda arealerna har beräknats på ett tillförlitligt sätt och det kvarvarande beloppet för finansiering av åtgärder för att främja användningen av linfibrer har fastställts till 0.
(19) För att utvärdera effekterna av de nya åtgärderna skall kommissionen lämna rapporter till Europaparlamentet och rådet dels under 2003 om de garanterade nationella kvantiteterna och den högsta halten av orenheter och ved i korta linfibrer och hampfibrer och dels under 2005 om konsekvenserna för producenterna och marknaderna av stödet till beredning och det kompletterande stödet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Den gemensamma organisationen av marknaderna för lin och hampa som odlas för fiberproduktion skall omfatta ett system för den inre marknaden och ett system för handel med tredje land. Den skall omfatta följande produkter:
%gt%Plats för tabell%gt%
2. I denna förordning avses med
a) jordbrukare: en jordbrukare enligt definitionen i artikel 10 a i rådets förordning (EG) nr 1259/1999 av den 17 maj 1999 om upprättande av gemensamma bestämmelser för system för direktstöd inom ramen för den gemensamma jordbrukspolitiken(15),
b) godkänd förste beredare: en fysisk eller juridisk person eller en sammanslutning av fysiska eller juridiska personer, oavsett vilken juridisk status sammanslutningen eller dess medlemmar har enligt nationell rätt, som har godkänts av den medlemsstats behöriga myndighet på vars territorium det beredningsföretag är beläget som skall producera linfibrer eller hampfibrer.
3. Denna förordning skall tillämpas utan att tillämpningen av förordning (EG) nr 1251/1999 påverkas.
AVDELNING I
Den inre marknaden
Artikel 2
1. Härmed införs ett stöd för beredning av linstrån och hampstrån avsedda för fiberproduktion.
Stödet skall beviljas en godkänd förste beredare för den kvantitet fibrer som faktiskt framställts av stråna och för vilken det har ingåtts ett köpe- och försäljningsavtal med en jordbrukare.
Dock
a) skall köpe- och försäljningsavtalet, om den godkände förste beredaren och jordbrukaren är en och samma person, ersättas av ett åtagande av den berörda personen att utföra beredningen själv,
b) skall stödet beviljas jordbrukaren om denne behåller stråna som han har låtit bereda genom kontrakt med en godkänd förste beredare och styrker att han har släppt ut de erhållna fibrerna på marknaden.
2. Stöd skall inte beviljas en godkänd förste beredare eller en jordbrukare om det konstateras att denne på ett konstlat sätt har uppfyllt de villkor som krävs för att få stödet och därmed får en förmån som inte är förenlig med målet för detta system.
3. Stödbeloppet för beredningsstödet skall fastställas enligt följande:
a) För långa linfibrer
- 100 euro/ton för regleringsåret 2001/2002,
- 160 euro/ton för regleringsåren 2002/2003, 2003/2004, 2004/2005 och 2005/2006,
- 200 euro/ton från och med regleringsåret 2006/2007.
b) För korta linfibrer och hampfibrer, innehållande högst 7,5 % orenheter och ved, skall stödbeloppet vara 90 euro/ton för regleringsåren 2001/2002-2005/2006.
Medlemsstaten får dock för regleringsåren 2001/2002-2003/2004 besluta att också bevilja stödet med hänsyn till de traditionella avsättningsmöjligheterna
- för korta linfibrer som innehåller 7,5-15 % orenheter och ved av lin,
- för hampfibrer som innehåller 7,5-25 % orenheter och ved.
I dessa fall skall medlemsstaten bevilja stödbeloppet för en kvantitet som motsvarar högst 7,5 % orenheter och ved i den producerade kvantiteten.
4. De fiberkvantiteter som berättigar till stöd skall begränsas till de arealer för vilka det finns ett avtal eller åtagande enligt punkt 1.
Medlemsstaterna skall fastställa de begränsningar som avses i första stycket så att de överensstämmer med de garanterade nationella kvantiteter som avses i artikel 3.
5. På den godkände förste beredarens begäran skall ett förskott betalas ut för den kvantitet fibrer som framställts.
Artikel 3
1. För långa linfibrer fastställs en garanterad maximikvantitet på 75250 ton per regleringsår som skall fördelas mellan alla medlemsstater i form av garanterade nationella kvantiteter. Kvantiteten skall fördelas på följande sätt:
- 13800 ton för Belgien,
- 300 ton för Tyskland,
- 50 ton för Spanien,
- 55800 ton för Frankrike,
- 4800 ton för Nederländerna,
- 150 ton för Österrike,
- 50 ton för Portugal,
- 200 ton för Finland,
- 50 ton för Sverige,
- 50 ton för Förenade kungariket.
2. För stödberättigade korta linfibrer och hampfibrer fastställs en garanterad maximikvantitet på 135900 ton per regleringsår. Denna kvantitet skall fördelas i form av
a) garanterade nationella kvantiteter för följande medlemsstater:
- 10350 ton för Belgien,
- 12800 ton för Tyskland,
- 20000 ton för Spanien,
- 61350 ton för Frankrike,
- 5550 ton för Nederländerna,
- 2500 ton för Österrike,
- 1750 ton för Portugal,
- 2250 ton för Finland,
- 2250 ton för Sverige,
- 12100 ton för Förenade kungariket.
b) 5000 ton som skall fördelas i garanterade nationella kvantiteter, för varje regleringsår, mellan Danmark, Grekland, Irland, Italien och Luxemburg. Denna fördelning skall baseras på de arealer för vilka ett av de avtal ingåtts eller det åtagande gjorts som avses i artikel 2.1.
De nationella garanterade kvantiteterna för korta linfibrer och hampfibrer, eventuellt nedsatta enligt punkt 5 i denna artikel, skall inte tillämpas från och med regleringsåret 2006/2007.
3. Om de fibrer som har framställts i en medlemsstat kommer från strån som producerats i en annan medlemsstat skall dessa kvantiteterna fibrer påföras den garanterade nationella kvantiteten i den medlemsstaten där stråna har skördats. Stödet skall utbetalas av den medlemsstat på vars garanterade nationella kvantitet fibrerna har påförts.
4. De medlemsstater som så önskar får en enda gång och före den 30 juni 2001 mellan sig överföra en del av sina garanterade nationella kvantiteter enligt punkt 1 eller punkt 2, eventuellt anpassade i enlighet med punkt 5. I detta fall skall de underrätta kommissionen som skall underrätta de övriga medlemsstaterna.
5. En medlemsstat får överföra en del av sin nationella garanterade kvantitet enligt punkt 1 till sin nationella garanterade kvantitet enligt punkt 2 och vice versa.
Vid de överföringar som avses i första stycket skall 1 ton långa linfibrer vara lika med 2,2 ton korta linfibrer och hampfibrer.
Stödbeloppen för beredningen skall beviljas för högst de kvantiteter som anges i punkt 1 respektive punkt 2, anpassade enligt de första två styckena i denna punkt och enligt punkt 4.
Artikel 4
Fram till och med regleringsåret 2005/2006 skall ett extra stöd beviljas till den förste godkände beredaren för de linarealer som befinner sig i de områden som beskrivs i bilagan och för vars stråproduktion
- sådana köpe- eller försäljningsavtal ingås eller ett sådant åtagande görs som avses i artikel 2.1, och
- till vilken ett stöd ges för beredning av långa fibrer.
Det extra stödbeloppet skall vara 120 euro per hektar i område I och 50 euro per hektar i område II.
AVDELNING II
Handel med tredje land
Artikel 5
1. Denna artikel skall inte påverka tillämpningen av mer restriktiva bestämmelser som medlemsstaterna kan ha antagit med beaktande av fördraget och av de åtaganden som följer av Världshandelsorganisationens avtal om jordbruk.
2. Vid all import av hampa med ursprung i tredje land skall det utfärdas ett intyg om att följande villkor är uppfyllda:
- Oberedd mjukhampa som omfattas av KN-nummer 5302 10 00 skall uppfylla de villkor som anges i artikel 5a i förordning (EG) nr 1251/1999.
- Olika sorters hampfrön avsedda för utsäde som omfattas av KN-nummer 1207 99 10 skall åtföljas av ett bevis om att tetrahydrocannabiolhalten inte överstiger den som fastställs i artikel 5a i förordning (EG) nr 1251/1999.
- Andra hampfrön än sådana som är avsedda för utsäde och som omfattas av KN-nummer 1207 99 91 får importeras endast genom av medlemsstaten godkända importörer för att säkerställa att de inte skall användas för utsäde.
Till gemenskapen importerade produkter enligt första och andra strecksatsen skall kontrolleras för att avgöra om de uppfyller villkoren enligt denna artikel.
Artikel 6
Om inte annat föreskrivs i denna förordning eller i en bestämmelse som antagits i enlighet därmed, skall följande vara förbjudet i handeln med tredje land:
- Uttag av en avgift som har motsvarande verkan som en tull.
- Tillämpning av kvantitativa begränsningar eller åtgärder med motsvarande verkan.
Artikel 7
1. Om gemenskapsmarknaden för en eller flera av de produkter som förtecknas i artikel 1.1 på grund av import eller export påverkas eller hotas av allvarliga störningar som sannolikt kommer att äventyra uppnåendet av de mål som anges i artikel 33 i fördraget, får lämpliga åtgärder vidtas i samband med handeln med tredje land till dess att sådan störning eller sådant hot om störning har upphört.
Rådet skall på kommissionens förslag och med kvalificerad majoritet anta allmänna tillämpningsföreskrifter för denna punkt och skall bestämma i vilka fall och inom vilka gränser medlemsstater får vidta skyddsåtgärder.
2. I det fall som avses i punkt 1 skall kommissionen på begäran av en medlemsstat eller på eget initiativ besluta om nödvändiga åtgärder; åtgärderna skall meddelas medlemsstaterna och skall tillämpas omedelbart. Om kommissionen mottar en begäran från en medlemsstat, skall den fatta beslut därom inom tre arbetsdagar från och med mottagandet av begäran.
3. Varje medlemsstat får hänskjuta kommissionens beslut till rådet inom tre arbetsdagar efter det att beslutet meddelades. Rådet skall sammanträda utan dröjsmål. Det får med kvalificerad majoritet ändra eller upphäva beslutet ifråga inom en månad efter den dag då det hänskjutits till rådet.
4. Denna artikel skall tillämpas med beaktande av de skyldigheter som följer av avtal som har ingåtts i enlighet med artikel 300.2 i fördraget.
AVDELNING III
Allmänna bestämmelser
Artikel 8
Om inte annat föreskrivs i denna förordning skall artiklarna 87, 88 och 89 i fördraget tillämpas på produktion av och handel med de produkter som anges i artikel 1.1 i denna förordning.
Artikel 9
De åtgärder som krävs för att genomföra denna förordning och som rör de frågor som anges nedan skall antas i enlighet med det förvaltningsförfarande som avses i artikel 10.2. Det gäller särskilt
- villkoren för godkännande av förste beredare,
- villkoren för en godkänd förste beredare när det gäller de köpe- eller försäljningsavtal och åtaganden som avses i artikel 2.1,
- villkoren för jordbrukarna i det fall som avses i artikel 2.1 b,
- kriterierna för dels långa linfibrer, dels korta linfibrer och hampfibrer,
- metoderna för beräkning av de stödberättigade kvantiteterna i de fall som avses i artikel 2.3 b andra stycket,
- villkoren för att bevilja stöd och förskott, och särskilt bevis för beredningen av strån,
- villkoren för att fastställa de begränsningar som avses i artikel 2.4,
- fördelningen av den kvantitet på 5000 ton som avses i artikel 3.2 b,
- villkoren för överföring mellan de garanterade nationella kvantiteter som avses i artikel 3.5,
- villkoren för beviljande av det extra stöd som avses i artikel 4.
Åtgärderna får även gälla alla kontroller som är nödvändiga för att skydda gemenskapens finansiella intressen mot bedrägeri och andra oegentligheter.
Artikel 10
1. Kommissionen skall biträdas av Förvaltningskommittén för naturfibrer (nedan kallad kommittén).
2. När det hänvisas till denna punkt skall artiklarna 4 och 7 i beslut 1999/468/EG tillämpas.
Den tid som avses i artikel 4.3 i beslut 1999/468/EG skall vara en månad.
3. Kommittén får behandla varje annan fråga som dess ordförande, antingen på eget initiativ eller på begäran av företrädaren för en medlemsstat, hänskjuter till den.
4. Kommittén skall själv anta sin arbetsordning.
Artikel 11
Förordning (EG) nr 1258/1999 och de bestämmelser som har fastställts för dess genomförande skall tillämpas för de produkter som anges i artikel 1.1 i den här förordningen.
AVDELNING IV
Övergångsbestämmelser och slutbestämmelser
Artikel 12
1. För regleringsåret 2000/2001 skall stödbeloppen för i gemenskapen producerad lin och hampa fastställas, senast den 31 oktober 2000, i enlighet med förfarandet i artikel 10.2.
Dessa belopp skall fastställas genom att på de belopp som gäller för regleringsåret 1999/2000 tillämpa en koefficient och som är lika med förhållandet mellan
- de genomsnittliga utgifterna per hektar som motsvarar 88 miljoner euro för den totala areal som framgår av skördedeklarationerna, och
- de beräknade genomsnittliga utgifterna på 721 euro per hektar för regleringsåret 1999/2000.
Stödbeloppen för regleringsåret 2000/2001 får under inga omständigheter överstiga de belopp som har fastställts för regleringsåret 1999/2000.
2. För regleringsåret 2000/2001 skall det belopp som tas ut på stödet till lin och som är avsett att finansiera de åtgärder som främjar användningen av linfibrer fastställas till 0 euro per hektar.
3. Regleringsåret 2000/2001 slutar den 30 juni 2001.
Artikel 13
Förordningarna (EEG) nr 1308/70, (EEG) nr 619/71, (EEG) nr 620/71, (EEG) nr 1172/71, (EEG) nr 1430/82 och (EEG) nr 2059/84 skall upphöra att gälla från och med den 1 juli 2001.
Artikel 14
Kommissionen skall i enlighet med förfarandet i artikel 10.2 besluta om
- de åtgärder som krävs för att underlätta övergången från bestämmelserna i förordningarna (EEG) nr 1308/70 och (EEG) nr 619/71 till dem som införs genom denna förordning,
- de åtgärder som krävs för att lösa särskilda praktiska problem. Under förutsättning att de är vederbörligen motiverade får sådana åtgärder avvika från vissa delar av denna förordning.
Artikel 15
1. Senast den 31 december 2003 skall kommissionen för Europaparlamentet och rådet lägga fram en rapport, eventuellt tillsammans med förslag, om produktionstendenserna i de olika medlemsstaterna och om konsekvenserna av reformen av den gemensamma organisationen av marknaden för sektorns avsättningsmöjligheter och ekonomiska livskraft. Den skall även behandla den maximala nivån orenheter och ved som skall gälla för korta linfibrer och hampfibrer.
Rapporten skall eventuellt utgöra grunden för en ny fördelning och för en möjlig ökning av de garanterade nationella kvantiteterna. Kommissionen skall särskilt ta hänsyn till produktionsnivån, beredningskapaciteten och avsättningsmöjligheterna på marknaden.
2. År 2005 skall kommissionen för Europaparlamentet och rådet lägga fram en rapport om beredningsstödet, eventuellt tillsammans med förslag.
Rapporten skall innehålla en bedömning av konsekvenserna av beredningsstödet, särskilt för
- producenternas situation när de gäller de odlade arealerna och de pris som de får,
- tendenserna på marknaderna för textilfibrer och utvecklingen av nya produkter,
- beredningsindustrin.
I rapporten skall det, med hänsyn till den alternativa produktionen, anges om industrin kan fungera enligt de fastställda riktlinjerna. Den skall även behandla möjligheten att permanent behålla beredningsstödet per ton korta linfibrer och hampfibrer och det extra stöd per hektar lin som avses i artikel 4 efter regleringsåret 2005/2006.
Artikel 16
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska gemenskapernas officiella tidning.
Artiklarna 1-11 skall tillämpas från och med regleringsåret 2001/2002.
Förordning (EEG) nr 1308/70 och förordning (EEG) nr 619/71 skall fortsätta att tillämpas när det gäller regleringsåren 1998/1999, 1999/2000 och 2000/2001.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens beslut
av den 27 december 2000
om ändring för fjärde gången av beslut 1999/467/EG om fastställande av officiellt tuberkulosfri status för nötkreatursbesättningarna i vissa medlemsstater eller regioner i medlemsstater
[delgivet med nr K(2000) 4144]
(Text av betydelse för EES)
(2001/26/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 64/432/EEG om djurhälsoproblem som påverkar handeln med nötkreatur och svin inom gemenskapen(1), senast ändrat genom direktiv 2000/20/EG(2), särskilt bilaga A.I.4 i detta, och
av följande skäl:
(1) Genom kommissionens beslut 1999/467/EG av den 15 juli 1999 om fastställande av officiellt tuberkulosfri status för nötkreatursbesättningarna i vissa medlemsstater eller regioner i medlemsstater och om upphävande av beslut 97/76/EG(3), senast ändrat genom beslut 2000/694/EG(4), förklarades vissa medlemsstater och regioner i medlemsstater vara officiellt tuberkulosfria.
(2) De behöriga myndigheterna i Frankrike har till kommissionen överlämnat belägg för att samtliga krav i bilaga A.I.4 till direktiv 64/432/EEG är uppfyllda, och framför allt kravet på att mer än 99,9 % av nötkreatursbesättningarna i Frankrike under de sex senaste åren skall ha varit officiellt fria från bovin tuberkulos på grundval av läget den 31 december varje år. De behöriga myndigheterna har också lagt fram belägg för att informationen i den databas som upprättades i december 1999 gör det möjligt att spåra nötkreatur som identifierats enligt gemenskapens lagstiftning.
(3) Det förefaller därför lämpligt att klassa Frankrike som officiellt fritt från bovin tuberkulos enligt ovannämnda direktiv.
(4) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga I till beslut 1999/467/EG skall ersättas med bilagan till det här beslutet.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Rådets beslut
av den 22 december 2000
om undertecknande och provisorisk tillämpning av det i Bryssel den 8 november 2000 paraferade avtalet mellan Europeiska gemenskapen och Republiken Kroatien om handel med textilprodukter
(2001/55/EG)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 133 jämförd med artikel 300.2 första stycket första meningen i detta,
med beaktande av kommissionens förslag, och
av följande skäl:
(1) Kommissionen har på gemenskapens vägnar förhandlat fram ett avtal med Republiken Kroatien om handel med textilprodukter.
(2) Avtalet paraferades den 8 november 2000.
(3) Avtalet bör undertecknas på gemenskapens vägnar, med förbehåll för att det senare ingås.
(4) Avtalet bör tillämpas provisoriskt från och med den 1 januari 2001 till dess att de relevanta förfarandena för det formella ingåendet har slutförts, under förutsättning att det tillämpas ömsesidigt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Rådets ordförande bemyndigas härmed att utse de personer som skall ha rätt att på gemenskapens vägnar underteckna avtalet mellan Europeiska gemenskapen och Republiken Kroatien om handel med textilprodukter, med förbehåll för att det senare ingås.
Artikel 2
Det avtal som avses i artikel 1 skall tillämpas provisoriskt från och med den 1 januari 2001 till dess att förfarandena för dess ingående har slutförts, under förutsättning att det tillämpas ömsesidigt.
Texten till avtalet bifogas detta beslut.
Rådets beslut
av den 22 januari 2001
om inrättande av Europeiska unionens militära stab
(2001/80/GUSP)
EUROPEISKA UNIONENS RÅD HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om Europeiska unionen, särskilt artikel 28.1 i detta,
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 207.2 i detta, och
av följande skäl:
(1) Inom ramen för den förstärkning av den gemensamma utrikes- och säkerhetspolitiken (GUSP), och särskilt den gemensamma europeiska säkerhets- och försvarspolitiken, som det föreskrivs om i artikel 17 i Fördraget om Europeiska unionen, uppnåddes vid mötet i Europeiska rådet i Nice den 7-11 december 2000 en överenskommelse om inrättande av Europeiska unionens militära stab, i vilken fastställs dennas uppdrag och uppgifter.
(2) Enligt Europeiska rådets riktlinjer bör den militära staben göras redo att inleda arbetet. HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Militär personal kommer att avdelas från medlemsstaterna till rådets generalsekretariat för att bilda Europeiska unionens militära stab (EUMS).
2. Den militära staben kommer att ingå i rådets generalsekretariat.
Artikel 2
Den militära stabens uppdrag och uppgifter fastställs i bilaga V till ordförandeskapets rapport som godkänts av Europeiska rådet i Nice och som återges i bilagan.
Artikel 3
Alla medlemmar i den militära staben skall vara medborgare i Europeiska unionens medlemsstater.
Artikel 4
1. Medlemmarna i den militära staben skall omfattas av regler som kommer att fastställas i ett rådsbeslut.
2. Tills det beslut som omnämns i punkt 1 träder i kraft skall rådets beslut 2000/178/GUSP av den 28 februari 2000 om de regler som skall gälla för utstationerade militära nationella experter vid rådets generalsekretariat under interimsperioden under den interimistiska perioden(1) förbli gällande.
Artikel 5
Detta beslut blir gällande samma dag som det antas.
Det skall tillämpas från och med ett datum som fastställs av generalsekreteraren/den höge representanten, efter samråd med Kommittén för utrikes- och säkerhetspolitik och med det interimistiska militära organet/den militära kommittén, och i princip före slutet av juni månad 2001.
Fram till datum för tillämpningen av detta beslut skall generaldirektören för den militära staben (DGEUMS), som kommer att tillträda sin tjänst den 1 mars 2001(2), fungera som chef för de militära experter som avdelats från medlemsstaterna till rådets sekretariat(3).
Artikel 6
Detta beslut skall offentliggöras i Officiella tidningen.
Europeiska centralbankens beslut
av den 6 december 2001
om fördelning av de monetära inkomsterna för de deltagande medlemsstaternas nationella centralbanker från och med räkenskapsåret 2002
(ECB/2001/16)
(2001/914/EG)
ECB-RÅDET HAR FATTAT DETTA BESLUT
med beaktande av Stadgan för Europeiska centralbankssystemet och Europeiska centralbanken (nedan kallad stadgan), särskilt artikel 32 i denna, och
av följande skäl:
(1) Enligt artikel 32.1 i stadgan är monetära inkomster sådana inkomster som uppkommer då de nationella centralbankerna fullgör monetära uppgifter. I enlighet med artikel 32.2 i stadgan skall summan av de monetära inkomsterna för varje nationell centralbank vara lika med centralbankens årliga inkomster av de tillgångar som den innehar som motvärden till sedlar i omlopp och till inlåning från kreditinstitut. Dessa tillgångar skall reserveras av de nationella centralbankerna i enlighet med ECB-rådets riktlinjer. Från och med räkenskapsåret 2003 skall de nationella centralbankerna reservera sådana tillgångar som uppkommit som ett resultat av att de nationella centralbankerna fullgör monetära uppgifter som tillgångar som de innehar som motvärden till sedlar i omlopp och till inlåning från kreditinstitut. Enligt artikel 32.4 i stadgan skall varje nationell centralbanks monetära inkomster minskas med ett belopp som motsvarar centralbankens räntebetalningar till följd av förpliktelser på grund av inlåning från kreditinstituten enligt artikel 19 i stadgan.
(2) Enligt artikel 32.5 i stadgan skall summan av de nationella centralbankernas monetära inkomster fördelas på de nationella centralbankerna i förhållande till deras inbetalda andelar av Europeiska centralbankens (ECB) kapital.
(3) Enligt artikel 32.6 och 32.7 i stadgan åligger det ECB-rådet att fastställa riktlinjer för hur ECB skall utföra avräkningen och betalningen av saldona från fördelningen av de monetära inkomsterna och att vidta alla övriga åtgärder som behövs för tillämpningen av artikel 32 i stadgan.
(4) Av artikel 10 i rådets förordning (EG) nr 974/98 av den 3 maj 1998 om införande av euron(1) framgår att ECB och de nationella centralbankerna (nedan kallade Eurosystemet) från och med den 1 januari 2002 skall sätta sedlar som anges i euro i omlopp. Enligt artikel 15 i nämnda förordning skall sedlar i nationell valuta behålla sin ställning som lagligt betalningsmedel under högst sex månader efter övergångsperiodens utgång. År 2002 måste därför betraktas som ett speciellt år, eftersom de sedlar som är i omlopp i nationella valutaenheter fortfarande kan utgöra en avsevärd del av det totala värdet på de sedlar som befinner sig i omlopp i Eurosystemet och olika mönster kan förekomma i olika medlemsstater. Denna situation är jämförbar med situationen mellan 1999-2001, varför man under räkenskapsåret 2002 skall beräkna monetära inkomster med en metod som motsvarar den som fastställdes i beslut ECB/2000/19 av den 3 november 1998 i dess ändrade lydelse enligt beslut av den 14 december 2000 om fördelningen av de monetära inkomsterna för de deltagande medlemsstaternas nationella centralbanker och ECB:s förluster för räkenskapsåren 1999-2001(2), så att det säkerställs att förändringar i det mönster enligt vilket sedlar befinner sig i omlopp inte medför väsentliga ändringar i de nationella centralbankernas relativa inkomstlägen. För 2002 kan ECB-rådet enligt artikel 32.3 besluta att de monetära inkomsterna, med avvikelse från artikel 32.2 i stadgan, skall beräknas enligt en annan metod.
(5) Enligt artikel 9.1 i riktlinje ECB/2001/1 av den 10 januari 2001 om antagande av vissa bestämmelser avseende utbytet av sedlar och mynt 2002(3) skall eurosedlar som förhandstilldelas kreditinstitut eller deras utsedda ombud debiteras respektive konto hos de nationella centralbankerna till nominella värdet enligt följande %quot%linjära modell%quot% för debitering: en tredjedel av det förhandstilldelade beloppet debiteras den 2 januari 2002, en tredjedel den 23 januari 2002 och den sista tredjedelen den 30 januari 2002. Vid beräkningen av monetära inkomster för 2002 måste hänsyn tas till denna %quot%linjära modell%quot% för debitering.
(6) Detta beslut har samband med beslut ECB/2001/15 av den 6 december 2001 om utgivningen av eurosedlar(4), där det stadgas att ECB och de nationella centralbankerna skall ge ut eurosedlar. Av beslut ECB/2001/15 framgår att tilldelningen av eurosedlar i omlopp till de nationella centralbankerna skall ske i förhållande till deras inbetalda andelar av ECB:s kapital. Enligt samma beslut skall ECB:s tilldelning av det sammanlagda värdet av eurosedlar i omlopp vara 8 procent. Fördelningen av eurosedlar bland Eurosystemets medlemmar kommer att medföra att olika saldon uppkommer inom Eurosystemet. Förräntningen av dessa saldon inom Eurosystemet för eurosedlar i omlopp får direkta inkomstkonsekvenser för var och en av Eurosystemets medlemmar och skall därför regleras genom detta beslut. ECB:s inkomster från avkastningen på de fordringar ECB har inom Eurosystemet på de nationella centralbankerna avseende dess andel av eurosedlar i omlopp skall i princip, i enlighet med ECB-rådets beslut, fördelas bland de nationella centralbankerna i förhållande till deras andel i fördelningsnyckeln för tecknat kapital under samma räkenskapsår som inkomsterna uppkommer.
(7) Nettosaldot av fordringar och skulder inom Eurosystemet för eurosedlar i omlopp skall förräntas enligt ett objektivt kriterium som motsvarar kapitalkostnaden. För detta ändamål bedöms räntan för de huvudsakliga refinansieringstransaktionerna som används inom Eurosystemet vid de huvudsakliga refinansieringstransaktionerna vara ändamålsenlig.
(8) Nettoskulderna inom Eurosystemet för eurosedlar i omlopp skall ingå i skuldbasen vid beräkningen av de nationella centralbankernas monetära inkomster enligt stadgans artikel 32.2, eftersom de motsvarar sedlar i omlopp. Avveckling av räntebetalningarna inom Eurosystemet för saldon avseende eurosedlar i omlopp kommer därför att leda till att en avsevärd del av Eurosystemets monetära inkomster kommer att fördelas mellan de nationella centralbankerna i förhållande till deras inbetalda andelar av ECB:s kapital. Dessa saldon inom Eurosystemet bör justeras så att de nationella centralbankernas balans- och resultaträkningar kan anpassas gradvis. Justeringarna bör baseras på värdet av de sedlar som varje nationell centralbank har i omlopp under en period innan eurosedlarna införs. Dessa justeringar bör ta hänsyn till de speciella omständigheterna under 2002, då medlemsstaterna har olika övergångsscenarier och kreditinstituten kommer att ha större innehav av kontanter än normalt, och bör tillämpas på årsbasis i enlighet med en fastställd formel under högst fem år därefter.
(9) Justeringarna av Eurosystemets saldon för eurosedlar i omlopp har beräknats så att de skall kompensera för varje väsentlig ändring i de nationella centralbankernas inkomstlägen som kan bli konsekvensen av att eurosedlarna införs och den därpå följande fördelningen av monetära inkomster. ECB-rådet har därför beslutat att inte göra något avsteg från stadgans artikel 32, vilket är tillåtet enligt stadgans artikel 51.
(10) Justeringarna av saldon inom Eurosystemet för eurosedlar i omlopp måste ta hänsyn till Storhertigdömet Luxemburgs speciella situation som har sin grund i landets monetära historia.
(11) ECB-rådet har antagit detta beslut med den avsikten att dess ekonomiska resultat, och den finansiella jämnvikt dessa ekonomiska resultat medför, skall förbli oförändrade under den tidsperiod artikel 4 i detta beslut tillämpas och ECB-rådet har därför åtagit sig att säkerställa att bestämmelserna i detta beslut upprätthålls till den 31 december 2007.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Definitioner
I detta beslut avses med
a) deltagande medlemsstater: de medlemsstater som har infört den gemensamma valutan i enlighet med Fördraget om upprättandet av Europeiska gemenskapen,
b) nationella centralbanker: de deltagande medlemsstaternas nationella centralbanker,
c) skuldbasen: summan av de i bilaga I till detta beslut angivna skuldposterna i varje nationell centralbanks balansräkning,
d) reserverade tillgångar: värdet av de i bilaga II till detta beslut angivna tillgångar som hålls som motvärden till skuldbasen i varje nationell centralbanks balansräkning,
e) Eurosystemets saldon för eurosedlar i omlopp: fordringar och skulder som uppkommer mellan en nationell centralbank och ECB samt mellan en nationell centralbank och övriga nationella centralbanker som resultat av att artikel 4 i beslut ECB/2001/15 av den 6 december 2001 om utgivningen av eurosedlar tillämpas,
f) fördelningsnyckel för tecknat kapital: procenttal som erhålls när man tillämpar vikten i den fördelningsnyckel som avses i artikel 29.1 i stadgan och som fastställs i beslut ECB/1998/13 av den 1 december 1998 om de nationella centralbankernas procentandelar i fördelningsnyckeln till Europeiska centralbankens kapital(5) på de nationella centralbankerna,
g) kreditinstitut: kreditinstitut som omfattas av kassakrav enligt förordning ECB/1998/15(6) angående tillämpningen av minimireserver (kassakrav), ändrad genom förordning ECB/2000/8(7),
h) den harmoniserade balansräkningen: den harmoniserade balansräkning som redovisas i bilaga IX till riktlinje ECB/2000/18 om den rättsliga ramen för redovisning och rapportering inom Europeiska centralbankssystemet, med de ändringar som gjordes den 15 december 1999 och den 14 december 2000(8),
i) referensräntan: den senaste tillgängliga marginalränta som Eurosystemet använt för sina huvudsakliga refinansieringstransaktioner enligt kapitel 3.1.2 i bilaga I till riktlinje ECB/2000/7 av den 31 augusti 2000 om Eurosystemets penningpolitiska instrument och förfaranden(9). Om mer än en refinansieringstransaktion genomförs med samma likviddag, skall ett enkelt genomsnitt av de parallella transaktionernas marginalränta användas.
Artikel 2
Eurosystemets saldon för eurosedlar i omlopp
1. Eurosystemets saldon för eurosedlar i omlopp skall beräknas månadsvis och bokföras hos ECB och de nationella centralbankerna den första öppethållandedagen i månaden med den föregående månadens sista öppethållandedag som valutadag.
Den första beräkningen av Eurosystemets saldon för eurosedlar i omlopp enligt föregående stycke skall göras för förhandstilldelade eurosedlar den 2 januari 2002 med valutadag den 1 januari 2002.
2. Eurosystemets saldon för eurosedlar i omlopp, inklusive sådana som uppkommer genom tillämpningen av artikel 4 i detta beslut, skall förräntas till referensräntan.
3. Den förräntning som avses i föregående punkt skall avvecklas genom kvartalsvisa betalningar via Target.
4. Med avvikelse från föregående punkt skall den förräntning som avses i punkt 2 för räkenskapsåret 2002 avvecklas vid årets slut.
Artikel 3
Metod för beräkning av monetära inkomster
1. Under 2002 skall de monetära inkomsterna för varje nationell centralbank beräknas enligt följande formel:
%gt%Hänvisning till %gt%,där:
MI är en nationell centralbanks monetära inkomster som skall läggas samman med motsvarande belopp för övriga nationella centralbanker,
LB är den nationella centralbankens skuldbas, och
RR är referensräntan.
2. Från och med 2003 skall varje nationell centralbanks monetära inkomster fastställas genom beräkning av de faktiska inkomsterna från de bokförda reserverade tillgångarna. Ett undantag från detta är guld, som inte skall anses generera några inkomster.
3. Om en nationell centralbanks reserverade tillgångar över- eller understiger värdet på dess skuldbas, skall mellanskillnaden kompenseras genom att man på mellanskillnadens värde tillämpar den genomsnittliga procentuella avkastningen från alla nationella centralbankers sammanlagda reserverade tillgångar.
Denna genomsnittliga procentuella avkastning skall beräknas på följande sätt. De nationella centralbankernas samtliga inkomster från reserverade tillgångar skall sammanräknas - exklusive sådana inkomster som är resultatet av nettofordringar inom Eurosystemet på grund av Target-transaktioner (punkt A 3 i bilaga II) och nettofordringar inom Eurosystemet från eurosedlar i omlopp inklusive sådana som är resultatet av tillämpningen av artikel 4 (punkt A 4 i bilaga II) - och divideras med det genomsnittliga beloppet på Eurosystemets samtliga reserverade tillgångar. Denna genomsnittliga procentsats skall tillämpas på basis av ett år om 360 dagar.
Artikel 4
Justering av saldon inom Eurosystemet
1. Vid beräkningen av de monetära inkomsterna skall varje nationell centralbanks saldon inom Eurosystemet för eurosedlar i omlopp justeras med ett utjämningsbelopp som beräknas enligt följande formel:
%gt%Hänvisning till %gt%,där:
CA är utjämningsbeloppet,
K är det belopp för varje nationell centralbank som erhålls om man använder fördelningsnyckeln för tecknat kapital på det genomsnittliga värdet av sedlar i omlopp under perioden 1 juli 1999 till och med 30 juni 2001,
A är det genomsnittliga beloppet för varje nationell centralbank av sedlar i omlopp under perioden 1 juli 1999 till och med 30 juni 2001,
C är följande koefficient för varje räkenskapsår:
%gt%Plats för tabell%gt%
2. Summan av de nationella centralbankernas utjämningsbelopp skall vara 0.
3. Utjämningsbeloppen och motposter till dessa utjämningsbelopp skall den första öppethållandedagen varje kalenderår bokföras på separata Eurosystem-konton hos varje nationell centralbank med valutadag den 1 januari. De bokföringsposter som används för att utjämna utjämningsbeloppen skall inte förräntas.
4. Om beloppet för de eurosedlar som Banque centrale du Luxembourg sätter i omlopp under 2002 överstiger det genomsnittliga beloppet för dess sedlar i omlopp under perioden 1 juli 1999 till och med 30 juni 2002 med 25 procent eller mer, skall bokstaven A i den formel som återfinns i punkt 1 för Banque centrale du Luxembourg vara det belopp för sedlar som Banque centrale du Luxembourg sätter i omlopp under 2002, dock högst 2,2 miljarder euro. Om detta undantag tillämpas skall alla de utjämningsbelopp som beräknats enligt artikel 4.1 justeras retroaktivt i slutet av 2002, så att överensstämmelse med punkt 2 säkerställs. Sådana retroaktiva justeringar skall ske proportionellt till fördelningsnyckeln för tecknat kapital.
5. Om det inträffar sådana speciella omständigheter som beskrivs i bilaga III till detta beslut rörande sedlarnas ändrade omloppsmönster skall, med avvikelse från punkt 1 ovan, varje nationell centralbanks saldo inom Eurosystemet för eurosedlar i omlopp justeras i enlighet med föreskrifterna i nämnda bilaga.
6. Föreskrifterna i denna artikel om justeringar av saldon inom Eurosystemet skall upphöra att gälla från och med den 1 januari 2008.
Artikel 5
Beräkning och fördelning av de monetära inkomsterna
1. ECB skall för varje dag beräkna de monetära inkomsterna för varje nationell centralbank. Beräkningen skall göras på grundval av de redovisningsuppgifter som de nationella centralbankerna rapporterar till ECB. ECB skall varje kvartal underrätta de nationella centralbankerna om de kumulerade beloppen.
2. De olika nationella centralbankernas monetära inkomster skall minskas med ett belopp som motsvarar upplupen eller erlagd ränta för skulder som ingår i skuldbasen och i enlighet med beslut som ECB-rådet fattar på grundval av artikel 32.4 andra stycket i stadgan.
3. Fördelningen av de nationella centralbankernas monetära inkomster proportionellt i förhållande till fördelningsnyckeln för tecknat kapital skall göras i slutet av varje räkenskapsår.
Artikel 6
Slutbestämmelser
1. Detta beslut träder i kraft den 1 januari 2002.
2. Detta beslut skall offentliggöras i Europeiska gemenskapernas officiella tidning.
Rådets gemensamma ståndpunkt
av den 27 december 2001
om tillämpning av särskilda åtgärder i syfte att bekämpa terrorism
(2001/931/GUSP)
EUROPEISKA UNIONENS RÅD HAR ANTAGIT FÖLJANDE GEMENSAMMA STÅNDPUNKT
med beaktande av Fördraget om Europeiska unionen, särskilt artiklarna 15 och 34 i detta, och
av följande skäl:
(1) Europeiska rådet förklarade vid sitt extra möte den 21 september 2001 att terrorismen är en verklig utmaning för världen och Europa och att kampen mot terrorismen skall vara ett prioriterat mål för Europeiska unionen.
(2) Den 28 september 2001 antog Förenta nationernas säkerhetsråd resolution 1373(2001), i vilken omfattande strategier läggs fram för att bekämpa terrorism och i synnerhet finansieringen av terrorism.
(3) Den 8 oktober 2001 bekräftade rådet unionens beslutsamhet att i nära samarbete med Förenta staterna angripa terrorismens finansieringskällor.
(4) I enlighet med FN:s säkerhetsråds resolution 1333(2000) antog rådet den 26 februari 2001 gemensam ståndpunkt 2001/154/GUSP(1), i vilken det bland annat föreskrivs att kapital som tillhör Usama Bin Ladin och med honom associerade individer och organ skall frysas. Följaktligen omfattas inte dessa individer och organ av denna gemensamma ståndpunkt.
(5) Europeiska unionen bör vidta ytterligare åtgärder för att genomföra FN:s säkerhetsråds resolution 1373/2001.
(6) Medlemsstaterna har till Europeiska unionen överlämnat den information som är nödvändig för att genomföra några av dessa extra åtgärder.
(7) Gemenskapens insatser är nödvändiga för att några av dessa extra åtgärder skall kunna genomföras, och det krävs även insatser från medlemsstaterna, särskilt när det gäller tillämpningen av former för polissamarbete och straffrättsligt samarbete.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Denna gemensamma ståndpunkt skall tillämpas i enlighet med bestämmelserna i följande artiklar på personer, grupper och enheter som deltar i terroristhandlingar och finns förtecknade i bilagan.
2. I denna gemensamma ståndpunkt avses med personer, grupper och enheter som deltar i terroristhandlingar:
- personer som begår eller försöker begå terroristhandlingar eller som deltar i eller underlättar genomförandet av terroristhandlingar,
- grupper och enheter som ägs eller kontrolleras direkt eller indirekt av sådana personer och personer, grupper eller enheter som agerar på sådana personers, gruppers eller enheters vägnar eller under deras ledning, inklusive kapital som härrör från eller uppstår genom egendom som direkt eller indirekt ägs eller kontrolleras av sådana personer och av associerade personer, grupper och enheter.
3. I denna gemensamma ståndpunkt avses med terroristhandling: en av följande avsiktliga handlingar som på grund av sin art eller sitt sammanhang allvarligt kan skada ett land eller en internationell organisation och som definieras som ett brott enligt nationell lagstiftning och begås i syfte att
i) injaga allvarlig fruktan hos en befolkning,
ii) otillbörligen tvinga ett offentligt organ eller en internationell organisation att utföra eller att avstå från att utföra en viss handling, eller
iii) allvarligt destabilisera eller förstöra de grundläggande politiska, konstitutionella, ekonomiska eller sociala strukturerna i ett land eller i en internationell organisation:
a) angrepp mot en persons liv som kan leda till döden,
b) allvarliga angrepp på en persons fysiska integritet,
c) människorov eller tagande av gisslan,
d) förorsakande av omfattande förstörelse av en regeringsanläggning eller offentlig anläggning, transportsystem, infrastruktur, inklusive datasystem, en fast plattform belägen på kontinentalsockeln, en offentlig plats eller privat egendom som sannolikt kommer att förorsaka att människoliv utsätts för fara eller leda till betydande ekonomiska förluster,
e) kapning av luftfartyg och fartyg eller andra kollektiva transportmedel eller godstransporter,
f) tillverkning, innehav, förvärv, transport, tillhandahållande eller användning av skjutvapen, sprängämnen eller kärnvapen, av biologiska eller kemiska vapen, samt, när det gäller biologiska och kemiska vapen, forskning och utveckling,
g) utsläpp av farliga ämnen eller orsakande av brand, explosioner eller översvämningar som kan förorsaka att människoliv utsätts för fara,
h) att störa eller avbryta försörjningen av vatten, elkraft eller andra grundläggande naturresurser som kan förorsaka att människoliv utsätts för fara,
i) hot om att utföra någon av de handlingar, som räknas upp i a-h,
j) att leda en terroristgrupp,
k) att delta i en terroristgrupps verksamhet, vari inbegrips att förse den med upplysningar eller ge den materiellt stöd eller bidra med vilken form av finansiering som helst av denna verksamhet, med kännedom om att deltagandet kommer att bidra till gruppens brottsliga verksamhet.
I denna punkt avses med %quot%terroristgrupp%quot% en strukturerad grupp, inrättad för en viss tid, bestående av mer än två personer som handlar i samförstånd för att begå terroristhandlingar. Med strukturerad grupp avses: en grupp som inte tillkommit slumpartat i det omedelbara syftet att begå en terroristhandling och som inte nödvändigtvis har formellt fastställda roller för medlemmarna, kontinuitet i sammansättningen eller en noggrant utarbetad struktur.
4. Förteckningen i bilagan skall upprättas på grundval av exakta uppgifter eller fakta i det relevanta ärendet som visar att ett beslut har fattats av en behörig myndighet beträffande de personer, grupper eller enheter som avses, oavsett om det gäller inledande av undersökningar eller rättsliga åtgärder i fråga om en terroristhandling, försök att begå, deltaga i eller underlätta en sådan handling, grundat på bevis eller allvarliga och trovärdiga indicier eller en dom för sådana handlingar. Personer, grupper och enheter som enligt FN:s säkerhetsråd är knutna till terrorism eller mot vilka säkerhetsrådet har utfärdat sanktioner kan ingå i förteckningen.
I denna punkt avses med behörig myndighet: en rättslig myndighet eller, om rättsliga myndigheter inte har behörighet på det område som omfattas av denna punkt, en likvärdig myndighet som är behörig på det området.
5. Rådet skall se till att namnen på fysiska eller juridiska personer, grupper eller enheter i förteckningen i bilagan förses med tillräckliga detaljer för att enskilda individer, juridiska personer, enheter eller organ med säkerhet skall kunna identifieras och att de som har samma eller liknande namn lättare skall kunna rentvås.
6. Namnen på de personer och enheter som finns i förteckningen i bilagan skall ses över med jämna mellanrum minst en gång var sjätte månad för att man skall försäkra sig om att det är berättigat att behålla dem i förteckningen.
Artikel 2
Europeiska gemenskapen, som handlar inom ramen för sina befogenheter enligt Fördraget om upprättandet av Europeiska gemenskapen, kommer att beordra att alla penningmedel och andra finansiella tillgångar eller ekonomiska resurser frysas för personer, grupper och enheter som finns i förteckningen i bilagan.
Artikel 3
Europeiska gemenskapen, som handlar inom ramen för sina befogenheter enligt Fördraget om upprättandet av Europeiska gemenskapen, skall se till att penningmedel, finansiella tillgångar eller ekonomiska resurser eller finansiella eller andra därmed besläktade tjänster varken direkt eller indirekt görs tillgängliga för personer, grupper och enheter som finns i förteckningen i bilagan.
Artikel 4
Medlemsstaterna skall genom polissamarbete och straffrättsligt samarbete inom ramen för avdelning VI i Fördraget om Europeiska unionen ge varandra största möjliga bistånd när det gäller att förhindra och bekämpa terroristhandlingar. Därför kommer de, med hänsyn till undersökningar och förfaranden som genomförs av deras myndigheter när det gäller någon av de personer, grupper och enheter som finns i förteckningen i bilagan, att på anmodan fullt ut utnyttja sina befintliga befogenheter i enlighet med Europeiska unionens rättsakter och andra internationella avtal, ordningar och konventioner som är bindande för medlemsstaterna.
Artikel 5
Denna gemensamma ståndpunkt får verkan samma dag som den antas.
Artikel 6
Denna gemensamma ståndpunkt skall ses över fortlöpande.
Artikel 7
Denna gemensamma ståndpunkt skall offentliggöras i Officiella tidningen.
Kommissionens direktiv 2001/2/EG
av den 4 januari 2001
om anpassning till den tekniska utvecklingen av rådets direktiv 1999/36/EG om transportabla tryckbärande anordningar
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 1999/36/EG av den 29 april 1999 om transportabla tryckbärande anordningar(1), särskilt artikel 14 i detta, och
av följande skäl:
(1) I artikel 3.1 i direktiv 1999/36/EG fastställs att nya kärl och nya tankar skall uppfylla de tillämpliga bestämmelserna i rådets direktiv 94/55/EG av den 21 november 1994 om tillnärmning av medlemsstaternas lagstiftning om transport av farligt gods på väg(2), senast ändrat genom Europaparlamentets och rådets direktiv 2000/61/EG(3), och att de skall uppfylla de tillämpliga bestämmelserna i rådets direktiv 96/49/EG av den 23 juli 1996 om tillnärmning av medlemsstaternas lagstiftning om transport av farligt gods på järnväg(4), senast ändrat genom Europaparlamentets och rådets direktiv 2000/62/EG(5).
(2) Bestämmelserna i europeiska överenskommelsen om internationell transport av farligt gods på väg (ADR) och reglementet om internationell järnvägsbefordran av farligt gods (RID)(6), och ändringarna av dessa, finns som bilagor till direktiv 94/55/EG och direktiv 96/49/EG. En ny version av ADR och RID kommer att träda i kraft den 1 juli 2001.
(3) I bilaga V till direktiv 1999/36/EG fastställs moduler för bedömning av överensstämmelse av nya kärl och tankar. Dessa bestämmelser överensstämmer inte längre med den nya versionen av ADR och RID. Följaktligen bör bilagan ändras.
(4) De ändringar som är nödvändiga för att anpassa bilagorna till direktiv 1999/36/EG skall antas i enlighet med artikel 14 i direktivet, i enlighet med förfarandet i artikel 15.
(5) De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från den kommitté som anges i artikel 15 i direktiv 1999/36/EG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till direktiv 1999/36/EG skall ersättas med bilagan till det här direktivet.
Artikel 2
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 1 juli 2001. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när det offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 3
Detta direktiv träder i kraft den sjunde dagen efter det att det har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
Europaparlamentets och rådets direktiv 2001/10/EG
av den 22 maj 2001
om ändring av rådets direktiv 91/68/EEG vad gäller scrapie
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 152.4 b i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
efter att ha hört med Regionkommittén,
i enlighet med förfarandet i artikel 251 i fördraget(3), och
av följande skäl:
(1) Djurhälsovillkoren i samband med scrapie, vilka reglerar avyttring av djur, fastställs i rådets direktiv 91/68/EEG av den 28 januari 1991 om djurhälsovillkor för handeln med får och getter inom gemenskapen(4).
(2) Kommissionen har erhållit vetenskapliga utlåtanden, framför allt från Vetenskapliga styrkommittén, om flera aspekter på transmissibel spongiform encefalopati (TSE). Bestämmelserna i direktiv 91/68/EEG bör omprövas mot bakgrund av dessa utlåtanden.
(3) Det bör fastställas bestämmelser för alla frågor i samband med TSE, särskilt de bestämmelser som skall tillämpas på framställning och avyttring av levande djur och animaliska produkter enligt artikel 1.1 i Europaparlamentets och rådets förordning (EG) nr 999/2001 av den 22 maj 2001 om fastställande av bestämmelser för förebyggande, kontroll och utrotning av vissa typer av transmissibel spongiform encefalopati(5).
(4) Detta direktiv avser direkt folkhälsan och hänför sig till den inre marknadens funktion. Följaktligen är det lämpligt att bibehålla artikel 152.4 b i fördraget som rättslig grund för bestämmelserna om förebyggande och bekämpning av vissa typer av transmissibel spongiform encefalopati.
(5) Direktiv 91/68/EEG bör ändras i enlighet med detta.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 91/68/EEG ändras på följande sätt:
1. I artikel 2.7 skall orden %quot%uppförd på förteckningen under avdelningarna I och II i bilaga B%quot% ersättas med orden %quot%uppförd på förteckningen i bilaga B, avdelning I%quot%.
2. Artikel 6 b skall utgå.
3. I artikel 7.1 skall orden %quot%som avses i bilaga B, avdelningarna II och III%quot% ersättas med orden %quot%som avses i bilaga B, avdelning III%quot%.
4. I artikel 8.1 skall orden %quot%som räknas upp i avdelningarna II och III i bilaga B%quot% ersättas med %quot%som räknas upp i bilaga B, avdelning III%quot%.
5. Avdelning II i bilaga B skall utgå.
Artikel 2
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 30 juni 2001. De skall genast underrätta kommissionen om detta.
De skall tillämpa dessa bestämmelser från och med den 1 juli 2001.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv. Kommissionen skall underrätta övriga medlemsstater om detta.
Artikel 3
Detta direktiv träder i kraft den tjugonde dagen efter det att det har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Artikel 4
Detta direktiv riktar sig till medlemsstaterna.
Kommissionens förordning (EG) nr 306/2001
av den 12 februari 2001
om klassificering av vissa varor i Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan(1), senast ändrad genom förordning (EG) nr 2559/2000(2), särskilt artikel 9 i denna, och
av följande skäl:
(1) För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovannämnda förordning, är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till denna förordning.
(2) I förordning (EEG) nr 2658/87 har allmänna regler fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
(3) Enligt dessa allmänna regler måste de varor som beskrivs i kolumn 1 i tabellen som är bifogad den här förordningen klassificeras enligt motsvarande KN-nummer i kolumn 2 med de motiveringar som ges i kolumn 3.
(4) Det är lämpligt att bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter avseende varuklassificeringen i Kombinerade nomenklaturen och som inte överensstämmer med de rättigheter som fastställs i denna förordning fortfarande kan åberopas av innehavaren enligt bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(3), senast ändrad genom Europaparlamentets och rådets förordning (EG) nr 2700/2000(4), under en period av tre månader.
(5) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Tullkodexkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 2
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
Artikel 3
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1370/2001
av den 5 juli 2001
om ändring av förordning (EG) nr 174/1999 om fastställande av särskilda tillämpningsföreskrifter till rådets förordning (EEG) nr 804/68 i fråga om exportlicenser och exportbidrag inom sektorn för mjölk och mjölkprodukter
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1255/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter(1), senast ändrad genom förordning (EG) nr 1670/2000(2), särskilt artikel 26.3 i denna, och
av följande skäl:
(1) I kommissionens förordning (EG) nr 174/1999(3), senast ändrad genom förordning (EG) nr 1202/2001(4), fastställs särskilda tillämpningsföreskrifter till rådets förordning (EEG) nr 804/68(5) i fråga om exportlicenser och exportbidrag inom sektorn för mjölk och mjölkprodukter. För att säkerställa en god förvaltning av ordningen med exportbidrag och minska risken för spekulation och störningar inom ordningen för vissa mjölkprodukter är det nödvändigt att höja den säkerhet som fastställs i nämnda förordning.
(2) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för mjölk och mjölkprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 9 i förordning (EG) nr 174/1999, skall ersättas med följande: %quot%Artikel 9
Beloppet för den säkerhet som avses i artikel 15.2 i kommissionens förordning (EG) nr 1291/2000(6) skall motsvara följande procentsats av det bidragsbelopp som fastställts för varje produktkod och som gäller på inlämningsdagen för ansökan om exportlicens:
a) 5 % för produkter enligt KN-nummer 0405,
b) 30 % för produkter enligt KN-nummer 0402 10,
c) 30 % för produkter enligt KN-nummer 0406,
d) 20 % för övriga produkter.
Säkerhetsbeloppet får emellertid aldrig underskrida 6 euro per 100 kg.
Det bidragbelopp som avses i första stycket skall vara det som beräknats för den totala mängden av den berörda produkten, förutom när det gäller mjölkprodukter med tillsats av socker.
För mjölkprodukter med tillsats av socker skall det bidragsbelopp som avses i första stycket beräknas genom att den sammanlagda mängden av hela den berörda produkten multipliceras med den bidragssats som gäller per kilo mjölkprodukt.%quot%
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Rådets förordning (EG) nr 1452/2001
av den 28 juni 2001
om specifika åtgärder för vissa jordbruksprodukter till förmån för de franska utomeuropeiska departementen, ändring av direktiv 72/462/EEG samt upphävande av förordning (EEG) nr 525/77 och förordning (EEG) nr 3763/91 (Poseidom)
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artiklarna 36 och 37 samt artikel 299.2 i detta,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande(1), och,
av följande skäl:
(1) På grund av de franska utomeuropeiska departementens avlägsna belägenhet och ökaraktär antog rådet genom beslut 89/687/EEG(2) ett särskilt åtgärdsprogram (Poseidom) för dessa departement inom ramen för gemenskapens politik till förmån för de yttersta randområdena. Syftet med programmet är att främja den ekonomiska och sociala utvecklingen i dessa områden och göra det möjligt för dem att dra nytta av fördelarna som erbjuds av den inre marknaden, som dessa områden tillhör, även om de befinner sig avsides både geografiskt och ekonomiskt. Programmet avser tillämpningen av den gemensamma jordbrukspolitiken i dessa områden och föreskriver att specifika åtgärder skall vidtas. Programmet föreskriver bland annat förbättring av möjligheterna till produktion och saluföring av de franska utomeuropeiska departementens jordbruksprodukter och lindring av de negativa effekterna av det speciella geografiska läget och övriga begränsningar, i enlighet med artikel 299.2 i fördraget.
(2) De franska utomeuropeiska departementens speciella geografiska läge i förhållande till försörjningskällorna för vissa basprodukter för bearbetning och som insatsvaror i jordbruket innebär ökade transportkostnader i dessa områden. Även andra faktorer som har samband med ökaraktären och läget i gemenskapens yttersta randområden begränsar ytterligare verksamheten för aktörer och producenter. Detta gäller särskilt försörjningen med spannmål, som knappast alls produceras och inte kan produceras i större mängder i dessa departement, som följaktligen är beroende av leveranser utifrån. Effekterna av dessa begränsningar kan lindras genom att priset på dessa basprodukter sänks. Således bör en särskild försörjningsordning införas för att garantera departementens försörjning genom den lokala produktionen och för att minska de merkostnader som uppstår till följd av områdenas avlägsna belägenhet, ökaraktär och läge i gemenskapens yttersta randområden.
(3) För detta ändamål, genom undantag från artikel 23 i fördraget, bör importen av produkter från tredje land befrias från tillämpliga importtullar.
(4) För att effektivt kunna uppnå målet att sänka priserna i de franska utomeuropeiska departementen samt lindra de merkostnader som uppstår till följd av den avlägsna belägenheten, ökaraktären och läget i gemenskapens yttersta randområden, men samtidigt bibehålla gemenskapsprodukternas konkurrenskraft, bör stöd beviljas för leverans av gemenskapsprodukter till departementen. Stödet kommer att ta hänsyn till ökade transportkostnader till departementen och exportpriser till tredje land samt, när det gäller insatsvaror i jordbruket eller produkter avsedda för bearbetning, till merkostnader till följd av departementens ökaraktär och läge i gemenskapens yttersta randområden.
(5) Eftersom de kvantiteter som omfattas av den särskilda försörjningsordningen är begränsade till de franska utomeuropeiska departementens försörjningsbehov stör systemet inte den inre marknadens funktion. De ekonomiska fördelarna med den särskilda försörjningsordningen bör inte leda till omläggning av handeln med de berörda produkterna. Det bör således vara förbjudet att vidaresända eller återexportera dessa produkter från departementen. Handelsflödena mellan departementen omfattas dock inte av detta förbud. Vid bearbetning gäller detta förbud på vissa villkor inte heller export till tredje länder för att främja regional handel eller traditionell export till den övriga gemenskapen.
(6) De ekonomiska fördelarna med den särskilda försörjningsordningen bör återverka på produktionskostnaderna ända fram till slutanvändaren. Stöd bör således beviljas endast på villkor att det har önskad effekt, och de nödvändiga kontrollerna bör genomföras.
(7) Med tanke på den senaste jordbruksutvecklingen i Franska Guyana har bestämmelser införts för att främja utvecklingen av risodlingen genom förordning (EEG) nr 3763/91(3). Bestämmelserna upphörde att gälla i slutet av regleringsåret 1996. Eftersom ingen förlängning har begärts av den berörda medlemsstaten har bestämmelserna upphävts. Det finns bestämmelser om avsättning och saluföring av en del av den lokala produktionen i Guadeloupe, Martinique och i övriga gemenskapen. Hela den lokala produktionen kan inte konsumeras på platsen, eftersom lagringsmöjligheterna är mycket begränsade och därför bör bestämmelserna, som är av yttersta vikt för balansen i den lokala produktions- och handelskedjan, bibehållas på samma villkor som i den gällande lagstiftningen.
(8) Traditionell animalieproduktion bör stödjas i syfte att tillgodose de lokala konsumtionsbehoven i de franska utomeuropeiska departementen. Undantag bör göras från vissa bestämmelser i de gemensamma organisationerna av marknaderna när det gäller begränsningar av produktionen så att hänsyn tas till utvecklingen och de särskilda lokala produktionsvillkoren som skiljer sig helt från den övriga gemenskapen. Detta mål kan understödjas genom finansiering av program för genetisk förbättring som omfattar inköp av renrasiga avelsdjur och inköp av raser som är bättre anpassade till de lokala förhållandena, genom beviljande av tillägg till am- och dikobidraget samt slaktbidraget, samt vid behov genom möjligheten att från tredje land importera handjur av nötkreatur för uppfödning under vissa villkor och bevilja undantag från tillämpningen av villkoren för import av djur och animaliska livsmedel.
(9) De bristfälliga villkoren för försörjning av den lokala marknaden i de franska utomeuropeiska departementen med färska mjölkprodukter, som nu för närvarande företrädesvis sker genom importerade produkter, bör åtgärdas. Detta mål kan genomföras, å ena sidan, genom fortsatt stöd till utvecklingen av komjölksproduktionen inom gränserna för de lokala konsumtionsbehoven vilka utvärderas inom ramen för en försörjningsbalans och, å andra sidan, genom att inte tillämpa systemet med tilläggsavgifter för producenterna av komjölk enligt förordning (EEG) nr 3950/92(4). De bristfälliga villkoren för försörjning som kännetecknar dessa yttersta randområden, helt annorlunda än de som råder i den övriga gemenskapen, liksom nödvändigheten att utveckla incitament till lokal produktion motiverar detta undantag.
(10) Ett gemenskapsbidrag har tillfälligt införts för perioden 1996-2000 för finansiering av regionala program på Martinique och Réunion för produktion och saluföring av lokala produkter inom djuruppfödnings- och mjölkproduktsektorerna. För de berörda sektorerna är täckningen av de lokala behoven fortsatt låg. Aktörernas möjlighet att utforma och genomföra strategier som är anpassade till de lokala förhållandena i fråga om ekonomisk utveckling, fysisk planering av produktionen och branschkunskaper förutsätter möjligheten att effektivt kunna uppbåda gemenskapsstöd. Stödet bör tillfälligt fortsätta så att produktionen kan utvecklas till en högkvalitativ och modern sektor. Denna bestämmelse bör utökas till att omfatta Franska Guyana och Guadeloupe under förutsättning att branschorganisationer etablerar sig lokalt.
(11) När det gäller frukt, grönsaker, växter och blommor har åtgärder vidtagits för att förbättra jordbruksföretagens produktivitet och produkternas kvalitet, strukturera sektorerna, utveckla produkter som bearbetas lokalt och för att stödja vissa traditionella produktioner (vanilj, oljor m.m.) till förmån för den lokala saluföringen av dessa produkter, samt bearbetning och extern saluföring av dem. Eftersom dessa åtgärder har gjort det möjligt att förstärka den lokala produktionens konkurrenskraft gentemot yttre konkurrens från tillväxtmarknader, bättre motsvara konsumenternas och nya distributionskedjors förväntningar och se till att dessa produkter marknadsförs i den övriga gemenskapen, bör dessa ansträngningar fortsätta.
(12) Genom förordning (EEG) nr 525/77(5) införs en stödordning för produktion av konserverad ananas som endast har tillämpats på Martinique. För att uppnå en harmoniserad lagstiftning och administration bör detta system, med beaktande av systemets och produktionsområdets särdrag, integreras i den här förordningen. Förordning (EEG) nr 525/77 bör således upphöra att gälla. Ananassektorn kan endast bevaras genom att alla sektorns aktörer medverkar. Ananasproduktionen är särskilt viktig för Martinique i både ekonomiskt och socialt hänseende. Med produktionen följer höga kostnader och de bearbetade produkterna utsätts för konkurrens från tredje land. Man bör se till att bearbetningsindustrin får fortsatt stöd, att de små jordbruksföretagen fortlever, att försörjningen av industrin säkerställs, att producentorganisationernas roll förstärks och samtidigt göra det möjligt att på medellång sikt styra produktionen mot bättre lönsamhet samt eventuellt mot saluföring av färska produkter.
(13) Rörsockersektorn är central för de franska utomeuropeiska departementens ekonomi. Departementens nackdelar är betydande (avlägsen belägenhet, ökaraktär, läge i gemenskapens yttersta randområden, bergsnatur, småskaliga och utspridda jordbruksföretag, litet antal fabriker, höga lokala transportkostnader, otillräckligt vägnät) och innebär merkostnader. Det finns också särskilda nackdelar jämfört med fastlandsproduktionen av sockerbetor, i synnerhet i fråga om insamlingen av sockerrör. För att se till att sektorn utvecklas på ett bra sätt och för att minska dessa svårigheter bör åtgärder vidtas för att delvis kompensera merkostnaderna i fråga om transport av sockerrören från fälten till uppsamlingscentralerna.
(14) Rom är en produkt vars ekonomiska betydelse och avsättningsmöjligheter är av yttersta vikt för de franska utomeuropeiska departementen. Ett gradvist avskaffande av de nuvarande förmåner som kommer romproduktionen till del skulle få allvarliga följder för producenternas inkomster. Främst bör åtgärder vidtas för stöd till sockerrörsodlingen och den direkta bearbetningen till jordbruksrom och sockerrörssaft i så måtto som detta har en positiv effekt för bibehållande av produktionen av sockerrör som levereras till destillerier, som på så sätt får möjlighet att planera och rationalisera investeringar i produktionsutrustning, påverka ersättningen till odlaren och uppmuntras att förbättra sin produktionsutrustning så att avkastningen och kvaliteten på de levererade sockerrören kan garanteras.
(15) Jordbruksproducenterna i de franska utomeuropeiska departementen bör uppmuntras att leverera kvalitetsprodukter, och avsättningen av dessa produkter bör stödjas. För detta ändamål kan gemenskapens grafiska symbol användas.
(16) Jordbruksproduktionen i de franska utomeuropeiska departementen har särskilda växtskyddsproblem som hänger samman med klimatförhållandena och med bristen på resurser för bekämpning. Det bör genomföras bekämpningsprogram mot skadliga organismer, även med biologiska metoder. Ett ekonomiskt stöd från gemenskapen bör fastställas för genomförandet av programmen.
(17) I förordning (EG) nr 1257/1999(6) fastställs de åtgärder för utveckling av landsbygden som kan berättiga till stöd från gemenskapen samt villkoren för att erhålla detta stöd.
(18) Denna förordning syftar till att kompensera för de ogynnsamma betingelser som har sin grund i de franska utomeuropeiska departementens avlägsna belägenhet och ökaraktär samt förbättra villkoren för produktion och saluföring av deras jordbruksprodukter.
(19) Vissa jordbruksföretag eller bearbetnings- och saluföringsföretag i de franska utomeuropeiska departementen uppvisar allvarliga strukturella brister, vilket leder till särskilda svårigheter. För vissa typer av investeringar bör undantag därför kunna beviljas från de bestämmelser som begränsar eller förhindrar beviljandet av vissa strukturstöd enligt förordning (EG) nr 1257/1999.
(20) Enligt artikel 29.3 i förordning (EG) nr 1257/1999 skall stödet till skogsbruk endast beviljas för skogar och arealer som ägs av privata ägare, deras sammanslutningar, eller av kommuner och sammanslutningar av kommuner. Större delen av skogarna och skogsarealerna i de franska utomeuropeiska departementen ägs av andra offentliga myndigheter än kommuner. Villkoren i nämnda artikel bör därför mjukas upp.
(21) Gemenskapens medfinansiering av tre av de kompletterande åtgärderna i artikel 35.1 i förordning (EG) nr 1257/1999 får uppgå till 85 % av den totala stödberättigande kostnaden i de yttersta randområdena. Enligt artikel 47.2 tredje strecksatsen i samma förordning skall däremot gemenskapens medfinansiering av de åtgärder för miljövänligt jordbruk som utgör den fjärde kompletterande åtgärden begränsas till 75 % för alla områden som omfattas av mål 1. Med tanke på den betydelse som miljövänligt jordbruk tillskrivs i samband med landsbygdsutvecklingen bör nivån på gemenskapens medfinansiering harmoniseras för alla kompletterande åtgärder i de yttersta randområdena.
(22) Varje plan, ram för gemenskapsstöd, operativt program eller samlat programdokument skall i enlighet med artikel 14 i förordning (EG) nr 1260/1999(7) omfatta en period på sju år, och programperioden skall inledas den 1 januari 2000. Av konsekvensskäl och för att undvika en diskriminering av stödmottagare som omfattas av samma program bör de undantag som föreskrivs i denna förordning i undantagsfall kunna tillämpas för hela denna programperiod.
(23) Ett undantag får beviljas från kommissionens bestämda politik att inte tillåta statligt stöd till driften inom produktionssektorn och till bearbetning och saluföring av jordbruksprodukter som omfattas av bilaga I till fördraget, för att lindra effekterna av de särskilda begränsningar som jordbruksproduktionen i de franska utomeuropeiska departementen utsätts för på grund av deras avlägsna belägenhet, ökaraktär, läge i gemenskapens yttersta randområden, ringa storlek, besvärliga terräng- och klimatförhållanden samt ekonomiska beroende av ett fåtal produkter.
(24) Övergångsbestämmelser bör kunna antas för att underlätta övergången från de ordningar som fastställs i förordning (EEG) nr 3763/91 och i förordning (EEG) nr 525/77 till den nya ordning som fastställs i den här förordningen och för att se till att det inte uppstår några avbrott vid en eventuell förlängning av de befintliga åtgärderna.
(25) De åtgärder som krävs för att genomföra denna förordning bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(8).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I denna förordning fastställs specifika åtgärder för att med avseende på vissa jordbruksprodukter avhjälpa de svårigheter som beror på de franska utomeuropeiska departementens avlägsna belägenhet, läge i gemenskapens yttersta randområden och ökaraktär.
AVDELNING I
SÄRSKILD FÖRSÖRJNINGSORDNING
Artikel 2
1. Härmed inrättas en särskild försörjningsordning för de jordbruksprodukter som finns förtecknade i bilaga I och som är nödvändiga i de franska utomeuropeiska departementen som livsmedel, för bearbetning och som insatsvaror i jordbruket.
2. Genom en prognostiserad försörjningsbalans skall de årliga försörjningsbehoven beräknas i fråga om produkterna i bilaga I. En separat prognos kan göras för att bedöma bearbetnings- och förpackningsindustrins behov av produkter för den lokala marknaden och för export, på vissa villkor till tredje länder eller traditionella sändningar till den övriga gemenskapen.
Artikel 3
1. Tullar skall inte tillämpas vid direktimport till de franska utomeuropeiska departementen av produkter som omfattas av den särskilda försörjningsordningen, och som kommer från tredje land, inom ramen för den kvantitetsbegränsning som fastställs i försörjningsbalansen.
2. För att säkerställa de behov som fastställts i enlighet med artikel 2 vad beträffar mängd, pris och kvalitet och för att bevara den del av försörjningen som kommer från gemenskapen skall ett stöd beviljas för försörjning av de franska utomeuropeiska departementen med produkter med ursprung i gemenskapen och som förvaras i offentliga interventionslager eller finns tillgängliga på gemenskapsmarknaden.
Stödbeloppet skall fastställas med hänsyn till merkostnaderna för transport till de franska utomeuropeiska departementen och exportpriser till tredje land samt, när det gäller produkter avsedda för bearbetning eller insatsvaror i jordbruket, till merkostnader till följd av departementens ökaraktär och läge i gemenskapens yttersta randområden.
3. Den särskilda försörjningsordningen skall genomföras på ett sätt som särskilt tar hänsyn till
- de franska utomeuropeiska departementens specifika behov och, när det gäller produkter avsedda för bearbetning eller insatsvaror i jordbruket, de speciella kvalitetskraven,
- handeln med den övriga gemenskapen,
- den ekonomiska aspekten av de planerade stöden.
4. Den särskilda försörjningsordningen skall tillämpas under förutsättning att de förmåner som följer av befrielsen från importtullar eller, när det gäller försörjning från den övriga gemenskapen, av stöd, faktiskt kommer slutanvändaren till godo.
5. De produkter som omfattas av den särskilda försörjningsordningen får inte återexporteras till tredje land eller sändas tillbaka till den övriga gemenskapen. Förbudet i denna punkt skall inte gälla handeln mellan de franska utomeuropeiska departementen.
Om produkterna bearbetas i departementen skall detta förbud inte gälla export till tredje länder eller traditionella sändningar till den övriga gemenskapen av de bearbetade produkterna, enligt villkor som skall fastställas av kommissionen i enlighet med förfarandet i artikel 23.2.
Inget exportbidrag skall beviljas.
6. Tillämpningsföreskrifter för denna avdelning skall fastställas i enlighet med förfarandet i artikel 23.2. De skall särskilt omfatta
- fastställande av stöden för försörjning från gemenskapen,
- bestämmelser för att säkerställa att förmånerna kommer slutanvändaren till godo,
- införande av ett system för import- eller leveranslicenser vid behov.
Kommissionen skall i enlighet med förfarandet i artikel 23.2 upprätta försörjningsbalanser; enligt samma förfarande får kommissionen se över dessa balanser samt förteckningen över produkter i bilaga I beroende på hur de franska utomeuropeiska departementens behov förändras.
Artikel 4
Inom ramen för en årlig kvantitet på 8000 ton skall den avgift som fastställs enligt artiklarna 10 och 11 i förordning (EEG) nr 1766/92(9) inte tillämpas på import till ön Réunion av vetekli enligt KN-nummer 2302 30 med ursprung i AVS-stater.
AVDELNING II
ÅTGÄRDER FÖR LOKAL PRODUKTION
KAPITEL I
RIS
Artikel 5
1. Gemenskapsstöd skall beviljas, inom ramen för en årlig volym om 12000 ton ris uttryckt som helt slipat ris, för ris skördat i Franska Guyana som är föremål för årskontrakt som avser avsättning och saluföring i Guadeloupe och Martinique samt i den övriga gemenskapen. För avsättning och saluföring i övriga gemenskapen skall stöd betalas ut för en volym på högst 4000 ton.
Sådana kontrakt skall ingås mellan producenter i Franska Guyana, å ena sidan, och fysiska eller juridiska personer som är etablerade i Guadeloupe, Martinique eller den övriga gemenskapen, å andra sidan.
Stödbeloppet skall uppgå till 10 % av värdet av den produktion som avsätts i Guadeloupe, Martinique eller den övriga gemenskapen, för en vara som levererats i den första lossningshamnen. Procentsatsen skall höjas till 13 % om den ena kontraktsparten är en sammanslutning eller en förening av producenter.
Stödet skall betalas ut till den köpare som saluför produkterna enligt årskontraktet.
2. Tillämpningsföreskrifter för denna artikel skall antas i enlighet med förfarandet i artikel 23.2. Enligt samma förfarande kan kommissionen se över den årliga volym om 12000 ton som avses i punkt 1 första stycket.
KAPITEL II
DJURUPPFÖDNING OCH MJÖLKPRODUKTER
Artikel 6
1. Inom djuruppfödningssektorn skall stöd beviljas för leverans till de franska utomeuropeiska departementen av renrasiga djur och raser för handelsbruk samt produkter med ursprung i gemenskapen.
2. Villkoren för beviljande av stöd skall fastställas främst med hänsyn till de franska utomeuropeiska departementens försörjningsbehov för att få igång produktion av olika slag, genetisk förbättring av djurbesättningar och raser som är bäst anpassade till de lokala förhållandena. Stödet skall betalas ut för leverans av varor som uppfyller gemenskapsbestämmelsernas krav.
3. Stöden skall fastställas med beaktande av
- försörjningsförhållandena för de franska utomeuropeiska departementen till följd av det geografiska läget, särskilt när det gäller kostnader,
- varornas priser på gemenskapsmarknaden och på världsmarknaden,
- om tullar tas ut vid import från tredje land eller ej,
- den ekonomiska aspekten av de planerade stöden.
4. Artikel 3.4 och 3.5 skall tillämpas på varor för vilka stöd beviljas enligt punkt 1 i den här artikeln.
5. Såväl tillämpningsföreskrifter för den här artikeln som förteckningen över de produkter och stödbelopp som avses i punkt 1 skall fastställas i enlighet med förfarandet i artikel 23.2.
Artikel 7
1. Till dess att det lokala beståndet av unga nötkreatur av hankön har blivit tillräckligt stort för att säkerställa utvecklingen av den lokala köttproduktionen, och inom den begränsning som avses i artikel 9, skall möjligheten införas att importera nötkreatur med ursprung i tredje land för uppfödning på plats och för konsumtion i de franska utomeuropeiska departementen, utan att de tullar som avses i artikel 30 i förordning (EG) nr 1254/1999(10) tillämpas.
Artikel 3.4 och 3.5 skall tillämpas på de djur som omfattas av den befrielse från tullar som avses i första stycket i den här punkten.
2. Antalet djur som omfattas av den befrielse från tullar som avses i punkt 1 skall, när importbehovet är motiverat, fastställas med hänsyn till utvecklingen av den lokala produktionen. Antalet djur samt tillämpningsföreskrifter för denna artikel, som bland annat skall omfatta en minimiperiod för uppfödning, skall fastställas i enlighet med förfarandet i artikel 23.2. Dessa djur är först och främst avsedda för producenter som innehar minst 50 % av göddjuren av lokalt ursprung.
Artikel 8
I direktiv 72/462/EEG(11) skall följande artikel införas: %quot%Artikel 31a
Utan att det påverkar tillämpningen av artikel 13 i direktiv 91/496/EEG(12) får kommissionen, i enlighet med förfarandet i artikel 29 i det här direktivet, göra undantag från bestämmelserna i det här direktivet när det gäller import till de franska utomeuropeiska departementen(13).
När sådana beslut som avses i första stycket antas skall de regler som skall tillämpas efter importen fastställas i enlighet med samma förfarande.%quot%
Artikel 9
1. För att främja traditionell verksamhet och kvalitetsförbättrande åtgärder inom nötköttsproduktionen inom ramen för konsumtionsbehoven i de franska utomeuropeiska departementen enligt beräkning i en regelbundet upprättad försörjningsbalans, skall stöd beviljas enligt punkterna a och b i andra stycket.
Försörjningsbalansen skall också omfatta djur som levererats med tillämpning av artiklarna 6 och 7.
a) Ett tillägg till am- och dikobidraget i artikel 6 i förordning (EG) nr 1254/1999 skall betalas ut till nötköttsproducenter. Detta tillägg skall uppgå till 50 euro för varje am- eller diko som producenten håller den dag ansökan lämnas in.
b) Ett tillägg till slaktbidraget i artikel 11 i förordning (EG) nr 1254/1999 skall betalas ut till nötköttsproducenter. Detta tillägg skall vara 25 euro per djur.
2. Bestämmelserna om
a) det regionala tak som införs genom artikel 4 i förordning (EG) nr 1254/1999, när det gäller det särskilda bidraget,
b) det individuella tak för sådana djur som hålls på företaget och som införs genom artikel 6 i förordning (EG) nr 1254/1999, när det gäller grundbidraget för am- och dikor,
c) det nationella tak som införs genom artikel 11 i förordning (EG) nr 1254/1999, när det gäller det särskilda grundbidraget för slakt,
d) den djurtäthetsfaktor på jordbruksföretag som införs genom artikel 12 i förordning (EG) nr 1254/1999,
skall inte tillämpas i de franska utomeuropeiska departementen, varken när det gäller det särskilda bidraget, grundbidraget för am- och dikor, grundbidraget för slakt eller de tilläggsbidrag som avses i punkt 1 a och b i den här artikeln.
3. De grund- och tilläggsbidrag som avses i punkt 1 skall varje år beviljas för högst 10000 handjur av nötkreatur, 35000 am- och dikor och 20000 slaktade djur.
4. Tillämpningsföreskrifter för denna artikel skall antas i enlighet med förfarandet i artikel 23.2. De skall innefatta upprättandet av de försörjningsbalanser som avses i punkt 1 i den här artikeln samt eventuell översyn till följd av utvecklingen av behoven.
a) För det särskilda bidraget för handjur av nötkreatur skall det i dessa föreskrifter anges
- en %quot%frysning%quot%, inom ett regionalt tak enligt artikel 4 i förordning (EG) nr 1254/1999, av det antal djur för vilka särskilt bidrag i de franska utomeuropeiska departementen beviljades år 1994,
- beviljande av bidrag, dock för högst nittio djur per åldersgrupp, kalenderår och företag.
b) För am- och dikobidraget skall det i föreskrifterna
- finnas bestämmelser för att, i den mån det behövs, säkerställa rättigheterna för de producenter som beviljats bidrag med tillämpning av artikel 6 i förordning (EG) nr 1254/1999,
- anges att en särskild reserv skall upprättas för de franska utomeuropeiska departementen samt anges särskilda villkor för tilldelning eller omfördelning av rättigheter, med hänsyn till de mål som eftersträvas för djuruppfödningen; reservens storlek skall bestämmas i förhållande till det tak som fastställs i punkt 3 och till det antal bidrag som beviljades år 1994.
c) För det särskilda slaktbidraget skall det föreskrivas
- en %quot%frysning%quot%, inom ett nationellt tak enligt artikel 38.1 i förordning (EG) nr 2342/1999(14), av det antal djur för vilka slaktbidrag beviljades år 2000.
Tillämpningsföreskrifterna kan innehålla ytterligare villkor för beviljande av tilläggsbidrag.
Kommissionen får enligt samma förfarande se över de tak som avses i punkt 3.
Artikel 10
1. Stöd för utveckling av komjölksproduktion skall beviljas inom ramen för de franska utomeuropeiska departementens behov av mjölkprodukter som livsmedel för varje regleringsår enligt beräkning i en försörjningsbalans. Mjölk som används för tillverkning av skummjölk till djurfoder är inte stödberättigande.
Stödet skall beviljas producenter eller producentgrupper för de mängder som levereras till mejerierna. Stödet skall betalas ut via mejerierna.
Stödet skall uppgå till 8,45 euro per 100 kilogram helmjölk.
Stödet skall betalas ut varje år för högst 40000 ton mjölk.
2. Den tilläggsavgift för producenter av komjölk som införs genom förordning (EEG) nr 3950/92 skall inte tillämpas i de franska utomeuropeiska departementen.
3. Kommissionen skall i enlighet med förfarandet i artikel 23.2 fastställa tillämpningsföreskrifter för denna artikel samt den försörjningsbalans som avses i punkt 1 i den artikeln.
Enligt samma förfarande får kommissionen se över den högsta kvantitet som avses i punkt 1 fjärde stycket.
Artikel 11
1. Under perioden 2001-2006 skall ett stöd beviljas för genomförandet av övergripande stödprogram för produktion och saluföring av lokala produkter inom djuruppfödnings- och mjölkproduktsektorerna i departementen Martinique och Réunion. Under 2001 skall stödet beviljas för årliga övergångsprogram. De övergripande programmen skall ha en varaktighet på fem år under perioden 2002-2006.
Programmen får omfatta stimulansåtgärder för förbättringar av kvalitet och hygien, saluföring, strukturering av sektorer, rationalisering av strukturer för produktion och saluföring, information på lokal nivå om kvalitetsprodukter och genomförande av tekniskt stöd. Programmen får inte omfatta beviljande av stöd utöver de bidrag som betalas ut med tillämpning av artiklarna 9 och 10.
Programmen skall utarbetas och genomföras i nära samråd mellan de behöriga myndigheter som medlemsstaten utsett och de erkända branschorganisationer som är mest representativa för de berörda ekonomiska sektorerna.
2. Tillämpningsföreskrifter för denna artikel skall fastställas i enlighet med förfarandet i artikel 23.2. De behöriga myndigheterna skall till kommissionen överlämna programprojekt med en varaktighet på högst fem år; kommissionen skall godkänna dem i enlighet med förfarandet i artikel 23.2. Enligt samma förfarande får kommissionen låta denna artikel omfatta departementen Guadeloupe och Franska Guyana, under förutsättning att branschorganisationer etablerar sig där.
3. De franska myndigheterna skall varje år lägga fram en rapport om genomförandet av programmen. Före utgången av 2005 skall kommissionen för Europaparlamentet och rådet lägga fram en utvärderingsrapport om tillämpningen av den åtgärd som avses i denna artikel, eventuellt tillsammans med lämpliga förslag.
KAPITEL III
FRUKT, GRÖNSAKER, VÄXTER OCH BLOMMOR
Artikel 12
1. Stöd skall beviljas för frukt, grönsaker, blommor och levande växter som anges i kapitlen 6, 7 och 8 i Kombinerade nomenklaturen, peppar enligt KN-nummer 0904 samt kryddor enligt KN-nummer 0910 vilka skördats i de franska utomeuropeiska departementen och är avsedda för försörjning av marknaderna i departementen. För Martinique och Guadeloupe skall detta stöd inte beviljas för andra bananer än mjölbananer enligt KN-nummer 0803 00 11.
Stödet skall beviljas för produkter som uppfyller de gemensamma normer som fastställs i gemenskapslagstiftningen eller, om sådana saknas, som överensstämmer med de detaljerade beskrivningar som ingår i leveransavtalen.
Stödet skall beviljas om leveransavtal för ett eller flera regleringsår ingåtts mellan å ena sidan enskilda producenter, producentgrupper eller de producentorganisationer som avses i artiklarna 11, 13 och 14 i förordning (EG) nr 2200/96(15) och å andra sidan aktörer inom distributions- eller restaurangsektorn eller sammanslutningar.
Stödet skall betalas ut till ovannämnda enskilda producenter, producentgrupper eller producentorganisationer inom ramen för de kvantiteter som årligen fastställs för varje produktkategori.
Stödbeloppet skall fastställas som ett schablonbelopp för varje produktkategori enligt de berörda produkternas medelvärde. Det skall differentieras beroende på om det gäller en av de producentorganisationer som avses i artiklarna 11, 13 och 14 i förordning (EG) nr 2200/96 eller någon annan stödmottagare.
2. Ett stöd om 6,04 euro per kilogram skall beviljas för produktion av grön vanilj enligt KN-nummer 0905 00 00 ämnad för produktion av torkad vanilj (svart) eller vaniljextrakt.
Stödet skall betalas ut för en årlig maximikvantitet om 75 ton.
3. Ett stöd om 44,68 euro per kilogram skall beviljas för produktion av pelargon- och vetiveriaoljor enligt KN-nummer 3301 21 respektive 3301 26.
Stödet skall betalas inom ramen för en årlig maximikvantitet om 30 ton pelargonolja och 5 ton vetiveriaolja.
4. Tillämpningsföreskrifter för denna artikel skall fastställas i enlighet med förfarandet i artikel 23.2. Samma förfarande skall användas för att fastställa de produktkategorier och stödbelopp som avses i punkt 1 i den här artikeln, och vid behov skall de maximikvantiteter som avses i punkterna 2 och 3 i den artikeln.
Artikel 13
1. Stöd skall beviljas för produktion av bearbetade frukter och grönsaker som framställts av produkter som skördats i de franska utomeuropeiska departementen.
Produktionsstödet skall betalas ut till bearbetningsföretag som åt producenten betalat minst ett minimipris för råvaran enligt avtal mellan å ena sidan producenterna eller deras erkända organisationer i enlighet med förordning (EG) nr 2200/96, och å andra sidan bearbetningsföretagen eller deras i laglig ordning stiftade föreningar eller sammanslutningar. Medlemsstaten skall fastställa ett minimipris för råvaran enligt produktionskostnaderna för denna.
2. Stödbeloppet skall fastställas som ett schablonbelopp för varje produktkategori på grundval av priset för den lokala råvara som används samt priset för import av samma råvara.
3. Stödet skall betalas ut inom ramen för den mängd som årligen fastställs för varje produktkategori.
4. En förteckning över bearbetade produkter för vilka stöd beviljas samt tillämpningsföreskrifter för denna artikel skall fastställas i enlighet med förfarandet i artikel 23.2. Samma förfarande skall användas för att fastställa de produktkategorier och stödbelopp som avses i punkt 2 i den här artikeln, samt de maximikvantiteter som avses i punkt 3.
Artikel 14
1. De franska myndigheterna skall för kommissionen lägga fram ett stödprogram för ananassektorn på Martinique.
Programmet skall omfatta stimulansåtgärder för förbättring av villkoren för produktion, saluföring och bearbetning av ananas och skall också bidra till att förstärka sektorns konkurrenskraft och understödja dess omstrukturering samt till att bevara småföretagen. Ananas som odlas på Martinique omfattas inte av stöd som betalas ut enligt artikel 13.
2. Programprojekten, som högst får pågå under fem år, skall läggas fram för kommissionen av de franska myndigheterna tillsammans med en genomföranderapport för föregående program, och de skall godkännas i enlighet med förfarandet i artikel 23.2.
Artikel 15
1. Stöd skall beviljas för ingående av årskontrakt om avsättning och saluföring av de produkter som avses i artikel 12.1. Detta stöd skall betalas ut inom ramen för en handelsvolym om högst 3000 ton per produkt, år och departement.
Avtalen skall ingås mellan å ena sidan de producenter eller producentorganisationer som avses i artiklarna 11, 13 och 14 i förordning (EG) nr 2200/96 och å andra sidan fysiska eller juridiska personer som är etablerade i den övriga gemenskapen.
2. Stödbeloppet skall vara 10 % av den saluförda produktionens värde, fritt bestämmelseorten.
3. Stödet skall beviljas uppköpare som förbinder sig att saluföra produkter från departementen som omfattas av sådana kontrakt som avses i punkt 1.
4. Om de åtgärder som avses i punkt 1 vidtas av gemensamma företag som har bildats av producenter, producentsammanslutningar eller producentföreningar i dessa departement, eller fysiska eller juridiska personer som är etablerade inom den övriga gemenskapen, i syfte att saluföra produkter som skördats i departementen, och om parterna förbinder sig att under en period om minst tre år gemensamt utnyttja det kunnande och den kompetens som krävs för att uppnå företagets mål, skall det stödbelopp som anges i punkt 2 höjas till 13 % av värdet av den produktion som gemensamt avsätts varje år.
5. Stöd enligt denna artikel skall också betalas ut, enligt villkor som fastställs i punkterna 1-4,
- för bearbetade produkter av frukt och grönsaker som skördats i departementen,
- för pelargon- och vetiveriaolja enligt KN-nummer 3301 21 respektive 3301 26,
- för torkad (svart) vanilj enligt KN-nummer ex 0905 00 00 samt för vaniljextrakt enligt KN-nummer 3301 90 90,
som är föremål för årskontrakt som avser avsättning och saluföring.
6. För meloner med KN-nummer ex 0807 19 00 och ananas med KN-nummer ex 0804 30 00 kan stöd dock beviljas i ett departement för en mängd som överstiger 3000 ton, om den totala stödberättigande mängden för samtliga departement inte överskrids.
7. Tillämpningsföreskrifter för denna artikel skall fastställas i enlighet med förfarandet i artikel 23.2.
KAPITEL IV
SOCKER OCH SEKTORN FÖR SOCKERRÖR, SOCKER OCH ROM
Artikel 16
1. Ett stöd för transport av sockerrör från skördeplatsen till uppsamlingscentralerna skall beviljas de producenter för vilka behöriga organ som skall utses av medlemsstaten har dokumenterat leveranser till bearbetningsindustrin.
2. Stödbeloppet skall fastställas enligt avstånd och andra objektiva kriterier som berör transporten; det får inte överskrida hälften av transportkostnaderna per ton som schablonmässigt har fastställts av de franska myndigheterna i varje departement.
Artikel 17
1. Stöd skall beviljas för direkt bearbetning av sockerrör som producerats i de franska utomeuropeiska departementen till sockerrörssaft eller jordbruksrom enligt definitionen i artikel 1.4 a 2 i förordning (EEG) nr 1576/89(16).
Stödet skall, beroende på situationen, betalas ut till producenten av sockerrörssaft eller till destillatören förutsatt att denne betalat sockerrörsproducenten ett lägsta pris som skall fastställas.
2. Stödet skall betalas ut
- beträffande produktion av sockerrörssaft, för en mängd om 250 ton årligen,
- beträffande produktion av jordbruksrom, för en total mängd om 75600 hektoliter ren alkohol.
Artikel 18
Tillämpningsföreskrifter för detta kapitel samt stödbeloppet och det lägsta pris som avses i artikel 17.1 skall fastställas i enlighet med förfarandet i artikel 23.2.
KAPITEL V
GRAFISK SYMBOL
Artikel 19
1. Branschorganisationerna skall föreslå bestämmelser för användningen av en grafisk symbol i syfte att öka kunskapen om och konsumtionen av obearbetade och bearbetade jordbruksprodukter av hög kvalitet som är karakteristiska för de franska utomeuropeiska departementen i deras egenskap av yttersta randområden. De franska myndigheterna skall vidarebefordra sådana förslag, tillsammans med sitt yttrande, till kommissionen för godkännande.
Användningen av symbolen skall kontrolleras av en offentlig myndighet eller ett organ som godkänts av de behöriga franska myndigheterna.
2. Tillämpningsföreskrifter för denna artikel skall vid behov fastställas i enlighet med förfarandet i artikel 23.2.
AVDELNING III
FYTOSANITÄRA ÅTGÄRDER
Artikel 20
1. De franska myndigheterna skall för kommissionen lägga fram program för bekämpning av skadegörare på växter och växtprodukter. I programmen skall särskilt anges de mål som skall uppnås, åtgärder som skall vidtas samt deras varaktighet och kostnad. De program som läggs fram i enlighet med denna artikel skall inte beröra skyddsåtgärder för bananer.
2. Gemenskapen skall bidra till finansieringen av dessa program på grundval av en teknisk analys av situationen inom den berörda regionen.
3. Gemenskapens medfinansiering och stödbeloppet skall fastställas i enlighet med förfarandet i artikel 23.2. De åtgärder som gemenskapen kan lämna bidrag till skall fastställas i enlighet med samma förfarande.
4. Medfinansieringen kan uppgå till högst 60 % av de stödberättigande utgifterna. Utbetalning skall ske på grundval av handlingar som tillhandahålls av de franska myndigheterna. Kommissionen kan vid behov initiera undersökningar, som genomförs för dess räkning av sådana sakkunniga som avses i artikel 21 i direktiv 2000/29/EG(17).
TITEL IV
UNDANTAG FRÅN STRUKTURÅTGÄRDER
Artikel 21
1. Trots bestämmelserna i artikel 7 i förordning (EG) nr 1257/1999 skall stödets totala värde, uttryckt i procent av den stödberättigande investeringsvolymen, begränsas till högst 75 % för de investeringar som bl.a. syftar till att främja diversifiering, omstrukturering eller omställning till hållbart jordbruk på jordbruksföretag med begränsade tillgångar som skall definieras i det programkomplement som avses i artikel 19.4 i förordning (EG) nr 1260/1999.
2. Trots bestämmelserna i artikel 28.2 i förordning (EG) nr 1257/1999 skall stödets totala värde, uttryckt i procent av den stödberättigande investeringsvolymen, begränsas till högst 65 % för investeringar i företag för bearbetning och saluföring av jordbruksprodukter som huvudsakligen härrör från lokal produktion och från sektorer som skall definieras i det programkomplement som avses i artikel 19.4 i förordning (EG) nr 1260/1999. För små och medelstora företag skall stödets totala värde på samma villkor begränsas till högst 75 %.
3. Den begränsning som föreskrivs i artikel 29.3 i förordning (EG) nr 1257/1999 skall inte gälla tropiska skogar och skogsarealer i de franska utomeuropeiska departementen.
4. Trots bestämmelserna i artikel 47.2 andra stycket tredje strecksatsen i förordning (EG) nr 1257/1999 skall gemenskapens medfinansiering av åtgärder för miljövänligt jordbruk enligt artiklarna 22, 23 och 24 i den förordningen uppgå till 85 %.
5. En kortfattad beskrivning av de åtgärder som planeras i enlighet med den här artikeln skall ingå i de samlade programdokument för dessa departement som avses i artikel 19 i förordning (EG) nr 1260/1999.
AVDELNING V
ALLMÄNNA BESTÄMMELSER OCH SLUTBESTÄMMELSER
Artikel 22
De åtgärder som krävs för att genomföra denna förordning skall antas i enlighet med förvaltningsförfarandet i artikel 23.2.
Artikel 23
1. Kommissionen skall biträdas av Förvaltningskommittén för spannmål, som inrättats genom artikel 22 i förordning (EEG) nr 1766/92, eller av förvaltningskommittéer som inrättats genom förordningar om den gemensamma organisationen av marknaderna för de berörda produkterna.
För de jordbruksprodukter som omfattas av förordning (EEG) nr 827/68(18) samt för de produkter som inte omfattas av någon av de gemensamma organisationerna av marknaden skall kommissionen biträdas av Förvaltningskommittén för humle som inrättats genom artikel 20 i förordning (EEG) nr 1696/71(19).
När det gäller den grafiska symbolen och i andra fall som omfattas av denna förordning skall kommissionen biträdas av Förvaltningskommittén för färsk frukt och färska grönsaker som inrättats genom förordning (EG) nr 2200/96.
För genomförandet av avdelning III skall kommissionen biträdas av Ständiga kommittén för växtskydd som inrättats genom beslut 76/894/EEG(20).
För genomförandet av avdelning IV skall kommissionen biträdas av kommittén för utveckling och omställning av regioner och kommittén för jordbrukets struktur och landsbygdens utveckling, som inrättats genom artikel 48 respektive artikel 50 i förordning (EG) nr 1260/1999.
2. När det hänvisas till denna punkt skall artiklarna 4 och 7 i beslut 1999/468/EG tillämpas.
När det gäller avdelning III skall dock förfarandet i artikel 18 i direktiv 2000/29/EG tillämpas.
Den tid som avses i artikel 4.3 i beslut 1999/468/EG skall vara en månad.
3. Kommittéerna skall själva anta sina arbetsordningar.
Artikel 24
För de jordbruksprodukter som omfattas av bilaga I till fördraget får kommissionen för de produkter som omfattas av artiklarna 87-89 i fördraget tillåta stöd till sektorerna för produktion, bearbetning och saluföring av dessa produkter för att lindra de särskilda begränsningar för jordbruksproduktionen i de franska utomeuropeiska departementen som har samband med den avlägsna belägenheten, ökaraktären och läget i gemenskapens yttersta randområden.
Artikel 25
De åtgärder som fastställs i denna förordning, med undantag av artikel 21, skall utgöra interventioner avsedda att stabilisera jordbruksmarknaderna i enlighet med artikel 2.2 i förordning (EG) nr 1258/1999(21).
Artikel 26
Medlemsstaterna skall vidta nödvändiga åtgärder för att se till att bestämmelserna i denna förordning iakttas, särskilt när det gäller kontrollåtgärder och administrativa sanktioner och informera kommissionen om detta.
Tillämpningsföreskrifter för denna artikel skall fastställas i enlighet med förfarandet i artikel 23.2.
Artikel 27
1. Frankrike skall lägga fram en årsrapport för kommissionen om genomförandet av de åtgärder som föreskrivs i denna förordning.
2. Senast vid slutet av det femte tillämpningsåret skall kommissionen till Europaparlamentet och rådet överlämna en allmän rapport med en redogörelse för verkningarna av de åtgärder som vidtagits i enlighet med denna förordning, eventuellt tillsammans med lämpliga förslag.
Artikel 28
Förordning (EEG) nr 3763/91 upphör härmed att gälla. Hänvisningar till förordning (EEG) nr 3763/91 skall tolkas som hänvisningar till denna förordning enligt jämförelsetabellen i bilaga II.
Förordning (EEG) nr 525/77 upphör härmed att gälla från och med regleringsåret 2002/2003.
Kommissionen får, i enlighet med förfarandet i artikel 23.2, vidta nödvändiga övergångsåtgärder för en smidig övergång från den ordning som gäller under år 2000 eller under regleringsåret 2000-2001 till den ordning som införs genom den här förordningen. Om de befintliga åtgärderna förlängs skall kommissionen se till att den nödvändiga kontinuiteten bevaras.
Artikel 29
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Den skall tillämpas från och med den dag den träder i kraft. Emellertid skall
- artikel 10 tillämpas från och med den 1 januari 2001,
- artikel 11 tillämpas från och med den 1 januari 2001,
- artikel 16 tillämpas på sockerrör som skördas från och med regleringsåret 2001/2002,
- artikel 21 tillämpas från och med den 1 januari 2000.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Rådets förordning (EG) nr 2157/2001
av den 8 oktober 2001
om stadga för europabolag
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättande av Europeiska gemenskapen, särskilt artikel 308 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2),
med beaktande av Ekonomiska och sociala kommitténs yttrande(3), och
av följande skäl:
(1) Genomförandet av den inre marknaden och den förbättring av den ekonomiska och sociala situationen i hela gemenskapen detta bör leda till kräver, förutom slopande av handelshindren, en omstrukturering av produktionsfaktorerna så att de anpassas till gemenskapens dimension. För att så skall kunna ske, är det av största vikt att de företag vilkas verksamhet inte begränsar sig till att tillgodose rent lokala behov kan utforma och fullfölja omorganisationen av sin verksamhet på gemenskapsnivå.
(2) En sådan omorganisering förutsätter att redan existerande företag i flera medlemsstater får möjlighet att genom fusionsåtgärder samla sin potential. Sådana åtgärder får dock vidtas endast under förutsättning att fördragets konkurrensregler efterlevs.
(3) Vid genomförandet av omstrukturerings- och samarbetsåtgärder som inbegriper företag i olika medlemsstater uppstår svårigheter av juridisk, psykologisk och skatteteknisk art. Åtgärderna för tillnärmning av medlemsstaternas bolagsrätt genom direktiv grundade på artikel 44 är ägnade att undanröja vissa av dessa svårigheter. Dessa åtgärder befriar dock inte företag som omfattas av olika lagstiftningar från skyldigheten att välja en bolagsform som regleras av en viss nationell lagstiftning.
(4) Den rättsliga ram inom vilken företagen i gemenskapen måste hålla sig och som fortfarande är huvudsakligen nationell överensstämmer således inte med den ekonomiska ram inom vilken de bör utvecklas för att möjliggöra genomförandet av de mål som anges i artikel 18 i fördraget. Detta förhållande är ägnat att avsevärt försvåra sammanslagning av bolag hemmahörande i olika medlemsstater.
(5) Medlemsstaterna är skyldiga att sörja för att de bestämmelser som skall tillämpas på europabolagen enligt denna förordning varken leder till diskriminering genom oberättigad särbehandling av europabolag i förhållande till aktiebolag eller till oproportionerliga inskränkningar i rätten att bilda ett europabolag eller att flytta dess säte.
(6) Det är nödvändigt att i största möjliga mån få till stånd överensstämmelse mellan det europeiska företagets ekonomiska och dess rättsliga enheter. Därför bör föreskrifter antas som gör det möjligt att, vid sidan av bolag som faller under en viss nationell lag, stifta bolag vilkas bildande och verksamhet regleras av en gemenskapsförordning som är direkt tillämplig i alla medlemsstater.
(7) Bestämmelserna i en sådan förordning kommer att göra det möjligt att bilda och driva bolag med en europeisk dimension, utan att olikheterna i och den begränsade territoriella tillämpningen av de nationella lagstiftningar som gäller för affärsdrivande bolag hindrar eller försvårar detta.
(8) Stadgan för europabolag (nedan kallade %quot%SE-bolag%quot%) tillhör de rättsakter som skulle antas av rådet före 1992 enligt kommissionens vitbok om den inre marknaden, vilken godkändes i juni 1985 av Europeiska rådet i Milano. Vid sitt möte i Bryssel 1987 uttryckte Europeiska rådet önskemålet att en sådan stadga snabbt skulle upprättas.
(9) Sedan kommissionen 1970 lade fram förslaget till förordning om stadga för europeiska aktiebolag, vilket ändrades 1975, har arbetet på en tillnärmning av den nationella bolagsrätten avancerat betydligt, varför det är möjligt att i stadgan för SE-bolag hänvisa till lagstiftningen om aktiebolag i den medlemsstat där SE-bolaget har sitt säte på de områden där dess verksamhet inte kräver enhetliga gemenskapsbestämmelser.
(10) Det huvudsakliga mål som eftersträvas i den rättsliga ordningen för SE-bolag kräver under alla omständigheter, utan att de ekonomiska behov som kan uppstå i framtiden åsidosätts, att ett SE-bolag kan bildas både för att tillåta bolag hemmahörande i olika medlemsstater att gå samman eller bilda ett holdingbolag och för att ge möjlighet åt bolag och andra juridiska personer med ekonomisk verksamhet hemmahörande i olika medlemsstater att bilda gemensamma dotterbolag.
(11) I samma syfte bör ett aktiebolag tillåtas att ombildas till SE-bolag med säte och huvudkontor i gemenskapen utan att bolaget först måste upplösas, om bolaget har ett dotterbolag i en annan medlemsstat än den där bolaget har sitt säte.
(12) De nationella bestämmelser som gäller för publika aktiebolag och för aktieaffärer bör även tillämpas när SE-bolag bildas i form av ett publikt bolag, liksom på SE-bolag som senare önskar bli publika.
(13) SE-bolaget självt bör bildas i form av ett aktiebolag, som är den rättsliga form som, både från finansierings- och förvaltningssynpunkt, bäst svarar mot behoven hos företag som bedriver verksamhet på europeisk nivå. För att säkerställa att sådana företag får ett lämpligt format bör det fastställas en lägsta gräns för aktiekapitalet så att bolagen förfogar över tillräckliga tillgångar, utan att det för den skull försvåras för små och medelstora företag (SMF) att bilda SE-bolag.
(14) Det är viktigt att möjliggöra att ett SE-bolag drivs effektivt samtidigt som en noggrann tillsyn över förvaltningen säkerställs. Hänsyn bör tas till att det för närvarande, vad beträffar administration av aktiebolag, förekommer två olika system inom gemenskapen. Samtidigt som SE-bolag bör tillåtas att välja mellan dessa båda system, bör dock en klar ansvarsfördelning göras mellan de personer som sköter bolagets förvaltning och dem som utövar tillsynen.
(15) Rättigheter och skyldigheter i fråga om skydd för minoritetsaktieägare och tredje man när ett företag utövar kontroll över ett annat företag som omfattas av en annan lagstiftning skall, enligt den internationella privaträttens allmänna regler och principer, regleras av den lag av vilken det kontrollerade företaget omfattas, utan att detta påverkar de skyldigheter som åvilar det kontrollerande företaget i kraft av de lagbestämmelser detta omfattas av, till exempel i fråga om koncernredovisning.
(16) Utan att det påverkar konsekvenserna av en framtida samordning av medlemsstaternas lagstiftningar, krävs för närvarande ingen särskild reglering avseende SE-bolag på detta område. Därför bör dessa allmänna regler och principer tillämpas både då SE-bolaget är det kontrollerande bolaget och då SE-bolaget är det kontrollerade bolaget.
(17) De regler som faktiskt är tillämpliga då SE-bolaget kontrolleras av ett annat företag bör preciseras, och det bör därvid hänvisas till den lag som är tillämplig på aktiebolag som omfattas av lagstiftningen i den medlemsstat där SE-bolaget har sitt säte.
(18) Varje medlemsstat måste vara förpliktad att vid överträdelser av bestämmelserna i denna förordning tillämpa de sanktioner som gäller för aktiebolag som omfattas av dess lagstiftning.
(19) Reglerna för arbetstagarinflytande i SE-bolag är föremål för rådets direktiv 2001/86/EG av den 8 oktober 2001 om komplettering stadgan för europabolag vad gäller arbetstagarinflytande(4). Dessa bestämmelser utgör ett oskiljbart komplement till denna förordning och måste tillämpas tillsammans med denna.
(20) Denna förordning omfattar inga andra rättsliga områden, såsom skatterätt, insolvensrätt, immaterial- eller konkursrätt. Följaktligen skall bestämmelserna i medlemsstaternas lagstiftning och i gemenskapsrätten tillämpas på de ovannämnda områdena samt på andra områden som inte omfattas av denna förordning.
(21) Direktiv 2001/86/EG syftar till att tillförsäkra arbetstagarna rätt till inflytande beträffande frågor och beslut som påverkar verksamheten och förhållandena i SE-bolagen. Övriga frågor av social- och arbetsrättslig art, särskilt arbetstagarnas rätt till information och samråd, såsom den är utformad i medlemsstaterna, regleras av de nationella bestämmelser som under samma omständigheter gäller för aktiebolag.
(22) Denna förordnings ikraftträdande måste uppskjutas så att varje medlemsstat i sin nationella lagstiftning kan införliva bestämmelserna i direktiv 2001/86/EG och i förväg inrätta den struktur som behövs för att bilda och driva SE-bolag med säten inom den statens territorium, så att förordningen och direktivet kan tillämpas samtidigt.
(23) Ett bolag som inte har sitt huvudkontor i gemenskapen bör få delta i bildandet av ett SE-bolag, om bolaget bildas i överensstämmelse med lagstiftningen i en medlemsstat, har sitt säte i den medlemsstaten och har faktisk och fortlöpande anknytning till ekonomin i den medlemsstaten enligt de principer som fastställs i 1962 års allmänna program för upphävande av begränsningar i etableringsfriheten. Sådan anknytning föreligger särskilt om bolaget har ett driftsställe i medlemsstaten och driver verksamhet därifrån.
(24) Ett SE-bolag bör ha möjlighet att flytta sitt säte till en annan medlemsstat. Ett adekvat skydd av intressena för de minoritetsaktieägare som motsätter sig flyttningen samt av borgenärers och andra rättsinnehavares intressen bör vara proportionerligt. Flyttningen bör inte påverka de rättigheter som har tillkommit före flyttningen.
(25) Denna förordning påverkar inte tillämpningen av någon bestämmelse som kan komma att införas i 1968 års Brysselkonvention eller i någon text som antas av medlemsstaterna eller rådet för att ersätta den konventionen och som avser de behörighetsregler som gäller när ett publikt aktiebolag flyttar sitt säte från en medlemsstat till en annan.
(26) Finansinstitutens verksamhet regleras av särskilda direktiv, och de nationella bestämmelserna för genomförande av dessa direktiv och andra nationella regler för denna verksamhet gäller fullt ut för SE-bolag.
(27) Med hänsyn till SE-bolagens särskilda gemenskapskaraktär påverkar den ordning för ett SE-bolags faktiska säte som antas genom denna förordning inte tillämpningen av medlemsstaternas lagstiftningar och åsidosätter inte de val som kan göras när det gäller andra gemenskapstexter om bolagsrätt.
(28) I fördraget anges inte några andra befogenheter för att anta denna förordning än de som finns i artikel 308.
(29) Eftersom målen för de föreslagna åtgärderna såsom de skisseras ovan inte i tillräcklig utsträckning kan uppnås av medlemsstaterna, eftersom det är fråga om att bilda SE-bolag på europeisk nivå och de därför på grund av åtgärdernas omfattning och effekter bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidaritetsprincipen i artikel 5 i fördraget. I enlighet med proportionalitetsprincipen i samma artikel går detta beslut inte utöver vad som är nödvändigt för att uppnå dessa mål.
HÄRIGENOM FÖRESKRIVS FÖLJANDE
AVDELNING I
ALLMÄNNA BESTÄMMELSER
Artikel 1
1. Ett bolag får bildas inom gemenskapens territorium i form av ett europeiskt publikt aktiebolag (Societas Europaea, nedan kallat %quot%SE-bolag%quot%) på de villkor och enligt de bestämmelser som fastställs i denna förordning.
2. Ett SE-bolag skall vara ett bolag vars aktiekapital är fördelat på aktier. Varje aktieägare skall vara ekonomiskt ansvarig endast för den del av aktiekapitalet som han har tecknat.
3. Ett SE-bolag skall vara en juridisk person.
4. Arbetstagarinflytandet i ett SE-bolag skall följa bestämmelserna i direktiv 2001/86/EG.
Artikel 2
1. Publika aktiebolag som anges i bilaga I som har bildats i överensstämmelse med lagstiftningen i en medlemsstat och som har sitt säte och sitt huvudkontor i gemenskapen, får bilda ett SE-bolag genom fusion, om minst två av bolagen omfattas av olika medlemsstaters lagstiftning.
2. Publika och privata aktiebolag i bilaga II vilka har bildats i överensstämmelse med lagstiftningen i en medlemsstat samt har sitt säte och sitt huvudkontor i gemenskapen får ta initiativ till bildandet av ett SE-holdingbolag, om minst två av bolagen
a) omfattas av olika medlemsstaters lagstiftning eller
b) sedan minst två år har ett dotterbolag som omfattas av lagstiftningen i en annan medlemsstat eller en filial belägen i en annan medlemsstat.
3. Bolag enligt artikel 48 andra stycket i fördraget samt andra offentligrättsliga eller privaträttsliga rättsliga enheter, som har bildats i överensstämmelse med lagstiftningen i en medlemsstat och har sitt säte och sitt huvudkontor i gemenskapen, får bilda ett SE-dotterbolag genom att teckna aktier i detta, om minst två av dem
a) omfattas av olika medlemsstaters lagstiftning eller
b) sedan minst två år har ett dotterbolag som omfattas av lagstiftningen i en annan medlemsstat eller en filial belägen i en annan medlemsstat.
4. Ett publikt aktiebolag som har bildats enligt lagstiftningen i en medlemsstat och som har sitt säte och huvudkontor i gemenskapen får ombildas till ett SE-bolag om det sedan minst två år har ett dotterbolag som omfattas av lagstiftningen i en annan medlemsstat.
5. En medlemsstat har rätt att föreskriva att ett bolag som inte har sitt huvudkontor i gemenskapen får delta i bildandet av ett SE-bolag, om bolaget är bildat i överensstämmelse med lagstiftningen i en medlemsstat, har sitt säte i den medlemsstaten och har faktisk och fortlöpande anknytning till ekonomin i en medlemsstat.
Artikel 3
1. Vid tillämpningen av artikel 2.1, 2.2. och 2.3 skall ett SE-bolag anses som ett publikt aktiebolag som omfattas av lagstiftningen i den medlemsstat där det har sitt säte.
2. Ett SE-bolag får självt bilda ett eller flera dotterbolag i form av SE-bolag. Sådana bestämmelser i den medlemsstat där ett SE-dotterbolag har sitt säte enligt vilka krävs att ett publikt aktiebolag skall ha fler än en aktieägare skall inte tillämpas på SE-dotterbolaget. De nationella bestämmelser som har antagits i enlighet med rådets tolfte direktiv 89/667/EEG av den 21 december 1989 på bolagsrättens område om enmansbolag med begränsat ansvar(5) skall i tillämpliga delar gälla för SE.
Artikel 4
1. Ett SE-bolags aktiekapital skall vara uttryckt i euro.
2. Det tecknade aktiekapitalet skall uppgå till minst 120000 euro.
3. Om det i lagstiftningen i en medlemsstat föreskrivs ett större tecknat aktiekapital för bolag med vissa typer av verksamhet, skall den lagstiftningen tillämpas på SE-bolag som har sitt säte i den medlemsstaten.
Artikel 5
Om inte annat följer av bestämmelserna i artikel 4.1 och 4.2, skall ett SE-bolags aktiekapital, aktiekapitalets bibehållande, ändringar av det samt SE-bolagets aktier, obligationer och andra jämförbara värdepapper regleras av de bestämmelser som skulle tillämpas på ett publikt aktiebolag med säte i den medlemsstat där SE-bolaget är registrerat.
Artikel 6
I denna förordning avses med ett SE-bolags bolagsordning både SE-bolagets stiftelseurkund och dess bolagsordning, om denna utgör ett separat dokument.
Artikel 7
Ett SE-bolags säte skall vara beläget inom gemenskapen i samma medlemsstat som huvudkontoret. En medlemsstat får dessutom föreskriva att SE-bolag som är registrerade inom dess territorium skall vara skyldiga att förlägga sitt huvudkontor och säte till samma plats.
Artikel 8
1. Ett SE-bolags säte får flyttas till en annan medlemsstat i enlighet med punkterna 2-13. En sådan flyttning skall inte medföra vare sig bolagets avveckling eller bildandet av en ny juridisk person.
2. Ett förslag om flyttning skall upprättas av lednings- eller förvaltningsorganet och offentliggöras i enlighet med artikel 13, utan att detta påverkar eventuella ytterligare former av offentliggörande som föreskrivs i den medlemsstat där bolaget har sitt säte. I förslaget skall SE-bolagets aktuella firma, säte och nummer anges, samt
a) det säte som föreslås för SE-bolaget,
b) den bolagsordning som föreslås för SE-bolaget och, i förekommande fall, bolagets nya firma,
c) eventuella följder som flyttningen kan få för arbetstagarinflytandet,
d) den tidsplan som föreslås för flyttningen,
e) eventuella rättigheter till skydd av aktieägare och/eller borgenärer.
3. Lednings- eller förvaltningsorganet skall avfatta en redogörelse där flyttningens juridiska och ekonomiska aspekter förklaras och motiveras och där det förklaras vilka följder flyttningen får för aktieägare, borgenärer och arbetstagare.
4. Senast en månad före den bolagsstämma vid vilken det skall beslutas om flyttningen skall ett SE-bolags aktieägare och borgenärer ha rätt att där bolaget har sitt säte granska förslaget om flyttning och den redogörelse som avfattats i enlighet med punkt 3 samt att på begäran kostnadsfritt få kopior av dessa dokument.
5. En medlemsstat får när det gäller SE-bolag som är registrerade inom dess territorium anta bestämmelser som är avsedda att säkerställa ett lämpligt skydd för de minoritetsaktieägare som motsätter sig flyttning.
6. Ett beslut om flyttning får inte fattas förrän två månader efter offentliggörandet av förslaget. Beslutet skall fattas enligt bestämmelserna i artikel 59.
7. Innan den behöriga myndigheten utfärdar det intyg som avses i punkt 8, skall SE-bolaget visa denna att, när det gäller sådana skulder som uppkommit före offentliggörandet av förslaget om flyttning, de intressen som borgenärer och innehavare av övriga rättigheter har gentemot SE-bolaget (inbegripet offentliga organs intressen) är skyddade på ett betryggande sätt i överensstämmelse med de krav som har fastställts av den medlemsstat där SE-bolaget har sitt säte före flyttningen.
En medlemsstat får utvidga tillämpningen av det första stycket till att omfatta skulder som uppkommer (eller kan uppkomma) före flyttningen.
Föregående stycken skall inte påverka tillämpningen på SE-bolag av medlemsstaternas nationella lagstiftning om erläggande eller säkring av betalningar till offentliga organ.
8. En domstol, notarie eller annan behörig myndighet i den medlemsstat där ett SE-bolag har sitt säte skall utfärda ett intyg som slutgiltigt bekräftar att vad som krävs i fråga om handlingar och formaliteter före flyttningen har fullgjorts.
9. Ny registrering får inte ske förrän det intyg som avses i punkt 5 har framlagts och det har styrkts att de formaliteter som krävs för registrering i det land där bolagets nya säte skall vara beläget har uppfyllts.
10. Flyttningen av ett SE-bolags säte samt den därav följande ändringen av bolagets bolagsordning skall bli gällande den dag då SE-bolaget i enlighet med artikel 12 registreras i registret där bolaget har sitt nya säte.
11. När SE-bolagets nya registrering har gjorts, skall en underrättelse om detta lämnas från det register där den nya registreringen gjorts till det register där den gamla registreringen fanns. Den gamla registreringen skall strykas vid mottagandet av denna underrättelse, men inte före detta.
12. Den nya registreringen och strykningen av den gamla skall offentliggöras i de berörda medlemsstaterna i enlighet med artikel 13.
13. I och med offentliggörandet av SE-bolagets nya registrering kan det nya sätet åberopas gentemot tredje man. Så länge strykningen ur registret av SE-bolagets registrering på dess föregående säte inte har offentliggjorts kan emellertid tredje man fortsätta att åberopa det föregående sätet, såvida inte SE-bolaget bevisar att tredje man hade kännedom om det nya sätet.
14. Genom lagstiftningen i en medlemsstat får det, i fråga om SE-bolag som är registrerade i den medlemsstaten, föreskrivas att en flyttning av bolagets säte som skulle medföra en ändring av tillämplig lag inte skall bli gällande om någon behörig myndighet i medlemsstaten motsätter sig flyttningen inom den tvåmånadersfrist som avses i punkt 6. Motsättandet får grundas endast på hänsyn till allmänintresset.
Om ett SE-bolag kontrolleras av en nationell finansiell tillsynsmyndighet enligt gemenskapens direktiv skall rätten att motsätta sig ändring av säte också gälla denna myndighet.
Överklagande till domstol skall vara möjligt.
15. Ett SE-bolag som har varit föremål för ett rättsligt förfarande rörande avveckling, likvidation, insolvens eller betalningsinställelse eller andra liknande förfaranden får inte flytta sitt säte.
16. Ett SE-bolag som har flyttat sitt säte till en annan medlemsstat skall, när det gäller rättsanspråk som kan uppkomma före den flyttning som avses i punkt 10 i denna artikel, anses ha sitt säte i den medlemsstat där SE-bolaget var registrerat före flyttningen, även om talan skulle väckas mot SE-bolaget efter flyttningen.
Artikel 9
1. Ett SE-bolag skall regleras
a) av bestämmelserna i denna förordning,
b) om denna förordning uttryckligen tillåter det, av bestämmelserna i bolagets bolagsordning,
eller
c) beträffande frågor som inte regleras i denna förordning eller - om en fråga endast delvis regleras i den - beträffande de aspekter som inte omfattas av denna förordning, av
i) de lagbestämmelser som har antagits av medlemsstaterna för att tillämpa gemenskapsåtgärder som specifikt avser SE bolag,
ii) de lagbestämmelser i medlemsstaterna som skulle gälla för ett publikt aktiebolag bildat i överensstämmelse med lagstiftningen i den medlemsstat där SE-bolaget har sitt säte,
iii) bestämmelserna i bolagsordningen på samma villkor som för ett publikt aktiebolag bildat i överensstämmelse med lagstiftningen i den medlemsstat där SE-bolaget har sitt säte.
2. De lagbestämmelser som antas av medlemsstaterna specifikt för SE-bolag måste stämma överens med de direktiv som är tillämpliga på de publika aktiebolag som anges i bilaga I.
3. Om det finns särskilda bestämmelser i nationell lagstiftning för den typ av verksamhet som ett SE-bolag bedriver skall dessa bestämmelser gälla fullt ut för SE-bolaget.
Artikel 10
Om inte annat följer av bestämmelserna i denna förordning, skall ett SE-bolag i varje medlemsstat behandlas som ett publikt aktiebolag bildat i överensstämmelse med lagstiftningen i den medlemsstat där SE-bolaget har sitt säte.
Artikel 11
1. SE-bolagets firma skall innehålla förkortningen %quot%SE%quot% före eller efter firman.
2. Endast SE-bolag får ha firmor som innehåller förkortningen %quot%SE%quot%.
3. Bolag eller andra juridiska personer som har registrerats i en medlemsstat före den dag då denna förordning träder i kraft och vilkas firmor innehåller förkortningen %quot%SE%quot% skall dock inte vara skyldiga att ändra sina firmor.
Artikel 12
1. Varje SE-bolag skall registeras i den medlemsstat där det har sitt säte i ett register som anges i lagstiftningen i denna medlemsstat i enlighet med artikel 3 i rådets direktiv 68/151/EEG av den 9 mars 1968 om samordning av de skyddsåtgärder som krävs i medlemsstaterna av de i artikel 58 andra stycket i fördraget avsedda bolagen i bolagsmännens och tredje mans intressen, i syfte att göra skyddsåtgärderna likvärdiga inom gemenskapen(6).
2. Ett SE-bolag får inte registeras om det saknas en överenskommelse om riktlinjer för arbetstagarinflytande enligt artikel 4 i direktiv 2001/86/EG eller ett beslut enligt artikel 3.6 i det direktivet eller om förhandlingsperioden enligt artikel 5 i det direktivet har löpt ut utan att en överenskommelse har träffats.
3. För att ett SE-bolag skall kunna registreras i en medlemsstat som har utnyttjat möjligheten i artikel 7.3 i direktiv 2001/86/EG, är det nödvändigt att ett avtal har slutits i enlighet med artikel 4 i det direktivet om en ordning för hur arbetstagarinflytande och -medverkan skall utformas, eller att inget av de bolag som ingår lyder under bestämmelser om medverkan före registreringen av SE-bolaget.
4. Ett SE-bolags bolagsordning får aldrig strida mot de riktlinjer för arbetstagarinflytande som har fastställts på detta sätt. Om nya riktlinjer som fastställts i enlighet med direktiv 2001/86/EG strider mot gällande bolagsordning, skall bolagsordningen ändras i nödvändig omfattning.
I detta fall skall SE-bolagets lednings- eller förvaltningsorgan ha rätt att vidta åtgärder för att ändra bolagsordningen utan något ytterligare beslut från bolagsstämman.
Artikel 13
De handlingar och uppgifter rörande ett SE-bolag som skall offentliggöras enligt denna förordning skall offentliggöras på det sätt som föreskrivs i lagstiftningen i den medlemsstat där SE-bolaget har sitt säte i enlighet med direktiv 68/151/EEG.
Artikel 14
1. Ett meddelande om registrering och avregistrering av ett SE-bolag skall offentliggöras för kännedom i Europeiska gemenskapernas officiella tidning när offentliggörande har skett i enlighet med artikel 13. Meddelandet skall innehålla uppgift om SE-bolagets namn, registreringsnummer, registreringsdatum och registreringsort, datum och ort för offentliggörandet, samt om bolagets säte och dess verksamhetsområde.
2. Vid flyttning av SE-bolagets säte enligt artikel 8 skall ett meddelande därom offentliggöras innehållande de uppgifter som avses i punkt 1 samt uppgifter om den nya registreringen.
3. De uppgifter som avses i punkt 1 skall översändas till Byrån för Europeiska gemenskapernas officiella publikationer inom en månad efter det offentliggörande som avses i artikel 13.
AVDELNING II
BILDANDE
Avsnitt 1
Allmänna bestämmelser
Artikel 15
1. Om inte annat följer av denna förordning, skall bildandet av ett SE-bolag regleras av den lag som gäller för publika aktiebolag i den stat dit SE-bolaget förlägger sitt säte.
2. Registrering av ett SE-bolag skall offentliggöras enligt artikel 13.
Artikel 16
1. Ett SE-bolag får status som juridisk person den dag då det registreras i det register som avses i artikel 12.
2. Om rättshandlingar har företagits i SE-bolagets namn före dess registrering enligt artikel 12 och om SE-bolaget efter registreringen inte påtar sig de skyldigheter som härrör från dessa rättshandlingar, skall de fysiska personer, bolag eller andra juridiska personer som företagit handlingarna vara solidariskt och obegränsat ansvariga för dessa, såvida inte annat överenskommits.
Avsnitt 2
Bildande av ett SE-bolag genom fusion
Artikel 17
1. Ett SE-bolag får bildas genom fusion i enlighet med artikel 2.1.
2. Fusionen kan genomföras
a) enligt förfarandet för fusion genom förvärv i artikel 3.1 i direktiv 78/855/EEG(7), eller
b) enligt förfarandet för fusion genom bildande av ett nytt bolag i artikel 4.1 i samma direktiv.
I fallet med fusion genom förvärv skall det övertagande bolaget anta bolagsformen SE-bolag samtidigt med fusionen. I fallet med fusion genom bildande av ett nytt bolag skall SE-bolaget vara det nybildade bolaget.
Artikel 18
Beträffande frågor som inte innefattas i detta avsnitt, eller - om en fråga endast delvis innefattas av detta - beträffande de aspekter som inte innefattas i avsnittet skall varje bolag som deltar i bildandet av ett SE-bolag genom fusion vara underställt de lagbestämmelser i den medlemsstat där det hör hemma som gäller för fusion av publika aktiebolag i enlighet med direktiv 78/855/EEG.
Artikel 19
Genom lagstiftningen i en medlemsstat får det föreskrivas att ett bolag som omfattas av lagstiftningen i den medlemsstaten inte får delta i bildandet av ett SE-bolag genom fusion, om en behörig myndighet i denna medlemsstat motsätter sig detta före utfärdandet av det intyg som avses i artikel 25.2.
Ett sådant motsättande får grundas endast på hänsyn till allmänintresset. Överklagande till domstol skall vara möjligt.
Artikel 20
1. Lednings- eller förvaltningsorganen i de fusionerande bolagen skall utarbeta ett fusionsförslag. Förslaget skall innehålla
a) uppgift om de fusionerande bolagens firma och säte samt om SE-bolagets planerade firma och säte,
b) uppgift om aktiernas utbytesförhållande och om eventuellt kompensationsbelopp,
c) uppgift om villkoren för tilldelning av aktier i SE-bolaget,
d) uppgift om från och med vilket datum innehav av aktier i SE-bolaget ger rätt till del i vinsten samt om eventuella särskilda villkor rörande denna rätt,
e) uppgift om från och med vilket datum de fusionerande bolagens transaktioner bokföringsmässigt skall behandlas som hörande till SE-bolaget,
f) uppgift om vilka rättigheter SE-bolaget tilldelar innehavare av aktier med speciella rättigheter och innehavare av andra värdepapper än aktier eller om vilka åtgärder som föreslås beträffande dem,
g) uppgift om eventuella särskilda förmåner som beviljas de experter som granskar fusionsförslaget samt ledamöterna av förvaltnings-, lednings-, tillsyns- eller kontrollorganen i de fusionerande bolagen,
h) SE-bolagets bolagsordning,
i) information om de förfaranden genom vilka riktlinjerna för arbetstagarinflytandet skall fastställas i enlighet med direktiv 2001/86/EG.
2. De fusionerande bolagen får ta med ytterligare uppgifter i fusionsförslaget.
Artikel 21
För vart och ett av de fusionerande bolagen skall, med förbehåll för eventuella ytterligare krav som åläggs av den medlemsstat under vars lagstiftning det aktuella bolaget faller, följande uppgifter offentliggöras i denna medlemsstats allmänna tidning:
a) Form, firma och säte för varje fusionerande bolag.
b) Det register till vilket de handlingar som avses i artikel 3.2 i direktiv 68/151/EEG har ingivits för vart och ett av de fusionerande bolagen samt registreringsnummer i detta register.
c) En uppgift om hur det aktuella bolagets borgenärer skall förfara för att utöva sina rättigheter enligt artikel 24 samt den adress där fullständig information om detta förfarande kostnadsfritt kan erhållas.
d) En uppgift om hur minoritetsaktieägarna i det berörda bolaget skall förfara för att utöva sina rättigheter enligt artikel 24 samt den adress där fullständig information om detta förfarande kostnadsfritt kan erhållas.
e) SE-bolagets planerade firma och säte.
Artikel 22
Som alternativ till experter som granskar förslaget för varje fusionerande bolags räkning får en eller flera oberoende experter, enligt artikel 10 i direktiv 78/855/EEG, utsedda för detta ändamål och på gemensam begäran av de fusionerande bolagen av en rättslig eller administrativ myndighet i den medlemsstat av vars lagstiftning något av de fusionerande bolagen eller det blivande SE-bolaget omfattas, granska fusionsförslaget och upprätta ett gemensamt yttrande avsett för samtliga aktieägare.
Experterna skall ha rätt att av vart och ett av de fusionerande bolagen begära de upplysningar som de anser vara nödvändiga för att de skall kunna slutföra sin uppgift.
Artikel 23
1. Bolagsstämman i vart och ett av de fusionerande bolagen skall godkänna fusionsförslaget.
2. Arbetstagarinflytandet i SE-bolaget skall fastställas i enlighet med direktiv 2001/86/EG och denna förordning. Bolagsstämman i vart och ett av de fusionerande bolagen får förbehålla sig rätten att ställa som villkor för registrering av SE-bolaget att den uttryckligen bekräftar de riktlinjer som har beslutats på detta sätt.
Artikel 24
1. Lagstiftningen i den medlemsstat under vars lagstiftning vart och ett av de fusionerande bolagen lyder skall, under beaktande av att fusionen är gränsöverskridande, tillämpas på samma sätt som vid fusion mellan publika aktiebolag vad beträffar skyddet av följande personers intressen:
a) De fusionerande bolagens borgenärer.
b) De fusionerande bolagens rättighetsinnehavare.
c) Innehavare av andra värdepapper än aktier, vilka är förenade med speciella rättigheter i de fusionerande bolagen.
2. En medlemsstat får, vad beträffar fusionerande bolag som faller under dess lagstiftning, anta bestämmelser avsedda att säkerställa lämpligt skydd för de minoritetsaktieägare som motsatt sig fusionen.
Artikel 25
1. Kontrollen av fusionens lagenlighet skall, beträffande den del av förfarandet som rör varje fusionerande bolag, ske i enlighet med den lag som tillämpas på fusion mellan publika aktiebolag i den medlemsstat under vars lagstiftning bolaget lyder.
2. I varje berörd medlemsstat skall domstol, notarie eller annan behörig myndighet utfärda ett intyg genom vilket slutgiltigt bekräftas att alla rättshandlingar och formaliteter inför fusionen har fullgjorts.
3. Om det i lagstiftningen i en medlemsstat under vars lagstiftning fusionerande bolaget lyder föreskrivs ett förfarande för kontroll och ändring av aktiernas utbytesförhållande eller för kompensation av minoritetsaktieägare utan att det hindrar fusionens registrering, skall dessa förfaranden gälla endast om övriga fusionerande bolag belägna i medlemsstater som inte ger utrymme för ett sådant förfarande vid godkännandet av fusionsförslaget i enlighet med artikel 23.1 uttryckligen godtar möjligheten för det fusionerande bolagets aktieägare att tillgripa detta förfarande. I sådana fall kan domstolen, notarien eller annan behörig myndighet utfärda intyg enligt punkt 2 även om ett sådant förfarande har inletts. I intyget skall dock anges att förfarandet är oavslutat. Beslutet som förfarandet leder fram till är bindande för det övertagande bolaget och dess aktieägare.
Artikel 26
1. Kontrollen av fusionens lagenlighet skall, beträffande den del av förfarandet som rör genomförandet av fusionen och bildandet av ett SE-bolag, utföras av domstol, notarie eller annan myndighet som i den medlemsstat där SE-bolaget kommer att ha sitt säte är behörig att kontrollera denna aspekt av lagenligheten vid fusion mellan publika aktiebolag.
2. Varje fusionerande bolag skall därför överlämna det intyg som avses i artikel 25.2 till denna myndighet inom sex månader från och med intygets utfärdande samt en kopia av det av bolaget godkända fusionsförslaget.
3. Den myndighet som avses i punkt 1 skall särskilt kontrollera att de fusionerande bolagen har godkänt ett fusionsförslag med samma lydelse och att riktlinjer för arbetstagarinflytande har fastställts i enlighet med direktivet.
4. Myndigheten skall vidare kontrollera att SE-bolaget har bildats i överensstämmelse med de villkor som fastställs i lagen i den medlemsstat där det enligt artikel 15 har sitt säte.
Artikel 27
1. Fusionen och det samtidiga bildandet av ett SE-bolag skall träda i kraft vid det datum då SE-bolaget registreras i enlighet med artikel 12.
2. Ett SE-bolag får inte registreras förrän alla de formaliteter som avses i artiklarna 25 och 26 har fullgjorts.
Artikel 28
Varje fusionerande bolag skall offentliggöra genomförandet av fusionen enligt bestämmelserna i varje medlemsstats lag i enlighet med artikel 3 i direktiv 68/151/EEG.
Artikel 29
1. Då fusionen genomförs enligt artikel 17.2 a skall följande rättsverkningar inträda samtidigt:
a) Varje överlåtande bolags samtliga tillgångar och skulder överförs till det övertagande bolaget.
b) Aktieägarna i det överlåtande bolaget blir aktieägare i det övertagande bolaget.
c) Det överlåtande bolaget upphör att existera.
d) Det övertagande bolaget antar den juridiska formen SE-bolag.
2. Då fusionen genomförs enligt artikel 17.2 b skall följande rättsverkningar inträda samtidigt:
a) De fusionerande bolagens samtliga tillgångar och skulder överförs till SE-bolaget.
b) Aktieägarna i de fusionerande bolagen blir aktieägare i SE-bolaget.
c) De fusionerande bolagen upphör att existera.
3. Om lagen i en medlemsstat vid fusion mellan publika aktiebolag kräver att särskilda formaliteter uppfylls för att de fusionerande bolagens överföring av vissa tillgångar, rättigheter och skyldigheter skall få rättsverkan gentemot tredje man, skall dessa formaliteter tillämpas och fullgöras antingen av de fusionerande bolagen eller av SE-bolaget efter dess registrering.
4. De deltagande bolagens rättigheter och skyldigheter i fråga om sådana anställningsvillkor som härrör från nationell lagstiftning, praxis och enskilda anställningskontrakt eller anställningsförhållanden och som föreligger vid tidpunkten för registreringen, skall med anledning av registreringen överföras till SE-bolaget när det registreras.
Artikel 30
När SE-bolaget har registrerats, kan en fusion som skett enligt bestämmelserna i artikel 2.1 inte ogiltigförklaras.
Utebliven kontroll av fusionens lagenlighet enligt artiklarna 25 och 26 kan utgöra en av grunderna för att avveckla ett SE-bolag.
Artikel 31
1. När en fusion enligt artikel 17.2 a genomförs av ett bolag som innehar samtliga aktier och övriga värdepapper som berättigar till rösträtt vid ett överlåtande bolags bolagsstämma, skall bestämmelserna i artiklarna 20.1 b, 20.1 c, 20.1 d, 22 och 29.1 b inte tillämpas. Dock skall de nationella bestämmelser under vilka vart och ett av de fusionerande bolagen lyder och som reglerar fusioner mellan publika aktiebolag i enlighet med artikel 24 i direktiv 78/855/EEG tillämpas.
2. När en fusion genom förvärv av ett annat bolags tillgångar och skulder genomförs av ett bolag som inte innehar samtliga men 90 % eller mer av de aktier och övriga värdepapper som berättigar till rösträtt i ett överlåtande bolags bolagsstämma, skall redogörelser från lednings- eller förvaltningsorganet, yttranden från en eller flera oberoende experter samt de handlingar som behövs för kontrollen endast erfordras i den mån detta föreskrivs i den nationella lag under vilken det övertagande bolaget faller eller av den nationella lag under vilken det överlåtande bolaget faller.
Medlemsstaterna får emellertid föreskriva att denna punkt kan gälla när ett bolag innehar aktier som berättigar till 90 % eller mer av rösterna, men inte till samtliga röster.
Avsnitt 3
Bildande av ett SE-holdingbolag
Artikel 32
1. Ett SE-bolag får bildas i enlighet med artikel 2.2.
Ett bolag som tar initiativet till bildande av ett SE-bolag i enlighet med artikel 2.2 upphör inte att existera.
2. Lednings- eller förvaltningsorganen i de bolag som tar initiativet till bildandet skall utarbeta ett likalydande förslag till bildande av ett SE-bolag. Förslaget skall innehålla en redogörelse där bolagsbildningens juridiska och ekonomiska aspekter förklaras och motiveras och där det anges vilka följder antagandet av bolagsformen SE-bolag får för aktieägare och för arbetstagare. Förslaget skall vidare innehålla de uppgifter som anges i artikel 20.1 a, b, c, f, g, h och i och fastställa den lägsta procentuella andel aktier i vart och ett av de bolag som tar initiativet till bildandet som måste tillskjutas av aktieägarna för att ett SE-bolag skall bildas. Denna andel skall bestå av aktier som berättigar till över 50 % av de ordinarie rösterna.
3. För vart och ett av de initiativtagande bolagen skall förslaget till bildande av SE-bolaget offentliggöras på det sätt som föreskrivs i varje medlemsstats lagstiftning, i enlighet med artikel 3 i direktiv 68/151/EEG, senast en månad före datum för den bolagsstämma vid vilken det skall beslutas om bildandet.
4. En eller flera oberoende experter i de initiativtagande bolagen, utsedda eller godkända enligt de nationella bestämmelser som antagits för att genomföra direktiv 78/855/EEG av en rättslig eller administrativ myndighet i den medlemsstat under vars lagstiftning vart och ett av bolagen faller, skall granska det enligt punkt 2 upprättade förslaget till bildande och avge ett skriftligt yttrande avsett för aktieägarna i varje bolag. Genom överenskommelse mellan de initiativtagande bolagen får ett skriftligt yttrande avges för aktieägarna i samtliga bolag av en eller flera oberoende experter utsedda eller godkända av en rättslig eller administrativ myndighet i den medlemsstat under vars lagstiftning av vilken något av de initiativtagande bolagen eller det blivande SE-bolaget omfattas enligt de nationella bestämmelser som antagits för att genomföra direktiv 78/855/EEG.
5. I yttrandet skall anges vilka särskilda problem värderingen har vållat och om aktiernas föreslagna utbytesförhållande är rättvist och rimligt, vilka metoder som använts för att fastställa det och om dessa metoder är adekvata i det aktuella fallet.
6. Bolagsstämman i vart och ett av de initiativtagande bolagen skall godkänna förslaget till bildande av ett SE-bolag.
Arbetstagarinflytandet i SE-bolaget skall avgöras i enlighet med direktiv 2001/86/EG och denna förordning. Bolagsstämman i vart och ett av de initiativtagande bolagen får förbehålla sig rätten att ställa som villkor för registrering av SE-bolaget att det uttryckligen bekräftar de riktlinjer som har beslutats på detta sätt.
7. Bestämmelserna i denna artikel skall i tillämpliga delar gälla för privata aktiebolag.
Artikel 33
1. Aktieägarna i de initiativtagande bolagen skall beredas tillfälle att inom tre månader meddela de initiativtagande bolagen om de har för avsikt att tillskjuta sina aktier för bildandet av SE-bolaget. Denna period skall börja samma dag som handlingen avseende bildandet av SE-bolaget har upprättats i enlighet med artikel 32.
2. SE-bolaget får bildas endast om aktie- eller andelsägarna i de initiativtagande bolagen inom den tid som anges i punkt 1 har tillskjutit den minimala procentuella andel aktier eller andelar i varje bolag som har fastställts i förslaget till bildande och om alla övriga villkor är uppfyllda.
3. Om samtliga villkor för bildandet av ett SE-bolag är uppfyllda i enlighet med punkt 2, skall detta offentliggöras för vart och ett av de initiativtagande bolagen enligt de bestämmelser i nationell lagstiftning för dessa bolag som antagits för att genomföra artikel 3 i direktiv 68/151/EEG.
De aktie- eller andelsägare i de initiativtagande bolag som inte inom den i punkt 1 angivna tiden har meddelat om de har för avsikt att ställa sina aktier till de initiativtagande bolagens förfogande för bildandet av ett SE-bolag skall beviljas en extra frist på en månad för att göra detta.
4. De aktieägare som har tillskjutit sina värdepapper för bildandet av SE-bolaget skall erhålla aktier i detta.
5. SE-bolaget får endast registreras mot intyg om att formaliteterna i artikel 32 och villkoren i punkt 2 ovan har uppfyllts.
Artikel 34
En medlemsstat får när det gäller de initiativtagande bolagen anta bestämmelser som avser att säkerställa skydd för minoritetsaktieägare som motsätter sig bildandet samt för borgenärer och arbetstagare.
Avsnitt 4
Bildande av ett SE-dotterbolag
Artikel 35
Ett SE-bolag får bildas i enlighet med artikel 2.3.
Artikel 36
För de bolag eller andra juridiska personer som deltar i bildandet gäller de bestämmelser som reglerar deras deltagande i bildandet av ett dotterbolag i form av ett publikt aktiebolag enligt nationell rätt.
Avsnitt 5
Ombildning av ett publikt aktiebolag till ett SE-bolag
Artikel 37
1. Ett SE-bolag kan bildas enligt artikel 2.4.
2. Utan att det påverkar tillämpningen av artikel 12 får ombildningen av ett publikt aktiebolag till ett SE-bolag inte innebära att bolaget avvecklas eller att en ny juridisk person skapas.
3. Bolagets säte får inte flyttas från en medlemsstat till en annan enligt artikel 8 i samband med ombildningen.
4. Det berörda bolagets lednings- eller förvaltningsorgan skall lämna ett förslag till ombildning och en redogörelse där juridiska och ekonomiska aspekter på ombildningen förklaras och motiveras och där det anges vilka verkningar antagandet av SE-bolagsformen får för aktieägarna och arbetstagarna.
5. Förslaget till villkor för ombildning skall offentliggöras på det sätt som föreskrivs i varje medlemsstats lagstiftning enligt artikel 3 i direktiv 68/151/EEG senast en månad före den bolagsstämma som sammankallas för att besluta om ombildningen.
6. Före den bolagsstämma som anges i punkt 7 skall en eller flera oberoende sakkunniga som, enligt de nationella bestämmelser som antagits för att tillämpa artikel 10 i direktiv 78/855/EEG, utsetts eller godkänts av en rättslig eller administrativ myndighet i den medlemsstat under vars lagstiftning bolaget under ombildning till SE-bolag lyder, med iakttagande av tillämpliga delar av rådets direktiv 77/91/EEG(8), intyga att bolaget förfogar över tillgångar som åtminstone motsvarar aktiekapitalet och de reserver som enligt lag eller enligt bolagsordningen inte får delas ut.
7. Bolagsstämman i det berörda bolaget skall godkänna förslaget till villkor för ombildningen samt SE-bolagets bolagsordning. Bolagsstämmans beslut skall godkännas genom omröstning på det sätt som föreskrivs i de nationella bestämmelser som antagits för att tillämpa artikel 7 i direktiv 78/855/EEG.
8. Medlemsstaterna kan göra ombildningen avhängig av kvalificerad röstmajoritet eller enhällighet i det organ i bolaget under ombildning inom vilket arbetstagarinflytandet organiseras.
9. Rättigheterna och skyldigheterna för bolaget under ombildning i fråga om sådana anställningsvillkor som omfattas av nationell lagstiftning, praxis och enskilda anställningskontrakt eller anställningsförhållanden och som föreligger vid tidpunkten för registreringen, skall med anledning av registreringen överföras till SE-bolaget.
AVDELNING III
SE-BOLAGS SAMMANSÄTTNING
Artikel 38
Ett SE-bolag skall enligt bestämmelserna i denna förordning bestå av
a) en bolagsstämma och
b) antingen ett tillsynsorgan och ett ledningsorgan (dualistiskt system) eller ett förvaltningsorgan (monistiskt system), beroende på vilket alternativ som fastställs i bolagsordningen.
Avsnitt 1
Dualistiskt system
Artikel 39
1. Ledningsorganet skall ansvara för SE-bolagets ledning och förvaltning. En medlemsstat kan föreskriva att en verkställande direktör eller verkställande direktörer skall ansvara för den löpande förvaltningen på samma villkor som gäller för publika aktiebolag med säte på denna medlemsstats territorium.
2. Ledamoten/ledamöterna i ledningsorganet skall väljas och entledigas av tillsynsorganet.
En medlemsstat får dock föreskriva eller ge möjlighet att i bolagsordningen föreskriva, att ledamoten/ledamöterna i ledningsorganet skall väljas och entledigas av bolagsstämman på samma sätt som sker i de publika aktiebolag som har sitt säte inom dess territorium.
3. Ingen får samtidigt vara ledamot i SE-bolagets ledningsorgan och dess tillsynsorgan. Dock får tillsynsorganet i händelse av vakans utse någon av sina ledamöter till ledamot i ledningsorganet. Under denna period upphävs tillfälligt dennes uppdrag som ledamot i tillsynsorganet. En medlemsstat får föreskriva att denna period skall vara tidsbegränsad.
4. Antalet ledamöter i ledningsorganet eller reglerna för hur detta antal skall bestämmas skall fastställas i SE-bolagets bolagsordning. Dock kan ett lägsta och/eller högsta antal fastställas av en medlemsstat.
5. En medlemsstat som saknar bestämmelser om ett dualistiskt system för publika aktiebolag med säte inom dess territorium får vidta lämpliga åtgärder rörande SE-bolag.
Artikel 40
1. Tillsynsorganet skall kontrollera ledningsorganets förvaltning. Det får inte för egen del ha några befogenheter att vidta förvaltningsåtgärder avseende SE-bolaget.
2. Ledamöterna i tillsynsorganet skall väljas av bolagsstämman. Dock får ledamöterna i det första tillsynsorganet utses i bolagsordningen. Denna bestämmelse gäller utan att detta påverkar tillämpningen av artikel 47.4 eller någon sådan ordning för arbetstagarnas medverkan som fastställs i enlighet med direktivet.
3. Bolagsordningen skall innehålla en bestämmelse om antalet ledamöter i tillsynsorganet eller regler för hur detta antal skall fastställas. En medlemsstat får dock föreskriva hur många ledamöter tillsynsorganet skall ha i de SE-bolag som är registrerade inom dess territorium eller hur många dessa minst och/eller högst skall vara.
Artikel 41
1. Ledningsorganet skall minst var tredje månad informera tillsynsorganet om SE-bolagets ekonomiska ställning och dess förutsebara framtida utveckling.
2. Utöver den periodiska informationen enligt punkt 1 skall ledningsorganet i god tid underrätta tillsynsorganet om alla händelser som kan ha påtagliga återverkningar på SE-bolaget.
3. Tillsynsorganet får från ledningsorganet begära in all den information som krävs för att det skall kunna utöva sin kontroll enligt artikel 40.1. En medlemsstat får föreskriva att även varje ledamot i tillsynsorganet skall ha denna möjlighet.
4. Tillsynsorganet får verkställa eller låta verkställa de kontroller som krävs för att det skall kunna fullgöra sitt uppdrag.
5. Var och en av ledamöterna av tillsynsorganet skall ha rätt att ta del av all information som tillställs detta organ.
Artikel 42
Tillsynsorganet skall välja en ordförande bland sina ledamöter. Om hälften av ledamöterna har utsetts av arbetstagarna, får endast en ledamot utsedd av bolagsstämman väljas till ordförande.
Avsnitt 2
Monistiskt system
Artikel 43
1. Förvaltningsorganet skall leda och förvalta SE-bolaget. En medlemsstat kan föreskriva att en verkställande direktör eller verkställande direktörer skall ansvara för den dagliga ledningen och förvaltningen på samma villkor som gäller för publika aktiebolag med säte på denna medlemsstats territorium.
2. Antalet ledamöter i förvaltningsorganet eller reglerna för hur detta antal skall bestämmas skall fastställas i SE-bolagets bolagsordning. Dock får en medlemsstat fastställa ett lägsta och, i förekommande fall, högsta antal ledamöter.
Detta förvaltningsorgan skall dock bestå av minst tre ledamöter, om arbetstagarnas medverkan är reglerad i enlighet med direktiv 2001/86/EG.
3. Ledamoten/ledamöterna i förvaltningsorganet skall väljas av bolagsstämman. Dock får ledamöterna av det första förvaltningsorganet utses i bolagsordningen. Dessa bestämmelser gäller utan att detta påverkar tillämpningen av artikel 47.4 eller någon sådan ordning för arbetstagarnas medverkan som fastställs i enlighet med direktiv 2001/86/EG.
4. Om det inte finns någon bestämmelse om ett monistiskt system beträffande publika aktiebolag med säte inom en medlemsstats territorium får denna medlemsstat anta lämpliga bestämmelser beträffande SE-bolag.
Artikel 44
1. Förvaltningsorganet skall sammanträda minst var tredje månad, med ett intervall som fastställs i bolagsordningen, för att diskutera SE-bolagets ekonomiska ställning och dess förutsebara framtida utveckling.
2. Var och en av ledamöterna i förvaltningsorganet skall ha rätt att ta del av all information som tillställs detta organ.
Artikel 45
Förvaltningsorganet skall välja en ordförande bland sina ledamöter. Om hälften av ledamöterna har utsetts av arbetstagarna, får endast en ledamot utsedd av bolagsstämman väljas till ordförande.
Avsnitt 3
Gemensamma regler för det monistiska och det dualistiska systemet
Artikel 46
1. Ledamöterna i organen skall utses för den period som fastställs i bolagsordningen och denna får inte vara längre än sex år.
2. Såvida inte bolagsordningen innehåller några inskränkningar, får ledamöterna omväljas en eller flera gånger för den period som fastställts enligt punkt 1.
Artikel 47
1. SE-bolagets bolagsordning får föreskriva att ett bolag eller en annan juridisk person skall ha rätt att vara ledamot i ett organ, såvida inte annat stadgas i den på publika aktiebolag tillämpliga lagen i den medlemsstat där SE-bolaget har sitt säte.
Bolaget eller annan juridisk person skall för utövandet av sina befogenheter i det aktuella organet utse en fysisk person till sin företrädare.
2. Till ledamöter i ett visst organ i ett SE-bolaget eller till företrädare för en ledamot enligt punkt 1 får inte väljas personer som
a) enligt lagen i den medlemsstat där SE-bolaget har sitt säte inte får ingå i motsvarande organ i ett publikt aktiebolag som faller under denna medlemsstats lagstiftning,
b) på grund av ett rättsligt eller administrativt avgörande meddelat i en medlemsstat inte får ingå i motsvarande organ i ett publikt aktiebolag som faller under lagstiftningen i en medlemsstat i gemenskapen.
3. SE-bolagets bolagsordning får, i likhet med vad som föreskrivs för publika aktiebolag i lagen i den medlemsstat där SE-bolaget har sitt säte, fastställa särskilda villkor för valbarhet beträffande de ledamöter som företräder aktieägarna.
4. Denna förordning påverkar inte tillämpningen av de nationella lagstiftningar som tillåter en minoritet av aktieägare eller andra personer eller myndigheter att välja en del av ledamöterna i organen.
Artikel 48
1. Ett SE-bolags bolagsordning skall innehålla en uppräkning av de kategorier av åtgärder för vilka tillsynsorganets medgivande måste inhämtas i det dualistiska systemet, eller för vilka det krävs ett uttryckligt beslut av förvaltningsorganet i det monistiska systemet.
Dock får en medlemsstat föreskriva att, i det dualistiska systemet, tillsynsorganet självt får besluta att dess medgivande skall inhämtas för vissa kategorier av åtgärder.
2. En medlemsstat får bestämma vilka kategorier av åtgärder som under alla omständigheter skall finnas upptagna i bolagsordningen för de SE-bolag som är registrerade på dess territorium.
Artikel 49
Ledamöterna av ett SE-bolags organ får inte, inte heller efter avslutat uppdrag, lämna någon information de innehar om SE-bolaget och vars röjande skulle kunna skada bolagets intressen, med undantag av de fall där ett sådant röjande krävs eller medges i bestämmelserna i den nationella lag som tillämpas på publika aktiebolag eller är av allmänt intresse.
Artikel 50
1. Utom i de fall då annat föreskrivs i denna förordning eller i bolagsordningen, skall de interna reglerna beträffande SE-organens beslutsförhet och beslutsfattande vara följande:
a) Beslutsförhet: minst hälften av ledamöterna skall vara närvarande eller företrädda.
b) Beslutsfattande: beslut fattas med majoriteten av de närvarande eller företrädda ledamöternas röster.
2. Om bolagsordningen inte innehåller några bestämmelser därom, skall varje organs ordförande ha utslagsröst vid lika röstetal. Dock får bolagsordningen inte innehålla några bestämmelser i strid härmed, om hälften av tillsynsorganets ledamöter företräder arbetstagarna.
3. Om arbetstagarmedverkan organiseras i enlighet med direktiv 2001/86/EG får en medlemsstat föreskriva att tillsynsorganets beslutsförhet och beslutsfattande, med undantag från punkt 1 och 2, skall regleras av de föreskrifter som under samma förhållanden gäller för publika aktiebolag som omfattas av den aktuella medlemsstatens lagstiftning.
Artikel 51
Ledamöterna i lednings-, tillsyns- eller förvaltningsorganet skall, i enlighet med de bestämmelser som gäller för publika aktiebolag i den medlemsstat där SE-bolaget har sitt säte, vara ansvariga för skada som tillfogas SE-bolaget till följd av att de har åsidosatt sina skyldigheter enligt lagen eller bolagsordningen eller andra skyldigheter som är förenade med deras uppdrag.
Avsnitt 4
Bolagsstämma
Artikel 52
Bolagsstämman skall besluta i de frågor som specifikt ankommer på stämman enligt
a) denna förordning,
b) bestämmelserna i lagstiftningen i den medlemsstat där SE-bolaget har sitt säte antagna med tillämpning av direktiv 2001/86/EG.
Vidare skall bolagsstämman besluta i de frågor för vilka bolagsstämman i ett publikt aktiebolag som faller under lagstiftningen i den medlemsstat där SE-bolaget har sitt säte är behörig, antingen enligt denna medlemsstats lag eller enligt den av samma lag reglerade bolagsordningen.
Artikel 53
Utan att det påverkar tillämpningen av reglerna i detta avsnitt, skall planeringen och genomförandet av bolagsstämman samt röstningsförfarandena regleras av lagstiftningen i den medlemsstat där SE-bolaget har sitt säte avseende publika aktiebolag.
Artikel 54
1. Bolagsstämman skall sammanträda minst en gång per kalenderår inom sex månader efter räkenskapsårets utgång, såvida inte lagstiftningen i den medlemsstat där SE-bolaget har sitt säte och som gäller för publika aktiebolag med samma typ av verksamhet som SE-bolag föreskriver tätare sammanträden. Dock får en medlemsstat föreskriva att den första bolagsstämman skall äga rum inom arton månader efter SE-bolagets bildande.
2. Bolagsstämman kan sammankallas när som helst av ledningsorganet, förvaltningsorganet, tillsynsorganet, eller av annat organ eller behörig myndighet i enlighet med den nationella lagen i den medlemsstat där SE-bolaget har sitt säte och som gäller för publika aktiebolag.
Artikel 55
1. Sammankallande av bolagsstämman och fastställande av dagordning får begäras av en eller flera aktieägare som tillsammans innehar aktier motsvarande minst 10 % av det tecknade aktiekapitalet, varvid en lägre procentsats får föreskrivas i bolagsordningen eller i den nationella lagen på samma villkor som gäller för publika aktiebolag.
2. I begäran om sammankallande skall anges vilka punkter som bör upptas på dagordningen.
3. Om efter den begäran som framställts enligt punkt 1 bolagsstämman inte hålls inom lämplig tid och i varje fall inte inom högst två månader, får den behöriga rättsliga eller administrativa myndigheten på den ort där SE-bolaget har sitt säte beordra att stämman skall sammankallas inom en bestämd tid och ge antingen de aktieägare som har begärt att så skall ske eller ett ombud för dessa rätt att sammankalla stämman. Detta påverkar inte tillämpningen av de nationella bestämmelser som eventuellt ger aktieägarna själva möjlighet att sammankalla bolagsstämman.
Artikel 56
En eller flera aktieägare som tillsammans innehar aktier motsvarande minst 10 % av det tecknade aktiekapitalet får begära att en eller flera nya punkter skall upptas på dagordningen för en bolagsstämma. De förfaranden och tidsfrister som gäller för denna begäran skall fastställas i den nationella lagen i den medlemsstat där SE-bolaget har sitt säte eller, om sådana bestämmelser saknas, i SE-bolagets bolagsordning. Den ovannämnda procentsatsen får sänkas i bolagsordningen eller i den nationella lagen på samma villkor som gäller för publika aktiebolag.
Artikel 57
Bolagsstämmans beslut skall fattas med majoriteten av de vederbörligen avgivna rösterna, såvida inte högre majoritet krävs enligt denna förordning eller, om den inte innehåller sådana bestämmelser, enligt den lag som gäller för publika aktiebolag i den medlemsstat där SE-bolaget har sitt säte.
Artikel 58
I de avgivna rösterna innefattas inte de som är knutna till aktier för vilka aktieägaren har underlåtit att delta i omröstningen eller har lagt ned sin röst eller röstat blankt eller avgivit ogiltig röst.
Artikel 59
1. För ändring av bolagsordningen krävs ett beslut av bolagsstämman fattat med en majoritet som inte får understiga två tredjedelar av de avgivna rösterna, såvida inte den lag som gäller för publika aktiebolag hemmahörande i den medlemsstat där SE-bolaget har sitt säte föreskriver eller medger högre majoritet.
2. Dock får en medlemsstat föreskriva att enkel majoritet av de i punkt 1 angivna rösterna skall räcka, när minst hälften av det tecknade aktiekapitalet är företrädd.
3. Ändringar av bolagsordningen för ett SE-bolag skall offentliggöras i enlighet med artikel 13.
Artikel 60
1. Då ett SE-bolag har två eller flera aktiekategorier, måste beslut av bolagsstämman föregås av en separat omröstning för varje kategori av aktieägare vilkas specifika rättigheter påverkas av beslutet.
2. Då bolagsstämmans beslut kräver den majoritet av rösterna som avses i artikel 59.1 och 59.2, skall denna majoritet också krävas för den separata omröstningen i varje kategori av aktieägare vilkas specifika rättigheter påverkas av beslutet.
AVDELNING IV
ÅRSBOKSLUT OCH KONCERNBOKSLUT
Artikel 61
Om inte annat följer av bestämmelserna i artikel 62 skall vad gäller upprättande av årsbokslut och, i förekommande fall, koncernbokslut, inbegripet den åtföljande verksamhetsberättelsen, samt revisionsberättelse och offentliggörande av boksluten SE-bolaget vara underkastat de regler som gäller för publika aktiebolag som omfattas av lagstiftningen i den medlemsstat där SE-bolaget har sitt säte.
Artikel 62
1. Ett SE-bolag som är kredit- eller finansinstitut skall i fråga om upprättande av årsbokslut och, i förekommande fall, koncernbokslut, inbegripet den åtföljande verksamhetsberättelsen, samt revisionsberättelse och offentliggörande av boksluten vara underkastade de regler som föreskrivs i den nationella lagen i den medlemsstat där SE-bolaget har sitt säte i enlighet med Europaparlamentets och rådets direktiv 2000/12/EG av den 20 mars 2000 om rätten att starta och driva verksamhet i kreditinstitut(9).
2. Ett SE-bolag som är försäkringsföretag skall i fråga om upprättande av årsbokslut och, i förekommande fall, koncernbokslut, inbegripet den åtföljande verksamhetsberättelsen, samt revisionsberättelse och offentliggörande av boksluten vara underkastade de regler som föreskrivs i den nationella lagen i den medlemsstat där SE-bolaget har sitt säte i enlighet med rådets direktiv 91/674/EEG av den 19 december 1991 om årsbokslut och sammanställd redovisning för försäkringsföretag(10).
AVDELNING V
AVVECKLING, LIKVIDATION, OBESTÅND OCH BETALNINGSINSTÄLLELSE
Artikel 63
Vad beträffar avveckling, likvidation, obestånd, betalningsinställelse och liknande förfaranden skall SE-bolaget vara underkastat bestämmelserna i den lag som skulle gälla för ett publikt aktiebolag bildat i enlighet med lagstiftningen i den medlemsstat där SE-bolaget har sitt säte, inbegripet bestämmelserna om bolagsstämmans beslutsfattande.
Artikel 64
1. Om ett SE-bolag inte längre uppfyller skyldigheten i artikel 7, skall den medlemsstat där SE-bolaget har sitt säte vidta lämpliga åtgärder för att få SE-bolaget att anpassa sig till gällande bestämmelser inom viss tid
a) antingen genom att flytta tillbaka sitt huvudkontor till den medlemsstat där det har sitt säte,
b) eller genom att flytta sitt säte enligt det förfarande som anges i artikel 8.
2. Den medlemsstat i vilken SE-bolagets huvudkontor är beläget skall vidta nödvändiga åtgärder för att säkerställa att ett SE-bolag som inte följer bestämmelserna i artikel 64.1 försätts i likvidation.
3. Den medlemsstat där SE-bolaget har sitt säte skall inleda ett rättsligt förfarande vid varje konstaterad överträdelse av bestämmelserna i artikel 7. Denna talan har suspensiv verkan på de förfaranden som avses i punkt 1 och 2.
4. Om det antingen på initiativ av myndigheterna eller på initiativ av en berörd part fastställs att ett SE-bolag har sitt huvudkontor i en medlemsstat i strid med artikel 7, skall myndigheterna i denna medlemsstat omgående underrätta den medlemsstat där SE-bolagets säte är förlagt.
Artikel 65
Inledande av ett avvecklings-, likvidations-, obestånds- eller betalningsinställelseförfarande samt avslutande av förfarandet och beslut att verksamheten får fortsätta skall offentliggöras i enlighet med artikel 13, utan att detta påverkar tillämpningen av sådana bestämmelser i den nationella lagstiftningen som föreskriver ytterligare åtgärder för offentliggörande.
Artikel 66
1. Ett SE-bolag får ombildas till ett publikt aktiebolag som faller under lagstiftningen i den medlemsstat där det har sitt säte. Beslutet om ombildning får inte fattas förrän två år efter SE-bolags registrering och inte förrän de första två årsredovisningarna har godkänts.
2. Ombildningen av ett SE-bolag till publikt aktiebolag innebär varken att det förra avvecklas eller att en ny juridiska person skapas.
3. Ett SE-bolags lednings- eller förvaltningsorgan skall upprätta ett förslag till ombildning och en redogörelse där ombildningens juridiska och ekonomiska aspekter förklaras och motiveras och där det anges vilka konsekvenser antagandet av bolagsformen SE-bolag får för aktieägare och arbetstagare.
4. Förslaget till ombildning skall offentliggöras på det sätt som föreskrivs i varje medlemsstats lagstiftning, i enlighet med artikel 3 i direktiv 68/151/EEG, senast en månad före datum för den bolagsstämma vid vilken fråga om godkännande av ombildningen skall behandlas.
5. Före den i punkt 6 avsedda bolagsstämman skall en eller flera oberoende experter, utsedda eller godkända enligt de nationella bestämmelser som antagits med tillämpning av artikel 10 i direktiv 78/855/EEG av en rättslig eller administrativ myndighet i den medlemsstat under vars lagstiftning det SE-bolag som skall ombildas till publikt aktiebolag lyder, intyga att bolaget förfogar över tillgångar som åtminstone motsvarar aktiekapitalet.
6. Ett SE-bolags bolagsstämma skall godkänna ombildningsförslaget samt det publika aktiebolagets bolagsordning. Bolagsstämmans beslut skall fattas på det sätt som föreskrivs i de nationella bestämmelser som antagits i enlighet med artikel 7 i direktiv 78/855/EEG.
AVDELNING VI
KOMPLETTERANDE BESTÄMMELSER OCH ÖVERGÅNGSBESTÄMMELSER
Artikel 67
1. Varje medlemsstat får, om och så länge som EMU:s tredje fas inte är tillämplig på staten i fråga, tillämpa samma bestämmelser på de SE-bolag som har sitt säte inom dess territorium som på de publika aktiebolag som faller under dess lagstiftning, vad beträffar i vilken valuta aktiekapitalet skall vara uttryckt. Ett SE-bolag får under alla omständigheter också uttrycka sitt aktiekapital i euro. I detta fall skall omräkningskursen mellan den nationella valutan och euron vara den som gäller den sista dagen i månaden före bildandet av SE-bolaget.
2. Om och så länge som EMU:s tredje fas inte är tillämplig på den medlemsstat där SE-bolaget har sitt säte, får emellertid SE-bolaget upprätta och offentliggöra sitt årsbokslut och, om så är lämpligt, sin koncernredovisning i euro. Medlemsstaten får kräva att SE-bolagets årsredovisning och, i förekommande fall, koncernredovisning upprättas och offentliggörs i nationell valuta på samma villkor som gäller för publika aktiebolag som omfattas av denna medlemsstats lagstiftning. Detta påverkar inte den möjlighet som ett SE-bolag har i enlighet med direktiv 90/604/EEG(11) att dessutom offentliggöra sin årsredovisning och, i förekommande fall, koncernredovisning i euro.
AVDELNING VII
SLUTBESTÄMMELSER
Artikel 68
1. Medlemsstaterna skall vidta alla lämpliga åtgärder för att säkerställa ett effektivt genomförande av denna förordning.
2. Varje medlemsstat skall utse de behöriga myndigheterna enligt artiklarna 8, 25, 26, 54, 55 och 64. Den skall underrätta kommissionen och de övriga medlemsstaterna om detta.
Artikel 69
Senast fem år efter det att denna förordning har trätt i kraft skall kommissionen förelägga rådet och Europaparlamentet en rapport om förordningens tillämpning och förslag om eventuella ändringar. Rapporten skall framför allt analysera lämpligheten av att
a) medge att ett SE-bolag har sitt huvudkontor och sitt säte i olika medlemsstater,
b) utvidga begreppet fusion i artikel 17.2 till att även tillåta andra typer av fusioner än de som anges i artiklarna 3.1 och 4.1 i direktiv 78/855/EEG,
c) se över klausulen om domstolsbehörighet i artikel 8.16 mot bakgrund av någon bestämmelse som kan ha införts i 1968 års Brysselkonvention eller i någon text som medlemsstaterna eller rådet antagit för att ersätta sådan konvention,
d) tillåta bestämmelser i ett SE-bolags bolagsordning genom lagar som en medlemsstat antar för att verkställa de befogenheter som medlemsstaterna har fått genom denna förordning, eller lagar som antas för att garantera en effektiv tillämpning av denna förordning på SE-bolag och som avviker från eller kompletterar dessa lagar, även när sådana bestämmelser inte är tillåtna i bolagsordningen för de publika aktiebolag som har sitt säte i medlemsstaten.
Artikel 70
Denna förordning träder i kraft den 8 oktober 2004.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 2430/2001
av den 12 december 2001
om komplettering av bilagan till förordning (EG) nr 2301/97 om att införa vissa benämningar i det %quot%register över skyddade särarter%quot% som föreskrivs i rådets förordning (EEG) nr 2082/92 om särartsskydd för jordbruksprodukter och livsmedel
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2082/92 av den 14 juli 1992 om särartsskydd för jordbruksprodukter och livsmedel(1), särskilt artikel 9.1 i denna, och
av följande skäl:
(1) Sverige har, i enlighet med artikel 7 i förordning (EEG) nr 2082/92, till kommissionen lämnat in en ansökan om att %quot%Falukorv%quot% skall registreras som särart.
(2) Det är endast för de benämningar som finns upptagna i registret som beteckningen %quot%garanterad traditionell specialitet%quot% får användas.
(3) Enligt artikel 8 i den förordningen framställdes ingen invändning till kommissionen till följd av offentliggörandet i Europeiska gemenskapernas officiella tidning(2) mot den beteckning som anges i bilagan till den här förordningen.
(4) Benämningen i bilagan förtjänar följaktligen att förtecknas i %quot%registret över skyddade särarter%quot% och därmed att skyddas enligt artikel 13.2 i förordning (EEG) nr 2082/92 som garanterad traditionell specialitet.
(5) Bilagan till den här förordningen kompletterar bilagan till kommissionens förordning (EG) nr 2301/97(3), senast ändrad genom förordning (EG) nr 1482/2000(4).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till förordning (EG) nr 2301/97 skall kompletteras med den benämning som anges i bilagan till den här förordningen och den skall förtecknas i %quot%registret över skyddade särarter%quot% enligt artikel 9.1 i förordning (EEG) nr 2082/92.
Den skall skyddas i enlighet med artikel 13.2 i den förordningen.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens beslut
av den 18 februari 2002
om en mall för föreläggande av en sammanfattning av nationella uppgifter om bränslekvalitet
[delgivet med nr K(2002) 508]
(2002/159/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets direktiv 98/70/EG av den 13 oktober 1998 om kvaliteten på bensin och dieselbränslen och om ändring av rådets direktiv 93/12/EEG(1), särskilt artikel 8.3 i detta, och
av följande skäl:
(1) För att uppfylla de miljöspecifikationer som anges i direktiv 98/70/EG och för att kunna se till att de åtgärder som vidtas för att minska utsläppen från motorfordon är effektiva, måste medlemsstaterna övervaka kvaliteten på bensin och dieselbränslen som saluförs på deras territorium.
(2) Det är nödvändigt att fastställa en gemensam mall för föreläggande av uppgifter om bränslekvalitet i enlighet med artikel 8.3 i direktiv 98/70/EG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Genom detta beslut fastställs en gemensam mall för föreläggande av nationella uppgifter om bränslekvalitet i enlighet med artikel 8 i direktiv 98/70/EG.
Artikel 2
Vid föreläggandet av uppgifter till kommissionen skall mallen i bilagan användas.
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 21 februari 2002
om ändring av bilaga D till rådets direktiv 90/426/EEG när det gäller test för diagnostisering av afrikansk hästpest
[delgivet med nr K(2002) 556]
(Text av betydelse för EES)
(2002/160/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 90/426/EEG av den 26 juni 1990 om djurhälsovillkor vid förflyttning och import av hästdjur från tredje land(1), senast ändrat genom direktiv 2001/298/EG(2), särskilt artikel 23 i detta, och
av följande skäl:
(1) I bilaga D till direktiv 90/426/EEG anges att komplementbindningstesten skall användas för diagnostisering av afrikansk hästpest.
(2) I november 2000 var gemenskapens referenslaboratorium i Algete i Spanien värd för det årliga mötet mellan medlemsstaternas nationella referenslaboratorier för afrikansk hästpest. Under mötet presenterades vetenskapliga rön som visar att komplementbindningstesten som för närvarande föreskrivs i bilaga D till direktiv 90/426/EEG har begränsningar av allvarlig art eftersom den endast lämpar sig för påvisande av antikroppar en kort tid efter infektion eller vaccination. Dessutom har testen i praktiken redan ersatts av moderna ELISA-tester vid nästan samtliga laboratorier i gemenskapen och även i de större exportländerna.
(3) Internationellt erkända laboratorietester för påvisande av antikroppar mot afrikansk hästpestvirus finns beskrivna i OIE:s (Internationella byrån för epizootiska sjukdomar) handbok för diagnostik och vaccination (Manual of Standards for Diagnosis and Vaccines)(3). I den nuvarande utgåvan anges emellertid bara en av de ELISA-tester som finns att tillgå.
(4) Bilaga D till direktiv 90/426/EEG bör därför ändras mot bakgrund av den tekniska utvecklingen och internationellt erkända normer.
(5) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga veterinärkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga D till direktiv 90/426/EEG skall ersättas med bilagan till detta beslut.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 18 december 2001
om genomförandebestämmelser för rådets beslut 2000/596/EG i fråga om förvaltnings- och kontrollsystem samt förfaranden för att genomföra finansiella korrigeringar beträffande åtgärder som medfinansieras av Europeiska flyktingfonden
[delgivet med nr K(2001) 4372]
(2002/307/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets beslut 2000/596/EG av den 28 september 2000 om inrättande av en europeisk flyktingfond(1), särskilt artikel 24 i detta,
efter samråd med den rådgivande kommitté som inrättats genom artikel 21.1 i beslut 2000/596/EG, och
av följande skäl:
(1) För att säkerställa en god finansiell förvaltning av de medel som beviljas genom Europeiska flyktingfonden (nedan kallad fonden) är det nödvändigt att medlemsstaterna upprättar riktlinjer för organisationen av de uppgifter som åligger den myndighet som ansvarar för genomförandet av medfinansierade åtgärder.
(2) För att gemenskapens resurser skall användas enligt principerna om en sund ekonomisk förvaltning måste medlemsstaternas förvaltnings- och kontrollsystem möjliggöra en tillfredsställande verifieringskedja, och medlemsstaterna måste lämna kommissionen allt nödvändigt bistånd vid genomförandet av kontroller, inbegripet stickprovskontroller.
(3) För att gemenskapens resurser skall användas på ett effektivt och korrekt sätt bör man fastställa enhetliga kriterier för de kontroller som medlemsstaterna genomför enligt artikel 18 i beslut 2000/596/EG.
(4) För att de utgiftsdeklarationer, för vilka betalning begärs enligt artikel 17.2 i beslut 2000/596/EG, skall kunna behandlas på ett enhetligt sätt bör ett standardformulär utarbetas för dessa deklarationer.
(5) För att möjliggöra återkrävande enligt artikel 18.1 i beslut 2000/596/EG av belopp som utbetalats på felaktiga grunder är det nödvändigt att föreskriva att uppdagade oegentligheter skall anmälas till kommissionen och att till anmälan skall fogas uppgifter om hur de administrativa eller rättsliga förfarandena har fortlöpt.
(6) Enligt artikel 19.1 i beslut 2000/596/EG skall medlemsstaterna genomföra finansiella korrigeringar i samband med enskilda eller systematiska oegentligheter genom att helt eller delvis dra in bidraget från gemenskapen. För att säkerställa att denna bestämmelse tillämpas på samma sätt i hela gemenskapen bör det fastställas bestämmelser om hur sådana korrigeringar skall beräknas och om rapportering till kommissionen.
(7) Om en medlemsstat inte uppfyller de krav som ställs på den enligt artikel 19.1 i beslut 2000/596/EG eller kraven i artikel 18 i beslutet, kan kommissionen själv göra de finansiella korrigeringarna med stöd av artikel 18.4 i beslutet. Det är lämpligt att beloppet för sådana korrigeringar alltid, när så är möjligt och genomförbart, beräknas utifrån handlingarna för det enskilda ärendet, och att det motsvarar de utgifter som felaktigt belastat fonden, varvid hänsyn skall tas till proportionalitetsprincipen. Om det inte är möjligt eller genomförbart att exakt kvantitativt fastställa värdet av de finansiella konsekvenserna av oegentligheten, eller om det skulle strida mot proportionalitetsprincipen att avföra samtliga de utgifter det gäller, bör kommissionen fastställa korrigeringen genom extrapolering eller genom att fastställa en klumpsumma utifrån den värdering som den gjort av omfattningen och de finansiella konsekvenserna av den oegentlighet som medlemsstaten har underlåtit att förebygga, påvisa eller korrigera.
(8) Det är nödvändigt att fastställa vissa former för genomförandet av de finansiella korrigeringar som avses i artikel 19.1 i beslut 2000/596/EG och att föreskriva att samma former skall tillämpas i de fall som avses i artikel 18.4 b i det beslutet.
(9) Det bör fastställas procentsatser för dröjsmålsräntan på belopp som blir föremål för återkrav och skall återbetalas till kommissionen enligt artikel 19.3 i beslut 2000/596/EG.
(10) Tillämpningen av detta beslut bör inte påverka bestämmelserna om återkrav av statligt stöd enligt artikel 14 i rådets förordning (EG) nr 659/1999 av den 22 mars 1999 om tillämpningsföreskrifter för artikel 93 i EG-fördraget(2).
(11) Tillämpningen av detta beslut bör inte påverka bestämmelserna i rådets förordning (Euratom, EG) nr 2185/96 av den 11 november 1996 om de kontroller och inspektioner på platsen som kommissionen utför för att skydda Europeiska gemenskapernas finansiella intressen mot bedrägerier och andra oegentligheter(3).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
KAPITEL I
TILLÄMPNINGSOMRÅDE OCH DEFINITIONER
Artikel 1
I detta beslut fastställs tillämpningsföreskrifter för rådets beslut 2000/596/EG när det gäller förvaltnings- och kontrollsystem för sådana bidrag från Europeiska flyktingfonden (nedan kallad fonden), som förvaltas av medlemsstaterna, samt förfarandet för tillämpliga finansiella korrigeringar av sådana bidrag.
Artikel 2
I detta beslut avses med
a) ansvarig instans: varje myndighet som utsetts av en medlemsstat i enlighet med artikel 7 i beslut 2000/596/EG,
b) förmedlande organ: alla offentliga förvaltningar eller icke-statliga organisationer till vilka en ansvarig instans delegerar genomförandeansvar i enlighet med artikel 7 i beslut 2000/596/EG.
KAPITEL II
FÖRVALTNINGS- OCH KONTROLLSYSTEM
Artikel 3
1. För tillämpningen av artikel 18.1 c i beslut 2000/596/EG skall varje medlemsstat meddela riktlinjer till den ansvariga instansen och till förmedlande organ som tilldelats delegerat ansvar för genomförandet.
Utan att detta skall påverka artikel 18.1 i beslut 2000/596/EG, skall riktlinjerna omfatta organisationen av de förvaltnings- och kontrollsystem som är nödvändiga för att säkerställa att ansökningarna om bistånd från gemenskapen är välgrundade, korrekta och berättigade till bidrag, och de skall utformas med beaktande av de allmänt erkända normer för god förvaltningssed som redovisas i bilaga 1.
2. För det fall då samtliga eller vissa av den ansvariga instansens uppgifter har delegerats till förmedlande organ skall det, i de riktlinjer som avses i punkt 1, bl.a. anges former för genomförandet av följande uppgifter:
a) Att klart definiera och fördela uppgifterna, bl.a. i fråga om förvaltning, utbetalning, kontroll och undersökning av överensstämmelsen med
i) de villkor som fastställs i kommissionens beslut om godkännande av de ansökningar om medfinansiering som avses i artikel 8 i beslut 2000/596/EG,
ii) de regler för stödberättigande för utgifter som anges i bilaga I till kommissionens beslut 2001/275/EG(4), och
iii) gemenskapens politik och åtgärder, bl.a. när det gäller konkurrensregler, offentlig upphandling, skydd och förbättring av miljön, avlägsnande av ojämlikhet och främjande av jämställdhet.
b) Att upprätta effektiva system för att säkerställa att de förmedlande organen utövar sina befogenheter på ett tillfredsställande sätt.
c) Att meddela upplysningar till den ansvariga instansen om det faktiska genomförandet av uppgifterna och redovisa de medel som använts för detta.
3. Enligt artikel 18.1 b i beslut 2000/596/EG skall varje medlemsstat senast två månader efter det att detta beslut trätt i kraft, och utöver upplysningarna i den första ansökningen om medfinansiering, överlämna en beskrivning av de inrättade förvaltnings- och kontrollsystemen samt av de förbättringar som planeras, särskilt med hänsyn till de allmänt erkända normer för god förvaltningssed som redovisas i bilaga 1.
Detta meddelande skall innehålla följande upplysningar beträffande varje ansvarig instans:
a) De uppgifter som instansen tilldelats.
b) Arbetsfördelningen, som inom den ansvariga instansen eller det förmedlande organet skall säkerställa att tillräcklig åtskillnad upprätthålls mellan förvaltnings-, utbetalnings- och kontrollfunktionerna för att en god finansiell förvaltning skall kunna garanteras.
c) Uppgifter om eventuella förmedlande organ.
d) Förfarandena vid mottagning, kontroll och godkännande av betalningsansökningarna samt för betalningsförordnande, utbetalning och utgiftsredovisning.
e) Bestämmelser om internrevision eller motsvarande förfaranden.
4. Kommissionen skall i samarbete med medlemsstaten granska förvaltnings- och kontrollsystemen och påvisa eventuella hinder som dessa medför för insynen i kontrollerna av fondens funktion och av att kommissionen fullgjort sitt ansvar enligt artikel 274 i fördraget.
Artikel 4
1. I medlemsstaternas förvaltnings- och kontrollsystem skall det finnas en tillfredsställande verifieringskedja.
2. En verifieringskedja skall anses tillfredsställande om den gör det möjligt att kontrollera
a) att de sammanlagda belopp som redovisats till kommissionen överensstämmer med enskilda utgiftsposter med tillhörande verifikationer som förvaras på de olika administrativa nivåerna och hos stödmottagarna, inbegripet de organ eller företag som ansvarar för genomförandet av projekten, och
b) hur de tillgängliga medlen från gemenskapen och de nationella medlen fördelas och överförs.
I bilaga II finns en vägledande beskrivning av de informationskrav som en tillfredsställande verifieringskedja skall uppfylla.
3. Den ansvariga instansen skall upprätta förfaranden som säkerställer att förvaringsplatsen för alla de dokument som avser enskilda utgifter inom det nationella genomförandeprogrammet finns registrerad, och att dessa dokument hålls tillgängliga för kontroll när så begärs av
a) personalen på den myndighet som ansvarar för behandlingen av betalningsansökningarna,
b) de nationella revisionsmyndigheterna, som skall utföra de kontroller som föreskrivs i artikel 5.1 i detta beslut,
c) den avdelning eller det organ inom den ansvariga instansen som ansvarar för den attestering av ansökningar om förskott eller slutbetalningar som avses i artikel 17 i beslut 2000/596/EG, och
d) bemyndigade tjänstemän och ombud från kommissionen och revisionsrätten.
De tjänstemän eller ombud som ansvarar för kontrollerna eller personer som givits sådana befogenheter får begära att kopior av de dokument som avses i den här punkten skall överlämnas till dem.
4. Under de fem år som följer efter kommissionens slutbetalning i samband med en åtgärd skall de ansvariga myndigheterna för kommissionen hålla tillgängliga samtliga verifikationer som rör utgifterna och kontrollerna för den berörda åtgärden, antingen i form av originalhandlingar eller i form av bestyrkta kopior på allmänt erkända datamedier. Rättsliga förfaranden eller en motiverad begäran från kommissionen skall ha suspensiv verkan på denna tidsfrist.
Artikel 5
1. Medlemsstaterna skall genomföra kontroller avseende ett lämpligt urval av projekt, särskilt för att
a) kontrollera att förvaltnings- och kontrollsystemen fungerar väl, och
b) selektivt, på grundval av en riskanalys, kontrollera de utgiftsdeklarationer som upprättats på olika berörda nivåer.
2. De kontroller som genomförs skall omfatta åtminstone 20 % av de totala stödberättigande utgifterna inom varje nationellt genomförandeprogram och grundas på ett representativt urval av godkända projekt med beaktande av bestämmelserna i punkt 3. Medlemsstaterna skall se till att sådana kontroller på lämpligt sätt hålls åtskilda från förfarandena för genomförande av insatser och därmed sammanhängande utbetalningar.
3. De utvalda projekten skall anges, urvalsmetoden beskrivas och en rapport sammanställas om resultaten av samtliga inspektioner och om åtgärder som vidtagits med anledning av konstaterade avvikelser och oegentligheter.
4. Urvalet av projekt för kontroll skall
a) omfatta projekt av tillräckligt varierande typ och omfattning,
b) beakta riskfaktorer som identifierats vid nationella kontroller eller gemenskapskontroller, och
c) ta hänsyn till om projekten koncentrerats till vissa stödmottagare, så att de mest betydande stödmottagarna kontrolleras åtminstone en gång innan varje slag av nationellt genomförandeprogram avslutas.
Artikel 6
Vid kontrollerna skall medlemsstaterna kontrollera följande:
a) Att förvaltnings- och kontrollsystemen fungerar effektivt.
b) Att det finns ett lämpligt antal relevanta redovisningshandlingar med tillhörande verifikationer hos de förmedlande organ som tilldelats visst ansvar för genomförandet av den ansvariga instansen, stödmottagarna och, i tillämpliga fall, de andra organ eller företag som genomför projekt.
c) Att det finns en tillfredsställande verifieringskedja.
d) Att typen av utgifter och de datum då de verkställdes uppfyller kraven i gemenskapens bestämmelser, de nationella bestämmelser som fastställts i samband med urvalsförfarandet och villkoren i avtalet eller handlingen om beviljande av stöd, samt att de avser faktiskt utförda insatser.
e) Att projektets faktiska eller planerade syften överensstämmer med de syften som beskrivs i det nationella genomförandeprogram som avses i artikel 8 i beslut 2000/596/EG.
f) Att gemenskapens finansiella bidrag ligger inom de gränser som anges i artikel 13 i beslut 2000/596/EG eller i andra tillämpliga gemenskapsbestämmelser, samt att de betalats ut till de slutliga stödmottagarna utan avdrag eller dröjsmål.
g) Att den nationella medfinansiering som krävs faktiskt har ställts till förfogande.
h) Att de medfinansierade insatserna har genomförts med iakttagande av bestämmelserna i artikel 4 och artikel 9.1 i beslut 2000/596/EG
Artikel 7
Genom kontrollerna skall det fastställas huruvida eventuella problem som förekommit är betingade av det tillämpade systemet och således innebär en risk för andra insatser som samma slutliga stödmottagare utför eller som administreras av samma förmedlande organ. De skall också identifiera orsakerna till sådana situationer, vilka ytterligare undersökningar som kan bli nödvändiga, samt nödvändiga korrigerande och förebyggande åtgärder.
Artikel 8
Medlemsstaterna skall årligen, genom den rapport som avses i artikel 20.2 i beslut 2000/596/EG, underrätta kommissionen om hur de under det föregående året har tillämpat artiklarna 5, 6 och 7 och därvid i tillämpliga fall komplettera eller uppdatera den beskrivning som avses i artikel 4.2.
Artikel 9
För insatser som mer än en medlemsstat deltar i eller som avser stödmottagare i mer än en medlemsstat skall de berörda medlemsstaterna och kommissionen komma överens om vilket administrativt bistånd som krävs för att säkerställa att kontrollerna håller erforderlig kvalitet.
KAPITEL III
UTGIFTSDEKLARATIONER
Artikel 10
1. Intyg om utgiftsdeklarationer skall upprättas enligt mallen i bilaga IV av en person eller enhet inom den ansvariga instansen som är oberoende av varje enhet som förordnar om utbetalningar.
2. Den ansvariga instansen skall i samband med varje utgiftsdeklaration avge en försäkran till kommissionen om att de nationella genomförandeprogrammen förvaltas i enlighet med all tillämplig gemenskapslagstiftning och att medlen används enligt principerna om en sund ekonomisk förvaltning. I denna deklaration skall intygas att ansökningen om medfinansiering inte avser andra slag av utgifter än sådana som
a) faktiskt betalats av stödmottagarna, enligt definitionen i artikel 2 d i beslut 2001/275/EG under den stödperiod som programmet avser enligt vad som anges i den relevanta artikeln i besluten om godkännande av medfinansieringsansökningar, och som
b) avser projekt som valts ut för medfinansiering inom det nationella genomförandeprogrammet enligt de fastställda urvalskriterierna och urvalsförfarandena och som har förvaltats i enlighet med gemenskapsbestämmelserna under hela den tid som utgifterna i fråga hänför sig till.
3. När ett program avslutas skall medlemsstaten inom sex månader överlämna en slutlig rapport enligt bilaga IV. Om ingen sådan sänds till kommissionen inom denna tidsfrist, avslutar kommissionen automatiskt programmet och de krediter som ingår i det.
4. Innan den ansvariga instansen sänder en ansökan till kommissionen, skall den förvissa sig om att tillräckliga kontroller har utförts. Det arbete som utförts skall redovisas ingående i den rapport som avses i artikel 20.3 i beslut 2000/596/EG. Kontrollerna skall avse såväl det praktiska genomförandet av projekten och graden av effektivitet som finansiella och redovisningsmässiga aspekter.
KAPITEL IV
FINANSIELLA KORRIGERINGAR SOM GÖRS AV MEDLEMSSTATERNA
Artikel 11
1. Vid oegentligheter som är betingade av systemets uppbyggnad skall undersökningen enligt artikel 19.1 i beslut 2000/596/EG omfatta samtliga transaktioner som kan vara berörda.
2. När gemenskapens bidrag helt eller delvis dras in, skall medlemsstaterna ta hänsyn till oegentligheternas art och omfattning samt till den ekonomiska förlusten för fonden.
3. Medlemsstaterna skall som bilaga till den rapport som avses i artikel 20.2 i beslut 2000/596/EG till kommissionen överlämna en förteckning över de förfaranden för indragande av stöd som inletts under det föregående året.
Artikel 12
1. När belopp skall återkrävas efter det att medfinansieringen dragits in enligt artikel 18.1 g i beslut 2000/596/EG, skall den behöriga avdelningen eller det behöriga organet inleda ett återkravsförfarande och rapportera detta till den ansvariga instansen. Kommissionen skall underrättas om återkraven, som skall redovisas i enlighet med artikel 13 i det här beslutet.
2. Medlemsstaterna skall i den rapport som avses i artikel 20.2 i beslut 2000/596/EG underrätta kommissionen om sina beslut eller förslag avseende ändrad tilldelning av de indragna beloppen.
Artikel 13
Den ansvariga instansen skall bokföra de belopp som skall återkrävas i fråga om redan utbetalat gemenskapsstöd, och de skall se till att dessa belopp återkrävs utan onödigt dröjsmål. Efter återkravet skall den ansvariga instansen i tillämpliga fall minska den följande utgiftsdeklarationen till kommissionen med ett belopp som motsvarar återkravet eller, om detta är otillräckligt, göra en återbetalning till gemenskapen. Utöver de belopp som skall återkrävas skall ränta betalas från förfallodagen med den procentsats som föreskrivs i artikel 94 i kommissionens förordning (EURATOM, EKSG, EG) nr 3418/93 av den 9 december 1993 om närmare bestämmelser för genomförandet av vissa bestämmelser i budgetförordningen av den 21 december 1977(5), senast ändrad genom förordning (EG) nr 1687/2001(6), för den första vardagen i den månad då fordringen förfaller till betalning.
När medlemsstaterna översänder den rapport som avses i artikel 20.2 i beslut 2000/596/EG, skall de bifoga en förteckning över påvisade oegentligheter med uppgift om belopp som återkrävts eller skall återkrävas samt i tillämpliga fall de administrativa och rättsliga förfaranden som inletts för återkrav av på felaktiga grunder utbetalda belopp.
KAPITEL V
FINANSIELLA KORRIGERINGAR SOM GÖRS AV KOMMISSIONEN
Artikel 14
1. Beloppen för de finansiella korrigeringar som görs av kommissionen enligt artikel 18.4 b i beslut 2000/596/EG för enskilda eller systematiska oegentligheter skall alltid när så är möjligt och praktiskt genomförbart fastställas på grundval av enskilda ärenden och motsvara de utgifter som felaktigt belastat fonderna, med beaktande av proportionalitetsprincipen.
2. Om det inte är möjligt eller praktiskt genomförbart att exakt bestämma det belopp som omfattas av en oegentlighet eller om det skulle vara oproportionerligt att helt dra in de berörda utgifterna, skall kommissionen grunda sina finansiella korrigeringar på antingen
a) en extrapolering, och därvid använda ett representativt urval av transaktioner med likartade egenskaper, eller
b) ett schablonbelopp, och därvid bedöma överträdelsens allvar samt omfattningen och de finansiella effekterna av den konstaterade oegentligheten.
3. När kommissionen grundar sitt ställningstagande på förhållanden som påvisats av utomstående revisorer, skall den själv bedöma de finansiella konsekvenserna av dessa efter att ha granskat de åtgärder som den berörda medlemsstaten vidtagit med tillämpning av artikel 18.1 i beslut 2000/596/EG.
4. Den tidsfrist inom vilken den berörda medlemsstaten skall besvara en förfrågan enligt artikel 18.3 i beslut 2000/596/EG skall vara två månader. I vederbörligen motiverade fall kan kommissionen bevilja en längre tidsfrist.
5. Om kommissionen föreslår en finansiell korrigering som fastställts genom extrapolering eller schablonmässigt, skall medlemsstaten ges möjlighet att med stöd av de berörda akterna visa, att oegentlighetens faktiska omfattning var mindre än enligt kommissionens bedömning. Efter överenskommelse med kommissionen får medlemsstaten begränsa omfattningen av undersökningen till en lämplig andel eller ett lämpligt urval av de berörda akterna. Utom i vederbörligen motiverade fall får förlängningen av tidsfristen för denna undersökning inte överskrida en ytterligare period av två månader efter den tvåmånadersperiod som anges i punkt 4. Kommissionen skall ta hänsyn till allt bevismaterial som medlemsstaterna tillhandahåller inom dessa tidsfrister.
6. Om kommissionen har inställt betalningar enligt artikel 19.2 i beslut 2000/596/EG och skälen till detta kvarstår vid utgången av den tidsfrist som anges i punkt 4, eller om den berörda medlemsstaten inte har underrättat kommissionen om de åtgärder som har vidtagits för att rätta till oegentligheterna, skall artikel 18.4 i beslut 2000/596/EG tillämpas.
7. Riktlinjer omfattande principerna och kriterierna samt vägledande skalor för kommissionens korrigeringar med schablonbelopp redovisas i bilaga III till detta beslut.
Artikel 15
1. Varje återbetalning till kommissionen enligt artikel 19.3 i beslut 2000/596/EG skall göras inom den tidsfrist som anges i ett föreläggande om återbetalning som upprättas enligt artikel 28 i budgetförordningen av den 21 december 1977(7). Utgången av denna tidsfrist skall vara slutet av den andra månaden efter det att föreläggandet utfärdades.
2. Varje försening av en återbetalning skall leda till att dröjsmålsränta tas ut från och med den förfallodag som anges i punkt 1 till och med den dag då beloppet faktiskt återbetalas. Tillämplig räntesats skall vara den som anges i artikel 13 i detta beslut.
3. En finansiell korrigering enligt artikel 19.2 i beslut 2000/596/EG skall inte påverka medlemsstatens skyldighet att återkräva medel enligt artikel 18.1 g i beslut 2000/596/EG och artikel 12.1 i detta beslut eller att återkräva statligt stöd enligt artikel 14 i förordning (EG) nr 659/1999.
KAPITEL VI
SLUTBESTÄMMELSER
Artikel 16
Detta beslut skall inte hindra medlemsstaterna från att tillämpa striktare nationella bestämmelser än de som fastställs genom detta beslut.
Artikel 17
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 17 juli 2002
om frågeformulär gällande rådets direktiv 96/82/EG om åtgärder för att förebygga och begränsa följderna av allvarliga olyckshändelser där farliga ämnen ingår
[delgivet med nr K(2002) 2656]
(2002/605/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 96/82/EG av den 9 december 1996 om åtgärder för att förebygga och begränsa följderna av allvarliga olyckshändelser där farliga ämnen ingår(1), särskilt artikel 19.4 i detta, och
av följande skäl:
(1) Enligt artikel 19.4 i direktiv 96/82/EG skall medlemsstaterna vart tredje år rapportera om genomförandet av detta direktiv.
(2) Rapporten skall upprättas på grundval av ett frågeformulär eller utkast som kommissionen utarbetat, i enlighet med det förfarande som anges i artikel 6 i direktiv 91/692/EEG av den 23 december 1991 om att standardisera och rationalisera rapporteringen om genomförandet av vissa direktiv om miljön(2).
(3) Treårsperioden bör omfatta åren 2003-2005.
(4) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från den kommitté som upprättats genom artikel 6 i direktiv 91/692/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Frågeformuläret i bilagan antas härmed.
Artikel 2
Medlemsstaterna skall utarbeta en rapport för perioden 2003-2005, i överensstämmelse med frågeformuläret i bilagan.
Artikel 3
Medlemsstaterna skall lämna treårsrapporten till kommissionen senast den 30 september 2006.
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
Rådets beslut
av den 22 juli 2002
om ingående på Europeiska gemenskapens vägnar av konventionen om bevarande och förvaltning av fiskeresurser i Sydostatlanten
(2002/738/EG)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 37 jämförd med artikel 300.2 första stycket första meningen och artikel 300.3 första stycket i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europaparlamentets yttrande(2), och
av följande skäl:
(1) Gemenskapen är behörig att i fråga om fiskeresurser anta bevarande- och förvaltningsåtgärder och att ingå avtal med andra länder eller internationella organisationer.
(2) Gemenskapen är avtalsslutande part i Förenta nationernas havsrättskonvention, enligt vilken samtliga medlemmar i det internationella samfundet skall samarbeta om bevarande och förvaltning av havets biologiska resurser.
(3) Gemenskapen har undertecknat avtalet om genomförande av bestämmelserna i Förenta nationernas havsrättskonvention av den 10 december 1982 om bevarande och förvaltning av gränsöverskridande och långvandrande fiskbestånd(3), men den har ännu inte avslutat ratifikationsförfarandet.
(4) Gemenskapen har sedan 1997 tillsammans med regionens kuststater och andra berörda parter deltagit aktivt i utarbetandet av en konvention om bevarande och förvaltning av fiskeresurser i Sydostatlanten. Gemenskapen undertecknade konventionen den 20 april 2001 under diplomatkonferensen i Windhoek, Namibia, i enlighet med det beslut som rådet fattat i detta syfte(4).
(5) Fiskare från gemenskapen bedriver fiske i det område som omfattas av konventionen. Det ligger följaktligen i gemenskapens intresse att bli fullvärdig medlem av den regionala fiskeriorganisation som skall upprättas genom konventionen. Gemenskapen bör därför godkänna konventionen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Konventionen om bevarande och förvaltning av fiskeresurser i Sydostatlanten godkänns härmed på gemenskapens vägnar.
Texten till konventionen åtföljer detta beslut.
Artikel 2
Rådets ordförande bemyndigas att utse den eller de personer som skall ha rätt att deponera instrumentet avseende godkännande hos generaldirektören för Förenta nationernas livsmedels- och jordbruksorganisation i enlighet med artikel 25.2 i konventionen.
Kommissionens beslut
av den 16 december 2002
om fortsatta jämförande försök och tester i gemenskapen när det gäller utsäde och förökningsmaterial av gramineae, Triticum aestivum, Vitis vinifera, Brassica napus och Allium ascalonicum inom ramen för rådets direktiv 66/401/EEG, 66/402/EEG, 68/193/EEG, 92/33/EEG, 2002/54/EG, 2002/55/EG, 2002/56/EG och 2002/57/EG
(Text av betydelse för EES)
(2002/984/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 66/401/EEG av den 14 juni 1966 om saluföring av utsäde av foderväxter(1), senast ändrat genom direktiv 2001/64/EG(2),
med beaktande av rådets direktiv 66/402/EEG av den 14 juni 1966 om saluföring av utsäde av stråsäd(3), senast ändrat genom direktiv 2001/64/EG,
med beaktande av rådets direktiv 68/193/EEG av den 9 april 1968 om saluföring av vegetativt förökningsmaterial av vinstockar(4), senast ändrat genom direktiv 2002/11/EG(5),
med beaktande av rådets direktiv 92/33/EEG av den 28 april 1992 om saluförande av annat föröknings- och plantmaterial av grönsaker än utsäde(6), senast ändrat genom kommissionens beslut 2002/111/EG(7),
med beaktande av rådets direktiv 2002/54/EG av den 13 juni 2002 om saluföring av betutsäde(8),
med beaktande av rådets direktiv 2002/55/EG av den 13 juni 2002 om saluföring av utsäde av köksväxter(9),
med beaktande av rådets direktiv 2002/56/EG av den 13 juni 2002 om saluföring av utsädespotatis(10),
med beaktande av rådets direktiv 2002/57/EG av den 13 juni 2002 om saluföring av utsäde av olje- och spånadsväxter(11), senast ändrat genom direktiv 2002/68/EG(12),
med beaktande av kommissionens beslut 2001/897/EG av den 12 december 2001 om villkor för gemenskapens jämförande försök och tester av utsäde och förökningsmaterial från vissa växter enligt rådets direktiv 66/400/EEG, 66/401/EEG, 66/402/EEG, 66/403/EEG, 68/193/EEG, 69/208/EEG, 70/458/EEG och 92/33/EEG(13), särskilt artikel 3 i detta, och
av följande skäl:
(1) I beslut 2001/897/EG fastställs villkor för gemenskapens jämförande försök och tester som skall genomföras i enlighet med rådets direktiv 66/401/EEG, 66/402/EEG, 68/193/EEG, 92/33/EEG, 2002/54/EG, 2002/55/EG, 2002/56/EG och 2002/57/EG fr.o.m. 2002 t.o.m. 2003.
(2) De försök och tester som genomfördes 2002 bör fortsätta under 2003.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Enda Artikel
Gemenskapens jämförande försök och tester som inleddes 2002 för utsäde och förökningsmaterial av gramineae, Triticum aestivum, Brassica napus, Allium ascalonicum och Vitis vinifera skall fortsätta under 2003 i enlighet med beslut 2001/897/EG.
Europaparlamentets och rådets beslut nr 1600/2002/EG
av den 22 juli 2002
om fastställande av gemenskapens sjätte miljöhandlingsprogram
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 175.3 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
med beaktande av Regionkommitténs yttrande(3),
i enlighet med förfarandet i artikel 251 i fördraget(4), på grundval av det gemensamma utkast som förlikningskommittén godkände den 1 maj 2002, och
av följande skäl:
(1) En ren och hälsosam miljö är en förutsättning för vårt samhälles välbefinnande och välfärd, men fortsatt tillväxt på global nivå kommer att medföra att miljön utsätts för fortsatt belastning.
(2) Gemenskapens femte miljöhandlingsprogram %quot%Mot en hållbar utveckling%quot% löpte ut den 31 december 2000, och har medfört en rad viktiga förbättringar.
(3) Fortsatta ansträngningar krävs för att uppfylla de miljömål som gemenskapen redan fastställt och det finns ett behov av det sjätte miljöhandlingsprogram (nedan kallat %quot%programmet%quot%) som fastställs genom detta beslut.
(4) Ett antal allvarliga miljöproblem återstår att lösa och nya håller på att framträda som kräver ytterligare insatser.
(5) Det krävs större koncentration på förebyggande och på tillämpning av försiktighetsprincipen när en strategi för skydd av människors hälsa och miljön skall utvecklas.
(6) Försiktig användning av naturresurserna och skydd av det globala ekosystemet utgör tillsammans med ekonomisk välfärd och en balanserad social utveckling förutsättningarna för hållbar utveckling.
(7) Programmet syftar till en hög skyddsnivå för miljön och för människors hälsa och till en allmän förbättring av miljön och livskvaliteten. Programmet anger vidare prioriteringar för miljödimensionen i strategin för hållbar utveckling, och bör beaktas när åtgärder läggs fram enligt strategin.
(8) Programmet syftar till att bryta sambandet mellan belastning på miljön och ekonomisk tillväxt samtidigt som det är förenligt med subsidiaritetsprincipen och respekterar de många skilda förutsättningar som råder i Europeiska unionens olika regioner.
(9) Genom programmet fastställs miljöprioriteringar för gemenskapens åtgärder med inriktning särskilt på klimatförändringar, natur och biologisk mångfald, miljö och hälsa och livskvalitet, samt naturresurser och avfall.
(10) För vart och ett av dessa områden anges övergripande mål och vissa delmål och ett antal åtgärder fastställs för att nå målen. Dessa mål och delmål utgörs av prestanda eller av resultat som skall eftersträvas.
(11) De mål, prioriteringar och åtgärder som anges i programmet bör bidra till en hållbar utveckling i kandidatländerna och vara uttryck för en strävan efter att säkerställa skyddet av naturvärdena i dessa länder.
(12) Lagstiftningen är av avgörande betydelse om miljömålen skall nås, och ett fullständigt och korrekt genomförande av gällande lagstiftning kommer därför att prioriteras. Andra möjligheter för att uppnå miljömål bör också övervägas.
(13) Programmet bör främja processen för integration av miljöhänsyn i all gemenskapspolitik och verksamhet i enlighet med artikel 6 i fördraget för att minska belastning på miljön från olika källor.
(14) Det krävs ett integrerat strategiskt tillvägagångssätt där nya former för samarbete med marknaden införs, som engagerar medborgarna, företagen och övriga intressenter för att få till stånd de nödvändiga förändringarna både i produktionen och i de offentliga och privata konsumtionsmönster som påverkar miljöns tillstånd och utveckling negativt. Detta tillvägagångssätt bör uppmuntra en hållbar användning och förvaltning av land och hav.
(15) Möjlighet att få tillgång till information i miljöfrågor och till överprövning samt allmänhetens deltagande i beslutsfattandet kommer att vara viktigt för programmets framgång.
(16) I de temainriktade strategierna kommer hänsyn att tas till det utbud av möjligheter och instrument som krävs för att behandla en rad komplicerade frågor som kräver ett öppet och flerdimensionellt synsätt, och nödvändiga åtgärder kommer att föreslås, och om så är lämpligt kommer Europaparlamentet och rådet att engageras.
(17) Inom vetenskapliga kretsar råder det enighet om att mänsklig verksamhet leder till ökade koncentrationer av växthusgaser, vilket i sin tur medför högre temperaturer globalt sett och störningar av klimatet.
(18) Följderna av klimatförändringar kan allvarligt påverka vårt samhälle och naturen och måste minskas. Åtgärder som leder till minskade utsläpp av växthusgaser kan genomföras utan att tillväxt- och välfärdsnivåerna sänks.
(19) Oavsett om insatserna för att minska påverkan lyckas eller inte, måste samhället anpassas till och förberedas för följderna av klimatförändringar.
(20) Sunda naturliga system som befinner sig i balans är en förutsättning för livet på vår jord.
(21) Mänsklig verksamhet medför betydande belastning på naturen och den biologiska mångfalden. Åtgärder krävs för att motverka belastning särskilt i form av föroreningar, införande av främmande arter, potentiella risker från utsättning av genetiskt modifierade organismer och det sätt på vilket land och hav exploateras.
(22) Mark är en begränsad resurs som står under miljöbelastning.
(23) Trots förbättringar av miljönormerna ökar sannolikheten för en koppling mellan miljöförstöring och vissa sjukdomar hos människor. Därför bör man ta itu med de potentiella risker som uppkommer till exempel från utsläpp och farliga kemikalier, bekämpningsmedel och buller.
(24) Det krävs större kunskaper om de potentiella negativa verkningarna av användning av kemikalier, och ansvaret för att utveckla kunskaperna bör ligga på tillverkarna, importörerna och användare i efterföljande led.
(25) Kemikalier som är farliga bör ersättas med säkrare kemikalier eller säkrare alternativ teknik som inte medför användning av kemikalier, i syfte att minska riskerna för människor och för miljön.
(26) Bekämpningsmedel bör användas på ett hållbart sätt så att riskerna för människors hälsa och för miljön minskas.
(27) Omkring 70 % av befolkningen lever i stadsmiljö och gemensamma ansträngningar behövs för att garantera bättre miljö och livskvalitet i städerna.
(28) Vår planets förmåga att motsvara de ökade kraven på resurser och att absorbera de utsläpp och det avfall som blir följden av resursanvändningen är begränsad och det finns tecken på att den nuvarande efterfrågan i många fall är högre än vad miljön kan bära.
(29) Gemenskapens avfallsvolym fortsätter att växa och en betydande mängd av detta avfall är farligt, vilket leder till förlust av resurser och ökade risker för förorening.
(30) Den ekonomiska globaliseringen innebär att miljöåtgärder allt oftare behövs på internationell nivå, däribland inom transportpolitiken, vilket kräver nya åtgärder från gemenskapen inom politikområden som handel, utveckling samt yttre förbindelser för att möjliggöra att hållbar utveckling eftersträvas i andra länder. God förvaltning bör bidra till att detta ändamål uppnås.
(31) Handel, internationella investeringsflöden och exportkrediter bör lämna ett större bidrag till miljöskydd och hållbar utveckling.
(32) Med tanke på frågornas komplexa natur måste beslutsfattandet på miljöområdet grundas på bästa tillgängliga vetenskapliga och ekonomiska bedömningar, och på kunskap om miljöns tillstånd och utvecklingstendenser i enlighet med artikel 174 i fördraget.
(33) Information till beslutsfattare, berörda parter och till allmänheten måste vara relevant, tydlig, aktuell och lättbegriplig.
(34) Framstegen i fråga om att nå miljömålen måste mätas och utvärderas.
(35) På grundval av en bedömning av miljöns tillstånd, med beaktande av den information som regelbundet lämnas av Europeiska miljöbyrån, bör efter halva programtiden de framsteg som gjorts ses över och en bedömning göras av huruvida programmets inriktning behöver ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Programmets räckvidd
1. Genom detta beslut upprättas ett program för gemenskapsåtgärder på miljöområdet, nedan kallat %quot%programmet%quot%. I programmet behandlas de huvudsakliga miljömålen och miljöprioriteringarna, vilka grundas på en bedömning av miljöförhållanden och aktuella trender, inklusive nyligen uppkomna problem, och som kräver ett initiativ från gemenskapens sida. Programmet skall främja integreringen av miljöhänsyn på alla gemenskapens politikområden och bidra till att en hållbar utveckling uppnås i hela den nuvarande och i den framtida utvidgade gemenskapen. Programmet skall vidare sörja för fortlöpande insatser för att de miljömål som redan fastställts av gemenskapen skall uppnås.
2. I programmet fastställs de huvudsakliga miljömål som skall uppnås. Där fastställs, där så är lämpligt, delmål och tidsplaner. Målen och delmålen bör uppnås innan programmet löper ut, om inte något annat anges.
3. Programmet skall omfatta en period på tio år från och med 22 juli 2002. I syfte att uppfylla målen skall lämpliga initiativ inom de olika politikområdena bestå av en rad åtgärder, som inbegriper lagstiftning och de strategier som beskrivs i artikel 3. Dessa initiativ bör läggas fram successivt, dock senast fyra år efter det att detta beslut har antagits.
4. Målen motsvarar de huvudsakliga miljöprioriteringarna för gemenskapen på områdena
- klimatförändringar,
- natur och biologisk mångfald,
- miljö och hälsa samt livskvalitet,
- naturresurser och avfall.
Artikel 2
Principer och övergripande syften
1. Programmet utgör en ram för gemenskapens miljöpolitik under programtiden i syfte att ge en hög skyddsnivå, varvid hänsyn skall tas till subsidiaritetsprincipen och till olikheterna i olika regioner inom gemenskapen, och att bryta sambandet mellan belastning på miljön och ekonomisk tillväxt. Det skall särskilt grundas på principen om att förorenaren skall betala, försiktighetsprincipen och principen om förebyggande åtgärder samt principen om åtgärdande av föroreningar vid källan.
Programmet skall utgöra grunden för miljödimensionen i strategin för hållbar utveckling i Europa och bidra till att miljöhänsyn införlivas i gemenskapens samtliga politikområden bland annat genom att ange miljöprioriteringar för strategin.
2. Programmet syftar till följande:
- Att betona att klimatförändringar kommer att vara en utomordentligt stor utmaning under de kommande tio åren och även därefter samt att bidra till det långsiktiga målet att uppnå en stabilisering av koncentrationerna av växthusgaser i atmosfären på en nivå som kan förhindra farlig antropogen inverkan på klimatsystemet. Därför skall ett långsiktigt mål på en maximal global temperaturhöjning på 2 °Celsius över de förindustriella nivåerna och en CO2-koncentration under 550 ppm styra programmet. På lång sikt kräver detta troligen en global minskning av utsläppen av växthusgaser med 70 % jämfört med 1990 års nivåer i enlighet med vad som har fastställts av Mellanstatliga panelen för klimatförändringar (IPCC).
- Att skydda, bevara, återställa och utveckla de naturliga systemens, de naturliga livsmiljöernas samt vilda växters och djurs sätt att fungera i syfte att hejda ökenspridningen och förlusten av biologisk mångfald, inklusive mångfalden av genetiska resurser, både i Europeiska unionen och globalt sett.
- Att bidra till hög livskvalitet och social välfärd för medborgarna genom att sörja för en miljö där föroreningsnivåerna inte leder till skadliga konsekvenser för människors hälsa eller för miljön och genom att stödja en hållbar stadsutveckling.
- Bättre resurseffektivitet, resurshushållning och avfallshantering för att säkerställa mer hållbara produktions- och konsumtionsmönster, så att resursanvändning och uppkomsten av avfall inte längre kopplas till graden av ekonomisk tillväxt och en strävan att säkerställa att användningen av förnybara och icke-förnybara resurser inte ställer större krav på miljön än vad denna förmår bära.
3. Programmet skall säkerställa att miljömålen, vilka bör inriktas på de miljöresultat som skall åstadkommas, uppnås genom de mest effektiva och lämpliga metoder som finns att tillgå, med beaktande av de principer som anges i punkt 1 och de strategier som beskrivs i artikel 3. Full hänsyn skall tas till säkerställandet av att gemenskapens miljöpolitiska beslut fattas på ett integrerat sätt och till alla till buds stående möjligheter och instrument, med beaktande av regionala och lokala olikheter samt ekologiskt känsliga områden och med tonvikten på
- utvecklandet av europeiska initiativ som syftar till att höja medvetenheten hos medborgarna och de lokala myndigheterna,
- en omfattande dialog med berörda parter, höjande av medvetenheten om miljöfrågor och allmänhetens medverkan,
- kostnads-nyttoanalys och hänsyn till behovet av att internalisera miljökostnaderna,
- bästa tillgängliga vetenskapliga data och förbättrade vetenskapliga kunskaper genom forskning och teknisk utveckling,
- data och information om miljöförhållanden och miljötrender.
4. Programmet skall främja en fullständig integrering av miljöskyddskrav i gemenskapens övriga politik och åtgärder genom att det där fastställs miljömål och, när så är lämpligt, delmål och tidsplaner, som skall beaktas inom de relevanta politikområdena.
Föreslagna och antagna åtgärder till förmån för miljön bör dessutom överensstämma med målen för den ekonomiska och sociala dimensionen av en hållbar utveckling och omvänt.
5. Programmet skall främja antagandet av politik och strategier som bidrar till att hållbar utveckling uppnås i de länder som är kandidater för anslutning (nedan kallade %quot%kandidatländerna%quot%) och som bygger på att gemenskapens regelverk överförs och genomförs. Utvidgningsprocessen bör stödja och skydda kandidatländernas miljövärden, till exempel rik biologisk mångfald, och bör bevara och stärka hållbara produktions- och konsumtions- samt markanvändningsmönster och miljömässigt sunda transportstrukturer genom
- integrering av miljöskyddskrav i gemenskapens program, inklusive sådana som har samband med utveckling av infrastrukturer,
- främjande av överföring av ren teknik till kandidatländerna,
- utvidgning av dialogen och utbytet av erfarenheter med kandidatländernas nationella och lokala förvaltningar om hållbar utveckling och bevarande av ländernas miljötillgångar,
- samarbete med det civila samhället, icke-statliga miljöorganisationer och näringsliv i kandidatländerna för att hjälpa till att öka allmänhetens medvetenhet och medverkan,
- uppmuntran till internationella finansinstitut och den privata sektorn att stödja genomförandet och efterlevnaden av gemenskapens regelverk på miljöområdet i kandidatländerna samt på lämpligt sätt beakta integrering av miljöhänsyn i den ekonomiska sektorns verksamhet.
6. Programmet skall stimulera
- Europeiska unionens positiva och konstruktiva roll som en ledande partner vid skyddet av den globala miljön och strävan efter att uppnå en hållbar utveckling,
- utvecklingen av ett globalt partnerskap för miljön och en hållbar utveckling,
- integrering av miljöhänsyn och miljömål i alla aspekter av gemenskapens yttre förbindelser.
Artikel 3
Strategier för att uppnå miljömålen
För att uppnå de syften och mål som fastställs i detta program skall bland annat följande medel användas:
1. Utarbetande av ny gemenskapslagstiftning och ändring av gällande lagstiftning, när så är lämpligt.
2. Främjande av ett effektivare genomförande och upprätthållande av gemenskapens miljölagstiftning, utan att det hindrar kommissionen att inleda överträdelseförfaranden. För detta krävs följande:
- Ökade åtgärder för att förbättra respekten för gemenskapens miljöskyddsregler och åtgärder för att ta itu med överträdelser av miljölagstiftningen.
- Främjande av bättre standarder för medlemsstaternas tillståndsgivning, inspektion, övervakning och verkställighet.
- En mer systematisk översyn av tillämpningen av miljölagstiftningen i samtliga medlemsstater.
- Förbättrat informationsutbyte om bästa metoder i fråga om genomförande, inklusive genom Europeiska nätverket för genomförande och upprätthållande av miljölagstiftning (Impel-nätverket) inom ramen för dess behörighet.
3. Ytterligare insatser behövs för att integrera miljöskyddskrav i förberedandet, fastställandet och genomförandet av gemenskapspolitik och gemenskapsverksamhet inom olika politikområden. Ytterligare insatser är nödvändiga inom olika sektorer, inklusive övervägande av särskilda miljömål, delmål, tidsplaner och indikatorer. För detta krävs
- säkerställande av att de integreringsstrategier som rådet utvecklar inom olika politikområden effektivt omsätts i praktiken och bidrar till genomförandet av programmets syften och mål för miljön,
- övervägande, innan åtgärder på det sociala och ekonomiska området antas, om huruvida dessa åtgärder bidrar till och stämmer överens med målen, delmålen och tidsramen för programmet,
- inrättande av lämpliga interna regelbundna mekanismer i gemenskapsinstitutionerna - varvid full hänsyn skall tas till behovet av att främja öppenhet och tillgång till information - för att säkerställa att miljöhänsyn fullt ut återspeglas i kommissionens politiska initiativ, inbegripet relevanta beslut och lagstiftningsförslag,
- regelbunden övervakning med hjälp av relevanta indikatorer, om möjligt framtagna på grundval av en gemensam metod för varje sektor, och rapportering om den sektoriella integreringsprocessen,
- ytterligare integrering av miljökriterier i gemenskapens finansieringsprogram, utan att redan befintliga kriterier påverkas,
- att miljökonsekvensbedömning och strategisk miljöbedömning används och genomförs fullt ut och effektivt,
- att hänsyn bör tas till målen i programmet i framtida översyner av budgetplanen för gemenskapens finansieringsorgan.
4. Främjande av hållbara produktions- och konsumtionsmönster genom effektivt genomförande av de principer som anges i artikel 2 i syfte att internalisera såväl de negativa som de positiva miljökonsekvenserna genom att utnyttja en kombination av styrmedel, inklusive marknadsbaserade och ekonomiska styrmedel. För detta krävs bland annat följande:
- Uppmuntra reformer av sådana subventioner som har avsevärda negativa miljökonsekvenser och är oförenliga med en hållbar utveckling, bland annat genom att senast vid halvtidsöversynen upprätta en förteckning över kriterier som gör det möjligt att registrera sådana subventioner som har negativ inverkan på miljön i syfte att avveckla dem stegvis.
- Analysera miljöeffektiviteten av överlåtbara miljötillstånd som ett allmänt styrmedel och handel med utsläppsrätter i syfte att främja och genomföra användningen av dessa när det är möjligt.
- Främja och uppmuntra skatteåtgärder såsom miljörelaterade skatter och incitament på lämplig nationell nivå eller på gemenskapsnivå.
- Främja integreringen av miljöskyddskrav i standardiseringsverksamheten.
5. Förbättrat samarbete och partnerskap med företag och deras representativa organ samt att engagera arbetsmarknadens parter, konsumenterna och deras organisationer i lämplig omfattning med syftet att förbättra företagens miljöprestanda och eftersträva hållbara produktionsmönster. För detta krävs
- främjande, genom hela programmet, av en integrerad produktpolitik, som uppmuntrar till beaktande av miljökraven genom produkternas hela livscykel och till en vidare tillämpning av miljövänliga processer och produkter,
- främjande av ett mer omfattande utnyttjande av gemenskapens miljölednings- och miljörevisionsordning (EMAS)(5) och utarbetande av sådana initiativ som uppmuntrar företagen att offentliggöra mycket noggranna rapporter som redogör för deras miljöprestanda eller deras insatser för en hållbar utveckling och som genomgått en oberoende granskning,
- införandet av ett stödprogram för hjälp med efterlevnaden, med särskilda stödåtgärder för små och medelstora företag,
- uppmuntra införandet av program för belöning av företags miljöprestanda,
- uppmuntran till innovation av produkter i syfte att göra marknaden mer miljöanpassad, bl.a. genom förbättrad spridning av resultaten av Life-programmet(6),
- främjande av frivilliga åtaganden och avtal för att uppnå tydliga miljömål, inklusive att bestämma vad som skall ske om dessa inte efterlevs.
6. Att bidra till att säkerställa att enskilda konsumenter, företag och offentliga organ i deras egenskap av köpare får tillgång till bättre information om vilka miljökonsekvenser olika processer och produkter har, i syfte att uppnå hållbara konsumtionsmönster. För detta krävs
- stöd till användande av miljömärkning och andra typer av miljöinformation och sådan märkning som ger konsumenterna möjlighet att jämföra miljöprestandan hos produkter av samma typ,
- stöd till användande av tillförlitliga miljöuppgifter från tillverkarna och förebyggande av missvisande uppgifter,
- främjande av en miljövänlig offentlig upphandlingspolitik, som gör det möjligt att ta hänsyn till miljöfaktorer och integrera miljöhänsyn i ett livscykelperspektiv, inklusive produktionsfasen, i upphandlingsförfarandena, dock i överensstämmelse med gemenskapens konkurrensregler och den inre marknaden, med riktlinjer för bästa metoder och inledande av en översyn av miljöanpassad upphandling i gemenskapsinstitutionerna.
7. Att stödja integrering av miljöhänsyn i den finansiella sektorn. För detta krävs
- övervägande av frivilliga initiativ tillsammans med den finansiella sektorn, som omfattar riktlinjer för införandet av uppgifter om miljökostnader i företagens årsredovisningar samt utbyte av bästa metoder mellan medlemsstater,
- uppmaning till Europeiska investeringsbanken att i större utsträckning integrera miljömål och miljööverväganden i låneverksamheten, särskilt i syfte att stödja en hållbar utveckling i kandidatländerna,
- stöd för integration av miljömål och miljöhänsyn i verksamheten i andra finansinstitut, t.ex. Europeiska banken för återuppbyggnad och utveckling (EBRD).
8. För att skapa en ansvarsordning för gemenskapen krävs bland annat
- lagstiftning om miljöansvar.
9. Främjande av den europeiska allmänhetens förståelse och engagemang för miljöfrågor och förbättrande av samarbete och partnerskap med konsumentgrupper och icke-statliga organisationer, kräver
- säkerställande av tillgång till information och deltagande samt till överprövning genom att gemenskapen och medlemsstaterna med det snaraste ratificerar Århuskonventionen(7),
- stöd för tillhandahållandet av lättillgänglig information till medborgarna om miljöförhållanden och miljötrender i förhållande till sociala och ekonomiska tendenser och hälsoutvecklingen,
- ett allmänt höjande av medvetenheten om miljöfrågor,
- utvecklande av allmänna regler och principer för god miljöförvaltning genom samrådsprocesser.
10. Effektiv och hållbar användning och förvaltning av land och hav med beaktande av miljöhänsyn skall uppmuntras och främjas. För detta krävs, samtidigt som subsidiaritetsprincipen efterlevs fullt ut, följande:
- Främjande av bästa metoder avseende hållbar markanvändning, varvid hänsyn skall tas till särskilda regionala omständigheter, med särskild betoning på programmet för integrerad förvaltning av kustområden.
- Främjande av bästa metoder och stödjande av nätverk som gynnar utbyte av erfarenheter av hållbar utveckling, vilket innefattar stadsområden, havs-, kust- och bergsområden, våtmarker och andra känsliga områden.
- Ökad användning, ökade resurser och större räckvidd för miljöåtgärder inom jordbruket inom ramen för den gemensamma jordbrukspolitiken.
- Uppmuntran till medlemsstaterna att överväga användningen av regional planering som ett instrument för att förbättra miljöskyddet för medborgarna och främja erfarenhetsutbytet om hållbar regional utveckling, särskilt när det gäller stadsområden och tättbefolkade områden.
Artikel 4
Temainriktade strategier
1. Åtgärder i enlighet med artiklarna 5-8 skall inbegripa utformning av temainriktade strategier och utvärdering av de befintliga strategier för prioriterade miljöproblem som kräver ett brett upplagt angreppssätt. Dessa strategier bör omfatta ett fastställande av vilka förslag som behövs för att målen i programmet skall uppnås samt de planerade förfarandena för antagandet. Dessa strategier skall tillställas Europaparlamentet och rådet och vid behov utformas som ett beslut av Europaparlamentet och rådet och skall antas i enlighet med förfarandet i artikel 251 i fördraget. Om inte annat följer av förslagets rättsliga grund skall de lagstiftningsförslag som bygger på dessa strategier antas i enlighet med förfarandet i artikel 251 i fördraget.
2. De temainriktade strategierna kan inbegripa sådana strategier som skisseras i artiklarna 3 och 9 samt relevanta kvalitativa och kvantitativa miljömål och tidsplaner, mot vilka de planerade åtgärderna kan mätas och utvärderas.
3. De temainriktade strategierna bör utarbetas och genomföras i nära samråd med relevanta parter, såsom icke-statliga organisationer, näringslivet, arbetsmarknadens övriga parter och offentliga myndigheter, och i förekommande fall bör det säkerställas att samråd med kandidatländerna ingår i denna process.
4. De tematiska strategierna bör presenteras för Europaparlamentet och rådets senast inom tre år efter det att programmet har antagits. Den halvtidsrapport i vilken kommissionen skall utvärdera de framsteg som har gjorts beträffande genomförandet av programmet skall omfatta en översyn av de temainriktade strategierna.
5. Kommissionen skall årligen rapportera till Europaparlamentet och rådet om framsteg i utarbetandet och genomförandet av strategierna samt om deras effektivitet.
Artikel 5
Mål och prioriterade områden för att hantera klimatförändringar
1. De syften som anges i artikel 2 bör tillgodoses genom att följande mål uppnås:
- Ratificering och ikraftträdande av Kyotoprotokollet till Förenta nationernas ramkonvention om klimatförändringar senast 2002 och uppfyllande av åtagandet enligt detta om att utsläppen för Europeiska gemenskapen som helhet senast 2008-2012 skall minskas med 8 % jämfört med 1990 års nivåer, i enlighet med varje enskild medlemsstats åtagande enligt rådets slutsatser av den 16-17 juni 1998.
- Påvisbara framsteg senast 2005 i fråga om uppfyllande av åtagandena enligt Kyotoprotokollet.
- Uppnående av en position som gör gemenskapen trovärdig i arbetet för ett internationellt avtal som fastställer mer långtgående mål om minskade utsläpp för den andra åtagandeperioden enligt Kyotoprotokollet. Målsättningen med detta avtal bör vara att minska utsläppen väsentligt, varvid full hänsyn bland annat skall tas till resultaten i den tredje utvärderingsrapporten från den mellanstatliga panelen för klimatförändringar (IPCC), och ta hänsyn till behovet av en global, rättvis fördelning av utsläppen av växthusgaser.
2. Dessa mål skall eftersträvas med hjälp av bland annat följande prioriterade åtgärder:
i) Genomförande av internationella klimatåtaganden, inklusive Kyotoprotokollet, genom
a) att studera resultaten av det europeiska klimatförändringsprogrammet och anta effektiva gemensamma och samordnade politiska riktlinjer och åtgärder för olika sektorer på grundval av detta, när det är lämpligt, för att komplettera nationella åtgärder i medlemsstaterna,
b) att verka för upprättandet av en gemenskapsram för att utveckla en fungerande handel med utsläppsrätter för CO2, vilken eventuellt kan utvidgas till att omfatta andra växthusgaser,
c) att förbättra övervakningen av växthusgaser och av hur medlemsstaterna lyckas uppfylla sina åtaganden enligt den interna överenskommelsen om bördefördelningen.
ii) Minskning av utsläppen av växthusgaser inom energisektorn:
a) Så snart som möjligt göra en genomgång och översyn av subventioner som motverkar en effektiv och hållbar energianvändning, i syfte att gradvis avveckla dem.
b) Uppmuntra användning av förnybara och fossila bränslen med lägre kolhalt för kraftproduktion.
c) Främja användningen av förnybara energikällor, inbegripet genom att vidta olika stimulansåtgärder, även på lokal nivå, i syfte att senast år 2010 uppnå det vägledande målet om 12 % av den totala energianvändningen.
d) Vidta stimulansåtgärder som främjar kraftvärme samt genomföra åtgärder för att fördubbla den totala andelen kraftvärme i gemenskapen som helhet, så att den uppgår till 18 % av den totala bruttoelproduktionen.
e) Förhindra och minska metanutsläpp från energiproduktion och energidistribution.
f) Främja energieffektivitet.
iii) Minskning av utsläppen av växthusgaser inom transportsektorn:
a) Fastställa och genomföra särskilda åtgärder för att minska utsläpp av växthusgaser från luftfarten, om man inte enas om sådana åtgärder inom ramen för Internationella civila luftfartsorganisationen (ICAO) senast 2002.
b) Fastställa och genomföra särskilda åtgärder för att minska utsläpp av växthusgaser från marin sjöfart, om man inte enas om sådana åtgärder inom Internationella sjöfartsorganisationen senast 2003.
c) Främja en övergång till effektivare och renare transportformer, inklusive bättre organisation och logistik.
d) Inom ramen för EU:s mål om en minskning med 8 % av utsläppen av växthusgaser uppmana kommissionen att före utgången av 2002 lägga fram ett meddelande om kvantifierade miljömål för ett hållbart transportsystem,
e) Fastställa och genomföra ytterligare särskilda åtgärder, inbegripet lämplig lagstiftning, för att minska utsläpp av växthusgaser, även N2O, från motorfordon.
f) Främja utveckling och användning av alternativa bränslen, samt fordon med låg bränsleförbrukning, i syfte att avsevärt och oavbrutet öka deras andel.
g) Främja åtgärder som återspeglar de totala miljökostnaderna i priset på transporttjänsterna.
h) Bryta kopplingen mellan ekonomisk tillväxt och efterfrågan på transporter i syfte att minska miljöpåverkan.
iv) Minskning av utsläppen av växthusgaser inom industriproduktionen:
a) Främja miljöeffektiva metoder och teknik inom industrin.
b) Ta fram metoder för att hjälpa små och medelstora företag att anpassa, förnya och förbättra sin verksamhet.
c) Stödja utvecklingen av miljömässigt sunda och tekniskt genomförbara alternativ, inbegripet fastställande av gemenskapsåtgärder, som syftar till att minska utsläppen, successivt avveckla produktionen där så är lämpligt och genomförbart samt minska användningen av fluorerade gaser HFC (vätefluorkolföreningar), FC (perfluorerade kolväten) och SF6 (svavelhexafluorid).
v) Minskning av utsläppen av växthusgaser inom andra sektorer:
a) Främja energieffektivitet, framför allt när det gäller uppvärmning, kylning och varmvattenförsörjning vid planering av byggnader.
b) Beakta behovet av att minska utsläppen av växthusgaser tillsammans med andra miljöhänsyn i den gemensamma jordbrukspolitiken och i gemenskapens strategi för avfallshantering.
vi) Användning av andra lämpliga styrmedel, t.ex. följande:
a) Främja tillämpningen av skatteåtgärder, inklusive att i rätt tid införa ett lämpligt ramverk för energibeskattning på gemenskapsnivå, för att uppmuntra till en övergång till effektivare energianvändning, renare energi och transporter och för att främja tekniska innovationer.
b) Främja miljöavtal med näringslivets sektorer om minskade utsläpp av växthusgaser.
c) Säkerställa att klimatförändringar blir ett tema av största vikt såväl i gemenskapens politik för forskning och teknisk utveckling som i nationella forskningsprogram.
3. Utöver att begränsa klimatförändringar bör gemenskapen förbereda insatser för anpassning till konsekvenserna av klimatförändringar, bland annat genom följande:
- Översyn av gemenskapspolitiken, i synnerhet de delar som berör klimatförändringar, så att behovet av anpassning beaktas tillräckligt i alla investeringsbeslut.
- Främjande av regionala klimatmodeller och bedömningar, både för att förbereda regionala anpassningsåtgärder, till exempel förvaltning av vattenresurser, bevarande av biologisk mångfald och förhindrande av ökenspridning och översvämningar, och för att bidra till att öka medborgarnas och näringslivets medvetenhet.
4. Det måste säkerställas att, vid gemenskapens utvidgning, hänsyn tas till den utmaning som klimatförändringarna innebär. Detta kommer bl.a. att kräva följande åtgärder beträffande kandidatländerna:
- Stödjande av kapacitetsuppbyggnad, för att nationella åtgärder skall kunna vidtas som möjliggör användning av Kyoto-mekanismerna samt förbättrad rapportering och övervakning av utsläppen.
- Främjande av en mer hållbar transport- och energisektor.
- Säkerställande av att samarbetet med kandidatländerna förstärks ytterligare när det gäller frågor om klimatförändringar.
5. Bekämpandet av klimatförändringar kommer att utgöra en integrerad del av Europeiska unionens politik i fråga om yttre förbindelser och utgöra en av prioriteringarna i unionens politik för en hållbar utveckling. Detta kommer att kräva gemensamma och samordnade insatser från gemenskapens och medlemsstaternas sida för att
- bygga upp kapacitet för att bistå utvecklingsländerna och länder med övergångsekonomier, till exempel genom att främja projekt under Kyotoprotokollets mekanismer för ren utveckling (CDM) och gemensamt genomförande (JI),
- bistå med tekniköverföring där behov identifieras, och
- bistå de berörda länderna i den utmaning som en anpassning till klimatförändringarna innebär.
Artikel 6
Mål och prioriterade områden för insatser avseende natur och biologisk mångfald
1. De syften som anges i artikel 2 bör tillgodoses genom att följande mål uppnås:
- Stoppa förlusten av biologisk mångfald i syfte att uppnå detta mål senast 2010, bl.a. genom att förhindra och mildra effekterna av främmande arter och främmande genotyper.
- Skydda mot skadliga föroreningar och på lämpligt sätt återställa natur och biologisk mångfald.
- Bevara, på lämpligt sätt återställa och på ett hållbart sätt nyttja havsmiljö, kuster och våtmarker.
- Bevara och på lämpligt sätt återställa särskilt natursköna områden, inklusive odlade och känsliga områden.
- Bevara arter och livsmiljöer, och särskilt förebygga fragmentering av livsmiljöer.
- Främja hållbart nyttjande av mark, med särskild uppmärksamhet på förebyggande av erosion, förstöring, förorening och ökenspridning.
2. Dessa mål skall uppnås bland annat med hjälp av följande prioriterade åtgärder, med beaktande av subsidiaritetsprincipen och på grundval av gällande globala och regionala konventioner och strategier och fullständigt genomförande av de relevanta gemenskapsrättsakterna. Den ekosystemansats som har antagits i konventionen om biologisk mångfald(8) bör alltid tillämpas när så är lämpligt.a) För biologisk mångfald:
- Säkerställa genomförandet och främjandet av övervakning och utvärdering av gemenskapens strategi för biologisk mångfald och därtill hörande handlingsplaner, bl.a. genom ett program för data- och informationsinsamling, framtagande av lämpliga indikatorer, och främjande av användningen av bästa tillgängliga teknik och bästa miljöpraxis.
- Främja forskning om biologisk mångfald, genetiska resurser, ekosystem och samspelet med mänsklig verksamhet.
- Utveckla åtgärder för att öka hållbart nyttjande, hållbar produktion och hållbara investeringar när det gäller biologisk mångfald.
- Främja en sammanhängande bedömning, ytterligare forskning och samarbete om hotade arter.
- På global nivå främja en rimlig och rättvis fördelning av vinster av nyttjandet av genetiska resurser för att genomföra artikel 15 i konventionen om biologisk mångfald och om tillgång till genetiska resurser med ursprung i tredje land.
- Utveckla åtgärder för att förhindra och kontrollera invaderande främmande arter, inklusive främmande genotyper.
- Upprätta Natura 2000-nätverket och genomföra nödvändiga tekniska och finansiella instrument och åtgärder för dess genomförande fullt ut och för skyddet utanför områdena för Natura 2000 av arter som skyddas enligt livsmiljö- och fågeldirektiven.
- Främja utvidgningen av Natura 2000-nätverket till att omfatta kandidatländerna.
b) För olyckor och katastrofer:
- Främja samordning inom gemenskapen av medlemsstaternas insatser i samband med olyckor och naturkatastrofer, genom att till exempel inrätta ett nätverk för utbyte av rutiner och verktyg för förebyggande åtgärder.
- Utveckla ytterligare åtgärder för att bidra till att förebygga risker för storolyckor, i synnerhet de som uppkommer på grund av rörledningar, gruvdrift och sjötransporter av farliga ämnen, samt utveckla åtgärder avseende avfall från gruvdrift.
c) En temainriktad strategi för markskydd genom att vidta förebyggande åtgärder mot bl.a. föroreningar, erosion, ökenspridning, markförstöring, markförbrukning och hydrogeologiska risker med beaktande av regional mångfald, inklusive bergsområdenas och de ofruktbara områdenas specifika karaktär.
d) Främja hållbar förvaltning av utvinningsindustrierna i syfte att minska deras miljöpåverkan.
e) Främja att bevarande och återställande av natursköna områden införlivas i övrig politik, till exempel turism, med beaktande av relevanta internationella instrument.
f) Främja integreringen av hänsynen till biologisk mångfald i jordbrukspolitiken och uppmuntra en hållbar utveckling av landsbygden, ett multifunktionellt och hållbart jordbruk genom följande åtgärder:
- Främja ett fullständigt utnyttjande av nuvarande möjligheter i den gemensamma jordbrukspolitiken och andra politiska åtgärder.
- Främja ett mer miljöansvarigt jordbruk, inbegripet när så är lämpligt extensiva produktionsmetoder, integrerade jordbruksmetoder, ekologiskt jordbruk och biologisk mångfald inom jordbruket, i kommande översyner av den gemensamma jordbrukspolitiken, med hänsyn till behovet av ett väl avvägt förhållningssätt till landsbygdssamhällenas multifunktionella roll.
g) Främja ett hållbart nyttjande av haven och bevarande av marina ekosystem, inklusive havsbottnar, områden kring flodmynningar och kustområden, med särskild hänsyn till platser med betydande biologisk mångfald, genom följande åtgärder:
- Främja en ökad integration av miljöhänsyn i den gemensamma fiskeripolitiken, varvid översynen av denna år 2002 skall utnyttjas.
- Utarbeta en temainriktad strategi för skydd och bevarande av havsmiljöer med beaktande av bland annat villkoren och genomförandeskyldigheterna i havskonventionerna samt behovet av att minska sjötransporters och andra havs- och landbaserade verksamheters utsläpp och miljöpåverkan.
- Främja en integrerad förvaltning av kustområden.
- Främja skyddet av havsområden ytterligare, framför allt genom Natura 2000-nätverket och genom andra genomförbara gemenskapsmedel.
h) I fråga om skogar genomföra och ytterligare utveckla strategier och åtgärder som är i linje med Europeiska unionens skogsstrategi, med beaktande av subsidiaritetsprincipen och hänsynen till biologisk mångfald, och där följande skall finnas med:
- Förbättra pågående gemenskapsåtgärder för skydd av skogar och genomföra en hållbar skogsförvaltning bland annat genom nationella skogsbruksprogram, i samband med planerna för landsbygdsutveckling, med ökad betoning på övervakning av skogens olika funktioner, i enlighet med rekommendationer som antagits av ministerkonferensen om skydd av skogarna i Europa samt FN:s skogsforum och konventionen om biologisk mångfald samt andra forum.
- Stödja effektiv samordning mellan alla politiska sektorer som berörs av skogsbruket, även den privata sektorn, samt samordning av alla intressenter som berörs av skogsbruksfrågor.
- Stimulera till större marknadsandelar för hållbart framställt trä, bland annat genom att uppmuntra certifiering av hållbar skogsförvaltning och uppmuntra märkning av berörda produkter.
- Fortsätta gemenskapens och medlemsstaternas aktiva medverkan i genomförandet av globala och regionala resolutioner och i diskussionerna och förhandlingarna om frågor som rör skogen.
- Undersöka möjligheterna att vidta aktiva åtgärder för att förhindra och bekämpa handeln med olagligt avverkad skog.
- Uppmuntra till diskussion om klimatförändringars verkningar på skogsbruket.
i) För genetiskt modifierade organismer:
- Utarbeta bestämmelser och metoder för riskbedömning, identifiering och märkning av genetiskt modifierade organismer och deras spårbarhet för att möjliggöra effektiv övervakning och kontroller av hälso- och miljöeffekter.
- Sträva efter att snarast ratificera och genomföra Cartagena-protokollet om biosäkerhet och stödja upprättandet av regelsystem i tredje land vid behov genom tekniskt och finansiellt bistånd.
Artikel 7
Mål och prioriterade områden för insatser avseende miljö, hälsa och livskvalitet
1. De syften som anges i artikel 2 bör tillgodoses genom att följande mål uppnås, med hänsyn till relevanta standarder, riktlinjer och program från Världshälsoorganisationen (WHO):
- Uppnå bättre kunskap om hoten mot miljön och människors hälsa i syfte att vidta åtgärder för att förebygga och minska hoten.
- Bidra till bättre livskvalitet genom ett integrerat förhållningssätt med fokus på stadsområden.
- Sträva efter att inom en generation (2020) åstadkomma att kemikalier produceras och används endast på sätt som inte har en betydande negativ inverkan på hälsan och miljön samt inse att den nuvarande bristen på kunskaper om egenskaper, användning, bortskaffande och exponering när det gäller kemikalier måste avhjälpas.
- Kemikalier som är farliga bör ersättas med säkrare kemikalier eller säkrare alternativa tekniker som inte innebär användning av kemikalier, så att riskerna för människan och miljön minskas.
- Minska påverkan av bekämpningsmedel för människors hälsa och miljön och, mer allmänt, åstadkomma en mer hållbar användning av bekämpningsmedel samt en betydande total minskning av riskerna och av användningen av bekämpningsmedel som är förenlig med ett tillräckligt skydd av grödor. De bekämpningsmedel som är beständiga eller anrikas i miljön eller är toxiska eller har andra negativa egenskaper bör ersättas med mindre farliga medel om det är möjligt.
- Uppnå en sådan kvalitet på grund- och ytvatten som inte leder till betydande konsekvenser och risker för människors hälsa eller miljön, och att se till att uttagen från vattenresurserna är hållbara på lång sikt.
- Uppnå en sådan luftkvalitet som inte leder till betydande negativa konsekvenser och risker för människors hälsa eller miljön.
- Avsevärt minska antalet personer som regelbundet utsätts för långsiktiga genomsnittliga bullernivåer, särskilt från trafiken, som enligt vetenskapliga undersökningar har skadliga effekter på människors hälsa och förbereda nästa steg i arbetet med bullerdirektivet.
2. Dessa mål skall uppnås med hjälp av följande prioriterade åtgärder:
a) Förstärkning av gemenskapens forskningsprogram och vetenskapliga expertis samt uppmuntran till internationell samordning av de nationella forskningsprogrammen i syfte att främja uppnåendet av fastställda mål inom området hälsa och miljö, och i synnerhet
- fastställa och rekommendera prioriterade områden för forskning och åtgärder, bland annat potentiella konsekvenser för hälsan från elektromagnetiska föroreningskällor och med särskild hänsyn till utvecklandet och valideringen av alternativa djurtestmetoder, i synnerhet på området för kemisk säkerhet,
- fastställa och utveckla hälso- och miljöindikatorer,
- undersöka på nytt, utveckla och uppdatera befintliga hälsostandarder och gränsvärden, och vid behov effekter på särskilt sårbara grupper, t.ex. barn och äldre, och olika förorenande ämnens synergier och deras ömsesidiga konsekvenser,
- granska utvecklingstendenser och tillhandahålla ett system för tidig varning vid nya eller framväxande problem.
b) För kemikalier:
- Lägga ansvaret på tillverkare, importörer och användare i efterföljande led för att utveckla kunskap om samtliga kemikalier (skyldighet att iaktta försiktighet) och bedöma riskerna med deras användning, också i produkter, samt materialåtervinning och bortskaffande.
- Utarbeta ett enhetligt system som grundar sig på ett angreppssätt som införs steg för steg, utom för kemiska ämnen som används i mycket små mängder, för testning, riskbedömning och riskhantering för nya och befintliga ämnen med testförfaranden som minimerar behovet av djurförsök samt utarbeta alternativa testmetoder.
- Se till att potentiellt skadliga kemiska ämnen omfattas av utökade riskhanteringsförfaranden och att potentiellt mycket skadliga kemiska ämnen, inbegripet cancerframkallande, arvsmassepåverkande och fortplantningsstörande ämnen när det gäller reproduktionsämnen och de som har POP-egenskaper (beständiga organiska föreningar), bara används i motiverade och klart definierade fall och att det krävs tillståndsgivning innan de får användas.
- Se till att resultaten av riskbedömningen av kemikalier till fullo beaktas i all gemenskapslagstiftning där kemikalier regleras och att undvika dubbelarbete.
- Tillhandahålla kriterier för att bland ämnen av mycket stor betydelse ta med sådana ämnen som är beständiga och bioackumulerande och toxiska, samt ämnen som är mycket beständiga och mycket bioackumulerande och överväga att ta med kända ämnen som kan orsaka en endokrin rubbning när överenskomna testmetoder och testkriterier fastställs.
- Se till att de viktigaste åtgärder som är nödvändiga med tanke på de fastställda målen utvecklas snabbt, så att de kan träda i kraft före halvtidsöversynen.
- Säkerställa allmänhetens tillgång till den icke-sekretessbelagda informationen i gemenskapens register över kemikalier (Reach-registret).
c) För bekämpningsmedel:
- Fullt genomförande och fullständig översyn av effektiviteten av den tillämpliga rättsliga ramen(9) för att säkerställa en hög skyddsnivå när den ändras. Denna översyn kan när så är lämpligt inbegripa en jämförande bedömning och utarbetande av tillståndsgivningsförfaranden på gemenskapsnivå för utsläppande på marknaden.
- En temainriktad strategi för hållbar användning av bekämpningsmedel som omfattar
i) en minimering av de risker för hälsa och miljö som användningen av bekämpningsmedel medför,
ii) förbättrade kontroller av användningen och spridningen av bekämpningsmedel,
iii) en minskning av halterna av skadliga aktiva ämnen också genom att ersätta de farligaste med säkrare, även kemikaliefria, alternativ,
iv) stöd till odling där mycket lite eller inget bekämpningsmedel behöver användas, bland annat genom att öka användarnas medvetenhet och främja användning av regler för god praxis och stödja diskussioner om eventuell tillämpning av finansiella styrmedel,
v) ett öppet system för att redogöra för och övervaka de framsteg som görs med att uppnå strategins mål, inklusive utarbetande av lämpliga indikatorer.
d) För kemikalier och bekämpningsmedel:
- Syfta till en snabb ratificering av Rotterdamkonventionen om förfarandet för ett förhandsgodkännande av vissa farliga kemikalier och bekämpningsmedel i internationell handel och Stockholmskonventionen om beständiga organiska föreningar (POP).
- Ändra rådets förordning (EEG) nr 2455/92 av den 23 juli 1992 om export och import av vissa farliga kemikalier(10) i syfte att anpassa denna till Rotterdamkonventionen, förbättra dess förfarandemekanismer och ge bättre information till utvecklingsländerna.
- Stödja förbättringen av hanteringen av kemikalier och bekämpningsmedel i utvecklings- och kandidatländerna, inklusive eliminering av lager av bekämpningsmedel som tagits ur bruk, bland annat genom att stödja projekt som syftar till sådan eliminering.
- Bidra till de internationella satsningarna på att utarbeta en strategi för internationell kemikaliehantering.
e) För hållbar vattenanvändning och hög vattenkvalitet:
- Säkerställa en hög skyddsnivå för ytvatten och grundvatten, förhindra förorening och främja hållbar vattenanvändning.
- Arbeta för fullständigt genomförande av ramdirektivet om vatten(11), vilket syftar till god ekologisk, kemisk och kvantitativ vattenstatus samt en sammanhängande och hållbar vattenförvaltning.
- Utveckla åtgärder för att eliminera utsläpp och spill av prioriterade farliga ämnen i linje med bestämmelserna i ramdirektivet om vatten.
- Säkerställa en hög skyddsnivå för badvatten, inklusive en översyn av badvattendirektivet(12).
- Säkerställa integrering av de koncept och tillvägagångssätt som fastställs i ramdirektivet för vatten och andra direktiv om vattenskydd i annan gemenskapspolitik.
f) För luftkvalitet: utvecklingen och genomförandet av åtgärderna i artikel 5 inom transport-, industri- och energisektorerna bör vara förenliga med och bidra till bättre luftkvalitet. Följande ytterligare åtgärder planeras:
- Förbättra övervakningen och bedömningen av luftkvaliteten och nedfallet av föroreningar och tillhandahålla information till allmänheten, bland annat genom att utarbeta och använda indikatorer.
- Utarbeta en temainriktad strategi för att stärka en konsekvent och integrerad politik när det gäller luftförorening, vilken omfattar prioriteringar för framtida åtgärder, översyn och uppdatering om så behövs av luftkvalitetsnormer och nationella utsläppstak i syfte att uppnå det långsiktiga målet att inte överskrida kritiska belastningsgränser och belastningsnivåer samt utveckla bättre system för insamling av information, modellering och prognosticering.
- Anta lämpliga åtgärder beträffande ozon och partiklar på marknivå.
- Undersöka inomhusluftens kvalitet och dess inverkan på människors hälsa, med rekommendationer för framtida åtgärder där så behövs.
- Spela en ledande roll i förhandlingarna och genomförandet av Montreal-protokollet om ämnen som bryter ned ozonskiktet.
- Spela en ledande roll vid förhandlingar om och stärkande av kopplingar och samverkan med sådana internationella processer som medverkar till ren luft i Europa.
- Vidareutveckla specifika gemenskapsinstrument för att minska utsläppen från relevanta kategorier av utsläppskällor.
g) För buller:
- Komplettera och ytterligare förbättra åtgärderna, till exempel lämpliga förfaranden för typgodkännande, mot bullerutsläpp från tjänster och produkter, särskilt motorfordon, inklusive åtgärder för att minska buller på grund av samspelet mellan däck och vägbana, vilka inte äventyrar trafiksäkerheten, samt från järnvägsvagnar, flygplan och stationära maskiner.
- Utveckla och införa instrument för att vid behov minska trafikbuller, exempelvis genom minskad efterfrågan på transporter, övergång till mindre bullersamma transportmedel, främjande av tekniska åtgärder och en hållbar transportplanering.
h) För stadsmiljö:
- Utarbeta en temainriktad strategi för att främja en integrerad horisontell lösning för gemenskapens alla politikområden och förbättra kvaliteten på stadsmiljön, med hänsyn till framstegen med genomförandet av den befintliga ramen för samarbete(13), och om så är nödvändigt se över denna strategi vilken omfattar
- främjande av lokal Agenda 21,
- minskning av sambandet mellan ekonomisk tillväxt och efterfrågan på passagerartransport,
- behovet att öka andelen kollektiv- och järnvägstrafik, trafik på inre vattenvägar, gång- och cykeltrafik,
- behovet att ta itu med de ökande trafikmängderna och att ta bort kopplingen mellan ökade transporter och BNP-tillväxt,
- behovet att främja användningen av miljövänliga fordon i kollektivtrafiken,
- övervägande av miljöindikatorer när det gäller städer.
Artikel 8
Mål och prioriterade områden för insatser avseende hållbar användning och förvaltning av naturresurser samt avfall
1. De syften som anges i artikel 2 bör tillgodoses genom att följande mål uppnås:
- Strävan efter att säkerställa att förbrukningen av resurser och dess följdeffekter inte överskrider vad miljön kan bära och att bryta sambandet mellan ekonomisk tillväxt och resursanvändning. I detta sammanhang erinras om det vägledande delmålet att i gemenskapen senast 2010 uppnå ett procenttal på 22 % när det gäller elproduktion från förnybara energikällor i syfte att drastiskt öka resurs- och energieffektiviteten.
- Uppnående av en betydande generell minskning av den mängd avfall som genereras genom initiativ för att förebygga avfall, bättre resurseffektivitet samt en övergång till mer hållbara produktions- och konsumtionsmönster.
- En betydande minskning av den mängd avfall som skall bortskaffas och mängden producerat farligt avfall, samtidigt som ökade utsläpp i luften, vattnet och marken undviks.
- Stöd till återanvändning och när det gäller avfall som fortfarande genereras: dess farlighetsgrad bör minskas och det bör medföra så liten risk som möjligt; företräde bör ges åt återvinning, särskilt materialåtervinning; mängden avfall som skall bortskaffas bör minimeras och bortskaffas på ett säkert sätt; avfall som är avsett att bortskaffas bör behandlas så nära uppkomstplatsen som möjligt, i den mån det inte leder till en minskning av effektiviteten i avfallshanteringen.
2. Målen skall nås med beaktande av strategin för en integrerad produktpolicy samt gemenskapsstrategin för avfallshantering(14) genom följande prioriterade åtgärder:
i) Utarbetande av en temainriktad strategi för hållbar användning och förvaltning av resurser, inbegripet bland annat
a) uppskattning av material- och avfallsflödena i gemenskapen, inklusive import och export, till exempel genom materialflödesanalys,
b) översyn av effektiviteten i de politiska åtgärderna och konsekvenserna av subventioner som rör naturresurser och avfall,
c) uppställande av mål för resurseffektivitet och en minskad användning av resurser för att bryta sambandet mellan ekonomisk tillväxt och negativa miljökonsekvenser,
d) främjande av utvinnings- och produktionsmetoder och teknik för att stödja ekoeffektivitet och en hållbar användning av råmaterial, energi, vatten och andra resurser,
e) utarbetande och genomförande av ett brett spektrum av instrument, däribland forskning, tekniköverföring, marknadsbaserade och ekonomiska instrument, program för bästa metoder samt indikatorer för resurseffektivitet.
ii) Utarbetande och genomförande av åtgärder för avfallsförebyggande och avfallshantering, bland annat genom att
a) sätta upp en rad kvantitativa och kvalitativa delmål för minskning som omfattar alla typer av relevant avfall, som skall uppnås på gemenskapsnivå senast 2010; kommissionen uppmanas att utarbeta ett förslag till sådana delmål senast 2002,
b) stödja miljövänlig och hållbar produktdesign,
c) öka medvetenheten om allmänhetens möjligheter att bidra till avfallsminskningen,
d) formulera operativa åtgärder för att stimulera förebyggande av uppkomsten av avfall, t.ex. genom att uppmuntra återanvändning och återvinning samt utfasning av vissa ämnen och material genom produktrelaterade åtgärder,
e) utarbeta ytterligare indikatorer inom avfallshanteringen.
iii) Utarbetande av en temainriktad strategi för avfallsåtervinning, vilken inbegriper bland annat
a) åtgärder för att ombesörja källsortering, insamling och materialåtervinning av prioriterade avfallsflöden,
b) ytterligare utveckling av producentansvar,
c) utarbetande och överföring av miljövänlig avfallsåtervinning och behandlingsteknik.
iv) Utveckling eller översyn av lagstiftningen om avfall, inbegripet bland annat bygg- och rivningsavfall, avloppsslam(15), biologiskt nedbrytbart avfall, förpackningar(16), batterier(17) samt avfallstransporter(18), klargörande av skillnaden mellan avfall och sådant som inte är avfall samt utarbetande av lämpliga kriterier för vidareutveckling av bilagorna IIA och IIB i ramdirektivet om avfall(19).
Artikel 9
Mål och prioriterade områden för åtgärder avseende internationella frågor
1. De syften som anges i artikel 2 avseende internationella frågor och internationella aspekter på de fyra prioriterade miljöområdena i detta program innehåller följande mål:
- Bedrivande av en ambitiös miljöpolitik på internationell nivå med särskild hänsyn till hur mycket den globala miljön kan bära.
- Ytterligare främjande av hållbara förbruknings- och produktionsmönster på internationell nivå.
- Framsteg mot säkerställande av att politik och åtgärder när det gäller handel och miljö ömsesidigt stöder varandra.
2. Dessa mål skall eftersträvas med hjälp av följande prioriterade åtgärder:
a) Integrering av miljöskyddskrav i all politik som rör gemenskapens yttre förbindelser, inklusive handels- och utvecklingssamarbete, för att uppnå en hållbar utveckling, bland annat genom utarbetande av riktlinjer.
b) Fastställande av ett antal samstämmiga miljö- och utvecklingsmål för antagande som en del av %quot%en ny global uppgörelse eller överenskommelse%quot% vid världstoppmötet om hållbar utveckling år 2002.
c) Strävan efter att förstärka den internationella miljöstyrningen genom ett gradvis stärkande av det multilaterala samarbetet och den institutionella ramen samt genom tilldelning av resurser.
d) Strävan efter snabb ratificering, faktisk efterlevnad och verkställighet av internationella konventioner och avtal om miljön där gemenskapen är part.
e) Främjande av hållbar miljöpraxis i samband med utlandsinvesteringar och exportkrediter.
f) Intensifierade ansträngningar på internationell nivå för att uppnå samsyn om metoder för bedömning av hälso- och miljörisker, samt om riskhanteringsförfaranden, inklusive försiktighetsprincipen.
g) Ömsesidigt stöd mellan handeln och miljöskyddsbehoven genom att vederbörlig hänsyn tas till miljödimensionen vid de konsekvensbedömningar av multilaterala handelsavtal ur hållbarhetssynvinkel som skall utföras i ett tidigt förhandlingsskede samt genom att efterleva resultaten av dessa.
h) Fortsatt stöd för ett världshandelssystem som fullt ut erkänner multilaterala eller regionala miljöavtal och försiktighetsprincipen och därigenom öka möjligheterna till handel med miljövänliga produkter och tjänster.
i) Främjande av gränsöverskridande miljösamarbete med grannländer och grannregioner.
j) Främjande av ökad konsekvens i politiken genom att det arbete som utförts inom ramen för de olika konventioner, inklusive en bedömning av sambanden mellan biologisk mångfald och klimatförändringar, kopplas till integreringen av hänsyn till den biologiska mångfalden i genomförandet av Förenta nationernas ramkonvention om klimatförändringar och av Kyotoprotokollet.
Artikel 10
Utformning av miljöpolitiken
De mål som fastställs i artikel 2 avseende utformning av miljöpolitiken, som grundar sig på delaktighet och på det främsta vetenskapliga kunnande som finns att tillgå och de strategiska metoder som anges i artikel 3, skall tillgodoses bland annat med hjälp av följande prioriterade åtgärder:
a) Utveckling av förbättrade mekanismer, allmänna regler och principer för god förvaltning som innebär ett omfattande och ingående samråd med berörda parter i alla skeden för att underlätta valet av de mest effektiva lösningarna och för att uppnå de bästa resultaten för miljön och en hållbar utveckling med avseende på kommande förslag till åtgärder.
b) Ökad medverkan av de icke-statliga miljöorganisationerna i dialogen, genom lämpligt stöd och gemenskapsfinansiering.
c) Bättre utformning av politiken genom
- utvärdering på förhand av de tänkbara konsekvenserna, i synnerhet miljökonsekvenserna, av en ny politik, inbegripet alternativet att inte vidta några åtgärder och av lagstiftningsförslagen samt offentliggörande av resultaten,
- utvärdering i efterhand av de befintliga åtgärdernas effektivitet när det gäller att nå miljömålen.
d) Se till att miljön och i synnerhet de prioriterade områden som identifieras i detta program utgör huvudprioriteringar i gemenskapens forskningsprogram. Regelbunden översyn av miljöforskningsbehov och prioriteringar bör göras inom gemenskapens ramprogram för forskning och teknisk utveckling. Säkerställa en bättre samordning av den miljörelaterade forskningen i medlemsstaterna, bl.a. för att förbättra tillämpningen av forskningsresultaten.
Bygga broar mellan miljöaktörer och andra aktörer inom områdena information, yrkesutbildning, forskning, utbildning och politik.
e) Se till att det från och med 2003 regelbundet tillhandahålls information som kan utgöra en grund för
- politiska beslut om miljö och hållbar utveckling,
- uppföljningen och översynen av sektoriella integreringsstrategier samt av strategin för en hållbar utveckling,
- information till den breda allmänheten.
Framställandet av denna information kommer att underlättas genom Europeiska miljöbyråns och andra relevanta organs regelbundna rapporter. Informationen skall främst utgöras av
- övergripande miljöindikatorer,
- indikatorer för miljöns aktuella tillstånd och utveckling,
- integreringsindikatorer.
f) Ompröva och regelbundet övervaka informations- och rapporteringssystemen för att få ett mer samstämmigt och effektivt system för att garantera enhetlig rapportering av högkvalitativ, jämförbar och relevant miljöinformation. Kommissionen uppmanas att så snart som möjligt vid behov lägga fram ett förslag i detta syfte. Kraven på övervakning, insamling av data och rapportering bör beaktas på ett effektivt sätt i framtida miljölagstiftning.
g) Förstärka utveckling och användning av system och verktyg för övervakning av jorden (t.ex. satellitteknik), som stöd för utformningen och genomförandet av politiken.
Artikel 11
Övervakning och utvärdering av resultaten
1. Under loppet av programmets fjärde år skall kommissionen utvärdera gjorda framsteg i programmets genomförande samt härmed förbundna tendenser och framtidsutsikter på miljöområdet. Detta bör göras på grundval av en övergripande uppsättning indikatorer. Kommissionen skall lägga fram denna rapport för Europaparlamentet och rådet efter halva tiden tillsammans med eventuella förslag till ändringar, som den anser lämpliga.
2. Kommissionen skall under loppet av programmets sista år till Europaparlamentet och rådet framlägga en slutbedömning av programmet och av tillståndet hos och utsikterna för miljön.
Artikel 12
Detta beslut skall offentliggöras i Europeiska gemenskapernas officiella tidning.
Europaparlamentets och rådets direktiv 2002/74/EG
av den 23 september 2002
om ändring av rådets direktiv 80/987/EEG om tillnärmning av medlemsstaternas lagstiftning om skydd för arbetstagarna vid arbetsgivarens insolvens
(Text av betydelse för EES)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 137.2 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Ekonomiska och sociala kommitténs yttrande(2),
efter att ha hört Regionkommittén,
i enlighet med förfarandet i artikel 251 i fördraget(3), och
av följande skäl:
(1) I punkt 7 i gemenskapens stadga om grundläggande sociala rättigheter för arbetstagare, som antogs den 9 december 1989, föreskrivs att förverkligandet av den inre marknaden måste leda till att levnad- och arbetsvillkoren för arbetstagare inom Europeiska gemenskapen förbättras samt att förbättringen, där så behövs, även måste medföra att vissa aspekter av anställningsreglerna utvecklas, såsom förfaranden vid kollektiva uppsägningar och konkurser.
(2) Direktiv 80/987/EEG(4) syftar till att garantera arbetstagarna ett minimiskydd vid arbetsgivarens insolvens. För detta ändamål är alla medlemsstater skyldiga att inrätta en institution som säkerställer att de berörda arbetstagarna får betalt för sina utestående fordringar.
(3) Rättsutvecklingen i medlemsstaterna avseende insolvens samt utvecklingen av den inre marknaden kräver en anpassning av vissa bestämmelser i ovannämnda direktiv.
(4) Av rättssäkerhetsskäl och för ökad insyn krävs dessutom preciseringar när det gäller tillämpningsområdet för och vissa definitioner i direktiv 80/987/EEG. Det är bl.a. lämpligt att i artikeldelen i direktivet precisera de möjligheter medlemsstaterna har att utesluta vissa kategorier, och som en följd därav upphäva bilagan till direktivet.
(5) För att säkerställa ett rättvist skydd för de berörda arbetstagarna bör man anpassa definitionen av insolvens till den nya utvecklingen av lagstiftningen i medlemsstaterna på detta område och genom detta begrepp även avse andra insolvensförfaranden än likvidationsförfaranden. I syfte att fastställa garantiinstitutionens betalningsskyldighet bör medlemsstaterna i detta sammanhang ha möjlighet att föreskriva att en insolvenssituation som leder till flera insolvensförfaranden skall hanteras som om det gällde ett enda insolvensförfarande.
(6) Det bör säkerställas att de arbetstagare som avses i rådets direktiv 97/81/EG av den 15 december 1997 om ramavtalet om deltidsarbete undertecknat av UNICE, CEEP och EFS(5), rådets direktiv 1999/70/EG av den 28 juni 1999 om ramavtalet om visstidsarbete undertecknat av EFS, UNICE och CEEP(6) och rådets direktiv 91/383/EEG av den 25 juni 1991 om komplettering av åtgärderna för att främja förbättringar av säkerhet och hälsa på arbetsplatsen för arbetstagare med tidsbegränsat anställningsförhållande eller tillfälligt anställningsförhållande(7) inte utesluts från tillämpningsområdet för detta direktiv.
(7) För att tillgodose arbetstagarnas rättssäkerhet när företag som bedriver verksamhet i flera medlemsstater blir insolventa och för att trygga arbetstagarnas rättigheter i enlighet med domstolens rättspraxis, är det nödvändigt att införa bestämmelser som uttryckligen fastställer vilken institution som är behörig att betala de utestående fordringarna till arbetstagarna i dessa fall och som fastställer målet för samarbetet mellan medlemsstaternas behöriga myndigheter att snarast möjligt reglera arbetstagarnas utestående fordringar. Det är vidare nödvändigt att föreskriva ett samarbete mellan behöriga administrativa myndigheter i medlemsstaterna för att se till att bestämmelserna på detta område tillämpas på rätt sätt.
(8) Medlemsstaterna kan införa begränsningar av garantiinstitutionernas ansvar. Begränsningarna bör vara förenliga med direktivets sociala mål, och vid införandet av dessa kan olika nivåer på fordringarna beaktas.
(9) För att underlätta fastställandet av insolvensförfaranden bl.a. i gränsöverskridande situationer bör det föreskrivas att medlemsstaterna skall informera kommissionen och övriga medlemsstater om de typer av insolvensförfaranden som ger anledning till åtgärd från garantiinstitutionen.
(10) Direktiv 80/987/EEG bör därför ändras i enlighet med detta.
(11) Eftersom målet för den föreslagna åtgärden, nämligen att ändra vissa bestämmelser i direktiv 80/987/EEG med anledning av att de verksamheter som bedrivs av företagen inom gemenskapen har förändrats, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna och de därför bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget. I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå detta mål.
(12) Kommissionen bör för Europaparlamentet och rådet lägga fram en rapport om genomförandet och tillämpningen av detta direktiv, särskilt med avseende på de nya anställningsformer som uppkommer i medlemsstaterna.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 80/987/EEG ändras på följande sätt:
1. Titeln skall ersättas med följande text: %quot%Rådets direktiv 80/987/EEG av den 20 oktober 1980 om skydd för arbetstagare vid arbetsgivarens insolvens.%quot%.
2. Avsnitt I skall ersättas med följande text: %quot%AVSNITT I
Tillämpningsområde och definitioner
Artikel 1
1. Detta direktiv skall tillämpas på fordringar som arbetstagare på grund av anställningsavtal eller anställningsförhållanden har gentemot arbetsgivare som är att anse som insolventa enligt artikel 2.1.
2. Medlemsstaterna får undantagsvis utesluta fordringar från vissa kategorier av arbetstagare från tillämpningsområdet för detta direktiv om det finns andra former av garanti som ger arbetstagarna ett skydd motsvarande det som följer av detta direktiv.
3. Medlemsstaterna får, om en sådan bestämmelse redan finns i deras nationella lagstiftning, fortsätta att utesluta följande kategorier från tillämpningsområdet för detta direktiv:
a) Arbetstagare i hushållet som är anställda av en fysisk person.
b) Fiskare som avlönas separat.
Artikel 2
1. I detta direktiv skall en arbetsgivare anses vara insolvent när en ansökan har inlämnats om att inleda ett kollektivt förfarande som grundas på arbetsgivarens insolvens i enlighet med respektive medlemsstats lagar och andra författningar och som innebär att arbetsgivarens tillgångar helt eller delvis tas i anspråk och att en förvaltare eller en person som utövar en liknande funktion utses, samt när den myndighet som är behörig enligt dessa lagar och andra författningar
a) har beslutat att inleda ett förfarande, eller
b) har fastställt att arbetsgivarens företag eller verksamheter definitivt har upphört och att befintliga tillgångar är otillräckliga för att motivera att förfarandet inleds.
2. Detta direktiv påverkar inte den definition som följer av nationell rätt beträffande termerna arbetstagare, arbetsgivare, lön, omedelbar rätt till och framtida rätt till.
Medlemsstaterna får från tillämpningsområdet för detta direktiv emellertid inte utesluta
a) deltidsanställda i den mening som avses i direktiv 97/81/EG,
b) visstidsanställda i den mening som avses i direktiv 1999/70/EG,
c) arbetstagare med ett tillfälligt anställningsförhållande i den mening som avses i artikel 1.2 i direktiv 91/383/EEG.
3. Medlemsstaterna får inte göra arbetstagarnas rätt enligt detta direktiv beroende av en minsta kvalifikationsperiod avseende anställningsavtal eller anställningsförhållande.
4. Detta direktiv hindrar inte medlemsstaterna från att utsträcka skyddet för arbetstagare till andra insolvenssituationer som fastställts genom andra förfaranden än de som nämns i punkt 1 och som föreskrivs i nationell lagstiftning, till exempel situationer där arbetsgivaren i praktiken inställt betalningarna permanent.
Sådana förfaranden skall dock inte leda till ett krav på garantier för institutionerna i de övriga medlemsstaterna i sådana fall som avses i avsnitt IIIa.%quot%
3. Artiklarna 3 och 4 skall ersättas med följande text: %quot%Artikel 3
Medlemsstaterna skall, om inte annat följer av artikel 4, vidta nödvändiga åtgärder för att tillförsäkra att garantiinstitutionerna säkerställer betalning av arbetstagarnas utestående fordringar som grundar sig på anställningsavtal eller anställningsförhållanden, inbegripet betalning av avgångsvederlag, förutsatt att nationell lagstiftning föreskriver det, när anställningsförhållandet upphör.
De utestående lönefordringar som garantiinstitutionen övertar avser en period före och/eller, i förekommande fall, efter ett datum som fastställts av medlemsstaterna.
Artikel 4
1. Medlemsstaterna får välja att begränsa garantiinstitutionernas betalningsansvar enligt artikel 3.
2. Om medlemsstaterna utnyttjar valmöjligheten enligt punkt 1, skall de fastställa den period för vilken garantiinstitutionen skall betala utestående fordringar. Denna period får dock inte vara kortare än en period som omfattar lönen för de tre senaste månaderna av anställningsförhållandet före och/eller efter det datum som avses i artikel 3. Medlemsstaterna får bestämma att denna minimiperiod på tre månader skall infalla under en referensperiod som inte får vara kortare än sex månader.
De medlemsstater som föreskriver en referensperiod på minst arton månader får begränsa den period för vilken garantiinstitutionen skall betala de utestående fordringarna till åtta veckor. I sådana fall skall de för arbetstagarna mest fördelaktiga perioderna användas vid beräkningen av minimiperioden.
3. Medlemsstaterna får dessutom fritt sätta övre gränser för garantiinstitutionens utbetalningar. Dessa gränser får inte vara lägre än en tröskel som är socialt förenlig med detta direktivs sociala målsättning.
Om medlemsstaterna utnyttjar denna valmöjlighet, skall de till kommissionen meddela vilka metoder de använder för att sätta denna övre gräns.%quot%
4. Följande avsnitt skall läggas till: %quot%AVSNITT IIIa
Bestämmelser om gränsöverskridande situationer
Artikel 8a
1. När ett företag som är verksamt på minst två medlemsstaters territorium är insolvent i den mening som avses i artikel 2.1, skall institutionen i den medlemsstat på vilkens territorium arbetstagarna normalt utför eller utförde sitt arbete vara behörig institution för betalningen av utestående fordringar till arbetstagarna.
2. Omfattningen av arbetstagarnas rättigheter skall fastställas i den lagstiftning som gäller för den behöriga garantiinstitutionen.
3. Medlemsstaterna skall vidta nödvändiga åtgärder för att säkerställa att, i de fall som avses i punkt 1, de beslut som fattas inom ramen för ett insolvensförfarande enligt artikel 2.1 som inletts i en annan medlemsstat beaktas för att fastställa arbetsgivarens insolvens i den mening som avses i detta direktiv.
Artikel 8b
1. För att genomföra artikel 8a skall medlemsstaterna föreskriva om utbyte av relevant information mellan de behöriga administrativa myndigheterna och/eller mellan de garantiinstitutioner som omnämns i artikel 3, vilket bland annat gör det möjligt att upplysa den behöriga garantiinstitutionen om arbetstagarnas utestående fordringar.
2. Medlemsstaterna skall till kommissionen och de andra medlemsstaterna lämna uppgifter om adress och telefon till sina behöriga administrativa myndigheter och/eller sina garantiinstitutioner. Kommissionen skall göra dessa upplysningar tillgängliga för allmänheten.%quot%
5. I artikel 9 skall följande stycke läggas till: %quot%Genomförandet av detta direktiv får under inga omständigheter utgöra skäl för att försämra den existerande situationen i medlemsstaterna och den allmänna skyddsnivån för arbetstagare inom det område som direktivet omfattar.%quot%
6. I artikel 10 skall följande punkt läggas till: %quot%c) vägra att ta på sig eller begränsa den betalningsskyldighet som avses i artikel 3 eller den garanterade förpliktelse som avses i artikel 7 i de fall då arbetstagaren ensam eller tillsammans med nära anförvanter var ägare till en väsentlig del av arbetsgivarens företag eller verksamhet och hade ett betydande inflytande över verksamheten.%quot%
7. Följande artikel skall läggas till: %quot%Artikel 10a
Medlemsstaterna skall till kommissionen och de övriga medlemsstaterna anmäla de typer av nationella insolvensförfaranden som omfattas av direktivets tillämpningsområde samt alla ändringar av dessa. Kommissionen skall offentliggöra dessa anmälningar i Europeiska gemenskapernas officiella tidning.%quot%
8. Bilagan skall utgå.
Artikel 2
1. Medlemsstaterna skall sätta i kraft de lagar och andra författningar som är nödvändiga för att följa detta direktiv före den 8 oktober 2005. De skall genast underrätta kommissionen om detta.
Medlemsstaterna skall tillämpa de bestämmelser som avses i första stycket på alla former av insolvens som drabbar en arbetsgivare efter den dag då dessa bestämmelser har trätt i kraft.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texten till de bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 3
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska gemenskapernas officiella tidning.
Artikel 4
Senast den 8 oktober 2010 skall kommissionen för Europaparlamentet och rådet lägga fram en rapport om genomförandet och tillämpningen av detta direktiv i medlemsstaterna.
Artikel 5
Detta direktiv riktar sig till medlemsstaterna.
Kommissionens förordning (EG) nr 141/2002
av den 25 januari 2002
om klassificering av vissa varor i Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan(1), senast ändrad genom förordning (EG) nr 2433/2001(2), särskilt artikel 9 i denna, och
av följande skäl:
(1) För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till ovannämnda förordning, är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till denna förordning.
(2) I förordning (EEG) nr 2658/87 har allmänna regler fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
(3) Enligt dessa allmänna regler måste de varor som beskrivs i kolumn 1 i tabellen som är bifogad den här förordningen klassificeras enligt motsvarande KN-nummer i kolumn 2 med de motiveringar som ges i kolumn 3.
(4) Det är lämpligt att bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter avseende varuklassificeringen i Kombinerade nomenklaturen och som inte överensstämmer med de rättigheter som fastställs i denna förordning fortfarande kan åberopas av innehavaren enligt bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(3) senast ändrad genom Europaparlamentets och rådets förordning (EG) nr 2700/2000(4), under en period av tre månader.
(5) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Tullkodexkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 2
Bindande tulltaxeupplysningar som meddelas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
Artikel 3
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 486/2002
av den 18 mars 2002
om ändring av förordning (EG) nr 2848/98 för tobakssektorn när det gäller fastställande av vissa tidsgränser
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2075/92 av den 30 juni 1992 om den gemensamma organisationen av marknaden för råtobak(1), senast ändrad genom förordning (EG) nr 1336/2000(2), särskilt artikel 11 i denna, och
av följande skäl:
(1) Eftersom det inte finns något rådsbeslut om kommissionens förslag(3) som avser att fastställa garantitrösklar för skördeåren 2002, 2003 och 2004 är det inte möjligt för medlemsstaterna att för 2002 års skörd iaktta tidsgränserna för att till producenterna utfärda kvotintyg och för att sluta odlingskontrakt enligt kommissionens förordning (EG) nr 2848/98 av den 22 december 1998 om tillämpningsföreskrifter till rådets förordning (EEG) nr 2075/92 när det gäller stödordningen, produktionskvoterna och det särskilda stöd som skall beviljas till producentsammanslutningar inom sektorn för råtobak(4), senast ändrad genom förordning (EG) nr 1441/2001(5). Dessa tidsgränser bör därför senareläggas.
(2) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för tobak.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 55 i förordning (EG) nr 2848/98 skall ersättas med följande: %quot%Artikel 55
1. För 2002 års skörd skall medlemsstaterna, genom undantag från artikel 22.3, till enskilda producenter som inte är medlemmar i någon organisation och till producentorganisationerna utfärda kvotintygen senast den 30 april 2002.
2. För 2002 års skörd skall odlingskontrakten, genom undantag från artikel 10.1, utom vid force majeure, slutas senast den 30 juni 2002.%quot%
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1889/2002
av den 23 oktober 2002
om genomförande av rådets förordning (EG) nr 448/98 om komplettering och ändring av rådets förordning (EG) nr 2223/96 om fördelning av indirekt mätta finansiella förmedlingstjänster (FISIM) inom ramen för det europeiska national- och regionalräkenskapssystemet (ENS)
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 448/98 av den 16 februari 1998 om komplettering och ändring av rådets förordning (EG) nr 2223/96 om fördelning av indirekt mätta finansiella förmedlingstjänster (FISIM) inom ramen för det europeiska national- och regionalräkenskapssystemet (ENS)(1), särskilt artikel 5.3 i denna, och
av följande skäl:
(1) Rådets förordning (EG) nr 2223/96 av den 25 juni 1996 om det europeiska national- och regionalräkenskapssystemet i gemenskapen(2), senast ändrad genom Europaparlamentets och rådets förordning (EG) nr 359/2002(3) (nedan kallat ENS 95) innehåller referensramen för de gemensamma standarder, definitioner, klassificeringar och räkenskapsregler som är avsedda att användas vid utarbetandet av medlemsstaternas räkenskaper för gemenskapens statistikbehov, för att sinsemellan jämförbara resultat skall erhållas från medlemsstaterna.
(2) Genom bilaga I till förordning (EG) nr 448/98 ändras bilaga A till förordning (EG) nr 2223/96 med syftet att i ENS 95-metodiken införa principen om fördelning av FISIM och fastställa försöksmetoder för fördelningen av FISIM vilka medlemsstaterna skulle testa för åren 1995 till 2001. Försöksperioden var tillräckligt lång för att göra det möjligt att pröva om denna fördelning ger mer tillförlitliga resultat för en korrekt mätning av ifrågavarande ekonomiska verksamhet än den nuvarande nollfördelningen.
(3) I enlighet med artikel 5.1 i förordning (EG) nr 448/98 lade kommissionen den 21 juni 2002 fram en slutrapport för Europaparlamentet och rådet med en kvalitativ och kvantitativ analys av konsekvenserna av försöksmetoderna för fördelning och beräkning av FISIM. Enligt slutsatserna i denna slutrapport är resultaten av försöksperioden positiva, eftersom det allmänt konstateras att fördelningen av FISIM skulle leda till avsevärda förbättringar av ENS 95-metodiken och mer exakta jämförelser av bruttonationalprodukten (BNP) inom Europeiska unionen.
(4) Eftersom slutsatserna i den slutliga utvärderingsrapporten är positiva i fråga om tillförlitligheten hos de resultat som erhållits under försöksperioden, måste den metod som skall användas för fördelningen av FISIM antas före den 31 december 2002 enligt artikel 5.3 i förordning (EG) nr 448/98.
(5) I sin slutrapport till Europaparlamentet och rådet anger kommissionen att det skulle vara ändamålsenligt om medlemsstaterna fick två år till på sig för att ytterligare förbättra de källor och metoder som använts för fördelningen av FISIM.
(6) Kommittén för valuta-, finans- och betalningsbalansstatistik, inrättad genom rådets beslut 91/115/EEG(4), ändrat genom beslut 96/174/EG(5), har hörts.
(7) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för det statistiska programmet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Medlemsstaterna skall göra följande beräkningar och fördelningar enligt de specificerade metoder som anges i bilaga III till rådets förordning (EG) nr 448/98:
a) Beräkningen och fördelningen av FISIM efter användarsektorer med hjälp av den referensränta som anges som %quot%Metod 1%quot% i punkt 1 b i bilaga III till rådets förordning (EG) nr 448/98.
b) Beräkningen och fördelningen av import och export av FISIM (inklusive FISIM mellan inhemska finansförmedlare och i utlandet etablerade finansförmedlare) med hjälp av den referensränta som anges som den %quot%externa%quot% referensräntan i punkt 1 b i bilaga III till rådets förordning (EG) nr 448/98.
c) Fördelningen av FISIM efter användande näringsgrenar baserat på stockarna för ut- och inlåning för varje näringsgren eller, om dessa uppgifter inte är tillförlitliga, på produktionen för varje näringsgren.
d) Beräkningen av FISIM till konstanta priser på basis av den formel som anges i punkt 3 i bilaga III till rådets förordning (EG) nr 448/98.
2. Medlemsstaterna skall till kommissionen översända resultaten av de beräkningar som görs enligt denna artikel som del av de sammanställningar som avses i artikel 3 i förordning (EG) nr 2223/96 (Leveransprogram för nationalräkenskapsdata), inklusive tillbakaskrivningar från 1995 och framåt.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Den skall tillämpas från och med den 1 januari 2005.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 2014/2002
av den 7 november 2002
om klassificering av vissa varor i Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan(1), senast ändrad genom kommissionens förordning (EG) nr 969/2002(2), särskilt artikel 9 i denna, och
av följande skäl:
(1) För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till förordning (EEG) nr 2658/87, är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till denna förordning.
(2) I förordning (EEG) nr 2658/87 har allmänna bestämmelser fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
(3) Enligt dessa allmänna bestämmelser måste de varor som beskrivs i kolumn 1 i tabellen som är bifogad den här förordningen klassificeras enligt motsvarande KN-nummer i kolumn 2 med de motiveringar som ges i kolumn 3.
(4) Det är lämpligt att bindande klassificeringsbesked som utfärdas av medlemsstaternas tullmyndigheter avseende varuklassificeringen i Kombinerade nomenklaturen och som inte överensstämmer med de rättigheter som fastställs i denna förordning fortfarande kan åberopas av innehavaren enligt bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(3), senast ändrad genom Europaparlamentets och rådets förordning (EG) nr 2700/2000(4), under en period av tre månader.
(5) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Tullkodexkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 2
Bindande klassificeringsbesked som utfärdas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 2147/2002
av den 2 december 2002
om ändring av förordning (EG) nr 1455/1999 om handelsnormer för paprika
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 2200/96 av den 28 oktober 1996 om den gemensamma organisationen av marknaden för frukt och grönsaker(1), senast ändrad genom förordning (EG) nr 545/2002(2), särskilt artikel 2.2 i denna, och
av följande skäl:
(1) I kommissionens förordning (EG) nr 1455/1999(3), ändrad genom förordning (EG) nr 2706/2000(4), fastställs bestämmelser om märkning och presentation av förpackningar med paprika.
(2) För att förbättra överskådligheten på världsmarknaden bör den ändring beaktas som nyligen gjordes av de handelsnormer för paprika som rekommenderats av Förenta nationernas ekonomiska kommission för Europa (ECE/FN) och som innebär att de förpackningar som innehåller paprika av olika färger inte nödvändigtvis behöver innehålla lika många paprikor av varje färg, förutsatt att märkningen på förpackningen är anpassad efter detta. Dessutom bör det föreskrivas att konsumentförpackningar bör få innehålla inte bara paprika av olika färg utan även paprika av olika typ.
(3) Bestämmelserna om märkning bör förtydligas på flera punkter, särskilt när det gäller märkningen av konsumentförpackningar som innehåller blandningar av paprikor av olika typ och/eller färg.
(4) Förordning (EG) nr 1455/1999 måste därför ändras.
(5) För att kunna tillämpa bestämmelserna i den här förordningen måste aktörerna genomföra vissa tekniska anpassningar, särskilt när det gäller förpackningsutrustningen. Den här förordningen bör därför börja tillämpas först sedan en tillräckligt lång period förflutit efter ikraftträdandet.
(6) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för färsk frukt och färska grönsaker.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till förordning (EG) nr 1455/1999 skall ändras i enlighet med bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Den skall tillämpas från och med den första dagen i den tredje månaden efter den månad då den träder i kraft.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Europeiska centralbankens beslut
av den 20 mars 2003
om valörer, tekniska specifikationer, reproducering, inlösen och indragning avseende eurosedlar
(ECB/2003/4)
(2003/205/EG)
ECB-RÅDET HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 106.1 i detta, och av artikel 16 i stadgan för Europeiska centralbankssystemet och Europeiska centralbanken, och
av följande skäl:
(1) Enligt artikel 106.1 i fördraget och artikel 16 i stadgan har Europeiska centralbanken (ECB) ensamrätt att tillåta sedelutgivning inom gemenskapen. Där anges även att ECB och de nationella centralbankerna får ge ut sådana sedlar. Enligt artikel 10 i rådets förordning (EG) nr 974/98 av den 3 maj 1998 om införande av euron(1) skall ECB och centralbankerna i de deltagande medlemsstaterna sätta eurosedlar i omlopp.
(2) Europeiska monetära institutet (EMI) förberedde framställningen och utgivningen av eurosedlar. Särskilt vad gäller utformningen av sedlarna underlättade EMI för användarna att känna igen och acceptera de nya sedlarnas valörer och tekniska specifikationer genom att beakta de olika visuella och tekniska krav som framfördes av europeiska sammanslutningar av professionella sedelanvändare.
(3) ECB har som EMI:s efterträdare övertagit upphovsrätten till mönstren för eurosedlarna från EMI. ECB och de nationella centralbankerna som företrädare för ECB får göra gällande denna upphovsrätt i fråga om reproduktioner som utgivits eller spritts och som innebär intrång i upphovsrätten, exempelvis reproduktioner som kan ha en negativ inverkan på förtroendet för eurosedlarna.
(4) Eftersom ECB och de nationella centralbankerna har rätt att ge ut eurosedlar inom gemenskapen har de även behörighet att vidta alla nödvändiga rättsliga åtgärder för att skydda eurosedlarnas ställning som betalningsmedel. ECB bör vidta åtgärder för att upprätta en lägsta skyddsnivå i alla deltagande medlemsstater, så att allmänheten kan skilja äkta eurosedlar från reproduktioner. Det är därför nödvändigt att gemensamt reglera i vilka fall reproducering av eurosedlar skall tillåtas.
(5) Bestämmelserna i detta beslut skall inte påverka tillämpningen av straffrättsliga bestämmelser, särskilt när det gäller penningförfalskning.
(6) Reproduktioner av eurosedlar i elektronisk form bör endast anses lagenliga om framställaren använder tekniska medel som förhindrar utskrifter i de fall allmänheten riskerar att förväxla reproduktionerna med äkta eurosedlar.
(7) Behörigheten att vidta åtgärder för att skydda eurosedlarnas ställning som betalningsmedel innefattar även behörighet att införa gemensamma regler, enligt vilka de nationella centralbankerna löser in skadade eurosedlar. I dessa regler anges vissa kategorier av eurosedlar som de nationella centralbankerna bör hålla kvar när de ges in för inlösen.
(8) För inlösen krävs att den del av en ursprunglig eurosedel som ges in skall ha en viss minsta storlek. För att undvika förvanskning av måtten, exempelvis om eurosedeln skadats genom krympning, skall storleken anges i procent av ytan på den ursprungliga eurosedeln, innan den skadades.
(9) För att förmå alla som yrkesmässigt handhar sedlar att använda stöldskyddsutrustningar på rätt sätt är det lämpligt att de får betala en avgift till de nationella centralbankerna, när de begär inlösen hos de nationella centralbankerna av eurosedlar som skadats av stöldskyddsutrustning. Avgiften skall kompensera för analyskostnader i samband med inlösen av eurosedlarna.
(10) Någon avgift skall inte tas ut om sedlarna skadats i samband med rån eller stöld eller försök till rån eller stöld. För att undvika obetydliga avgiftsbelopp skall avgift endast tas ut om ett visst, minsta antal skadade eurosedlar ges in för inlösen.
(11) Stora partier av eurosedlar som skadats genom användning av stöldskyddsutrustning bör ges in för inlösen i satser om ett visst, minsta antal eurosedlar.
(12) ECB:s ensamrätt att tillåta utgivning av eurosedlar inom gemenskapen innefattar behörighet att dra in eurosedlar och att införa gemensamma regler för hur ECB och de nationella centralbankerna skall genomföra dessa indragningar.
(13) Av tydlighets- och rättssäkerhetsskäl är det nödvändigt att kodifiera beslut ECB/2001/7 av den 30 augusti 2001 om valörer och tekniska specifikationer för, och reproducering, inlösen och indragning av, eurosedlar(2), ändrat genom beslut ECB/2001/14(3), och att förtydliga ECB:s och de nationella centralbankernas uppgifter med avseende på de regler som gäller för reproducering, inlösen och indragning av eurosedlar.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Valörer och tekniska specifikationer
1. De första serierna eurosedlar skall omfatta sju valörer mellan 5 euro och 500 euro på temat %quot%epoker och stilar i Europa%quot%, med följande grundläggande tekniska specifikationer:
%gt%Plats för tabell%gt%
2. De sju olika valörerna av eurosedlarna skall ha avbildningar av portar och fönster på framsidan (recto) och broar på baksidan (verso). De sju valörerna skall vara typiska för de olika perioder i den europeiska konsthistorien som nämns ovan. På sedlarna skall dessutom finnas symbolen för Europeiska unionen, valutans namn skrivet med romerska och grekiska bokstäver, ECB:s initialer i de olika officiella språkversionerna, symbolen ©, som anger att ECB innehar upphovsrätten, samt ECB-ordförandens underskrift.
Artikel 2
Regler för reproducering av eurosedlar
1. Med reproduktioner avses alla fysiska och icke fysiska bilder som hämtar material från hela eurosedlar eller delar därav, enligt specifikationerna i artikel 1, eller från delar av sedlarnas enskilda mönsterelement, såsom färger, mått, bokstäver eller symboler, och som kan likna eller erinra om en eurosedel, oberoende av
a) bildens storlek,
b) de material eller tekniker som använts för att framställa den,
c) om beståndsdelar eller bilder tillagts som inte kommer från sedlar, eller
d) om mönstret på eurosedlarna, exempelvis bokstäver eller symboler, har ändrats.
2. Reproduktioner som allmänheten kan förväxla med äkta eurosedlar skall anses vara icke lagenliga.
3. Reproduktioner som uppfyller följande krav skall anses lagenliga, eftersom det inte föreligger någon risk för att allmänheten kan förväxla dem med eurosedlar:
a) Reproduktioner som återger endast ena sidan av en eurosedel, enligt specifikationerna i artikel 1, under förutsättning att reproduktionens mått uppgår till minst 125 % av såväl längden som bredden eller högst 75 % av såväl längden som bredden på respektive eurosedel, enligt specifikationerna i artikel 1.
b) Reproduktioner som återger båda sidorna av en eurosedel, enligt specifikationerna i artikel 1, under förutsättning att reproduktionens mått uppgår till minst 200 % av såväl längden som bredden eller högst 50 % av såväl längden som bredden på respektive eurosedel, enligt specifikationerna i artikel 1.
c) Reproduktioner som återger enskilda mönsterelement på en eurosedel, enligt specifikationerna i artikel 1, under förutsättning att dessa mönsterelement inte avbildas mot en sedelliknande bakgrund.
d) Reproduktioner som återger endast en del av antingen framsidan eller baksidan av en eurosedel, under förutsättning att denna del är mindre än en tredjedel av eurosedelns ursprungliga framsida eller baksida, enligt specifikationerna i artikel 1.
e) Reproduktioner som görs av material som är helt olikt papper, och som ser påtagligt annorlunda ut än det material som används för sedlar.
f) Icke fysiska reproduktioner som görs tillgängliga elektroniskt på webbplatser, på trådbunden eller trådlös väg eller på annat sätt, och till vilka allmänheten har tillgång från en plats och vid en tidpunkt som de själva väljer, under förutsättning
- att ordet SPECIMEN är skrivet diagonalt över reproduktionen i Arial eller ett typsnitt jämförbart med Arial, att längden på ordet SPECIMEN är minst 75 % av längden på reproduktionen och höjden på ordet SPECIMEN minst 15 % av bredden på reproduktionen samt att det är utfört i ogenomskinlig färg som kontrasterar med den dominerande färgen på respektive eurosedel, enligt specifikationerna i artikel 1, och
- att upplösningen på den elektroniska reproduktionen i dess originalstorlek inte överstiger 72 dpi.
4. Efter skriftlig ansökan skall ECB och de nationella centralbankerna intyga att även reproduktioner som inte uppfyller kraven i punkt 3 är lagenliga, för såvitt allmänheten inte kan förväxla dem med äkta eurosedlar enligt specifikationerna i artikel 1. Om en reproduktion framställs på endast en deltagande medlemsstats territorium skall ansökan enligt ovan göras hos den nationella centralbanken i den medlemsstaten. I övriga fall skall ansökan göras hos ECB.
5. Reglerna för reproducering av eurosedlar gäller även i förhållande till eurosedlar som i enlighet med det här beslutet dragits in eller upphört att vara lagliga betalningsmedel.
Artikel 3
Inlösen av skadade eurosedlar
1. De nationella centralbankerna skall på begäran, och i enlighet med villkoren i punkt 2, lösa in skadade, äkta, giltiga eurosedlar i följande fall:
a) om mer än 50 % av eurosedeln ges in, eller
b) om 50 % eller mindre av eurosedeln ges in och inlämnaren kan visa att återstoden av sedeln har förstörts.
2. Utöver vad som anges i punkt 1 gäller följande för inlösen av skadade, giltiga eurosedlar:
a) Om det finns tvivel avseende inlämnarens rätt till eurosedlarna eller om deras äkthet skall inlämnaren identifiera sig.
b) När färgfläckade, förorenade eller infärgade sedlar ges in, skall inlämnaren ge en skriftlig förklaring avseende typen av färg, förorening eller infärgning.
c) När eurosedlar missfärgats på grund av att stöldskyddsutrustning har utlösts, skall en skriftlig förklaring lämnas om varför, och på vilket sätt, sedlarna blivit obrukbara i de fall eurosedlarna ges in av yrkesmässigt verksamma inrättningar enligt artikel 6.1 i rådets förordning (EG) nr 1338/2001 av den 28 juni 2001 om fastställande av nödvändiga åtgärder för skydd av euron mot förfalskning(4).
d) Om stora mängder av eurosedlar skadats genom användning av stöldskyddsutrustning skall de ges in i satser om 100 eurosedlar, när det antal eurosedlar som ges in är tillräckligt för att bilda sådana satser.
3. Trots vad som sägs ovan skall
a) de nationella centralbankerna vägra att lösa in eurosedlar som de vet eller har tillräckliga skäl att anta har skadats avsiktligt, samt hålla kvar eurosedlarna så att dessa inte åter sätts i omlopp eller ges in för inlösen i en annan nationell centralbank. De nationella centralbankerna skall emellertid lösa in de skadade eurosedlarna om de vet eller har tillräckliga skäl att anta att inlämnarna är i god tro, eller om inlämnarna kan visa att de är i god tro. Eurosedlar som endast skadats i mindre utsträckning, exempelvis genom att anteckningar, siffror eller korta fraser anbringats på dem, skall i princip inte anses utgöra avsiktligt skadade eurosedlar,
b) de nationella centralbankerna vägra att lösa in, och mot kvitto hålla kvar, skadade eurosedlar som bevis, om de vet, eller har tillräckliga skäl att anta, att ett brott har begåtts, samt ge in dem till de behöriga myndigheterna så att utredning kan inledas eller sedlarna kan användas som underlag i en pågående utredning. Såvida inte de behöriga myndigheterna beslutar annat, skall sedlarna vid utredningens slut återlämnas till inlämnaren och därefter kunna lösas in.
Artikel 4
Avgift för inlösen av skadade eurosedlar
1. De nationella centralbankerna skall ta ut en avgift av dem som yrkesmässigt handhar sedlar när dessa, i enlighet med artikel 3, begär att de nationella centralbankerna skall lösa in giltiga eurosedlar som skadats genom stöldskyddsutrustning.
2. Avgiften skall vara 10 cent för varje skadad eurosedel.
3. Avgift skall endast tas ut om 100 eller fler skadade eurosedlar löses in. Avgift skall tas ut för samtliga inlösta eurosedlar.
4. Någon avgift skall inte tas ut om eurosedlar skadats i samband med rån eller stöld eller försök till rån eller stöld.
Artikel 5
Indragning av eurosedlar
Indragning av en typ eller serie av eurosedlar skall regleras genom beslut av ECB-rådet, som offentliggörs för allmän kännedom i Europeiska unionens officiella tidning och i andra medier. Ett sådant beslut skall minst omfatta följande uppgifter:
- Den typ eller serie av eurosedlar som skall tas ur omlopp.
- Inlösenperiodens längd.
- Det datum då typen eller serien av eurosedlar upphör att vara lagliga betalningsmedel.
- Behandlingen av eurosedlar som lämnas in efter det att indragningsperioden upphört eller de förlorat sin ställning som lagliga betalningsmedel.
Artikel 6
Slutbestämmelser
1. Beslut ECB/2001/7 och ECB/2001/14 skall upphöra att gälla.
2. Hänvisningar till beslut ECB/1998/6(5), ECB/1999/2(6), ECB/2001/7 och ECB/2001/14 skall gälla som hänvisningar till det här beslutet.
3. Detta beslut träder i kraft dagen efter det att det offentliggörs i Europeiska unionens officiella tidning.
Rådets beslut
av den 16 december 2002
om likvärdighet av fältbesiktningar av utsädesodlingar i tredje land och om likvärdighet av utsäde producerat i tredje land
(Text av betydelse för EES)
(2003/17/EG)
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 66/401/EEG av den 14 juni 1966 om saluföring av utsäde av foderväxter(1), särskilt artikel 16.1 i detta,
med beaktande av rådets direktiv 66/402/EEG av den 14 juni 1966 om saluföring av utsäde av stråsäd(2), särskilt artikel 16.1 i detta,
med beaktande av rådets direktiv 2002/54/EG av den 13 juni 2002 om saluföring av betutsäde(3), särskilt artikel 23.1 i detta,
med beaktande av rådets direktiv 2002/57/EG av den 13 juni 2002 om saluföring av utsäde av olje- och spånadsväxter(4), särskilt artikel 20.1 i detta,
med beaktande av kommissionens förslag, och
av följande skäl:
(1) Enligt reglerna för officiell utsädeskontroll i Argentina, Australien, Bulgarien, Kanada, Chile, Tjeckien, Estland, Kroatien, Ungern, Israel, Lettland, Marocko, Nya Zeeland, Polen, Rumänien, Slovenien, Slovakien, Turkiet, Förenta staterna, Uruguay, Jugoslavien och Sydafrika skall en officiell fältbesiktning utföras under den tid då utsäde produceras.
(2) Enligt dessa regler får utsäde i princip certifieras officiellt och sädesförpackningar förslutas officiellt i enlighet med OECD:s system för sortkontroll av utsäde som är avsett för internationell handel. Reglerna innebär dessutom att provtagning och undersökning skall utföras i enlighet med Internationella frökontrollorganisationens (ISTA) metoder, eller i tillämpliga fall enligt AOSA:s (Association of Official Seed Analysts) regler.
(3) En granskning av dessa regler och tillämpningen av dem i nämnda tredje länder har visat att fältbesiktningarna av utsädesodlingar uppfyller de villkor som fastställs i direktiven 66/401/EEG, 66/402/EEG, 2002/54/EG och 2002/57/EG. De nationella bestämmelserna för utsäde som skördas och kontrolleras i dessa länder när det gäller utsädets egenskaper, möjligheterna till undersökning av utsädet, till säkerställande av utsädets identitet, till märkning och till kontroll, ger samma garantier som de bestämmelser som gäller för utsäde som skördas och kontrolleras inom gemenskapen, under förutsättning att ytterligare villkor för utsädesodlingar och för det producerade utsädet, i synnerhet när det gäller märkningen av förpackningarna, är uppfyllda.
(4) Genom rådets beslut 95/514/EG av den 29 november 1995 om likvärdighet av fältbesiktningar av utsädesodlingar i tredje land och om likvärdighet av utsäde producerat i tredje land(5) föreskrivs det att fältbesiktningar av utsädesodlingar av vissa arter i vissa tredje länder under en begränsad period är likvärdiga med fältbesiktningar som utförs enligt gemenskapens lagstiftning och att utsäde av vissa arter som producerats i de länderna är likvärdigt med utsäde som producerats enligt gemenskapens lagstiftning.
(5) Eftersom beslut 95/514/EG löper ut den 31 december 2002 bör ett nytt beslut antas och dess räckvidd utvidgas, särskilt genom att Estland, Lettland och Jugoslavien inkluderas.
(6) Det är önskvärt att begränsa erkännandet av denna likvärdighet enligt detta beslut till fem år.
(7) Det är lämpligt att i detta beslut inkludera specifika regler för ommärkning och återförslutning i gemenskapen genom att införliva regler motsvarande dem som föreskrivs i beslut 86/110/EEG(6), vilket inte längre är tillämpligt.
(8) Gällande lagstiftning föreskriver redan en skyldighet att för utsäde som saluförs inom gemenskapen, inklusive inte slutgiltigt certifierat utsäde, ange om utsädet är kemiskt behandlat eller om sorten är genetiskt modifierad. Det är lämpligt att fastställa detaljerade bestämmelser för hur detta skall anges på etiketten för sådant certifierat utsäde som importeras enligt detta beslut. Det är lämpligt att dessa bestämmelser återspeglar bestämmelserna i beslut 95/514/EG. Det är lämpligt att i framtiden uppdatera bilagorna till det här beslutet för att säkerställa att importerat utsäde omfattas av krav som är likvärdiga med alla nya bestämmelser som kan införas, särskilt för inte slutgiltigt certifierat utsäde.
(9) Vissa ändringar i bilagorna till detta beslut bör antas enligt rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(7).
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Sådana fältbesiktningar som avser utsädesodlingar av arterna i bilaga I och som utförs i de tredje länder som anges i samma bilaga, med undantag för utsäde från generationer som föregår basutsädet, skall anses likvärdiga med fältbesiktningar utförda enligt direktiven 66/401/EEG, 66/402/EEG, 2002/54/EG och 2002/57/EG på följande villkor:
a) De skall utföras officiellt av de myndigheter som förtecknas i bilaga I eller under dessa myndigheters officiella överinseende.
b) Villkoren i punkt A i bilaga II skall vara uppfyllda.
Artikel 2
Utsäde av de arter som anges i bilaga I, vilket producerats i de tredje länder som anges i samma bilaga och officiellt certifierats av de myndigheter som anges i denna bilaga, med undantag av utsäde från generationer som föregår basutsädet, skall betraktas som likvärdigt med utsäde som uppfyller villkoren i direktiven 66/401/EEG, 66/402/EEG, 2002/54/EG och 2002/57/EG, om det uppfyller de villkor som fastställs i punkt B i bilaga II.
Artikel 3
1. När likvärdiga utsädespartier har märkts om och återförslutits i gemenskapen enligt OECD:s system för sortkontroll av utsäde som är avsett för internationell handel, skall bestämmelserna i direktiven 66/401/EEG, 66/402/EEG, 2002/54/EG och 2002/57/EG för återförslutning av förpackningar som producerats i gemenskapen tillämpas på motsvarande sätt.
Första stycket skall inte påverka tillämpningen av de OECD-regler som omfattar sådana åtgärder.
2. När det är nödvändigt att märka om och återförsluta likvärdiga utsädespartier i gemenskapen, skall EG-märkning användas endast om
a) det utsäde som produceras i medlemsstaterna och det utsäde av samma sort och kategori som produceras i tredje land blandas för att förbättra grobarheten, under förutsättning att
- blandningen är homogen, och
- varje produktionsland anges på etiketten, eller
b) för EG-småförpackningar enligt direktiv 66/401/EEG eller 2002/54/EG.
Artikel 4
Ändringar i bilagorna skall, med undantag för dem som gäller kolumn 1 i tabellen i bilaga I, antas enligt förfarandet i artikel 5.2.
Artikel 5
1. Kommissionen skall biträdas av Ständiga kommittén för utsäde och uppförökningsmateriel för jordbruk, trädgårdsnäring och skogsbruk.
2. När det hänvisas till denna punkt skall artiklarna 4 och 7 i beslut 1999/468/EG tillämpas.
Den tid som avses i artikel 4.3 i beslut 1999/468/EG skall vara en månad.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 6
Detta beslut skall tillämpas från och med den 1 januari 2003 till och med den 31 december 2007.
Artikel 7
Detta beslut riktar sig till medlemsstaterna.
Rådets beslut
av den 19 december 2002
om ingående av ett protokoll om anpassning av handelsaspekterna i Europaavtalet om upprättande av en associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Rumänien, å andra sidan, för att beakta resultaten av förhandlingarna mellan parterna om nya ömsesidiga jordbruksmedgivanden
(2003/18/EG)
EUROPEISKA UNIONENS RÅD HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 133 jämförd med artikel 300.2 första stycket första meningen i detta,
med beaktande av kommissionens förslag, och
av följande skäl:
(1) I Europaavtalet om upprättande av en associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan och Rumänien å andra sidan(1), föreskrivs om vissa ömsesidiga handelsmedgivanden för vissa produkter.
(2) I artikel 21.5 i Europaavtalet föreskrivs att gemenskapen och Rumänien skall undersöka möjligheterna, produkt för produkt och på en ordnad ömsesidig grundval, att bevilja varandra ytterligare koncessioner.
(3) De första förbättringarna av förmånsordningen i Europaavtalet med Rumänien gjordes genom protokollet om anpassning av handelsaspekterna i Europaavtalet för att beakta Republiken Österrikes, Republiken Finlands och Konungariket Sveriges anslutning till Europeiska unionen och resultaten av förhandlingarna inom Uruguayrundan, däribland förbättringarna av den befintliga förmånsordningen, godkänt genom rådets beslut 98/626/EG(2).
(4) Förhandlingarna om liberalisering av jordbrukshandeln som avslutades 2000 ledde också till förbättringar av förmånsordningen. För gemenskapens del trädde förbättringarna i kraft den 1 juli 2000 genom rådets förordning (EG) nr 2435/2000 av den 17 oktober 2000 om vissa medgivanden i form av gemenskapstullkvoter för vissa jordbruksprodukter och om anpassning, som en autonom övergångsåtgärd, av vissa jordbruksmedgivanden enligt Europaavtalet med Rumänien(3). Denna andra anpassning av förmånsordningen har ännu inte integrerats med Europaavtalet som ett tilläggsprotokoll till detta.
(5) Förhandlingar för ytterligare förbättringar av förmånsordningen i Europaavtalet med Rumänien avslutades den 18 juni 2002.
(6) Det nya protokollet till Europaavtalet om anpassning av handelsaspekterna i Europaavtalet mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Rumänien, å andra sidan (nedan kallat %quot%protokollet%quot%) bör antas med sikte på en konsolidering av alla medgivanden inom jordbrukshandeln mellan de två parterna, inklusive resultaten av de förhandlingar som avslutades 2000 och 2002.
(7) I kommissionens förordning (EEG) nr 2454/93 av den 2 juli 1993 om tillämpningsföreskrifter för rådets förordning (EEG) nr 2913/92 om inrättandet av en tullkodex för gemenskapen(4) fastställs förvaltningsföreskrifterna för de tullkvoter som skall användas i kronologisk ordning efter tulldeklarationernas datum. Vissa tullkvoter som fastställs i det här beslutet bör därför förvaltas i enlighet med de föreskrifterna.
(8) De åtgärder som är nödvändiga för att genomföra detta beslut bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(5).
(9) Till följd av ovannämnda förhandlingar har förordning (EG) nr 2435/2000 blivit överflödig och bör därför upphöra att gälla.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Protokollet om anpassning av handelsaspekterna i Europaavtalet om upprättande av en associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Rumänien, å andra sidan, för att beakta resultaten av förhandlingarna mellan parterna om nya ömsesidiga jordbruksmedgivanden godkänns härmed på gemenskapens vägnar.
Artikel 2
1. Rådets ordförande bemyndigas härmed att utse den person som skall ha rätt att underteckna protokollet på gemenskapens vägnar med bindande verkan för denna.
2. Rådets ordförande skall på gemenskapens vägnar lämna den underrättelse om godkännande som det föreskrivs om i artikel 3 i protokollet.
Artikel 3
1. När detta beslut träder i kraft skall den ordning som föreskrivs i bilagan till protokollet som åtföljer detta beslut ersätta den ordning som avses i bilagorna XI och XII till vilka hänvisning görs i artikel 21.2 och 21.4, i deras ändrade lydelse, i Europaavtalet om upprättande av en associering mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Rumänien, å andra sidan.
2. Kommissionen skall anta tillämpningsföreskrifter för detta protokoll i enlighet med förfarandet i artikel 5.2.
Artikel 4
1. De löpnummer som gäller inom tullkvoterna i bilagan till detta beslut får ändras av kommissionen i enlighet med förfarandet i artikel 5.2. Tullkvoter med löpnummer över 09.5100 skall förvaltas av kommissionen i enlighet med artikel 308a, 308b och 308c i förordning (EEG) nr 2454/93.
2. De kvantiteter varor som omfattas av tullkvoter och övergår till fri omsättning från och med den 1 juli 2002 enligt de medgivanden som föreskrivs i bilaga A.b till förordning (EG) nr 2435/2000 skall till fullo räknas av mot de kvantiteter som det föreskrivs om i fjärde kolumnen bilaga A.b till bifogat protokoll, utom när det gäller kvantiteter för vilka importlicens utfärdades före den 1 juli 2002.
Artikel 5
1. Kommissionen skall biträdas av den förvaltningskommitté för spannmål som inrättades genom artikel 23 i rådets förordning (EEG) nr 1766/92(6) eller, i tillämpliga fall, den kommitté som inrättats genom tillämpliga bestämmelser i andra förordningar om den gemensamma organisationen av jordbruksmarknader.
2. När det hänvisas till denna punkt, skall artiklarna 4 och 7 i beslut 1999/468/EG tillämpas.
Den tid som avses i artikel 4.3 i beslut 1999/468/EG skall vara en månad.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 6
Förordning (EG) nr 2435/2000 skall upphöra att gälla samma dag som protokollet träder i kraft.
Kommissionens beslut
av den 30 december 2002
om att utveckla ett integrerat veterinärdatasystem
[delgivet med nr K(2002) 5496]
(2003/24/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 90/425/EEG av den 26 juni 1990 om veterinära och avelstekniska kontroller i handeln med vissa levande djur och varor inom gemenskapen med sikte på att förverkliga den inre marknaden(1), senast ändrat genom direktiv 118/20/EEG(2), särskilt artikel 20.3 i detta,
med beaktande av rådets beslut 92/438/EEG av den 13 juli 1992 om datorisering av veterinära förfaranden vid import (Shift-projektet), om ändring av direktiven 90/675/EEG, 91/496/EEG, 91/628/EEG och beslut 90/424/EEG och om upphävande av beslut 88/192/EEG(3), senast ändrat genom rådets beslut 95/1/EG(4), särskilt artikel 12 i detta,
med beaktande av rådets beslut 90/424/EEG av den 26 juni 1990 om utgifter inom veterinärområdet(5), senast ändrat genom beslut 2001/572/EG(6), särskilt artikel 37 och artikel 37a i detta, och
av följande skäl:
(1) Europaparlamentets och rådets direktiv 1999/93/EG av den 13 december 1999 om ett gemenskapsramverk för elektroniska signaturer(7) syftar till att göra elektronisk kommunikation säker och förtroendeingivande och att göra den lättare att använda av de nationella förvaltningarna och gemenskapens förvaltningar, både sinsemellan och vid kontakter med unionens medborgare och ekonomiska aktörer.
(2) Genom kommissionens beslut 92/563/EEG av den 19 november 1992 om den databas inom Shift-projektet som skall innehålla gemenskapens importbestämmelser(8), åläggs kommissionen att utveckla de relevanta databaserna.
(3) Genom kommissionens beslut 92/398 av den 19 juli 1991 om ett datoriserat nätverk som länkar samman veterinärmyndigheterna (Animo)(9) fastställs principerna för det kommunikationsnätverk som skall binda samman de veterinära enheterna.
(4) Flera arbeten som har utförts på gemenskapsnivå inom ramen för studier och seminarier har kommit till slutsatsen att det är nödvändigt att göra en översyn av Animo-nätets uppbyggnad för att införa ett veterinärsystem som integrerar olika datortillämpningar.
(5) I Europaparlamentets resolution A5-0396/2000 om revisionsrättens särskilda rapport nr 1/2000(10) om klassisk svinpest begärs att Animo-nätet skall förvaltas och utformas helt och hållet under kommissionens överinseende och att ändringar skall genomföras enligt revisionsrättens synpunkter.
(6) För att funktioner och användargränssnitt skall bli så bra som möjligt bör medlemsstaterna vara direkt engagerade i arbetet med att utveckla ett integrerat veterinärdatasystem.
(7) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Gemenskapen skall snarast möjligt införa ett datasystem som innebär att funktionerna i Animo- och Shift-systemen integreras i samma arkitektur. De tekniska specifikationerna anges i bilagan.
Artikel 2
1. Under det första steget skall kommissionen utarbeta specifikationer för det nya Animo-systemet, analysera det och lägga fram en prototyp.
Kommissionen disponerar 200000 euro för detta ändamål.
2. Under det andra steget skall kommissionen utarbeta Animo-systemet och ställa databasen till medlemsstaternas förfogande.
3. Kommissionen skall också se till att Shift-systemet utvecklas och integreras i det nya datasystemet, och särskilt de funktioner som krävs för att understödja beslutsfattandet vid gränskontroller, både när det gäller regelverket och när det gäller riskanalyser.
Artikel 3
Generaldirektören vid Generaldirektoratet för hälsa och konsumentskydd bemyndigas att på Europeiska kommissionens vägnar underteckna de avtal som är nödvändiga för att genomföra detta beslut.
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 18 mars 2003
om offentliggörande av referensnumret för standarden EN 613:2000 %quot%Gasutrustningar - Gaseldade konvektorer%quot% i enlighet med rådets direktiv 90/396/EEG
[delgivet med nr K(2003) 710]
(Text av betydelse för EES)
(2003/189/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 90/396/EEG av den 29 juni 1990 om tillnärmning av medlemsstaternas lagstiftning om anordningar för förbränning av gasformiga bränslen(1), ändrat genom direktiv 93/68/EEG(2), särskilt artikel 6.1 i detta,
med beaktande av yttrandet från den ständiga kommitté som inrättats med stöd av artikel 5 i Europaparlamentets och rådets direktiv 98/34/EG av den 22 juni 1998 om ett informationsförfarande beträffande tekniska standarder och föreskrifter samt föreskrifter för informationssamhällets tjänster(3), ändrat genom direktiv 98/48/EG(4), och
av följande skäl:
(1) I artikel 2 i direktiv 90/396/EEG föreskrivs att anordningar för förbränning av gasformiga bränslen får släppas ut på marknaden och tas i bruk endast om de, vid normal användning, inte äventyrar säkerheten för personer, husdjur eller egendom.
(2) I enlighet med artikel 5 i direktiv 90/396/EEG förutsätts de grundläggande krav för anordningar för förbränning av gasformiga bränslen som åsyftas i artikel 3 i direktivet vara uppfyllda när anordningarna följer de tillämpliga nationella standarder som överför de harmoniserade standarder vars referensnummer har offentliggjorts i Europeiska unionens officiella tidning.
(3) Medlemsstaterna skall offentliggöra referensnumren för de nationella standarder som överför de harmoniserade standarder vars referensnummer har offentliggjorts i Europeiska unionens officiella tidning.
(4) Förenade kungariket har protesterat formellt mot den harmoniserade standarden EN 613:2000 %quot%Gasutrustningar - Gaseldade konvektorer%quot%, som den europeiska standardiseringsorganisationen (CEN) antog den 13 juli 2000 och vars referensnummer offentliggjordes i Europeiska gemenskapernas officiella tidning den 18 juli 2001(5), med motiveringen att den inte helt uppfyller de grundläggande kraven i direktiv 90/396/EEG, särskilt inte dem som nämns i 2.1 och 3.2.2 i bilaga 1, och eftersom konstruktionskraven för gaseldade brasor med front av dekorationsglas inte är tillräckliga för att säkerställa en hög säkerhetsnivå. Förenade kungariket befarar i synnerhet att en farlig situation kan uppstå i förbindelse med sådana produkter vid en eventuell gasansamling, eftersom den samlade oförbrända gasen kan antändas och vålla allvarlig skada.
(5) På grundval av den information som har framkommit vid samråd med nationella myndigheter, CEN och den kommitté som inrättats med stöd av direktiv 98/34/EG har det inte framkommit några bevis till stöd för denna risk för gasansamling eller gasexplosion. Följaktligen saknas det belägg för att den harmoniserade standarden EN 613:2000 inte uppfyller de grundläggande kraven i direktiv 90/396/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Referensnumret för standarden EN 613:2000 %quot%Gasutrustningar - Gaseldade konvektorer%quot%, som den europeiska standardiseringsorganisationen (CEN) antog den 13 juli 2000 och som offentliggjordes i Europeiska gemenskapernas officiella tidning den 18 juli 2001, skall inte strykas från den förteckning över standarder som offentliggjorts i Europeiska unionens officiella tidning. Standarden innebär därför även fortsättningsvis att överensstämmelse med de relevanta bestämmelserna i direktiv 90/396/EEG kan förutsättas.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Rådets beslut
av den 13 juni 2003
om ändring av bilaga 12 till de gemensamma konsulära anvisningarna och bilaga 14 a till den gemensamma handboken vad gäller viseringsavgifter
(2003/454/EG)
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA BESLUT
med beaktande av rådets förordning (EG) nr 789/2001 av den 24 april 2001 om att förbehålla rådet genomförandebefogenheter avseende vissa detaljerade bestämmelser och praktiska förfaranden för behandlingen av ansökningar om visering(1),
med beaktande av rådets förordning (EG) nr 790/2001 av den 24 april 2001 om att förbehålla rådet genomförandebefogenheter avseende vissa detaljerade bestämmelser och praktiska förfaranden för genomförandet av gränskontroller och övervakning(2),
med beaktande av Republiken Greklands initiativ, och
av följande skäl:
(1) I rådets beslut 2002/44/EG av den 20 december 2001 om ändring av del VII i och bilaga 12 till de gemensamma konsulära anvisningarna samt av bilaga 14 a till den gemensamma handboken(3) fastställdes det att de avgifter som tas ut i samband med en ansökan om visering skall motsvara de administrativa kostnaderna. De gemensamma konsulära anvisningarna och den gemensamma handboken bör därför ändras i enlighet härmed.
(2) Avgiftsbeloppen bör ses över regelbundet.
(3) I enlighet med artiklarna 1 och 2 i det till Fördraget om Europeiska unionen och Fördraget om upprättandet av Europeiska gemenskapen fogade protokollet om Danmarks ställning deltar Danmark inte i antagandet av detta beslut, som inte är bindande för eller tillämpligt i Danmark. Eftersom detta beslut bygger på Schengenregelverket enligt bestämmelserna i avdelning IV i tredje delen av Fördraget om upprättandet av Europeiska gemenskapen, skall Danmark, i enlighet med artikel 5 i nämnda protokoll, inom en tid av sex månader efter det att rådet har antagit detta beslut besluta huruvida landet skall genomföra det i sin nationella lagstiftning.
(4) När det gäller Island och Norge utgör detta beslut i enlighet med avtalet mellan Europeiska unionens råd och Republiken Island och Konungariket Norge om dessa staters associering till genomförandet, tillämpningen och utvecklingen av Schengenregelverket(4), en utveckling av bestämmelser i Schengenregelverket vilka omfattas av det område som avses i artikel 1 punkt A i rådets beslut 1999/437/EG av den 17 maj 1999 om vissa tillämpningsföreskrifter för det avtalet(5).
(5) Detta beslut utgör en utveckling av bestämmelser i Schengenregelverket i vilka Förenade kungariket inte deltar i enlighet med rådets beslut 2000/365/EG av den 29 maj 2000 om en begäran från Förenade konungariket Storbritannien och Nordirland om att få delta i vissa bestämmelser i Schengenregelverket(6). Förenade kungariket deltar därför inte i antagandet av detta beslut, som inte är bindande för eller tillämpligt i Förenade kungariket.
(6) Detta beslut utgör en utveckling av bestämmelser i Schengenregelverket i vilka Irland inte deltar i enlighet med rådets beslut 2002/192/EG av den 28 februari 2002 om Irlands begäran om att få delta i vissa bestämmelser i Schengenregelverket(7). Irland deltar därför inte i antagandet av detta beslut, som är inte bindande för eller tillämpligt i Irland.
(7) Detta beslut utgör en rättsakt som bygger vidare på Schengenregelverket eller som på annat sätt har samband med det i den mening som avses i artikel 3.2 i 2003 års anslutningsakt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Tabellen i bilaga 12 till de gemensamma konsulära anvisningarna och tabellen i bilaga 14 a till den gemensamma handboken skall ersättas med följande tabell:
%quot%Avgifter motsvarande de administrativa kostnaderna för att behandla en ansökan om visering
%gt%Plats för tabell%gt%%quot%
Artikel 2
Detta beslut skall tillämpas senast från och med den 1 juli 2004.
Medlemsstaterna får tillämpa detta beslut före den 1 juli 2004, förutsatt att de meddelar rådets generalsekretariat från och med vilket datum de är i stånd att göra det.
Artikel 3
Detta beslut riktar sig till medlemsstaterna i enlighet med Fördraget om upprättandet a
Europaparlamentets och rådets direktiv 2003/25/EG
av den 14 april 2003
om särskilda stabilitetskrav för ro-ro-passagerarfartyg
(Text av betydelse för EES)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 80.2 i detta,
med beaktande av kommissionens förslag(1),
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande(2),
efter att ha hört Regionkommittén,
i enlighet med förfarandet i artikel 251 i fördraget(3), och
av följande skäl:
(1) Inom ramen för den gemensamma transportpolitiken bör ytterligare åtgärder vidtas för att öka säkerheten vid passagerartransporter till sjöss.
(2) Gemenskapen vill med alla lämpliga medel undvika att det inträffar olyckor till sjöss i vilka ro-ro-passagerarfartyg är inblandade och som resulterar i förluster av människoliv.
(3) Ro-ro-passagerarfartygens överlevnadsförmåga efter en kollisionsskada, som beror på den standard de håller när det gäller läckstabilitet, är en viktig faktor för passagerarnas och besättningens säkerhet och är särskilt betydelsefull vid räddningsinsatser. Det allvarligaste problemet för ett ro-ro-passagerarfartyg med slutet ro-ro-däck efter en kollisionsskada är effekten av den stora mängd vatten som samlas på det däcket.
(4) Passagerarna och besättningen ombord på ro-ro-passagerarfartyg i hela gemenskapen bör ha rätt att begära att fartyget håller samma höga säkerhetsnivå, oavsett i vilket område det går i trafik.
(5) Med tanke på den betydelse som passagerartransporter till sjöss har för den inre marknaden, är åtgärder på gemenskapsnivå det effektivaste sättet att fastställa en gemensam lägsta säkerhetsnivå för fartyg i hela gemenskapen.
(6) Åtgärder på gemenskapsnivå är det bästa sättet att säkerställa ett harmoniserat genomförande av de principer som överenskommits inom Internationella sjöfartsorganisationen (IMO), samtidigt som därigenom en snedvridning av konkurrensen mellan olika operatörer av ro-ro-passagerarfartyg som går i trafik i gemenskapen kan undvikas.
(7) Allmänna stabilitetskrav för ro-ro-passagerarfartyg i skadat skick fastställdes på internationell nivå genom 1990 års konferens om säkerheten för människoliv till sjöss (SOLAS 90) och infördes i regel II-1/B/8 i SOLAS-konventionen (SOLAS 90-kriterierna). Dessa krav gäller i hela gemenskapen, genom att SOLAS-konventionen är direkt tillämplig på internationella resor och genom att rådets direktiv 98/18/EG av den 17 mars 1998 om säkerhetsbestämmelser och säkerhetsnormer för passagerarfartyg(4) tillämpas på inrikes resor.
(8) Skadestabilitetskriterierna i SOLAS 90 omfattar underförstått effekten av vatten som tränger in på ro-ro-däcket under sjöförhållanden med ungefär 1,5 meters signifikant våghöjd.
(9) Genom IMO-resolution 14 från 1995 gav SOLAS IMO-medlemmar rätt att ingå regionala överenskommelser om de anser att de rådande sjöförhållandena och andra lokala förhållanden kräver särskilda stabilitetskrav i ett visst område.
(10) I Stockholm den 28 februari 1996 kom åtta nordeuropeiska länder, däribland sju medlemsstater, överens om att införa strängare stabilitetskriterier för ro-ro-passagerarfartyg i skadat skick för att hänsyn skall tas till effekten av vatten som samlas på ro-ro-däcket och för att fartygen skall kunna överleva under svårare sjöförhållanden än enligt kriterierna i SOLAS 90 och klara signifikanta våghöjder på upp till 4 meter.
(11) Enligt denna överenskommelse, den s.k. Stockholmsöverenskommelsen, beror de särskilda stabilitetskriterierna på det fartområde där fartyget går i trafik och närmare bestämt på den signifikanta våghöjd som registrerats i detta område. Den signifikanta våghöjden i det område där fartyget går i trafik bestämmer vattennivån på bildäcket efter en olycka där fartyget skadas.
(12) Vid avslutningen av den konferens där Stockholmsöverenskommelsen antogs, konstaterade kommissionen att överenskommelsen inte är tillämplig i andra delar av gemenskapen och förklarade att den hade för avsikt att undersöka de rådande lokala förhållandena i europeiska farvatten där ro-ro-passagerarfartyg går i trafik och att vidta lämpliga åtgärder.
(13) Vid sitt 2074:e möte den 17 mars 1998 avgav rådet en förklaring i vilken det betonades att det var nödvändigt att se till att alla passagerarfartyg som går i trafik under liknande förhållanden håller samma säkerhetsnivå, oavsett om de används för internationella eller inrikes resor.
(14) I sin resolution av den 5 oktober 2000 om den grekiska färjan Saminas förlisning(5) förklarade Europaparlamentet att det inväntar kommissionens utvärdering av Stockholmsöverenskommelsens effektivitet och av andra åtgärder för att förbättra passagerarfartygs stabilitet och säkerhet.
(15) En expertundersökning som kommissionen har låtit genomföra visar att våghöjderna i sydeuropeiska farvatten är ungefär desamma som i de nordeuropeiska farvattnen. Även om väderförhållandena i allmänhet är gynnsammare i söder, baseras de stabilitetskriterier som fastställs i Stockholmsöverenskommelsen enbart på den signifikanta våghöjden och på hur den påverkar ansamlingen av vatten på ro-ro-däcket.
(16) Tillämpningen av gemenskapens säkerhetskriterier i fråga om stabilitetskrav för ro-ro-passagerarfartyg är mycket viktig för säkerheten ombord på dessa fartyg, och sådana kriterier måste ingå i det gemensamma ramverket om säkerheten till sjöss.
(17) För att förbättra säkerheten och undvika en snedvridning av konkurrensen bör de gemensamma säkerhetskriterierna i fråga om stabilitet tillämpas på alla ro-ro-passagerarfartyg som är i reguljär trafik till eller från en hamn i en medlemsstat i internationell trafik, oavsett vilken flagg de för.
(18) Fartygssäkerheten är huvudsakligen flaggstaternas ansvar, och varje medlemsstat bör därför se till att de ro-ro-passagerarfartyg som för dess flagg uppfyller de tillämpliga säkerhetskraven.
(19) Medlemsstaterna bör också omfattas i egenskap av värdstater. De befogenheter som de utövar i denna egenskap bygger på särskilda hamnstatsbefogenheter som fullt ut överensstämmer med Förenta nationernas havsrättskonvention från 1982 (UNCLOS).
(20) De särskilda stabilitetskrav som införs genom detta direktiv bör baseras på en metod som fastställs i bilagorna till Stockholmsöverenskommelsen, enligt vilken vattennivån på ro-ro-däcket efter en kollisionsskada beräknas utifrån två grundläggande parametrar: fartygets restfribord och den signifikanta våghöjden i det fartområde där fartyget går i trafik.
(21) Medlemsstaterna bör bestämma och offentliggöra de signifikanta våghöjderna i de fartområden som korsas av ro-ro-passagerarfartyg i reguljär trafik till eller från deras hamnar. För internationella rutter bör, i tillämpliga fall och då så är möjligt, de stater där trafikens ändpunkter är belägna komma överens om vilken signifikant våghöjd som skall gälla. Signifikanta våghöjder för trafik som bedrivs i samma område under vissa delar av året kan också fastställas.
(22) Alla ro-ro-passagerarfartyg som omfattas av detta direktiv bör uppfylla de stabilitetskrav som gäller med hänsyn till de signifikanta våghöjder som fastställts för det område där fartyget går i trafik. De bör inneha ett certifikat om överensstämmelse som utfärdats av flaggstatens administration och som godtas av alla andra medlemsstater.
(23) Kriterierna i SOLAS 90 ger en säkerhetsnivå som motsvarar de särskilda stabilitetskrav som fastställs genom detta direktiv för fartyg som går i trafik i fartområden där den signifikanta våghöjden är 1,5 meter eller lägre.
(24) Med tanke på de ombyggnader av existerande ro-ro-passagerarfartyg som kan vara nödvändiga för att de skall uppfylla de särskilda stabilitetskraven, bör dessa krav införas successivt under ett antal år, så att den del av branschen som berörs får tillräckligt med tid att uppfylla kraven. En tidtabell för infasning av existerande fartyg bör därför fastställas. Denna tidtabell för infasning bör inte påverka tillämpningen av de särskilda stabilitetskraven i de fartområden som omfattas av bilagorna till Stockholmsöverenskommelsen.
(25) I artikel 4.1 e i rådets direktiv 1999/35/EG av den 29 april 1999 om ett system med obligatoriska besiktningar för en säker drift av ro-ro-passagerarfartyg och höghastighetspassagerarfartyg i reguljär trafik(6) föreskrivs att värdstaterna skall kontrollera att ro-ro-passagerarfartyg och höghastighetspassagerarfartyg uppfyller de särskilda stabilitetskrav som antagits på regional nivå och överförts till deras nationella lagstiftning, när de i den regionen bedriver trafik som omfattas av den nationella lagstiftningen.
(26) Det bör inte krävas att höghastighetspassagerarfartyg enligt definitionen i regel 1 i kapitel X i SOLAS-konventionen, med senare ändringar, skall uppfylla bestämmelserna i detta direktiv, under förutsättning att de fullt ut uppfyller bestämmelserna i IMO:s internationella säkerhetskod för höghastighetsfartyg, med senare ändringar.
(27) De åtgärder som är nödvändiga för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter(7).
(28) Eftersom målet med den föreslagna åtgärden, nämligen att slå vakt om säkerheten för människoliv till sjöss genom att öka ro-ro-passagerarfartygs överlevnadsförmåga efter en skada, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna och de därför på grund av åtgärdens omfattning och verkningar bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget. I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå detta mål.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Syfte
Syftet med detta direktiv är att fastställa en enhetlig nivå för de särskilda stabilitetskraven för ro-ro-passagerarfartyg, vilket kommer att förbättra överlevnadsförmågan för denna fartygstyp efter en kollisionsskada och säkerställa en hög säkerhetsnivå för passagerare och besättning.
Artikel 2
Definitioner
I detta direktiv används följande beteckningar med de betydelser som här anges:
a) ro-ro-passagerarfartyg: ett fartyg som medför fler än tolv passagerare och har ro-ro-lastutrymmen eller lastutrymmen av särskild kategori enligt definitionen i regel II-2/3 i SOLAS-konventionen med senare ändringar.
b) nytt fartyg: fartyg vars köl har sträckts eller som befinner sig på ett motsvarande byggnadsstadium den 1 oktober 2004 eller senare. Ett motsvarande byggnadsstadium avser det stadium på vilket
i) byggande som kan hänföras till ett visst fartyg har påbörjats, och
ii) sammanfogning av fartyget har påbörjats omfattande minst 50 ton eller 1 % av den beräknade mängden byggnadsmaterial, varvid den lägsta angivelsen skall gälla.
c) existerande fartyg: ett fartyg som inte är ett nytt fartyg.
d) passagerare: alla personer med undantag av befälhavaren och medlemmarna av besättningen eller andra personer som i någon egenskap är anställda eller sysselsatta ombord för fartygets behov med undantag av barn under ett år.
e) internationella konventioner: 1974 års internationella konvention om säkerheten för människoliv till sjöss (SOLAS-konventionen) och 1966 års internationella lastlinjekonvention samt därtill hörande protokoll och ändringar som är i kraft.
f) reguljär trafik: en rad överfarter med ro-ro-passagerarfartyg som går i trafik mellan samma två eller flera hamnar, antingen
i) enligt en offentliggjord tidtabell, eller
ii) med så regelbundna eller ofta förekommande överfarter att de utgör en igenkännlig systematisk serie.
g) Stockholmsöverenskommelsen: den överenskommelse som ingicks i Stockholm den 28 februari 1996 i enlighet med resolution 14 från 1995 års SOLAS-konferens, %quot%Regionala överenskommelser om särskilda stabilitetskrav för ro-ro-passagerarfartyg%quot%, antagen den 29 november 1995.
h) flaggstatens administration: de behöriga myndigheterna i den stat vars flagg ro-ro-passagerarfartyget har rätt att föra.
i) värdstat: en medlemsstat till eller från vars hamnar ett ro-ro-passagerarfartyg går i reguljär trafik.
j) internationell resa: en resa till sjöss från en hamn i en medlemsstat till en hamn utanför den medlemsstaten, eller omvänt.
k) särskilda stabilitetskrav: de stabilitetskrav som anges i bilaga I.
l) signifikant våghöjd (hs): den genomsnittliga höjden för den högsta tredjedel våghöjder som har iakttagits under en bestämd period.
m) restfribord (fr): det minsta avståndet mellan det skadade ro-ro-däcket och flytvattenlinjen efter skada, vid skadans placering på fartyget, utan att den ytterligare effekten av mängden vatten på det skadade ro-ro-däcket tas med i beräkningen.
Artikel 3
Räckvidd
1. Detta direktiv skall tillämpas på alla ro-ro-passagerarfartyg, oberoende av flagg, i reguljär trafik till eller från en medlemsstats hamn när de används på internationella resor.
2. Varje medlemsstat skall i egenskap av värdstat säkerställa att ro-ro-passagerarfartyg som för ett tredje lands flagg till fullo uppfyller kraven i detta direktiv innan de får användas på resor till eller från hamnar i den medlemsstaten i enlighet med bestämmelserna i artikel 4 i direktiv 1999/35/EG.
Artikel 4
Signifikanta våghöjder
De signifikanta våghöjderna (hs) skall användas för att bestämma vattennivån på bildäcket då de särskilda stabilitetskraven i bilaga I tillämpas. Värdena på de signifikanta våghöjderna skall vara de som inte överskrids med en sannolikhet på mer än 10 procent på en årlig basis.
Artikel 5
Fartområden
1. Värdstaterna skall senast den 17 maj 2004 upprätta en förteckning över de fartområden som korsas av ro-ro-passagerarfartyg i reguljär trafik till eller från deras hamnar samt motsvarande värden för de signifikanta våghöjderna i dessa områden.
2. Fartområdena och de signifikanta våghöjder som skall tillämpas i dessa områden skall fastställas i samråd mellan de medlemsstater eller, när det är tillämpligt och möjligt, mellan de medlemsstater och tredje länder, där trafikens ändpunkter är belägna. Om fartygets rutt korsar mer än ett fartområde, skall fartyget uppfylla de särskilda stabilitetskraven för den högsta signifikanta våghöjd som fastställts för dessa områden.
3. Förteckningen skall anmälas till kommissionen och offentliggöras i en offentlig databas som skall finnas tillgänglig på den behöriga sjöfartsmyndighetens webbplats. Kommissionen skall underrättas om var denna information finns att tillgå och om eventuella uppdateringar av förteckningen och skälen därtill.
Artikel 6
Särskilda stabilitetskrav
1. Utan att det påverkar tillämpningen av kraven i regel II-1/B/8 i SOLAS-konventionen (SOLAS 90-kriterier), beträffande vattentäta indelningar och stabilitet i skadat skick, skall alla ro-ro-passagerarfartyg som avses i artikel 3.1 uppfylla de särskilda stabilitetskraven i bilaga I till detta direktiv.
2. För ro-ro-passagerarfartyg som uteslutande går i trafik i fartområden där den signifikanta våghöjden är 1,5 meter eller lägre, skall uppfyllandet av kraven i den regel som avses i punkt 1 anses motsvara uppfyllandet av de särskilda stabilitetskrav som anges i bilaga I.
3. Vid tillämpning av kraven i bilaga I skall medlemsstaterna använda riktlinjerna i bilaga II, i den mån detta är praktiskt möjligt och lämpligt med hänsyn till det berörda fartygets konstruktion.
Artikel 7
Införande av de särskilda stabilitetskraven
1. Nya ro-ro-passagerarfartyg skall uppfylla de särskilda stabilitetskraven i bilaga I.
2. Existerande ro-ro-passagerarfartyg, med undantag av fartyg som omfattas av artikel 6.2, skall uppfylla de särskilda stabilitetskraven i bilaga I senast den 1 oktober 2010.
Existerande ro-ro-passagerarfartyg som den 17 maj 2003 uppfyller kraven i den regel som avses i artikel 6.1 skall uppfylla de särskilda stabilitetskraven enligt bilaga I senast den 1 oktober 2015.
3. Denna artikel skall inte påverka tillämpningen av artikel 4.1 e i direktiv 1999/35/EG.
Artikel 8
Certifikat
1. Alla nya och existerande ro-ro-passagerarfartyg som för en medlemsstats flagg skall inneha ett certifikat som visar att de särskilda stabilitetskrav som anges i artikel 6 och i bilaga I är uppfyllda.
Av detta certifikat, som skall utfärdas av flaggstatens administration och som kan kombineras med andra liknande certifikat, skall det framgå upp till vilken signifikant våghöjd fartyget kan uppfylla de särskilda stabilitetskraven.
Certifikatet skall vara giltigt så länge fartyget går i trafik i ett område med samma eller lägre signifikanta våghöjder.
2. Varje medlemsstat skall i egenskap av värdstat erkänna certifikat som utfärdats av en annan medlemsstat i enlighet med detta direktiv.
3. Varje medlemsstat skall i egenskap av värdstat godta certifikat som utfärdats av tredje land och som visar att fartyget uppfyller de särskilda stabilitetskrav som fastställts.
Artikel 9
Trafik under vissa delar av året och trafik under kortare tidsperioder
1. Om ett rederi som bedriver reguljär trafik året runt önskar införa ytterligare ro-ro-passagerarfartyg som skall nyttjas i samma trafik under en kortare period, skall det underrätta värdstatens eller värdstaternas behöriga myndigheter om detta senast en månad innan dessa fartyg börjar nyttjas i denna trafik. Om det emellertid på grund av oförutsedda omständigheter är nödvändigt att snabbt sätta in ett ro-ro-passagerarfartyg som ersättning för att säkerställa kontinuitet i trafiken skall direktiv 1999/35/EG tillämpas.
2. Om ett rederi önskar bedriva reguljär säsongstrafik under kortare tidsperioder som inte överstiger sex månader per år, skall det underrätta värdstatens eller värdstaternas behöriga myndighet om detta senast tre månader innan denna trafik börjar bedrivas.
3. Om sådan trafik bedrivs under förhållanden med lägre signifikant våghöjd än den som fastställts för samma fartområde vid trafik året runt, får den behöriga myndigheten, vid tillämpning av de särskilda stabilitetskraven i bilaga I, använda den signifikanta våghöjd som är tillämplig under denna kortare tidsperiod för att bestämma vattennivån på däck. Den signifikanta våghöjd som är tillämplig under denna kortare tidsperiod skall överenskommas mellan de medlemsstater eller, när så är tillämpligt och möjligt, de medlemsstater och tredje länder där trafikens ändpunkter är belägna.
4. När värdstatens eller värdstaternas behöriga myndighet har gett sitt samtycke till sådan trafik som avses i punkterna 1 och 2, skall ro-ro-passagerarfartyg som används i sådan trafik inneha ett certifikat enligt artikel 8.1 vilket visar att det uppfyller kraven i detta direktiv.
Artikel 10
Anpassning
Bilagorna får ändras i enlighet med förfarandet i artikel 11.2 för att hänsyn skall tas till den internationella utvecklingen, särskilt inom Internationella sjöfartsorganisationen (IMO) samt för att detta direktiv skall bli mer effektivt mot bakgrund av de erfarenheter som gjorts och den tekniska utvecklingen.
Artikel 11
Kommitté
1. Kommissionen skall biträdas av den genom artikel 3 i förordning (EG) nr 2099/2002(8) inrättade Kommittén för sjösäkerhet och förhindrande av förorening från fartyg.
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av artikel 8 i det beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara åtta veckor.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 12
Påföljder
Medlemsstaterna skall fastställa regler om de påföljder som skall gälla vid överträdelser av de nationella bestämmelser som har antagits enligt detta direktiv och skall vidta alla åtgärder som är nödvändiga för att se till att de verkställs. Påföljderna skall vara effektiva, proportionerliga och avskräckande.
Artikel 13
Genomförande
Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv före den 17 november 2004. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
Artikel 14
lkraftträdande
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska unionens officiella tidning.
Artikel 15
Adressater
Detta direktiv riktar sig till medlemsstaterna.
Kommissionens direktiv 2003/77/EG
av den 11 augusti 2003
om ändring av Europaparlamentets och rådets direktiv 97/24/EG och 2002/24/EG om typgodkännande av två- och trehjuliga motorfordon
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets direktiv 2002/24/EG av den 18 mars 2002 om typgodkännande av två- och trehjuliga motorfordon och om upphävande av rådets direktiv 92/61/EEG(1), särskilt artikel 17 i detta,
med beaktande av Europaparlamentets och rådets direktiv 97/24/EG av den 17 juni 1997 om vissa komponenter och karakteristiska egenskaper hos två- eller trehjuliga motorfordon(2), senast ändrat genom direktiv 2002/51/EG(3), särskilt artikel 7 i detta, och
av följande skäl:
(1) Direktiv 97/24/EG är ett av särdirektiven inom ramen för förfarandet för EG- typgodkännande i direktiv 92/61/EEG(4) som skall upphävas den 9 november 2003 genom direktiv 2002/24/EG.
(2) Genom Europaparlamentets och rådets direktiv 2002/51/EG av den 19 juli 2002 om minskning av de förorenande utsläppen från två- och trehjuliga motorfordon och om ändring av direktiv 97/24/EG infördes nya gränsvärden för utsläpp från tvåhjuliga motorcyklar. Dessa gränsvärden skall tillämpas i två steg, varav det första, som gäller alla fordonstyper, från och med den 1 april 2003, och det andra, som gäller nya typer, från och med den 1 januari 2006. I det andra steget grundas mätningen av utsläppen av föroreningar från tvåhjuliga motorcyklar på användningen av den grundläggande körcykeln för stadstrafik i enlighet med FN-ECE-föreskrift nr 40 och körcykeln för landsvägstrafik enligt rådets direktiv 70/220/EEG av den 20 mars 1970 om tillnärmning av medlemsstaternas lagstiftning om åtgärder mot luftförorening genom utsläpp från motorfordon(5), senast ändrat genom kommissionens direktiv 2002/80/EG(6).
(3) I direktiv 97/24/EG, i sin ändrade lydelse enligt direktiv 2002/51/EG, specificeras det typ I-prov som skall mäta utsläpp av föroreningar från två- och trehjuliga motorfordon. Det provet bör kompletteras av kommissionen genom Kommittén för anpassning till teknisk utveckling som inrättats genom artikel 13 i direktiv 70/156/EEG och tillämpas från och med 2006.
(4) Det är nödvändigt att förtydliga vissa sidor av provningsuppgifterna av typ II för den årliga trafiksäkerhetsprovningen enligt direktiv 2002/51/EG och att fastställa regler för registrering av dessa provningsuppgifter enligt bilaga VII till direktiv 2002/24/EG.
(5) Direktiven 97/24/EG och 2002/24/EG bör därför ändras.
(6) De åtgärder som föreskrivs i detta direktiv är förenliga med yttrandet från Kommittén för anpassning till teknisk utveckling.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga II till kapitel 5 i direktiv 97/24/EG skall ändras i enlighet med bilaga I till detta direktiv.
Artikel 2
Bilaga VII till direktiv 2002/24/EG skall ändras i enlighet med bilaga II till detta direktiv.
Artikel 3
1. Medlemsstaterna skall senast den 4 september 2004 anta och offentliggöra de lagar och andra författningar som är nödvändiga för att följa detta direktiv. De skall genast överlämna texterna till dessa bestämmelser till kommissionen tillsammans med en jämförelsetabell för dessa bestämmelser och bestämmelserna i detta direktiv.
De skall tillämpa dessa bestämmelser från och med den 4 september.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texten till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 4
Detta direktiv träder i kraft den tjugonde dagen efter det att det har offentliggjorts i Europeiska unionens officiella tidning.
Artikel 5
Detta direktiv riktar sig till medlemsstaterna.
Kommissionens förordning (EG) nr 47/2003
av den 10 januari 2003
om ändring av bilaga I till rådets förordning (EG) nr 2200/96
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 2200/96 av den 28 oktober 1996 om den gemensamma organisationen av marknaden för frukt och grönsaker(1), senast ändrad genom förordning (EG) nr 545/2002(2), särskilt artikel 2.3 i denna, och
av följande skäl:
(1) I bilaga I till förordning (EG) nr 2200/96 finns en förteckning över produkter som är avsedda att levereras i färskt tillstånd till konsumenten och som underkastas normer.
(2) Detaljhandelsförpackningar som innehåller flera olika arter av frukt och grönsaker blir allt vanligare på marknaden, vilket är en följd av att vissa konsumenter efterfrågar den typen av produkter.
(3) God affärssed innebär att färsk frukt och färska grönsaker som säljs i samma förpackning skall vara av samma kvalitet. Detta innebär att förteckningen över produkter som omfattas av handelsnormer måste utvidgas till att omfatta produkter som i detaljhandelsförpackningar blandas med produkter som redan finns med i förteckningen.
(4) Bilaga I till förordning (EG) nr 2200/96 bör därför ändras.
(5) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för färsk frukt och färska grönsaker.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I bilaga I till förordning (EG) nr 2200/96 skall följande läggas till:
%quot%Andra produkter enligt artikel 1 som ingår i blandningar, i detaljhandelsförpackningar med en nettovikt under 3 kg, som innehåller minst en av de produkter som förtecknas i denna bilaga.%quot%
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska gemenskapernas officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Rådets förordning (EG) nr 561/2003
av den 27 mars 2003
om ändring, när det gäller undantag från frysning av penningmedel och ekonomiska resurser, av förordning (EG) nr 881/2002 om införande av vissa särskilda restriktiva åtgärder mot vissa med Usama bin Ladin, nätverket al-Qaida och talibanerna associerade personer och enheter
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artiklarna 60, 301 och 308 i detta,
med beaktande av gemensam ståndpunkt 2002/402/GUSP av den 27 maj 2002 om restriktiva åtgärder mot Usama bin Ladin, medlemmar av al Qaida-organisationen, talibanerna och andra personer, grupper, företag och enheter associerade med dem och om upphävande av gemensamma ståndpunkterna 96/746/GUSP, 1999/727/GUSP, 2001/154/GUSP och 2001/771/GUSP(1),
med beaktande av gemensam ståndpunkt 2003/140/GUSP av den 27 februari 2003 om undantag från de restriktiva åtgärder som införts genom gemensam ståndpunkt 2002/402/GUSP(2),
med beaktande av kommissionens förslag(3),
med beaktande av Europaparlamentets yttrande(4), och
av följande skäl:
(1) Enligt gemensam ståndpunkt 2002/402/GUSP skall Europeiska gemenskapen bland annat vidta vissa restriktiva åtgärder, exempelvis frysning av penningmedel och ekonomiska resurser, i enlighet med FN:s säkerhetsråds resolution nr 1267 (1999), 1333 (2000) och 1390 (2002).
(2) Frysning av penningmedel och ekonomiska resurser har genomförts genom rådets förordning (EG) nr 881/2002(5).
(3) Genom sin resolution nr 1452 (2002) av den 20 december 2002 har säkerhetsrådet tillåtit vissa undantag när det gäller frysning av penningmedel och ekonomiska resurser enligt resolutionerna nr 1267 (1999), 1333 (2000) och 1390 (2002).
(4) Med hänsyn till resolution 1452 (2002) är det nödvändigt att anpassa de åtgärder som införts av gemenskapen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Följande artikel skall införas i förordning (EG) nr 881/2002:
%quot%Artikel 2a
1. Artikel 2 skall inte vara tillämplig på penningmedel eller ekonomiska resurser om
a) någon av medlemsstaternas behöriga myndigheter enligt förteckningen i bilaga II på begäran av en berörd fysisk eller juridisk person har fastställt att dessa penningmedel eller ekonomiska resurser
i) är nödvändiga för att täcka grundläggande utgifter, inbegripet betalning av livsmedel, hyra, amorteringar och räntor på bostadskrediter, mediciner och läkarvård, skatter, försäkringspremier och avgifter för samhällstjänster,
ii) endast är avsedda för betalning av rimliga arvoden och ersättning av utgifter i samband med tillhandahållande av juridiska tjänster,
iii) endast är avsedda för betalning av avgifter eller serviceavgifter för rutinmässig hantering eller förvaltning av frysta penningmedel eller frysta ekonomiska resurser, eller
iv) är nödvändiga för extraordinära kostnader, och
b) ett sådant fastställande har meddelats sanktionskommittén, och
c) i) när det gäller ett fastställande enligt punkt a i, a ii eller a iii ovan, sanktionskommittén inte har framfört några invändningar mot fastställandet inom 48 timmar efter det att meddelandet lämnats, eller
ii) när det gäller ett fastställande enligt punkt a iv ovan, sanktionskommittén har godkänt fastställandet.
2. Varje person som önskar utnyttja de bestämmelser som anges i punkt 1 skall rikta sin begäran till den relevanta behöriga myndigheten i medlemsstaten enligt förteckningen i bilaga II.
Den behöriga myndigheten enligt förteckningen i bilaga II skall skyndsamt skriftligen meddela den person som framställt begäran samt varje person, organ eller enhet som veterligen berörs direkt huruvida begäran har beviljats.
Den behöriga myndigheten skall också informera andra medlemsstater huruvida begäran om ett sådant undantag har beviljats.
3. Penningmedel som frigörs eller överförs inom gemenskapen för att ombesörja kostnader eller som erkänns enligt denna artikel skall inte omfattas av ytterligare restriktiva åtgärder enligt artikel 2.
4. Artikel 2.2 skall inte avse kreditering av frysta konton med
a) ränta eller andra intäkter på dessa konton, eller
b) betalningar enligt avtal, överenskommelser eller förpliktelser som uppstod före den dag då dessa konton kom att omfattas av bestämmelserna i FN:s säkerhetsråds resolutioner som successivt genomfördes genom förordning (EG) nr 337/2000(6), förordning (EG) nr 467/2001(7) eller denna förordning.
I likhet med det konto som krediteras skall sådan ränta, sådana andra intäkter och sådana betalningar också frysas.%quot%
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 627/2003
av den 4 april 2003
om klassificering av vissa varor i Kombinerade nomenklaturen
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2658/87 av den 23 juli 1987 om tulltaxe- och statistiknomenklaturen och om Gemensamma tulltaxan(1), senast ändrad genom kommissionens förordning (EG) nr 2176/2002(2), särskilt artikel 9 i denna, och
av följande skäl:
(1) För att säkerställa en enhetlig tillämpning av Kombinerade nomenklaturen, som är en bilaga till förordning (EEG) nr 2658/87, är det nödvändigt att anta bestämmelser för klassificering av de varor som avses i bilagan till denna förordning.
(2) I förordning (EEG) nr 2658/87 har allmänna bestämmelser fastställts för tolkningen av Kombinerade nomenklaturen och dessa regler gäller också för varje annan nomenklatur som helt eller delvis grundar sig på denna eller som tillfogar underuppdelningar till denna och som har upprättats genom särskilda gemenskapsbestämmelser för tillämpningen av tulltaxebestämmelser eller andra åtgärder för varuhandeln.
(3) Enligt dessa allmänna bestämmelser måste de varor som beskrivs i kolumn 1 i tabellen som är bifogad den här förordningen klassificeras enligt motsvarande KN-nummer i kolumn 2 med de motiveringar som ges i kolumn 3.
(4) Det är lämpligt att bindande klassificeringsbesked som utfärdas av medlemsstaternas tullmyndigheter avseende varuklassificeringen i Kombinerade nomenklaturen och som inte överensstämmer med de rättigheter som fastställs i denna förordning fortfarande kan åberopas av innehavaren enligt bestämmelserna i artikel 12.6 i rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om inrättandet av en tullkodex för gemenskapen(3), senast ändrad genom Europaparlamentets och rådets förordning (EG) nr 2700/2000(4), under en period av tre månader.
(5) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Tullkodexkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De varor som beskrivs i kolumn 1 i den bifogade tabellen skall i Kombinerade nomenklaturen klassificeras enligt motsvarande KN-nummer i kolumn 2 i samma tabell.
Artikel 2
Bindande klassificeringsbesked som utfärdas av medlemsstaternas tullmyndigheter och som inte stämmer överens med de rättigheter som fastställs i denna förordning kan fortfarande åberopas enligt bestämmelserna i artikel 12.6 i förordning (EEG) nr 2913/92 under en period av tre månader.
Artikel 3
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 808/2003
av den 12 maj 2003
om ändring av Europaparlamentets och rådets förordning (EG) nr 1774/2002 om hälsobestämmelser för animaliska biprodukter som inte är avsedda att användas som livsmedel
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 1774/2002 av den 3 oktober 2002 om hälsobestämmelser för animaliska biprodukter som inte är avsedda att användas som livsmedel(1), särskilt artiklarna 12.5 och 32.1 i denna, och
av följande skäl:
(1) Vetenskapliga styrkommittén lämnade den 16-17 januari 2003 ett yttrande om säkerheten avseende TSE i samband med användning av förbränningsanläggningar med låg kapacitet samt samförbränningsanläggningar för förbränning av animaliskt material som kan vara smittat med TSE.
(2) För att kunna beakta detta yttrande är det lämpligt att ändra bestämmelserna i förordning (EG) nr 1774/2002 avseende användningen av förbränningsanläggningar med låg kapacitet och samförbränningsanläggningar för att bortskaffa slaktkroppar av vissa djur.
(3) Dessutom bör ett antal tekniska ändringar göras i bilagorna till förordning (EG) nr 1774/2002 för att få dem att bättre överensstämma med förordningens artiklar och för att klargöra de bestämmelser som skall tillämpas på ett antal ytterligare produkter.
(4) Det bör fastställas ytterligare bestämmelser för hanteringen av avloppsvatten från anläggningar där det kan förekomma risk för mikrobiologisk eller annan smitta till följd av hantering av kategori 1- eller kategori 2-material.
(5) Det sakfel som gäller de tekniska kraven för bearbetning av biprodukter efter bearbetning med metod nr 2 bör också korrigeras.
(6) Samtidigt som det foderförbud som fastställs i rådets beslut 2000/766/EG(2) kvarstår bör mindre strikta bearbetningskrav tillämpas på bearbetat däggdjursprotein eftersom sådant material på grund av förbudet enbart kan klassificeras som avfall.
(7) Förordning (EG) nr 1774/2002 bör ändras i enlighet med ovanstående.
(8) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Ändring av förordning (EG) nr 1774/2002
Förordning (EG) nr 1774/2002 ändras på följande sätt:
1. Artikel 12.3 a skall ersättas med följande:
%quot%a) användas endast för bortskaffande av döda sällskapsdjur och sådana animaliska biprodukter som avses i artikel 4.1 b och artiklarna 5.1 och 6.1 och som inte omfattas av direktiv 2000/76/EG,%quot%
2. I artikel 12.3 skall följande punkt h läggas till:
%quot%h) uppfylla kraven i kapitel VII i bilaga IV när den används för att bortskaffa sådana animaliska biprodukter som avses i artikel 4.1 b,%quot%
3. Bilagorna I-IX skall ändras i enlighet med bilagan till denna förordning.
Artikel 2
Ikraftträdande
Denna förordning träder i kraft den samma dag som det att den har offentliggjorts i Europeiska unionens officiella tidning.
Den skall tillämpas från och med den 1 maj 2003.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1184/2003
av den 2 juli 2003
om ändring för tjugonde gången av rådets förordning (EG) nr 881/2002 beträffande införande av vissa särskilda restriktiva åtgärder mot vissa med Usama bin Ladin, nätverket al-Qaida och talibanerna associerade personer och enheter och om upphävande av rådets förordning (EG) nr 467/2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 881/2002 av den 27 maj 2002 om införande av vissa särskilda restriktiva åtgärder mot vissa med Usama bin Ladin, nätverket al-Qaida och talibanerna associerade personer och enheter och om upphävande av rådets förordning (EG) nr 467/2001 om förbud mot export av vissa varor och tjänster till Afghanistan, skärpning av flygförbudet och förlängning av spärrandet av tillgångar och andra finansiella medel beträffande talibanerna i Afghanistan(1), senast ändrad genom kommissionens förordning (EG) nr 1012/2003(2), särskilt artikel 7.1 första strecksatsen i denna, och
av följande skäl:
(1) I bilaga I till förordning (EG) nr 881/2002 anges de personer, grupper och enheter som omfattas av det spärrande av tillgångar och ekonomiska resurser som införs genom den förordningen.
(2) Den 25 juni 2003 beslutade sanktionskommittén att ändra förteckningen över de personer, grupper och enheter som bör omfattas av spärrandet av tillgångar och ekonomiska resurser, och bilaga I bör därför ändras i enlighet därmed.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga I till rådets förordning (EG) nr 881/2002 skall ändras i enlighet med bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1458/2003
av den 18 augusti 2003
om öppnande och förvaltning av tullkvoter för griskött
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2759/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för griskött(1), senast ändrad genom förordning (EG) nr 1365/2000(2), särskilt artikel 8.2, artikel 11.1 och artikel 22, andra stycket, i denna,
med beaktande av rådets förordning (EG) nr 1095/96 av den 18 juni 1996 om genomförande av medgivandena i lista CXL som fastställts sedan förhandlingarna enligt GATT artikel XXIV.6 avslutats(3), särskilt artikel 1 i denna, och
av följande skäl:
(1) Kommissionens förordning 1486/95 av den 28 juni 1995 om öppnande och förvaltning av tullkvoter för griskött(4) har ändrats på ett genomgripande sätt(5). För att skapa klarhet och överskådlighet bör den förordningen kodifieras.
(2) Inom ramen för de multilaterala handelsförhandlingarna i Uruguayrundan förhandlade gemenskapen fram olika avtal, särskilt ett jordbruksavtal. Enligt det protokollet fastställs bland annat tillgången till den gemensamma marknaden för vissa grisköttsprodukter med ursprung i tredje land. Det är därför lämpligt att fastställa särskilda tillämpningsföreskrifter för import inom grisköttssektorn.
(3) Enligt avtalet krävs att de rörliga importavgifterna upphävs och att samtliga importrestriktioner i fråga om jordbruksprodukter förvandlas till tullar.
(4) Förvaltningen av detta system bör säkerställas genom importlicenser. För detta ändamål bör särskilt bestämmelserna för licensansökningar och de uppgifter som dessa och licenserna skall innehålla definieras, med undantag från artikel 8 i kommissionens förordning (EEG) nr 1291/2000 av den 9 juni 2000 om gemensamma tillämpningsföreskrifter för systemet med import- och exportlicenser och förutfastställelselicenser för jordbruksprodukter(6), senast ändrad genom förordning (EG) nr 325/2003(7). Utfärdandet av licenser bör ske efter en viss betänketid och eventuellt bör en enhetlig procentsats för godkännande tillämpas på dessa. I aktörernas intresse bör det föreskrivas att licensansökan får dras tillbaka efter fastställandet av en godkännandekoefficient.
(5) För tydlighetens skull är det lämpligt att fastställa att en importlicens krävs för all import som sker inom ramen för en kvot. Den högsta kvantitet som tillåter aktörerna att dra tillbaka licensansökan efter tillämpning av den enhetliga procentsatsen för godkännande bör fastställas.
(6) För att underlätta handel mellan Europeiska gemenskapen och tredje land är det nödvändigt att tillåta import av grisköttsprodukter utan krav på import från ursprungslandet, av statistiska skäl måste dock detta skrivas in i fält 8 i importlicensen.
(7) I syfte att säkerställa en regelbunden import är det nödvändigt att dels definiera vilka produkter som omfattas av importsystemet, dels fördela de kvantiteter som anges i bilaga I till denna förordning under perioden 1 juli-30 juni.
(8) I syfte att säkerställa att systemet förvaltas effektivt är det lämpligt att fastställa 20 euro per 100 kg som säkerhet för importlicenser enligt detta system. Risken för spekulation inom grisköttssektorn gör det lämpligt att aktörernas tillgång till systemet omfattas av vissa preciserade villkor.
(9) Det är lämpligt att fästa aktörernas uppmärksamhet på att licenserna får användas endast för produkter som uppfyller samtliga gällande hygienkrav inom gemenskapen.
(10) För att garantera en god förvaltning av importordningarna behöver kommissionen få exakta uppgifter från medlemsstaterna om de kvantiteter som faktiskt importeras. För tydlighetens skull får medlemsstaterna bara använda en enda modell för att meddela kvantiteterna till kommissionen.
(11) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för griskött.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De importtullkvoter som anges i bilaga I skall öppnas årligen för de produktgrupper och på de villkor som anges i bilagan.
Artikel 2
I denna förordning avses med produkter enligt KN-nummer ex 0203 19 55 och ex 0203 29 55 i grupp G 2 och G 3 i bilaga I:
- benfria styckningsdelar: benfria styckningsdelar, med undantag av filé, med eller utan svål och sidfläsk,
- filé: den styckningsdel som omfattar muskelköttet musculus major psoas och musculus minor psoas, med eller utan huvud, även berett.
Artikel 3
De tullkvoter som anges i bilaga I skall fördelas i kvartalsandelar på 25 %, tillämpliga från och med den 1 juli, 1 oktober, 1 januari respektive 1 april.
Artikel 4
De importlicenser för tullkvoterna som avses i bilaga I skall omfattas av följande bestämmelser:
a) Den som ansöker om importlicens skall vara en fysisk eller juridisk person som vid tidpunkten för inlämnande av ansökan på ett tillfredsställande sätt kan visa medlemsstaternas behöriga myndigheter att han under minst de senaste 12 månaderna utövar handelsverksamhet med tredje land inom grisköttssektorn. Detaljhandel och restauranger som säljer sina produkter direkt till konsumenter skall inte omfattas av systemet.
b) I licensansökan skall endast ett av de gruppnummer som anges i bilaga I till denna förordning anges. Ansökan kan avse flera produkter som omfattas av olika KN-nummer och med ursprung i ett enda land. I detta fall skall alla KN-nummer och varuslag anges i fält 16 respektive 15 i ansökan. För grupp G 2 skall licensansökan avse minst 20 ton och högst 10 % av den disponibla kvantiteten för den period som anges i artikel 3. För de övriga grupperna skall licensansökan avse minst 1 ton och högst 10 % av den disponibla kvantiteten för den period som anges i artikel 3.
c) Fält 8 i licensansökningen och licensen skall innehålla uppgift om ursprungsland.
d) I licensansökan och licensen i fält 20 skall ett av följande anges:
- Reglamento (CE) n° 1458/2003
- Forordning (EF) nr. 1458/2003
- Verordnung (EG) Nr. 1458/2003
- Κανονισμός (ΕΚ) αριθ. 1458/2003
- Regulation (EC) No 1458/2003
- Règlement (CE) n° 1458/2003
- Regolamento (CE) n. 1458/2003
- Verordening (EG) nr. 1458/2003
- Regulamento (CE) n.o 1458/2003
- Asetus (EY) N:o 1458/2003
- Förordning (EG) nr 1458/2003
e) På licensen skall i fält 24 anges: %quot%tullavgift fastställd i ... med tillämpning av%quot% samt något av följande:
- Reglamento (CE) n° 1458/2003
- Forordning (EF) nr. 1458/2003
- Verordnung (EG) Nr. 1458/2003
- Κανονισμός (ΕΚ) αριθ. 1458/2003
- Regulation (EC) No 1458/2003
- Règlement (CE) n° 1458/2003
- Regolamento (CE) n. 1458/2003
- Verordening (EG) nr. 1458/2003
- Regulamento (CE) n.o 1458/2003
- Asetus (EY) N:o 1458/2003
- Förordning (EG) nr 1458/2003.
Artikel 5
1. Licensansökningarna får bara lämnas in under de sju första dagarna under den månad som föregår de perioder som anges i artikel 3.
2. Licensansökan skall inte godtas om den sökande inte skriftligen har förpliktat sig att under den berörda perioden inte lämna in en annan ansökan om produkter ur samma grupp enligt bilaga I i den medlemsstat där ansökan lämnas in eller i en annan medlemsstat.
Om en sökande lämnar in mer än en ansökan för produkter ur samma grupp enligt bilaga I skall ingen av ansökningarna godtas. Varje sökande får dock lämna in flera ansökningar om importlicens för produkter ur samma grupp enligt bilaga I om dessa produkter har sitt ursprung i olika länder.
3. Ansökningar som var och en anger endast ett ursprungsland skall lämnas in samtidigt till medlemsstatens behöriga myndighet. I fråga om den högsta kvantitet som anges i artikel 4 b och vid tillämpningen av bestämmelsen i punkt 2, andra stycket i denna artikel behandlas dessa som en enda ansökan.
4. En säkerhet på 20 euro per 100 kg skall ställas för ansökningar om importlicens för alla de produkter som anges i bilaga I.
5. Medlemsstaterna skall den tredje arbetsdagen efter utgången av perioden för inlämnande av ansökningar underrätta kommissionen om inlämnade ansökningar för var och en av de berörda produktgrupperna. Denna underrättelse skall innehålla en förteckning över de sökande och uppgift om begärda kvantiteter.
Samtliga underrättelser, inbegripet underrättelser om att inga ansökningar lämnats in, skall göras per telex eller telefax på den angivna arbetsdagen i enlighet med den mall som återges i bilaga II om ingen ansökan har lämnats in eller i enlighet med mallarna i bilagorna II och III om ansökningar har lämnats in.
6. Kommissionen skall snarast möjligt besluta i vilken omfattning den kan godkänna de ansökningar som avses i artikel 4.
Om de kvantiteter för vilka licenser har ansökts överstiger tillgängliga kvantiteter skall kommissionen fastställa en enhetlig procentandel för godkännande av begärda kvantiteter. I de fall då procentandelen är lägre än 5 % får kommissionen avslå ansökningarna; säkerheten skall frisläppas omedelbart.
7. Aktören kan dra tillbaka sin licensansökan inom tio arbetsdagar från det att den enhetliga procentsatsen för godkännande har offentliggjorts i Europeiska unionens officiella tidning, om tillämpning av denna procentsats leder till fastställandet av en kvantitet som är mindre än 20 ton för grupp G 2 och mindre än ett ton för de övriga grupperna. Medlemsstaterna skall inom fem dagar underrätta kommissionen om att licensansökan dragits tillbaka och skall omedelbart frisläppa säkerheten.
8. Kommissionen skall fastställa den resterande kvantitet som skall överföras till den tillgängliga kvantiteten för efterföljande period inom den tidsfrist som anges i artikel 1.
9. Licenserna skall utfärdas snarast möjligt efter det att kommissionen fattat sitt beslut.
10. Licenserna får inte användas för andra produkter än sådana som uppfyller samtliga gällande hygienkrav inom gemenskapen.
11. Före slutet av den fjärde månaden efter varje årlig period, från 1 juli till 30 juni, skall medlemsstaterna till kommissionen anmäla de kvantiteter som faktiskt importerats under perioden i fråga enligt denna förordning.
Alla anmälningar, även anmälningar om att inget har importerats, skall ske enligt den modell som anges i bilaga IV.
Artikel 6
1. Vid tillämpningen av artikel 23.2 i förordning (EG) nr 1291/2000 skall importlicensernas giltighetstid vara 150 dagar från och med utfärdandedagen.
Licensernas giltighetstid får dock inte i något fall utsträckas till efter den 30 juni under utfärdandeåret.
2. De importlicenser som utfärdas i enlighet med denna förordning får inte överlåtas.
Artikel 7
Bestämmelserna i förordning (EG) nr 1291/2000 skall tillämpas utan att det påverkar bestämmelserna i den här förordningen.
Med undantag från artikel 8.4 i förordning (EG) nr 1291/2000 får den kvantitet som importeras i enlighet med den här förordningen inte överstiga den kvantitet som anges i fält 17 och 18 på importlicensen. För detta ändamål skall siffran %quot%0%quot% anges i fält 19 på licensen.
Artikel 8
Förordning (EG) nr 1486/95 skall upphöra att gälla.
Hänvisningar till den upphävda förordningen skall anses som hänvisningar till denna förordning och skall läsas enligt jämförelsetabellen i bilaga VI.
Artikel 9
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 2011/2003
av den 14 november 2003
om ändring av bilagorna I och III i rådets förordning (EEG) nr 2377/90 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2377/90 av den 26 juni 1990 om inrättandet av ett gemenskapsförfarande för att fastställa gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung(1), senast ändrad genom kommissionens förordning (EG) nr 1873/2003(2), särskilt artiklarna 6, 7 och 8 i denna, och
av följande skäl:
(1) I enlighet med förordning (EEG) nr 2377/90 måste gränsvärden för högsta tillåtna restmängder successivt fastställas för samtliga farmakologiskt verksamma substanser som används inom gemenskapen i veterinärmedicinska läkemedel som är avsedda att ges till livsmedelsproducerande djur.
(2) Gränsvärden bör fastställas först efter det att Kommittén för veterinärmedicinska läkemedel har granskat all relevant information beträffande säkerheten med restmängder av ämnet i fråga för den som konsumerar livsmedel med animaliskt ursprung samt restmängdernas påverkan på den industriella bearbetningen av livsmedel.
(3) Vid fastställandet av gränsvärden för högsta tillåtna restmängder av veterinärmedicinska läkemedel i livsmedel med animaliskt ursprung är det nödvändigt att ange de djurarter i vilka restmängder kan förekomma, vilka mängder som kan förekomma i var och en av de relevanta vävnaderna från det behandlade djuret (målvävnad) samt vilket slag av restmängd som är relevant vid övervakningen av restmängder (restmarkör).
(4) För kontroll av resthalter bör enligt tillämplig gemenskapslagstiftning gränsvärden vanligtvis fastställas för målvävnaderna lever eller njure. I den internationella handeln avlägsnas dock ofta lever och njure från slaktkroppen, och gränsvärden bör därför alltid fastställas även för muskel- eller fettvävnader.
(5) För veterinärmedicinska läkemedel som är avsedda för äggläggande fåglar, mjölkdjur eller honungsbin, måste gränsvärden även fastställas för ägg, mjölk eller honung.
(6) Alfacypermetrin och Metamizol skall införas i bilaga I till förordning (EEG) nr 2377/90.
(7) För att möjliggöra komplettering av vetenskapliga studier Foxim skall införas i bilaga III till förordning (EEG) nr 2377/90.
(8) En tillräckligt lång tidsfrist bör fastställas innan denna förordning träder i kraft så att medlemsstaterna kan göra de nödvändiga anpassningarna till bestämmelserna i denna förordning av tillstånden att släppa ut de berörda veterinärmedicinska läkemedlen på marknaden, vilka beviljats enligt Europaparlamentets och rådets direktiv 2001/82/EG(3).
(9) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för veterinärmedicinska läkemedel.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagorna I och III till förordning (EEG) nr 2377/90 skall ändras i enlighet med bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Den skall tillämpas från och med den sextionde dagen efter att den har offentliggjorts.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 2314/2003
av den 29 december 2003
om inledande av en stående anbudsinfordran för försäljning på gemenskapsmarknaden av råg som innehas av det tyska interventionsorganet
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 1766/92 av den 30 juni 1992 om den gemensamma organisationen av marknaden för spannmål(1), särskilt artikel 5 i denna, och
av följande skäl:
(1) I kommissionens förordning (EEG) nr 2131/93 av den 28 juli 1993 om förfarandet vid och villkoren för försäljning av spannmål som innehas av interventionsorgan(2), föreskrivs bland annat att det spannmål som innehas av interventionsorgan skall försäljas genom anbudsinfordran och enligt sådana prisförhållanden att marknadsstörningar undviks.
(2) Tyskland förfogar fortfarande över interventionslager av råg.
(3) På grund av svåra klimatförhållanden i en stor del av gemenskapen minskade spannmålsproduktionen kraftigt under regleringsåret 2003/2004. Denna situation har lokalt medfört högre priser, vilket orsakar särskilda problem för uppfödare och för foderindustrin, som får svårigheter att göra inköp till konkurrenskraftiga priser.
(4) De lager av råg som innehas av det tyska interventionsorganet bör göras tillgängliga för den inre marknaden. Tidsfristen för inlämnande av anbud för den sista delanbudsinfordran enligt förordning (EG) nr 1510/20033(3) upphörde att gälla den 18 december 2003; det är lämpligt att inleda en ny stående anbudsinfordran.
(5) För att få överblick över situationen på gemenskapsmarknaden är det lämpligt att kommissionen fastställer villkoren för anbudsinfordran. Dessutom bör en tilldelningskoefficient fastställas för de anbud som ligger på samma nivå som det lägsta försäljningspriset.
(6) Det är viktigt att bevara anbudsgivarnas anonymitet i det tyska interventionsorganets anmälan till kommissionen.
(7) För att modernisera hanteringen är det också lämpligt att föreskriva att de uppgifter som kommissionen behöver skall förmedlas via e-post.
(8) Förvaltningskommittén för spannmål har inte avgivit något yttrande inom den tid som dess ordförande har bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Det tyska interventionsorganet skall inleda försäljning genom stående anbudsinfordran på gemenskapens inre marknad av 1139000 ton råg som det förfogar över.
Artikel 2
Försäljningen enligt artikel 1 skall ske enligt villkoren i förordning (EEG) nr 2131/93.
Genom undantag från den förordningen skall emellertid
a) anbuden utformas på grundval av den faktiska kvaliteten hos det parti som anbudet avser,
b) lägsta försäljningspris fastställas på en sådan nivå att det inte orsakar störningar på marknaderna för spannmål.
Artikel 3
Genom undantag från artikel 13.4 i förordning (EEG) nr 2131/93 skall säkerheten för anbudet fastställas till 10 euro per ton.
Artikel 4
1. Tidsfristen för inlämnande av anbud för den första delanbudsinfordran är den 8 januari 2004, kl. 9.00 (lokal tid, Bryssel).
Tidsfristen för inlämnande av anbud för de följande omgångarna skall löpa ut varje torsdag kl. 9.00 (lokal tid, Bryssel), med undantag av den 8 april och den 20 maj 2004.
Tidsfristen för inlämnande av anbud för den sista delanbudsinfordran skall löpa ut den 27 maj 2004, kl. 9.00 (lokal tid, Bryssel).
2. Anbuden skall lämnas in till det tyska interventionsorganet: Bundesanstalt für Landwirtschaft und Ernährung (BLE) Adickesallee 40 D - 60322 Frankfurt am Main Fax (00-49) 691 56 49 62
Artikel 5
Det tyska interventionsorganet skall underrätta kommissionen om de inkomna anbuden senast två timmar efter det att tidsfristen för inlämnande av anbud löpt ut. Anbuden skall skickas med elektronisk post och med hjälp av formuläret i bilagan.
Artikel 6
Kommissionen skall enligt förfarandet i artikel 23 i förordning (EG) nr 1766/92 fastställa det lägsta försäljningspriset eller besluta att avvisa de inlämnade anbuden. I de fall där anbud avser samma parti och en total kvantitet som överskrider den disponibla kvantiteten får fastställandet ske separat för varje parti.
När det gäller anbud som ligger på samma nivå som det lägsta försäljningspriset får en tilldelningskoefficient fastställas för de kvantiteter för vilka anbud har lämnats.
Artikel 7
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens beslut
av den 11 februari 2004
om att inte uppta fention i bilaga I till rådets direktiv 91/414/EEG och om återkallande av godkännande för växtskyddsmedel som innehåller detta verksamma ämne
[delgivet med nr K(2004) 313]
(Text av betydelse för EES)
(2004/140/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande av växtskyddsmedel på marknaden(1), senast ändrat genom kommissionens direktiv 2003/119/EG(2), särskilt artikel 8.2 tredje och fjärde stycket i detta,
med beaktande av kommissionens förordning (EEG) nr 3600/92 av den 11 december 1992 om närmare bestämmelser för genomförandet av den första etappen i det arbetsprogram som avses i artikel 8.2 i rådets direktiv 91/414/EEG om utsläppande av växtskyddsprodukter på marknaden(3), senast ändrad genom förordning (EG) nr 2266/2000(4), särskilt artikel 7.3a b i denna, och
av följande skäl:
(1) Enligt artikel 8.2 i direktiv 91/414/EEG skall kommissionen påbörja ett arbetsprogram som syftar till att undersöka de verksamma ämnen som används i växtskyddsprodukter som redan fanns på marknaden den 25 juli 1993. I förordning (EEG) nr 3600/92 fastställs närmare bestämmelser för genomförandet av programmet.
(2) Genom kommissionens förordning (EG) nr 933/94 av den 27 april 1994 om fastställande av verksamma ämnen i växtskyddsmedel och om val av rapporterande medlemsstater för genomförandet av kommissionens förordning (EEG) nr 3600/92(5), senast ändrad genom förordning (EG) nr 2230/95(6), fastställdes de verksamma ämnen som skulle bedömas inom ramen för förordning (EEG) nr 3600/92, fastställdes en medlemsstat som skulle fungera som rapporterande medlemsstat när det gällde bedömningen av varje verksamt ämne och fastställdes det vilka producenter av varje verksamt ämne som hade lämnat in en anmälan inom tidsfristen.
(3) Fention är ett av de 89 verksamma ämnen som anges i förordning (EG) nr 933/94.
(4) I enlighet med artikel 7.1 c i förordning (EEG) nr 3600/92 överlämnade Grekland, som utsetts till rapporterande medlemsstat, den 4 april 1996 en rapport till kommissionen om sin utvärdering av de uppgifter som anmälarna överlämnat i enlighet med artikel 6.1 i den förordningen.
(5) Efter att ha mottagit rapporten från den rapporterande medlemsstaten inledde kommissionen samråd med både medlemsstaternas experter och huvudanmälaren Bayer CropScience, i enlighet med artikel 7.3 i förordning (EEG) nr 3600/92.
(6) Kommissionen anordnade två trepartsmöten med den huvudsaklige uppgiftslämnaren och den rapporterande medlemsstaten för detta verksamma ämne den 18 april 1997 och den 11 februari 2003.
(7) Medlemsstaterna och kommissionen har granskat Greklands utvärderingsrapport inom ramen för Ständiga kommittén för livsmedelskedjan och djurhälsa. Resultatet av denna granskning presenterades den 4 juli 2003 i form av en kommissionsrapport om fention.
(8) Dokumentationen och resultatet av granskningen överlämnades också till Vetenskapliga kommittén för växter. Kommittén ombads att göra ett utlåtande om upprättande av nivåer för acceptabelt dagligt intag och godtagbar användarexponering. Grundat på slutsatser från riskbedömningarna avseende människor och miljö ansåg kommittén i sitt första yttrande av den 2 oktober 1998 att det inte är möjligt att sammanställa en fullständig bedömning i avsaknad av bevis för att ens en begränsad användning som bete på oliv- och citrusfruktodlingar var säker för folkhälsan och miljön. Kommittén noterade särskilt den mycket höga akuta risken för fåglar. I det yttrandet medgav kommittén att utveckling av en innovativ teknik för tillämpning, nämligen en typ av bete som innefattar fention och lockmedel på endast en del av grödan, skulle kunna vara intressant när det gäller att uppnå begränsad exponering av människor och miljö. Kommittén noterade att särskilda studier skulle behövas av en sådan tillämpning innan någon färdig utvärdering skulle kunna göras. Ytterligare uppgifter, särskilt när det gäller användningen som bete, har senare lämnats in av Bayer CropScience och utvärderats. Dessa ytterligare uppgifter och deras utvärdering har överlämnats till Vetenskapliga kommittén för växter. I sitt yttrande av den 17 december 2002 drog kommittén slutsatsen att risken för fåglar av de föreslagna användningarna av fention fortfarande är oklar. Följaktligen förblir frågorna i det tidigare yttrandet avseende möjliga risker för fåglar obesvarade.
(9) Resultatet av de utvärderingar som har gjorts på grundval av inlämnade uppgifter har inte visat att de växtskyddsmedel som innehåller fention, med de förslagna användningsföreskrifterna, allmänt uppfyller de krav som anges i artikel 5.1 a och 5.1 b i direktiv 91/414/EEG, särskilt inte när det gäller dess möjliga effekter på fåglar.
(10) Fention bör därför inte upptas i bilaga I till direktiv 91/414/EEG.
(11) Åtgärder bör vidtas för att se till att befintliga godkännanden för växtskyddsmedel med fention dras tillbaka inom en föreskriven period och inte förnyas samt att inga nya godkännanden beviljas för sådana produkter.
(12) Mot bakgrund av uppgifter som inkommit till kommissionen tycks det som om det, i avsaknad av effektiva alternativ för vissa begränsade användningar i vissa medlemsstater, finns behov för vidare användning av det verksamma ämnet så att alternativ kan utvecklas. Det är under rådande omständigheter således motiverat att under strikta förhållanden i syfte att minimera riskerna föreskriva en förlängd period för tillbakadragande av gällande godkännanden för de begränsade användningar som anses av behövas då det för närvarande inte existerar några alternativ för bekämpning av skadliga organismer.
(13) En övergångsperiod under vilken kvarvarande lager av de växtskyddsmedel som innehåller fention som är tillåtna av medlemsstaterna får omhändertas, lagras, släppas ut på marknaden och användas, skall begränsas till högst tolv månader för att kvarvarande lager inte skall användas mer än under en ytterligare växtodlingssäsong.
(14) Detta beslut påverkar inte de eventuella åtgärder som kommissionen kan komma att vidta i ett senare skede avseende detta verksamma ämne, inom ramen för rådets direktiv 79/117/EEG av den 21 december 1978 om förbud mot att växtskyddsprodukter som innehåller vissa verksamma ämnen släpps ut på marknaden och används(7), senast ändrat genom förordning (EG) nr 807/2003(8).
(15) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Fention skall inte upptas som ett verksamt ämne i bilaga I till rådets direktiv 91/414/EEG.
Artikel 2
Medlemsstaterna skall säkerställa följande:
1. Godkännanden av växtskyddsmedel med fention skall dras in senast den 11 augusti 2004.
2. Från och med den 17 februari 2004 får inga godkännanden av växtskyddsmedel som innehåller fention beviljas eller förnyas enligt det undantag som anges i artikel 8.2 i direktiv 91/414/EEG.
3. När det gäller de användningar som anges i kolumn B i bilagan får medlemsstaterna i kolumn A behålla godkännanden för växtskyddsmedel med fention t.o.m. den 30 juni 2007 under följande förutsättningar:
a) Medlemsstaten ser till att sådana växtskyddsmedel som finns kvar på marknaden får en ny märkning som motsvarar de skärpta villkoren för användning.
b) Medlemsstaten vidtar alla lämpliga lindrande åtgärder för att minska eventuella risker för att sörja för att människors och djurs hälsa samt miljön är väl skyddade.
c) Medlemsstaten skall se till att seriösa försök görs för att finna alternativa produkter eller metoder för sådana användningar, med hjälp av handlingsplaner.
Den berörda medlemsstaten skall underrätta kommissionen senast den 31 december 2004 om tillämpning av denna punkt och i synnerhet om åtgärder som vidtagits i enlighet med leden a-c, och varje år översända uppskattningar om hur mycket fention som använts i enlighet med den här artikeln.
Artikel 3
Alla anstånd som beviljas av medlemsstaterna i enlighet med artikel 4.6 i direktiv 91/414/EEG skall vara så korta som möjligt och får
a) för de användningar vilkas godkännanden skall återkallas senast den 11 augusti 2004, inte gälla längre än till och med den 11 augusti 2005,
b) för de användningar vilkas godkännanden skall återkallas senast den 30 juni 2007, inte gälla längre än till och med den 31 december 2007.
Artikel 4
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 18 november 2004
om tillåtelse för Slovakien att tillämpa det undantag som anges i artikel 3.2 i rådets direktiv 92/102/EEG om identifikation och registrering av djur
(delgivet med nr K(2004) 4382)
(Endast den slovakiska texten är giltig)
(Text av betydelse för EES)
(2004/775/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 92/102/EEG av den 27 november 1992 om identifikation och registrering av djur [1], särskilt artikel 3.2 i detta, och
av följande skäl:
(1) Enligt artikel 3.2 i direktiv 92/102/EEG kan medlemsstaterna få tillstånd att från den förteckning som avses i artikel 3.1 i direktivet undanta jordbruksföretag som håller högst tre får eller getter, för vilka de inte gör anspråk på särskilt stöd, eller ett svin, om dessa djur är avsedda för egen användning eller konsumtion, under förutsättning att djuren före eventuell flyttning underkastas de kontroller som beslutas om i direktivet.
(2) De slovakiska myndigheterna har begärt att tillståndet skall gälla till och med slutet av juni 2005 och har lämnat lämpliga garantier för veterinärmedicinska kontroller.
(3) Slovakien bör därför få tillstånd att tillämpa undantaget till och med den 30 juni 2005.
(4) De åtgärder som anges i detta beslut är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Slovakien ges härmed tillstånd att tillämpa det undantag som anges i artikel 3.2 i direktiv 92/102/EEG.
Artikel 2
Detta beslut skall tillämpas till och med den 30 juni 2005 och riktar sig till Republiken Slovakien.
Kommissionens beslut
av den 9 november 2004
om fastställelse av formulär för ansökningar om rättshjälp enligt rådets direktiv 2003/8/EG om förbättring av möjligheterna till rättslig prövning i gränsöverskridande tvister genom fastställande av gemensamma minimiregler för rättshjälp i sådana tvister
(delgivet med nr K(2004) 4285)
(2004/844/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 2003/8/EG av den 27 januari 2003 om förbättring av möjligheterna till rättslig prövning i gränsöverskridande tvister genom fastställande av gemensamma minimiregler för rättshjälp i sådana tvister [1], särskilt artikel 16.1 i detta,
efter samråd med den rådgivande kommitté som upprättats enligt artikel 17.1 i direktiv 2003/8/EG, och
av följande skäl:
(1) I artikel 16.1 i direktiv 2003/8/EG föreskrivs att kommissionen skall fastställa ett standardformulär för ansökningar om rättshjälp och för översändande av sådana ansökningar.
(2) Standardformuläret för översändande av ansökningar om rättshjälp mellan medlemsstaternas rättsliga myndigheter har fastställts genom kommissionens beslut K(2004) 1829 [2].
(3) Själva standardformuläret för ansökningar om rättshjälp skall, i kraft av artikel 16.2 andra stycket i direktiv 2003/8/EG, utarbetas senast den 30 november 2004. Formuläret bör följaktligen fastställas genom detta beslut.
(4) I överensstämmelse med artiklarna 1 och 2 i det protokoll om Danmarks ställning som är fogat till Fördraget om Europeiska unionen och Fördraget om upprättandet a
Rådets beslut
av den 25 oktober 2004
om ingående av ett avtal genom skriftväxling mellan Europeiska gemenskapen och Konungariket Norge om protokoll 2 till det bilaterala frihandelsavtalet mellan Europeiska ekonomiska gemenskapen och Konungariket Norge
(Text av betydelse för EES)
(2004/859/EG)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 133 jämförd med artikel 300.2 första meningen i första stycket i detta,
med beaktande av kommissionens förslag, och
av följande skäl:
(1) I protokoll 2 till det bilaterala frihandelsavtalet mellan Europeiska ekonomiska gemenskapen och Konungariket Norge [1], å ena sidan, och protokoll 3 till EES-avtalet, ändrat genom Gemensamma EES-kommitténs beslut nr 140/2001 [2], å andra sidan, fastställs handelsordningen mellan avtalsparterna när det gäller vissa jordbruksprodukter och bearbetade jordbruksprodukter.
(2) När beslut nr 140/2001 antogs förklarade Europeiska gemenskapen och Norge i ett gemensamt uttalande att den icke-jordbruksrelaterade delen av tullen på produkterna i tabell I i protokoll 3 skulle tas bort. På grundval av detta avslutades diskussionerna mellan tjänstemän från kommissionen och Norge den 11 mars 2004. De nya tullmedgivandena kommer att genomföras genom ett beslut av Gemensamma EES-kommittén om ändring av protokoll 3 till EES-avtalet.
(3) Ett avtal genom skriftväxling mellan Europeiska gemenskapen och Konungariket Norge om protokoll 2 till det bilaterala frihandelsavtalet mellan Europeiska ekonomiska gemenskapen och Konungariket Norge har också förhandlats fram för att beakta resultaten av dessa diskussioner.
(4) De åtgärder som är nödvändiga för att genomföra detta beslut bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter [3].
(5) Avtalet bör godkännas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Avtalet genom skriftväxling mellan Europeiska gemenskapen och Konungariket Norge om protokoll 2 till det bilaterala frihandelsavtalet mellan Europeiska ekonomiska gemenskapen och Konungariket Norge godkänns härmed på gemenskapens vägnar.
Texten till avtalet åtföljer detta beslut.
Artikel 2
Rådets ordförande bemyndigas att utse den person som skall ha rätt att underteckna det avtal med bindande verkan för gemenskapen.
Artikel 3
De åtgärder som är nödvändiga för att genomföra detta beslut skall antas i enlighet med förfarandet i artikel 4.2.
Artikel 4
1. Kommissionen skall biträdas av den förvaltningskommitté för övergripande frågor rörande handel med bearbetade jordbruksprodukter som avses i artikel 16 i rådets förordning (EG) nr 3448/93 [4] (nedan kallad "kommittén").
2. När det hänvisas till denna punkt skall artiklarna 4 och 7 i beslut 1999/468/EG tillämpas.
Den tid som avses i artikel 4.3 i beslutet skall fastställas till en månad.
3. Kommittén skall själv anta sin arbetsordning.
Rådets rekommendation
av den 14 oktober 2004
om genomförandet av medlemsstaternas sysselsättningspolitik
(2004/741/EG)
EUROPEISKA UNIONENS RÅD UTFÄRDAR DENNA REKOMMENDATION
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 128.4 i detta,
med beaktande av kommissionens rekommendation,
med beaktande av Sysselsättningskommitténs yttrande, och
av följande skäl:
(1) Den europeiska sysselsättningsstrategin är central för genomförandet av sysselsättnings- och arbetsmarknadsmålen i Lissabonstrategin. För att Lissabonagendan skall kunna genomföras framgångsrikt måste medlemsstaternas sysselsättningspolitik på ett balanserat sätt främja tre mål som kompletterar och ömsesidigt stödjer varandra, nämligen full sysselsättning, kvalitet och produktivitet i arbetet samt social sammanhållning och integration. För att dessa mål skall uppnås krävs ytterligare strukturreformer som inriktas på tio specifika prioriteringsområden samt bättre styrelseformer.
(2) Genom den reformerade europeiska sysselsättningsstrategin från 2003 har tonvikten lagts vid ett perspektiv på medellång sikt och vid betydelsen av att alla politiska åtgärder som rekommenderas i riktlinjerna för sysselsättningen genomförs. En komplett översyn av riktlinjerna för sysselsättningen bör därför endast göras vart tredje år. Under de mellanliggande åren bör de bara uppdateras i mycket begränsad omfattning.
(3) Rådet antog utan ändringar riktlinjerna för medlemsstaternas sysselsättningspolitik 2004 genom beslut 2004/740/EG [1].
(4) Rådet antog den 22 juli 2003 en rekommendation om genomförandet av medlemsstaternas sysselsättningspolitik [2]. Genomgången av medlemsstaternas nationella handlingsplaner för sysselsättning i den gemensamma rapporten om sysselsättningen 2003-2004 visar att medlemsstaterna och arbetsmarknadens parter bara i begränsad utsträckning har följt dessa rekommendationer från rådet.
(5) Den europeiska specialgruppen för sysselsättningsfrågor har rekommenderat att EU bör skärpa rekommendationerna till medlemsstaterna. Framför allt bör åtgärder vidtas för att öka anpassningsförmågan hos arbetstagare och företag, förmå fler människor att komma in och stanna kvar på arbetsmarknaden och se till att arbete lönar sig för alla, få till stånd fler och bättre riktade investeringar i humankapital och livslångt lärande, samt säkerställa ett effektivt genomförande av reformer genom bättre styrelseformer. Rådet och kommissionen delar denna bedömning och har integrerat de politiska budskap som framförs i specialgruppens rapport i den gemensamma rapporten om sysselsättningen.
(6) Analysen av genomförandet av riktlinjerna och rådets rekommendationer från 2003 i den gemensamma rapporten om sysselsättningen samt de generella och landspecifika politiska budskapen i rapporten från specialgruppen för sysselsättningsfrågor ligger till grund för EU:s rekommendationer till nationell sysselsättningspolitik 2004.
(7) Riktlinjerna för sysselsättningen gäller de nya medlemsstaterna sedan anslutningen. Alla nya medlemsstater har under de senaste åren avlagt rapport om genomförandet av de gemensamma utvärderingarna avseende riktlinjerna för sysselsättningen. De flesta nya medlemsstater måste tillsammans med arbetsmarknadens parter intensifiera sitt arbete med att modernisera sysselsättningspolitiken för att den pågående omstruktureringen av deras ekonomier skall kunna genomföras fullt ut. Det är mycket viktigt att det skapas en ny balans mellan flexibilitet och trygghet samt att öka sysselsättningen och investeringarna i humankapital genom ett livslångt lärande. Arbetskraftens hälsa måste också förbättras. För att uppnå en fullständig och effektiv användning a
Rådets direktiv 2004/113/EG
av den 13 december 2004
om genomförande av principen om likabehandling av kvinnor och män när det gäller tillgång till och tillhandahållande av varor och tjänster
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 13.1,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande [1],
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande [2],
med beaktande av Regionkommitténs yttrande [3], och
av följande skäl:
(1) Enligt artikel 6 i fördraget om Europeiska unionen bygger unionen på principerna om frihet, demokrati och respekt för de mänskliga rättigheterna och de grundläggande friheterna och på rättsstatsprincipen, vilka principer är gemensamma för medlemsstaterna, och unionen skall som allmänna principer för gemenskapsrätten respektera de grundläggande rättigheterna, såsom de garanteras i Europeiska konventionen om skydd för de mänskliga rättigheterna och de grundläggande friheterna och såsom de följer av medlemsstaternas gemensamma konstitutionella traditioner.
(2) Rätten till likställdhet inför lagen och skydd mot diskriminering för alla och envar är grundläggande rättigheter som erkänns i den allmänna förklaringen om de mänskliga rättigheterna, i FN:s konvention om avskaffandet av all slags diskriminering av kvinnor, i den internationella konventionen om avskaffandet av alla former av rasdiskriminering samt i FN:s konventioner om medborgerliga och politiska rättigheter och om ekonomiska, sociala och kulturella rättigheter samt genom Europeiska konventionen om skydd för de mänskliga rättigheterna och de grundläggande friheterna, vilka har undertecknats av alla medlemsstater.
(3) Samtidigt som diskriminering förbjuds är det viktigt att andra grundläggande fri- och rättigheter respekteras, bland annat skyddet för privat- och familjeliv och transaktioner som utförs i det sammanhanget samt religionsfrihet.
(4) Jämställdhet mellan kvinnor och män är en grundläggande princip för Europeiska unionen. Artiklarna 21 och 23 i Europeiska unionens stadga om de grundläggande rättigheterna förbjuder all könsdiskriminering och föreskriver att jämställdhet mellan kvinnor och män skall säkerställas på alla områden.
(5) Enligt artikel 2 i Fördraget om upprättandet av Europeiska gemenskapen är det en av gemenskapens grundläggande uppgifter att främja sådan jämställdhet. I artikel 3.2 i fördraget föreskrivs också att gemenskapen i all verksamhet skall syfta till att undanröja bristande jämställdhet mellan kvinnor och män och att främja jämställdhet mellan dem.
(6) Kommissionen aviserade i sitt meddelande om den socialpolitiska agendan att den hade för avsikt att lägga fram ett förslag till direktiv mot könsdiskriminering på områden utanför arbetsmarknaden. Ett sådant förslag är helt i enlighet med rådets beslut 2001/51/EG av den 20 december 2000 om inrättande av gemenskapens handlingsprogram avseende gemenskapens strategi för jämställdhet mellan kvinnor och män (2001–2005) [4], som omfattar samtliga av gemenskapens politikområden och syftar till att främja jämställdhet mellan kvinnor och män genom en anpassning av dessa politikområden och vidtagande av konkreta åtgärder för att förbättra situationen för kvinnor och män i samhället.
(7) Europeiska rådet uppmanade vid sitt möte i Nice den 7 och 9 december 2000 kommissionen att förstärka rättigheterna i fråga om likabehandling genom att anta ett förslag till direktiv för att främja jämställdhet mellan kvinnor och män inom andra områden än sysselsättning och yrkesverksamhet.
(8) Gemenskapen har antagit en rad rättsinstrument för att förebygga och motverka könsdiskriminering på arbetsmarknaden. Dessa instrument har visat hur viktig lagstiftning är för kampen mot diskriminering.
(9) Könsdiskriminering, inklusive trakasserier och sexuella trakasserier, förekommer även på andra områden än arbetsmarknaden. Denna diskriminering kan få lika stora negativa konsekvenser och hindra kvinnor och män från att i full utsträckning integreras väl i det ekonomiska och sociala livet.
(10) Dessa problem är särskilt tydliga när det gäller tillgång till och tillhandahållande av varor och tjänster. Könsdiskriminering bör därför förhindras och undanröjas på detta område. Precis som i fråga om rådets direktiv 2000/43/EG av den 29 juni 2000 om genomförandet av principen om likabehandling av personer oavsett deras ras eller etniska ursprung [5] kan detta mål uppnås bättre med hjälp av gemenskapslagstiftning.
(11) Sådan lagstiftning bör förbjuda könsdiskriminering när det gäller tillgång till och tillhandahållande av varor och tjänster. Med varor bör avses varor enligt bestämmelserna i fördraget om upprättandet av Europeiska gemenskapen i fråga om fri rörlighet för varor. Med tjänster bör avses tjänster enligt artikel 50 i det fördraget.
(12) För att förhindra diskriminering på grund av kön bör detta direktiv tillämpas på såväl direkt som indirekt diskriminering. Direkt diskriminering uppstår endast då en person på grund av kön behandlas sämre än en annan person i en jämförbar situation. Olika behandling av kvinnor och män när det gäller hälso- och sjukvård som grundar sig på fysiska skillnader mellan könen, till exempel, gäller inte jämförbara situationer och utgör därför inte diskriminering.
(13) Diskrimineringsförbudet bör gälla personer som tillhandahåller varor och tjänster som är tillgängliga för allmänheten och som erbjuds utanför området för privat- och familjeliv och transaktioner i samband med detta. Det bör inte gälla medie- och reklaminnehåll och inte heller offentlig eller privat utbildning.
(14) Alla individer har rätt att fritt sluta avtal inbegripet rätt att välja avtalspart för en transaktion. En individ som tillhandahåller varor eller tjänster kan ha ett antal subjektiva skäl till val av avtalspart. Så länge som valet av avtalspart inte grundar sig på denna persons kön bör inte detta direktiv påverka individens frihet att välja avtalspart.
(15) Det finns redan ett antal rättsliga instrument för genomförande av principen om likabehandling mellan kvinnor och män när det gäller frågor som rör arbetslivet. Detta direktiv bör därför inte gälla frågor som rör detta område. Samma princip gäller för egenföretagande i den mån detta omfattas av befintliga rättsliga instrument. Direktivet bör endast gälla försäkringar och pensioner som är privata, frivilliga och åtskilda från anställningsförhållandet.
(16) Skillnader i behandling kan endast godtas om de motiveras av ett berättigat syfte. Ett berättigat syfte kan till exempel vara skydd av offer för könsrelaterat våld (som vid upprättande av skyddat boende för enbart det ena könet), skäl som rör privatliv och anständighet (som då en person upplåter en bostad i en del av sitt hem), främjande av jämställdhet eller kvinnors eller mäns intressen (till exempel frivilligorganisationer för enbart det ena könet), föreningsfrihet (som medlemskap i privata klubbar för enbart det ena könet) samt anordnande av idrottsaktiviteter (som idrottsarrangemang för enbart det ena könet). Varje begränsning bör dock vara lämplig och nödvändig i enlighet med de kriterier som härrör ur Europeiska gemenskapernas domstols praxis.
(17) Principen om likabehandling beträffande tillgång till varor och tjänster innebär inte något krav på att kvinnor och män alltid skall erbjudas varor och tjänster på samma sätt, under förutsättning att de inte tillhandahålls på ett fördelaktigare sätt till det ena könet.
(18) Användningen av könsspecifika försäkringstekniska faktorer är utbredd i samband med att försäkringstjänster och andra liknande finansiella tjänster tillhandahålls. För att säkra likabehandling av kvinnor och män bör användningen av kön som en försäkringsteknisk faktor inte leda till skillnader i enskildas premier och ersättningar. För att marknaden inte skall utsättas för alltför plötsliga förändringar bör genomförandet av denna regel endast gälla nya avtal som ingås efter utsatt tidsfrist för införlivande av detta direktiv.
(19) Vissa riskkategorier kan variera mellan könen. I vissa fall är kön en men inte nödvändigtvis den enda avgörande faktorn vid bedömningen av de försäkrade riskerna. Beträffande avtal för försäkring av dessa risktyper får medlemsstaterna besluta att tillåta undantag från regeln om könsneutrala premier och ersättningar så länge de kan garantera att de bakomliggande försäkringstekniska och statistiska uppgifter som utgör grund för beräkningarna är tillförlitliga, regelbundet uppdateras och är tillgängliga för allmänheten. Undantag medges endast om den könsneutrala regeln inte redan tillämpas i den nationella lagstiftningen. Fem år efter införlivandet av detta direktiv bör medlemsstaterna på nytt granska motiveringen till dessa undantag med beaktande av de senaste försäkringstekniska och statistiska uppgifterna och en rapport från kommissionen tre år efter tidpunkten för införlivandet av detta direktiv.
(20) Mindre förmånlig behandling av kvinnor på grund av graviditet och moderskap bör anses vara en form av direkt könsdiskriminering och följaktligen förbjuden i försäkringstjänster och liknande finansiella tjänster. Kostnader som har samband med risk för graviditet och moderskap bör därför inte läggas på enbart de som tillhör det ena könet.
(21) Personer som har utsatts för könsdiskriminering bör tillförsäkras ett lämpligt rättsligt skydd. För att ett effektivare skydd skall tillhandahållas bör föreningar, organisationer och andra rättsliga enheter också ges befogenhet att, på det sätt medlemsstaterna bestämmer, engagera sig, antingen på den utsatta personens vägnar eller för att stödja denne, utan att detta påverkar tillämpningen av de nationella regler som rör ombud och försvar vid domstol.
(22) För att principen om likabehandling skall kunna tillämpas effektivt bör reglerna om bevisbördan anpassas på så sätt att bevisbördan övergår till svaranden när det föreligger ett prima facie-fall av diskriminering.
(23) För att principen om likabehandling skall kunna genomföras i praktiken krävs ett lämpligt rättsligt skydd mot repressalier.
(24) Medlemsstaterna bör i syfte att främja principen om likabehandling uppmuntra dialogen med berörda intressenter som i enlighet med nationell lagstiftning och praxis har ett berättigat intresse av att bidra till att motverka könsdiskriminering när det gäller tillgång till och tillhandahållande av varor och tjänster.
(25) Skyddet mot könsdiskriminering bör stärkas genom att det i varje medlemsstat finns ett eller flera organ med behörighet att analysera problemen, undersöka tänkbara lösningar och ge praktiskt stöd till människor som utsätts för diskriminering. Dessa organ kan vara desamma som de som på nationell nivå har till uppgift att tillvarata de mänskliga rättigheterna eller enskildas rättigheter eller som har till uppgift att genomföra principen om likabehandling.
(26) I detta direktiv fastställs minimikrav, vilket ger medlemsstaterna möjlighet att behålla eller införa mer förmånliga bestämmelser. Genomförandet av detta direktiv bör inte åberopas som skäl till inskränkningar i det skydd som för närvarande finns i varje medlemsstat.
(27) Medlemsstaterna bör föreskriva effektiva, proportionerliga och avskräckande påföljder för åsidosättande av skyldigheterna enligt detta direktiv.
(28) Eftersom målen för detta direktiv, nämligen att säkra en enhetlig och hög nivå av skydd mot diskriminering i alla medlemsstater, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna och de därför, på grund av den planerade åtgärdens omfattning och verkningar, bättre kan uppnås på gemenskapsnivå, får gemenskapen enligt subsidiaritetsprincipen i artikel 5 i fördraget vidta åtgärder. I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå dessa mål.
(29) I enlighet med punkt 34 i det interinstitutionella avtalet om bättre lagstiftning [6] uppmanas medlemsstaterna att för egen del och i gemenskapens intresse upprätta egna tabeller som så vitt det är möjligt visar överensstämmelsen mellan direktivet och införlivandeåtgärderna samt att offentliggöra dessa tabeller.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
KAPITEL I
ALLMÄNNA BESTÄMMELSER
Artikel 1
Syfte
Syftet med detta direktiv är att fastställa en ram för bekämpning av könsdiskriminering när det gäller tillgång till och tillhandahållande av varor och tjänster, för att i medlemsstaterna genomföra principen om likabehandling av kvinnor och män.
Artikel 2
Definitioner
I detta direktiv avses med
a)direkt diskriminering när en person på grund av kön behandlas mindre förmånligt än en annan person behandlas, har behandlats eller skulle ha behandlats i en jämförbar situation,b)indirekt diskrimineringnär en skenbart neutral bestämmelse eller ett skenbart neutralt kriterium eller förfaringssätt särskilt missgynnar personer av ett visst kön jämfört med personer av det andra könet, om inte bestämmelsen, kriteriet eller förfaringssättet objektivt kan motiveras av ett berättigat mål och medlen för att uppnå detta mål är lämpliga och nödvändiga,c)trakasseriernär ett oönskat beteende som har samband med en persons kön syftar till eller leder till att en persons värdighet kränks och att en hotfull, fientlig, förnedrande, förödmjukande eller kränkande stämning skapas,d)sexuella trakasseriernär ett oönskat beteende av sexuell natur, som tar sig fysiska, verbala eller icke-verbala uttryck, syftar till eller leder till att en persons värdighet kränks, särskilt då en hotfull, fientlig, förnedrande, förödmjukande eller kränkande stämning skapas.
Artikel 3
Tillämpningsområde
1. Inom ramen för gemenskapens befogenheter skall detta direktiv tillämpas på alla personer som tillhandahåller varor och tjänster som är tillgängliga för allmänheten oberoende av den berörda personen, såväl inom den offentliga som den privata sektorn, inklusive offentliga organ, och som erbjuds utanför området för privat- och familjeliv och transaktioner som utförs i det sammanhanget.
2. Detta direktiv påverkar inte individens frihet att välja avtalspart så länge som valet inte grundar sig på avtalspartens kön.
3. Detta direktiv skall inte gälla medie- och reklaminnehåll eller utbildning.
4. Detta direktiv skall inte gälla frågor som rör arbetslivet, inklusive verksamhet som egenföretagare, i den utsträckning dessa frågor omfattas av andra rättsakter i gemenskapslagstiftningen.
Artikel 4
Principen om likabehandling
1. I detta direktiv skall principen om likabehandling av kvinnor och män innebära att
a) ingen direkt könsdiskriminering får förekomma, inklusive mindre förmånlig behandling av kvinnor på grund av graviditet och moderskap,
b) ingen indirekt könsdiskriminering får förekomma.
2. Detta direktiv skall inte påverka tillämpningen av förmånligare bestämmelser om skydd av kvinnor i samband med graviditet och moderskap.
3. Trakasserier och sexuella trakasserier i den mening som avses i detta direktiv skall anses vara könsdiskriminering och skall därför förbjudas. Det förhållandet att en person avvisar eller låter bli att reagera mot ett sådant beteende får inte ligga till grund för ett beslut som gäller denna person.
4. En instruktion att direkt eller indirekt diskriminera personer på grund av kön skall anses vara diskriminering enligt detta direktiv.
5. Detta direktiv utesluter inte skillnader i behandling, om tillhandahållandet av varor och tjänster uteslutande eller främst till personer av ett kön motiveras av ett berättigat mål och medlen för att uppnå detta mål är lämpliga och nödvändiga.
Artikel 5
Försäkringstekniska faktorer
1. Medlemsstaterna skall se till att i alla nya kontrakt som ingås senast efter den 21 december 2007, användningen av kön som en faktor vid beräkningen av premier och ersättningar i samband med försäkringar och därmed sammanhängande finansiella tjänster inte resulterar i att skillnader uppstår i enskilda personers premier och ersättningar.
2. Trots vad som anges i punkt 1, får medlemsstaterna besluta att före den 21 december 2007 tillåta proportionerliga skillnader i enskildas personers premier och ersättningar om användningen av kön är en avgörande faktor vid en riskbedömning som grundas på relevanta och korrekta försäkringstekniska och statistiska uppgifter. Berörda medlemsstater skall underrätta kommissionen och se till att korrekta uppgifter som är relevanta för användningen av kön som en avgörande försäkringsteknisk faktor sammanställs, offentliggörs och regelbundet uppdateras. Dessa medlemsstater skall se över sitt beslut fem år efter den 21 december 2007 med beaktande av den rapport från kommissionen som nämns i artikel 16, och skall översända resultaten av denna översyn till kommissionen.
3. Kostnader som har samband med graviditet och moderskap skall i inget fall leda till skillnader i enskilda personers premier och ersättningar.
Medlemsstaterna får skjuta upp genomförandet av de åtgärder som krävs för att följa denna punkt i högst två år efter den 21 december 2007. I sådana fall skall den berörda medlemsstaten omedelbart underrätta kommissionen.
Artikel 6
Positiv särbehandling
I syfte att säkerställa full jämställdhet mellan kvinnor och män i praktiken får principen om likabehandling inte hindra en medlemsstat från att behålla eller besluta om särskilda åtgärder för att förhindra eller kompensera könsrelaterat missgynnande.
Artikel 7
Minimikrav
1. Medlemsstaterna får införa eller behålla bestämmelser som är mer fördelaktiga när det gäller att upprätthålla principen om likabehandling mellan kvinnor och män än de som anges i detta direktiv.
2. Genomförandet av detta direktiv får under inga omständigheter utgöra skäl för att inskränka det skydd mot diskriminering som redan finns i medlemsstaterna på de områden som omfattas av detta direktiv.
KAPITEL II
RÄTTSMEDEL OCH SÄKERSTÄLLANDE AV EFTERLEVNADEN AV BESTÄMMELSERNA
Artikel 8
Tillvaratagande av rättigheter
1. Medlemsstaterna skall säkerställa att alla som anser sig förfördelade på grund av att principen om likabehandling inte har tillämpats på dem har tillgång till rättsliga och/eller administrativa förfaranden, inbegripet, när de anser det lämpligt, förlikningsförfaranden, för att säkerställa efterlevnaden av skyldigheterna enligt detta direktiv, även efter det att den situation i vilken diskrimineringen uppges ha förekommit har upphört.
2. Medlemsstaterna skall i sina nationella rättsordningar införa nödvändiga bestämmelser för att säkerställa en faktisk och effektiv kompensation eller gottgörelse, enligt vad medlemsstaterna bestämmer, för den förlust och skada som lidits av den person som drabbats av diskriminering i den mening som avses i detta direktiv, på ett sätt som är avskräckande och står i proportion till den skada som lidits. En på förhand fastställd övre gräns får inte begränsa denna gottgörelse eller kompensation.
3. Medlemsstaterna skall säkerställa att föreningar, organisationer eller andra juridiska personer, som i enlighet med de kriterier som fastställs i deras nationella lagstiftning har ett berättigat intresse av att säkerställa att bestämmelserna i detta direktiv efterlevs får, på den klagande personens vägnar eller för att stödja denne och med hans eller hennes tillstånd engagera sig i de rättsliga och/eller administrativa förfaranden som finns för att säkerställa efterlevnaden av skyldigheterna enligt detta direktiv.
4. Punkterna 1 och 3 påverkar inte tillämpningen av nationella regler om tidsfrister för att väcka talan som rör principen om likabehandling.
Artikel 9
Bevisbörda
1. Medlemsstaterna skall, i enlighet med sina nationella rättssystem, vidta nödvändiga åtgärder för att säkerställa att det, när personer, som anser sig kränkta genom att principen om likabehandling inte har tillämpats på dem, inför domstol eller annan behörig myndighet lägger fram fakta som ger anledning att anta att det har förekommit direkt eller indirekt diskriminering, skall åligga svaranden att bevisa att det inte föreligger något brott mot principen om likabehandling.
2. Punkt 1 skall inte hindra att medlemsstaterna inför bevisregler som är fördelaktigare för käranden.
3. Punkt 1 skall inte tillämpas på straffrättsliga förfaranden.
4. Punkterna 1, 2 och 3 skall också tillämpas på förfaranden som inleds enligt artikel 8.3.
5. Medlemsstaterna kan avstå från att tillämpa punkt 1 på förfaranden där det åligger domstolen eller annan behörig myndighet att utreda fakta i målet.
Artikel 10
Repressalier
Medlemsstaterna skall i sina rättsordningar införa nödvändiga bestämmelser för att skydda personer mot ogynnsam behandling eller ogynnsamma följder på grund av klagomål eller rättsliga förfaranden som syftar till att se till att principen om likabehandling följs.
Artikel 11
Dialog med berörda intressenter
Medlemsstaterna skall i syfte att främja principen om likabehandling främja en dialog med berörda intressenter som i enlighet med nationella lagar och praxis har ett berättigat intresse av att motverka könsdiskriminering när det gäller tillgången till och tillhandahållande av varor och tjänster.
KAPITEL III
ORGAN FÖR FRÄMJANDE AV LIKABEHANDLING
Artikel 12
1. Medlemsstaterna skall utse och genomföra de nödvändiga förberedelserna för ett eller flera organ för främjande, analys och kontroll av samt till stöd för likabehandling av alla personer utan åtskillnad på grund av kön. Dessa organ får utgöra en del av myndigheter som på nationell nivå har till uppgift att tillvarata de mänskliga rättigheterna eller enskildas rättigheter eller att genomföra principen om likabehandling.
2. Medlemsstaterna skall säkerställa att behörigheten för de organ som avses i punkt 1 omfattar följande:
a) Att på ett oberoende sätt bistå personer som utsatts för diskriminering genom att driva klagomål om diskriminering, utan att det påverkar de rättigheter för personer som har blivit diskriminerade eller för föreningar, organisationer eller andra rättsliga enheter som avses i artikel 8.3.
b) Att genomföra oberoende undersökningar om diskriminering.
c) Att offentliggöra oberoende rapporter om och lämna rekommendationer i frågor som rör sådan diskriminering.
KAPITEL IV
SLUTBESTÄMMELSER
Artikel 13
Efterlevnad
Medlemsstaterna skall vidta nödvändiga åtgärder för att säkerställa att principen om likabehandling respekteras när det gäller tillgång till och tillhandahållande av varor och tjänster inom tillämpningsområdet för detta direktiv och i synnerhet att
a) lagar och andra författningar som strider mot principen om likabehandling upphävs,
b) avtalsbestämmelser, interna regler för företag och regler för vinstdrivande eller icke-vinstdrivande föreningar som strider mot principen om likabehandling, förklaras eller kan förklaras ogiltiga eller ändras.
Artikel 14
Påföljder
Medlemsstaterna skall föreskriva påföljder för överträdelser av nationella bestämmelser som har utfärdats enligt detta direktiv och skall vidta de åtgärder som krävs för att se till att dessa sanktioner tillämpas. Påföljderna, som kan bestå av skadestånd till den utsatta personen, skall vara effektiva, proportionerliga och avskräckande. Medlemsstaterna skall anmäla dessa bestämmelser till kommissionen senast den 21 december 2007, och alla senare ändringar som gäller dem så snart som möjligt.
Artikel 15
Informationsspridning
Medlemsstaterna skall se till att på lämpligt sätt och på hela sitt territorium informera berörda personer om de bestämmelser som antas enligt detta direktiv och om relevanta bestämmelser som redan gäller.
Artikel 16
Rapporter
1. Medlemsstaterna skall senast den 21 december 2009, och därefter vart femte år, till kommissionen lämna över all tillgänglig information om tillämpningen av detta direktiv.
Kommissionen skall utarbeta en sammanfattande rapport som skall innefatta en översikt över medlemsstaternas nuvarande förfaranden med avseende på artikel 4 när det gäller kön som en faktor vid beräkningen av premier och ersättningar. Den skall lägga fram denna rapport för Europaparlamentet och rådet senast den 21 december 2010. Vid behov skall kommissionen till sin rapport foga förslag till ändring av direktivet.
2. Kommissionen skall i sin rapport ta hänsyn till synpunkter från berörda intressenter.
Artikel 17
Införlivande
1. Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 21 december 2007. De skall genast överlämna texterna till dessa bestämmelser till kommissionen.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texten till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 18
Ikraftträdande
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska unionens officiella tidning.
Artikel 19
Adressater
Detta direktiv riktar sig till medlemsstaterna.
Kommissionens förordning (EG) nr 50/2004
av den 9 januari 2004
om ändring av förordning (EG) nr 2535/2001 om tillämpningsföreskrifter för rådets förordning (EG) nr 1255/1999 när det gäller ordningen för import av mjölk och mjölkprodukter och om öppnande av tullkvoter, och om undantag från förordning (EG) nr 2535/2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1255/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter(1), särskilt artiklarna 26.3 och 29.1 i denna, och
av följande skäl:
(1) Kapitel III i kommissionens förordning (EG) nr 2535/2001(2) innehåller bestämmelser om en årlig kvot smör som inte har fördelats under året. För att göra det möjligt att fördela importen inom denna kvot jämnt över kvotåret med syftet att på det sättet säkerställa tillräckliga leveranser till den inre marknaden bör den aktuella kvoten delas upp i en del per halvår med hänsyn tagen till den historiska utvecklingen av importen av produkten i fråga under kvotperioden.
(2) I kapitel I i kommissionens förordning (EG) nr 2535/2001 ges bestämmelser om kvoter som under januari och juli varje år fördelas på grundval av halvårskvoter. Med anledning av de tio nya medlemsstaternas anslutning den 1 maj 2004 bör det utformas föreskrifter som gör det möjligt för aktörerna i dessa länder att få del av gemenskapens kvoter från detta datum. Det är av det skälet lämpligt att begränsa de kvoter som öppnas i januari 2004 till de kvantiteter som motsvarar perioden januari-april 2004. Denna fördelning bör dock inte tillämpas på kvoter för hela kalenderåret, om de kännetecknas av underutnyttjande under den föregående perioden.
(3) I förordning (EG) nr 2535/2001 fastställs det inom sektorn för mjölk och mjölkprodukter bland annat tillämpningsföreskrifter för importordningar mellan gemenskapen och dess medlemsstater å ena sidan och vissa central- och östeuropeiska länder å andra sidan. För att de medgivanden skall kunna verkställas som föreskrivs i rådets beslut 2003/452/EG av den 26 maj 2003 om ingående av ett protokoll om anpassning av handelsaspekterna i Europaavtalet om upprättandet av en associering mellan Europeiska gemenskaperna och deras medlemsstater, som handlar inom ramen för Europeiska unionen, å ena sidan, och Republiken Slovenien, å andra sidan, för att beakta resultaten av förhandlingarna mellan parterna om nya ömsesidiga jordbruksmedgivanden(3) bör vissa redan befintliga kvoter ökas.
(4) För att det skall gå att följa utvecklingen när det gäller ostimportens sammansättning i de olika kvoterna föreskrivs det i artikel 19 i förordning (EG) nr 2535/2001 att aktörerna skall ange vissa halter på importdeklarationen. Om de angivna halterna överskrider de halter som anges i bilaga XIII till den nämnda förordningen skall de behöriga myndigheterna informera kommissionen. De meddelanden som har nått kommissionen, sedan detta krav infördes, vittnar om en viss stabilitet i sammansättningen av ostimporten, när det gäller ostens typ och ursprung. Meddelandena skapar en avsevärd arbetsbörda för tullmyndigheterna och för kommissionen och en betydande mängd dokument överförs, under det att större delen av fallen av överskridanden av bashalterna inte är särskilt omfattande. Meddelandena bör därför fortsättningsvis kunna begränsas till de fall där halterna är onormalt höga genom en anpassning av halterna i bilaga XIII. Det har vidare visat sig att intresset för att få information när halterna enligt bilaga XIII överskrids för vissa ostsorter är försumbart, eftersom variationen i halterna är begränsad till intervallet mellan de övre och undre gränserna för dessa produkter enligt KN. Kravet på meddelanden om dessa produkter bör upphävas.
(5) Nya Zeeland har skickat in uppgifter till kommissionen om ett nytt utfärdande organ. Bilaga XII till förordning (EG) nr 2535/2001 bör alltså uppdateras.
(6) Med anledning av nyanslutningarna den 1 maj 2004 bör giltighetstiden för de importlicenser som används för import från de nya medlemsstaterna begränsas till den 30 april 2004. Därför bör ett undantag göras från artikel 16.3 i förordning (EG) nr 2535/2001.
(7) Uppdelningen i halvårsdelar av smörkvoten enligt kapitel 3 i förordning (EG) nr 2535/2001 påverkar arbetsrytmen när det gäller att utfärda IMA 1-intyg för de utfärdande organen i de berörda tredjeländerna. För att ge möjlighet för de behöriga myndigheterna i dessa länder och för de berörda aktörerna att ta del av denna förändring innan den börjar gälla och för att uppfylla gemenskapens internationella förpliktelser bör det föreskrivas en tidsfrist mellan offentliggörandet och ikraftträdandet av uppdelningen av den nämnda kvoten som är tillräckligt lång. Eftersom IMA 1-intygen för 2004 kan utfärdas redan från 1 november 2003 av tredjeländernas utfärdande organ, bör godkännande ges för att utfärda importlicenser för alla IMA 1-intyg som har utfärdats fram till och med dagen före det datum då uppdelningen av kvoten träder i kraft.
(8) Förordning (EG) nr 2535/2001 bör alltså ändras och undantag göras från den.
(9) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för mjölk och mjölkprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 2535/2001 ändras på följande sätt:
1) Artikel 24.2 skall ersättas med följande:
%quot%2. De rättigheter som gäller och de största kvantiteter som får importeras under kvotperioden för den import som avses i punkt 1 a, anges i bilaga III.%quot%
2) I artikel 26.2 skall följande stycke läggas till:
%quot%IMA 1-intyg får dock utfärdas för kvot nr 09.4589
a) från och med den 1 november varje år och vara giltiga från och med den 1 januari följande år för kvantiteter som inte överskrider den maximala kvantiteten för den första kvotperioden för året enligt bilaga III.A; ansökningar om importlicenser får dock tidigast lämnas in den första arbetsdagen i januari,
b) från och med 1 maj varje år och gälla från och med närmast följande 1 juli för återstoden av den årskvot som avses i bilaga III.A; ansökningar om importlicenser får dock tidigast lämnas in den första arbetsdagen i juli.%quot%
3) Bilaga I skall ändras på följande sätt:
a) Del I.A skall ersättas med texten i bilaga I till den här förordningen.
b) I del I.B skall punkterna 5, 6, och 10 ersättas med bilaga II till den här förordningen.
c) Delarna I.F och I.H skall ersättas med bilaga III till den här förordningen.
4) I bilaga III.A skall de uppgifter som avser kvot nr 09.4589 ersättas med bilaga IV till den här förordningen.
5) I bilaga XII skall de uppgifter som avser det utfärdande organet för Nya Zeeland ersättas med följande:
%quot%%gt%Plats för tabell%gt%%quot%
6) Bilaga XIII skall ersättas med bilaga V till den här förordningen.
Artikel 2
Genom undantag från artikel 16.3 i förordning (EG) nr 2535/2001 skall licensernas giltighet löpa ut den 30 april för
a) import enligt de kvoter som avses i bilaga I.B, punkterna 1-4 och 7-10,
b) import från de nya medlemsstaterna enligt den kvot som avses i bilaga I.A.
Artikel 3
Genom undantag från artikel 24.2 och artikel 26.2 får importlicenser för 2004 avseende kvot nr 09.4589 utfärdas vid uppvisande av IMA 1-intyg som har utfärdats fram till och med dagen närmast före den dag då de bestämmelser träder i kraft som avses i artikel 1.1-1.2.
Artikel 4
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska unionens officiella tidning.
Artikel 1.1, 1.2 och 1.4 samt artikel 3 skall gälla från och med den tjuguförsta dagen efter det datum då den här förordningen har offentliggjorts i Europeiska unionens officiella tidning.
Artikel 1.3, 1.5 och 1.6 samt artikel 2 skall gälla från och med den 1 januari 2004.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Rådets förordning (EG) nr 57/2004
av den 27 oktober 2003
om ändring av kommissionens beslut 2002/602/EKSG om förvaltning av vissa importbegränsningar för vissa stålprodukter från Ryska federationen
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättande av Europeiska gemenskapen, särskilt artikel 133 i detta,
med beaktande av kommissionens förslag, och
av följande skäl:
(1) Avtalet om partnerskap och samarbete som upprättar ett partnerskap mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Ryska federationen, å andra sidan(1), trädde i kraft den 1 december 1997.
(2) I artikel 21 i avtalet om partnerskap och samarbete fastställs det att handel med produkter som omfattas av Fördraget om Europeiska kol- och stålgemenskapen (nedan kallad %quot%EKSG%quot%) skall regleras genom bestämmelserna i avdelning III, med undantag av artikel 15, och genom bestämmelserna i ett avtal.
(3) EKSG och Ryska federationens regering ingick den 9 juli 2002 ett sådant avtal om handel med vissa stålprodukter(2), vilket godkändes på EKSG:s vägnar genom kommissionens beslut 2002/603/EKSG(3).
(4) Fördraget om upprättandet av Europeiska kol- och stålgemenskapen upphörde att gälla den 23 juli 2002. I enlighet med artikel 10.2 i avtalet om handel med vissa stålprodukter enades parterna om att avtalet borde fortsätta att gälla och att alla rättigheter och skyldigheter borde bibehållas efter det att fördraget upphört att gälla. (5) Ryska federationens regering har i enlighet med artikel 3.3 i avtalet begärt överföring av vissa kvantiteter av de kvantitativa begränsningarna som inte utnyttjats under 2002. Följande överföringar har godkänts för varje produktgrupp: 2186980 kilogram för SA1, 10802830 kilogram för SA1a, 4200000 kilogram för SA2, 2505046 kilogram för SA3, 0 för SA4, 272850 kilogram för SB1, 4200000 för SB2 och 11550000 för SB3.
(6) Ryska federationens regering har i enlighet med artikel 3.4 i avtalet begärt att 4000 ton från produktgrupp SB2 och 6000 ton från produktgrupp SB3 skall överföras till produktgrupp SA1a.
(7) Parterna har inlett samråd enligt godkänt protokoll nr 2 till det ovannämnda avtalet och dragit slutsatsen att avtalets produkttäckning måste utvidgas så att även produktgrupperna SA5 och SA6 omfattas; detta genom ett nytt avtal som ändrar det tidigare avtalet.
(8) Gemenskapen godkände ingåendet av det nya avtalet, vilket trädde i kraft samma dag som det undertecknades(4).
(9) Kommissionens beslut 2002/602/EKSG om förvaltning av vissa importbegränsningar för vissa stålprodukter från Ryska federationen(5) måste därför ändras i syfte att beakta begäran om överföring av outnyttjade kvantiteter, begäran om överföring till en annan produktgrupp och det nya avtalet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Beslut 2002/602/EKSG ändras på följande sätt: 1. Bilaga I skall ersättas med texten i bilaga I till den här förordningen.
2. Bilaga IV skall ersättas med texten i bilaga II till den här förordningen.
Artikel 2
För import till gemenskapen av produkter som omfattas av produktgrupperna SA5 och SA6 och som åtföljs av ett kontrolldokument(6) utfärdat före dagen för ikraftträdandet av denna förordning skall det inte krävas ett sådant importtillstånd som anges i beslut 2002/602/EKSG, särskilt i artikel 2 i detta.
Artikel 3
Import till gemenskapen från Ryska federationen av produkter som omfattas av produktgrupperna SA5 och SA6, enligt definitionen i bilaga I, skall från och med den 1 januari 2003 dras av från de kvantitativa begränsningar för dessa produktgrupper för år 2003 som fastställs i bilaga II.
Artikel 4
Denna förordning träder i kraft den tionde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 592/2004
av den 30 mars 2004
om ändring av Europarlamentets och rådets förordning (EG) nr 998/2003 när det gäller förteckningarna över länder och territorier
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 998/2003 av den 26 maj 2003 om djurhälsovillkor som skall tillämpas vid transporter av sällskapsdjur utan kommersiellt syfte och om ändring av rådets direktiv 92/65/EEG(1), särskilt artiklarna 10 och 21 i denna, och
av följande skäl:
(1) I förordning (EG) nr 998/2003 fastställs de djurhälsovillkor som skall vara uppfyllda vid transporter av sällskapsdjur utan kommersiellt syfte samt de regler som skall gälla för kontroll av sådana transporter.
(2) I enlighet med förordning (EG) 998/2003 skall en förteckning upprättas över tredje länder före den 3 juli 2004. För att kunna upptas i förteckningen skall ett tredje land styrka sin rabiesstatus samt att det uppfyller vissa bestämmelser rörande anmälan, övervakning, veterinärmyndigheter, förebyggande och kontroll av rabies och föreskrifter gällande vacciner.
(3) För att inte i onödan störa transporterna av sällskapsdjur och för att ge tredje länder tid att lämna ytterligare garantier där detta är nödvändigt, är det lämpligt att upprätta en provisorisk förteckning över tredje länder. Förteckningen bör baseras på uppgifter från Internationella byrån för epizootiska sjukdomar (OIE), resultat från inspektioner utförda av kommissionens kontor för livsmedels- och veterinärfrågor i de berörda tredje länderna och information som samlats in av medlemsstaterna.
(4) Den provisoriska förteckningen över tredje länder bör omfatta länder som är rabiesfria och länder för vilka det har konstaterats att risken att rabies förs in till gemenskapen som en följd av transport från deras territorier inte är högre än riskerna i samband med transporter mellan medlemsstaterna.
(5) Förordning (EG) nr 998/2003 bör följaktligen ändras. För tydlighetens skull bör den förteckning över länder och territorier som anges i den förordningen ersättas i sin helhet.
(6) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga II till förordning (EG) nr 998/2003 skall ersättas med bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Den skall tillämpas från den 3 juli 2004.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1891/2004
av den 21 oktober 2004
om fastställande av tillämpningsföreskrifter för rådets förordning (EG) nr 1383/2003 om tullmyndigheternas ingripande mot varor som misstänks göra intrång i vissa immateriella rättigheter och om vilka åtgärder som skall vidtas mot varor som gör intrång i vissa immateriella rättigheter
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1383/2003 av den 22 juli 2003 om tullmyndigheternas ingripande mot varor som misstänks göra intrång i vissa immateriella rättigheter och om vilka åtgärder som skall vidtas mot varor som gör intrång i vissa immateriella rättigheter [1] särskilt artikel 20 i denna, och
av följande skäl:
(1) Genom förordning (EG) nr 1383/2003 införs gemensamma regler som har till syfte att förbjuda införsel, övergång till fri omsättning, utförsel, export, återexport, hänförande till ett suspensivt arrangemang eller uppläggning i en frizon eller ett frilager av varumärkesförfalskade och pirattillverkade varor och att effektivt bekämpa olaglig saluföring av sådana varor utan att för den skull hindra den lagliga handeln.
(2) Eftersom förordning (EG) nr 1383/2003 har ersatt rådets förordning (EG) nr 3295/94 av den 22 december 1994 om fastställande av vissa åtgärder avseende införsel till gemenskapen samt export och återexport från gemenskapen av varor som gör intrång i viss immateriell äganderätt [2] bör kommissionens förordning (EG) nr 1367/95 [3] om tillämpningsföreskrifter till förordning (EG) nr 3295/94 ersättas.
(3) För varje immateriell rättighet bör det fastställas vilka fysiska och juridiska personer som kan företräda rättighetshavaren eller varje annan person som är bemyndigad att använda denna rättighet.
(4) Det bör fastställas vilka former av handlingar som styrker att sökanden är rättighetshavare till en immateriell rättighet som krävs enligt artikel 5.5 andra stycket i förordning (EG) nr 1383/2003.
(5) I syfte att harmonisera och förenhetliga innehållet i och formen för formulären för ansökan om ingripande och de uppgifter som skall anges i formulären för de ansökningar om ingripande som avses i artikel 5.1 och 5.4 i förordning (EG) nr 1383/2003 bör en förlaga upprättas för dessa. Dessutom bör det närmare anges vilka språk som skall användas för den ansökan om ingripande som avses i artikel 5.4 i förordning (EG) nr 1383/2003.
(6) I syfte att underlätta för tullmyndigheterna att identifiera varor som kan göra intrång på en immateriell rättighet bör det fastställas vilka uppgifter som skall anges i ansökan om ingripande.
(7) Det bör fastställas vilken slags förklaring om rättighetshavarens ansvarsskyldighet som måste åtfölja ansökan om ingripande.
(8) I syfte att skapa ett klart rättsläge bör det fastställas när de tidsfrister som avses i artikel 13 i förordning (EG) nr 1383/2003 börjar.
(9) Förfaranden för informationsutbyte mellan medlemsstaterna och kommissionen bör fastställas dels för att göra det möjligt för kommissionen att övervaka tillämpningen av det förfarande som fastställs i förordning (EG) nr 1383/2003, vid lämplig tidpunkt utarbeta den rapport som avses i artikel 23 i den förordningen och försöka göra en kvantitativ och kvalitativ analys av de typer av bedrägerier som förekommer, dels för att medlemsstaterna skall kunna införa en lämplig riskanalys.
(10) Denna förordning bör tillämpas från och med samma dag som förordning (EG) nr 1383/2003 träder i kraft.
(11) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Tullkodexkommittén.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Med avseende på tillämpningen av artikel 2.2 b i förordning (EG) nr 1383/2003 (nedan kallad %quot%grundförordningen%quot%) kan rättighetshavaren eller varje annan person som bemyndigats att använda rättigheten företrädas av fysiska och juridiska personer.
De personer som avses i första stycket kan bl.a. vara upphovsrättsorganisationer vars enda eller huvudsakliga uppgift är att förvalta upphovsrätter och därmed sammanhängande rättigheter, sammanslutningar, eller företrädare för dessa, som lämnat en ansökan om registrering av en skyddad ursprungsbeteckning eller en skyddad geografisk beteckning, samt växtförädlare.
Artikel 2
1. I det fall en ansökan om ingripande enligt artikel 5.1 i grundförordningen lämnas av rättighetshavaren själv skall de styrkande handlingar som avses i artikel 5.5 andra stycket i grundförordningen utgöras av följande:
a) För rättigheter som har registrerats eller för vilka det inlämnats en ansökan fordras ett registreringsbevis utfärdat av berörd myndighet eller bevis för att ansökan inlämnats.
b) För upphovsrätter och därmed sammanhängande rättigheter och för mönsterskydd som inte registrerats eller för vilka det inte inlämnats någon ansökan fordras bevis för att den berörda personen är upphovsmannen eller den ursprunglige rättighetshavaren.
Som bevis enligt första stycket i punkt a, räknas en kopia av registreringen i databas hos en nationell myndighet eller ett internationellt organ.
För skyddade ursprungsbeteckningar och skyddade geografiska beteckningar skall beviset enligt första stycket punkt a dessutom innefatta ett bevis att rättighetsinnehavaren är producenten eller sammanslutningen och ett bevis för att ursprungsbeteckningen eller den geografiska beteckningen är registrerad. Detta gäller även i tillämpliga delar för viner och spritdrycker.
2. I det fall ansökan om ingripande lämnas av en annan person som bemyndigats att använda en rättighet enligt artikel 2.1 i grundförordningen skall de styrkande handlingarna, utöver de bevis som avses i punkt 1, utgöras av det dokument genom vilket den berörda personen bemyndigas att använda rättigheten i fråga.
3. I det fall ansökan om ingripande lämnas av en företrädare för rättighetshavaren eller en annan person som bemyndigats att använda en rättighet enligt artikel 2.2 i grundförordningen skall de styrkande handlingarna, utöver de bevis som avses i punkt 1 i denna artikel, utgöras av ett bevis om bemyndigandet att agera i rättighetshavarens ställe.
Företrädaren enligt första stycket skall uppvisa den förklaring som avses i artikel 6 i grundförordningen, vilken skall vara undertecknad av de personer som avses i punkterna 1 och 2 i denna artikel, eller ett dokument genom vilket han bemyndigas att i deras namn bära alla de kostnader som följer av tullmyndigheternas ingripande i deras namn i enlighet med artikel 6 i grundförordningen.
Artikel 3
1. Formuläret för de ansökningar om ingripande som avses i artikel 5.1 och 5.4 i grundförordningen, de beslut som avses i punkterna 7 och 8 i den artikeln och den förklaring som avses i artikel 6 i grundförordningen skall följa de förlagor som är bifogade den här förordningen.
Formulären skall ifyllas på elektronisk eller mekanisk väg alternativt för hand, under förutsättning att det är läsligt. Om det fylls i för hand skall formuläret fyllas i med bläck och med tryckbokstäver. Oavsett vilken metod som väljs accepteras inte raderingar, överskrivningar eller andra ändringar. När det gäller formulär som fylls i på elektronisk väg skall dessa finnas tillgängliga för dem som ansöker om formulär i digital form på minst en offentlig webbplats. Det är tillåtet att med hjälp av privat tryckningsutrustning flerfaldiga ett formulär som hämtats i elektronisk form.
I det fall det görs bruk av de extrablad som avses i fälten 8, 9, 10 och 11 i formuläret för den ansökan om ingripande som avses i artikel 5.1 i grundförordningen eller i fälten 7, 8, 9 och 10 i formuläret för den ansökan om ingripande som avses i artikel 5.4 i den förordningen skall dessa anses utgöra en integrerad del av formuläret.
2. Formulär som avser en ansökan enligt artikel 5.4 i grundförordningen skall tryckas och fyllas i på ett officiellt gemenskapsspråk som fastställs av de behöriga myndigheterna i den medlemsstat där ansökan om ingripande, och eventuella översättningar av denna, skall inlämnas.
3. Formuläret skall utfärdas i två exemplar:
a) Ett exemplar, märkt med nr 1, avsett för den medlemsstat i vilken ansökan lämnas in.
b) Ett exemplar, märkt med nr 2, avsett för rättighetshavaren.
Det ifyllda och undertecknade formuläret jämte ett antal utdrag ur detta motsvarande det antal medlemsstater som anges i ruta 6 i formuläret, samt styrkande handlingar som anges i rutorna 8, 9 och 10 skall uppvisas för behörig tullmyndighet och efter godkännandet bevaras av denna under minst ett år utöver formulärets giltighetstid.
Endast i det fall utdraget ur ett beslut om beviljande av ansökan om ingripande är ställd till en eller flera medlemsstater i enlighet med artikel 5.4 i grundförordningen skall den medlemsstat som mottar utdraget omgående fylla i dagen för mottagandet i det fält som är avsett för detta och återsända en kopia av utdraget till den behöriga myndighet som anges i ruta 2 i formuläret.
Rättighetshavaren kan så länge hans ansökan om gemenskapsingripande är giltig i den medlemsstat där ansökan ursprungligen lämnades, ansöka om ingripande i en ny medlemsstat som inte tidigare nämnts i ansökan. I detta fall skall giltighetstiden för den nya ansökan vara lika med den period som återstår av den ursprungliga ansökans giltighetstid och får förlängas i enlighet med de villkor som gäller för den ursprungliga ansökan.
Artikel 4
Med avseende på artikel 5.6 i grundförordningen kan den myndighet som tar emot och behandlar ansökningarna om ingripande begära uppgifter om tillverkningsorten, distributionsnätet, namnet på licensinnehavarna samt andra uppgifter i syfte att underlätta den tekniska analysen av de berörda varorna.
Artikel 5
I det fall en ansökan om ingripande lämnas i enlighet med artikel 4.1 i grundförordningen innan tidsfristen på tre arbetsdagar löpt ut skall de tidsfrister som avses i artiklarna 11 och 13 i grundförordningen börja löpa först dagen efter mottagandet av ansökan om ingripande, som godkänts av den tullmyndighet som utsetts för det ändamålet.
Om tullmyndigheten i enlighet med artikel 4.1 underrättar deklaranten eller varuinnehavaren om att frigörandet av varor uppskjutits eller att varor kvarhållits därför att de misstänks göra intrång på en immateriell rättighet, skall tidsfristen på tre arbetsdagar räknas först från och med den dag då rättighetshavaren delges underrättelsen.
Artikel 6
När det gäller lättfördärvliga varor skall förfarandet för uppskjutande av frigörandet av varorna eller för kvarhållande av varorna inledas i första hand för varor för vilka det redan inlämnats en ansökan om ingripande.
Artikel 7
1. Vid tillämpning av artikel 11.2 i grundförordningen skall rättighetshavaren underrätta tullmyndigheten om att det har inletts ett förfarande för att fastställa huruvida det gjorts intrång i en immateriell rättighet enligt den nationella lagstiftningen. Om den återstående tidsfristen enligt artikel 13.1 första stycket i grundförordningen inte är tillräcklig för att inleda ett sådant förfarande kan denna tidsfrist, utom när det gäller lättfördärvliga varor, förlängas enligt artikel 13.1 andra stycket i grundförordningen.
2. Om en förlängning med tio arbetsdagar redan beviljats i enlighet med artikel 11 i grundförordningen kan en förlängning i enlighet med artikel 13 i grundförordningen inte beviljas.
Artikel 8
1. Varje medlemsstat skall så snart som möjligt lämna uppgifter till kommissionen om den enhet vid tullmyndigheten som enligt artikel 5.2 i grundförordningen skall vara behörig att ta emot och behandla ansökningar om ingripande från rättighetshavaren.
2. Varje medlemsstat skall i slutet av varje kalenderår förelägga kommissionen en förteckning över samtliga skriftliga ansökningar om ingripande enligt artikel 5.1 och 5.4 i grundförordningen och uppge rättighetshavarens namn, adress och telefonnummer och vilken slags rättighet ansökan avser samt inge en kortfattad varubeskrivning. Även ansökningar som inte beviljats skall redovisas.
3. Månaden efter utgången av varje kvartal skall medlemsstaterna förelägga kommissionen en förteckning för varje produkttyp som skall innehålla närmare uppgifter om de fall där frigörandet av varorna har uppskjutits eller där varorna har kvarhållits. Förteckningen skall innehålla följande uppgifter:
a) Rättighetshavarens namn, varubeskrivning och, om detta är känt, ursprung, avsändarland och bestämmelseort för varorna och namnet på den immateriella rättighet som det gjorts intrång i.
b) Antalet varor av varje produkt för vilka frigörandet uppskjutits eller som kvarhållits, dessa varors tullstatus, den typ av immateriell rättighet som det gjorts intrång i och transportsätt.
c) Huruvida det rör sig om kommersiell trafik eller passagerartrafik, och huruvida det rör sig om ett förfarande som inletts till följd av en ansökan om ingripande eller ett förfarande som inletts på tullmyndigheternas initiativ. 4. Medlemsstaterna får underrätta kommissionen om det verkliga eller förmodade värdet på de varor för vilka frigörandet har uppskjutits eller som kvarhållits.
5. Kommissionen skall i slutet av varje år översända de uppgifter den erhållit i enlighet med punkterna 1-4 till medlemsstaterna.
6. Kommissionen skall i Europeiska unionens officiella tidning, C-serien, offentliggöra en förteckning över de behöriga tullmyndigheter som avses i artikel 5.2 i grundförordningen.
Artikel 9
Ansökningar om ingripande som lämnats in före den 1 juli 2004 är giltiga till dess att de rättsligen upphör att gälla och kan inte förlängas. De måste emellertid kompletteras med den förklaring som avses i artikel 6 i grundförordningen, varav en förlaga återfinns i bilagan till denna förordning. Genom denna förklaring frigörs de garantier som eventuellt skall erläggas i medlemsstaterna.
Om ett förfarande för avgörande i sakfrågan har inletts vid den behöriga myndigheten före den 1 juli 2004 och detta ännu inte har avslutats vid det datumet kommer garantin att frigöras först när förfarandet har avslutats.
Artikel 10
Förordning (EG) nr 1367/95 skall upphöra att gälla. Hänvisningar till den upphävda förordningen skall betraktas som hänvisningar till den här förordningen.
Artikel 11
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska unionens officiella tidning.
Den skall tillämpas från och med den 1 juli 2004.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 2140/2004
av den 15 december 2004
om tillämpningsföreskrifter för förordning (EG) nr 1245/2004 när det gäller ansökningar om fiskelicenser i vatten under Grönlands exklusiva ekonomiska zon
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1245/2004 av den 28 juni 2004 om ingående av protokollet om ändring av det fjärde protokollet om villkor för det fiske som föreskrivs i avtalet om fiske mellan Europeiska ekonomiska gemenskapen, å ena sidan, och Danmarks regering och Grönlands lokala regering, å andra sidan [1], särskilt artikel 4 andra stycket i denna, och
av följande skäl:
(1) I förordning (EG) nr 1245/2004 föreskrivs det att ägare till gemenskapsfartyg som får en licens för ett fartyg med rätt att fiska i vatten under Grönlands exklusiva ekonomiska zon skall betala en licensavgift enligt artikel 11.5 i det fjärde protokollet.
(2) I artikel 11.5 i det fjärde protokollet föreskrivs det att de tekniska genomförandevillkoren för tilldelningen av licenserna skall fastställas genom en administrativ överenskommelse mellan parterna.
(3) Grönlands regering och Europeiska gemenskapen har fört förhandlingar för att fastställa de formella reglerna för licensansökningarna och deras utfärdande, och förhandlingarna ledde fram till att en administrativ överenskommelse paraferades den 30 september 2004.
(4) Bestämmelserna i denna administrativa överenskommelse bör därför tillämpas.
(5) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Kommittén för fiske och vattenbruk.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De formella reglerna för ansökningar om fiskelicens och deras utfärdande enligt artikel 4 i förordning (EG) nr 1245/2004 fastställs i den administrativa överenskommelse som återges i bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft den sjunde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Den skall tillämpas från och med den 1 januari 2005.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Rådets förordning (EG) nr 2257/2004
av den 20 december 2004
om ändring av förordningarna (EEG) nr 3906/89, (EG) nr 1267/1999, (EG) nr 1268/1999 och (EG) nr 2666/2000 för att ta hänsyn till Kroatiens ställning som kandidatland
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 181a.2,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets yttrande, och
av följande skäl:
(1) Europeiska rådet beslutade vid sitt möte i Bryssel den 17 och 18 juni 2004 att Kroatien skulle få status som kandidatland för medlemskap och uppmanade kommissionen att utarbeta en föranslutningsstrategi för Kroatien inklusive nödvändiga finansiella instrument.
(2) För att kunna ge föranslutningsstöd till Kroatien bör landet tas upp bland stödmottagarna enligt rådets förordningar (EEG) nr 3906/89 av den 18 december 1989 om ekonomiskt stöd till vissa länder i Central- och Östeuropa (Phare) [1], rådets förordning (EG) nr 1267/1999 av den 21 juni 1999 om upprättande av ett strukturpolitiskt föranslutningsinstrument [2] (ISPA) och rådets förordning (EG) nr 1268/1999 av den 21 juni 1999 om gemenskapsstöd för föranslutningsåtgärder för jordbruket och landsbygdens utveckling i kandidatländerna i Central- och Östeuropa under föranslutningsperioden [3] (Sapard).
(3) I avdelning III i stabiliserings- och associeringsavtalet mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Republiken Kroatien, å andra sidan, undertecknat den 29 oktober 2001, uppmanas Kroatien att aktivt främja regionalt samarbete på västra Balkan.
(4) Den regionala aspekten av gemenskapsbiståndet till västra Balkan får särskild uppmärksamhet i rådets förordning (EG) nr 2666/2000 av den 5 december 2000 om bistånd till Albanien, Bosnien och Hercegovina, Kroatien, Förbundsrepubliken Jugoslavien och f.d. jugoslaviska republiken Makedonien [4] (Cards) vars syfte är att stärka det regionala samarbetet och Kroatien bör även fortsättningsvis vara berättigat till stöd för projekt och program som har regionala aspekter.
(5) I beslut 2004/648/EG [5] fastställs principerna, prioriteringarna och villkoren för det europeiska partnerskapet med Kroatien.
(6) Samförståndsavtalet rörande utvecklingen av sydöstra Europas huvudnätverk för regional transport bör underlätta förfarandet för att välja ut prioriterade åtgärder i syfte att utveckla ett alleuropeiskt transportnät under föranslutningsperioden.
(7) I och med ikraftträdandet av förordning (EG, Euratom) 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget [6] krävs vissa anpassningar av förordningarna i fråga för att få terminologi och nuvarande förfaranden förenliga med den.
(8) De nya medlemsstaterna nämns inte i denna förordning, men enligt artikel 33 i 2003 års anslutningsakt skall rådets förordningar (EG) nr 3906/89 och (EG) nr 1267/1999 tillämpas på dessa medlemsstater under en övergångsperiod.
(9) Kommissionen har antagit förordningarna (EG) nr 1419/2004 [7] och (EG) nr 447/2004 [8] som utgör den rättsliga grunden för finansieringen av åtgärder inom Sapard för åtaganden som på anslutningsdagen ännu inte var avslutade. De beslut som kommissionen kan behöva fatta innan dessa åtaganden har slutförts och som inte kan grundas på de båda nämnda förordningarna kan fortfarande grundas på förordning (EG) nr 1268/1999, eftersom den var i kraft innan den förordningen ändrades genom denna förordning.
(10) Förordningarna (EEG) nr 3906/89, (EG) nr 1267/1999, (EG) nr 1268/1999 och (EG) nr 2666/2000 bör ändras i enlighet med detta.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Rådets förordning (EEG) nr 3906/89 ändras på följande sätt:
1. Artikel 3 skall ändras på följande sätt:
a) Punkt 3 skall ersättas med följande:
"3. För ansökarländer som har ingått partnerskap för anslutning med Europeiska unionen skall finansieringen inom ramen för Phareprogrammet inriktas på de huvudsakliga prioriteringarna för antagandet av gemenskapens regelverk, det vill säga förstärkning av den administrativa och institutionella kapaciteten i ansökarländerna samt investeringar, med undantag av den typ av investeringar som finansieras i enlighet med rådets förordningar (EG) nr 1267/1999 av den 21 juni 1999 om upprättande av ett strukturpolitiskt föranslutningsinstrument [9] och (EG) nr 1268/1999 av den 21 juni 1999 om gemenskapsstöd för föranslutningsåtgärder för jordbruket och landsbygdens utveckling i kandidatländerna i Central- och Östeuropa under föranslutningsperioden [10], förutsatt att villkoren för finansiering enligt dessa båda förordningar är uppfyllda. Även åtgärder på områdena miljö, transport och jordbruk samt landsbygdsutveckling, vilka utgör en underordnad men nödvändig del av integrerade program som genomförs för omstrukturering av industrin eller regional utveckling, kan finansieras inom ramen för Phareprogrammet.
b) Följande punkter skall läggas till:
"4. Stödet får användas för att täcka utgifter vid mottagarländernas deltagande enligt denna förordning i regionalt, gränsöverskridande och, i tillämpliga fall, transnationellt och interregionalt samarbete dem emellan och mellan dem och EU:s medlemsstater.
5. I tillämpliga fall får stödet också användas för att täcka utgifter vid ett mottagarlands deltagande i regionala program inom ramen för andra rättsliga instrument."
2. I artikel 8 skall följande punkt läggas till:
"Inom de begränsningar som fastställs i artikel 54 i rådets förordning (EG, Euratom) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget [11] får kommissionen besluta att överlåta uppgifter som omfattar myndighetsutövning, särskilt uppgifter för genomförande av budgeten, till de organ som anges i artikel 54.2 i den förordningen. De organ som anges i artikel 54.2 c i förordning (EG, Euratom) nr 1605/2002 får anförtros uppgifter som omfattar myndighetsutövning om de har erkänt internationellt anseende, är uppfyller kraven i internationellt erkända förvaltnings- och kontrollsystem och övervakas av en offentlig myndighet.
3. Förteckningen i bilagan skall ersättas med följande:
"Bulgarien
Kroatien
Rumänien"
Artikel 2
Förordning (EG) nr 1267/1999 ändras på följande sätt:
1. Artikel 1.1 skall ersättas med följande:
"1. Ett strukturpolitiskt föranslutningsinstrument (nedan kallat "ISPA") skall upprättas.
Genom ISPA skall stöd ges för att bidra till Bulgariens, Kroatiens och Rumäniens (nedan kallade "de stödmottagande länderna") förberedelser inför anslutningen till Europeiska unionen på området ekonomisk och social sammanhållning, närmare bestämt med avseende på miljö- och transportpolitiken i enlighet med bestämmelserna i denna förordning."
2. Följande stycke skall läggas till i slutet av artikel 3:
"Oaktat vad som anges ovan skall gemenskapens stöd till Kroatien beviljas under perioden 2005–2006."
3. Följande stycke skall läggas till i slutet av artikel 4:
"Genom undantag från första och andra meningen i denna artikel skall tilldelningen till Kroatien för åren 2005 och 2006 från detta instrument fastställas av kommissionen på grundval av en bedömning av detta stödmottagande lands förmåga att administrera stödet och dess anslutningsrelaterade investeringsbehov."
4. I artikel 9.1 a skall orden "från och med den 1 januari 2000, och i alla händelser senast den 1 januari 2002," utgå.
Artikel 3
Förordning (EG) nr 1268/1999 ändras på följande sätt:
1. Artikel 1.1 skall ersättas med följande:
"1. Genom denna förordning upprättas en ram för gemenskapsstöd för ett hållbart jordbruk och en hållbar landsbygdsutveckling under föranslutningsperioden för Bulgarien, Kroatien och Rumänien. Förordningen skall också fortsätta att tillämpas för att avsluta de program som inletts i enlighet med denna i Estland, Lettland, Litauen, Polen, Slovakien, Slovenien, Tjeckien och Ungern före deras anslutning till Europeiska unionen."
2. Följande stycke skall läggas till i slutet av artikel 4.2:
"Genom avvikelse från första stycket skall planen för Kroatien, på samma villkor som anges i första stycket, omfatta en period på högst två år från och med år 2005."
3. Följande mening skall läggas till i slutet av artikel 5.1:
"När det gäller Kroatien skall programmen emellertid inte bedömas efter halva tiden."
4. Artikel 7 skall ändras på följande sätt:
a) Punkt 1 skall ersättas med följande:
"1. Gemenskapsstöd enligt denna förordning skall beviljas under perioden 2000–2006, med undantag av gemenskapsstödet för Kroatien som skall beviljas under perioden 2005–2005. Budgetmyndigheten skall godkänna de årliga anslagen inom ramen för budgetplanen."
b) Följande stycke skall läggas till i slutet av punkt 3:
"För Kroatien skall emellertid den årliga ekonomiska tilldelningen fastställas separat."
5. Artikel 11 skall ersättas med följande:
"Artikel 11
Kommissionen skall med avseende på genomförandet av artikel 7.2 fördela de tillgängliga resurserna till ansökarländerna. Inom tre månader efter beslutet att ett land skall vara berättigat till stöd enligt denna förordning skall kommissionen informera det ansökarlandet om sitt beslut om den vägledande finansiella fördelningen inom den nuvarande budgetplanen."
Artikel 4
Förordning (EG) nr 2666/2000 ändras på följande sätt:
1. Följande mening skall läggas till i slutet av artikel 1.1:
"Från och med år 2005 skall Kroatien som mottagarland endast ha tillgång till projekt och program med en regional dimension, såsom de som anges i artikel 2.2. Trots föregående mening skall Kroatien även fortsättningsvis vara berättigat till stöd för projekt och program enligt beslut 1999/311/EG."
2. Artikel 7 skall ändras på följande sätt:
a) Punkt 1 skall ersättas med följande:
"1. Kommissionen skall genomföra gemenskapsbiståndet i enlighet med rådets förordning (EG) nr 1605/2002 av den 25 juni 2002 med budgetförordning för Europeiska gemenskapernas allmänna budget [12].
b) Följande punkt skall införas:
"2a. Inom de begränsningar som fastställs i artikel 54 i förordning (EG) nr 1605/2002 får kommissionen besluta att överlåta uppgifter som omfattar myndighetsutövning, särskilt uppgifter för genomförande av budgeten, till de organ som anges i artikel 54.2 i den förordningen. De organ som anges i artikel 54.2 c i den förordningen får anförtros uppgifter som omfattar myndighetsutövning om de har erkänt internationellt anseende, uppfyller kraven i internationellt erkända förvaltnings- och kontrollsystem och övervakas av en offentlig myndighet."
Artikel 5
För genomförandet av föranslutningsinstrumenten och för genomförandet av rådets förordning (EG) nr 1266/1999 av den 21 juni 1999 om samordning av stödet till kandidatländerna inom ramen för föranslutningsstrategin [13] skall hänvisningen till anslutningspartnerskapet [14] och Europaavtalet för Kroatiens vidkommande förstås som en hänvisning till det europeiska partnerskapet [15] och till stabiliserings- och associeringsavtalet.
Artikel 6
Denna förordning träder i kraft den tredje dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Rådets yttrande
av den 8 mars 2005
om Sloveniens uppdaterade konvergensprogram för 2004–2007
(2005/C 177/06)
EUROPEISKA UNIONENS RÅD HAR AVGETT FÖLJANDE YTTRANDE
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1466/97 av den 7 juli 1997 om förstärkning av övervakningen av de offentliga finanserna samt övervakningen och samordningen av den ekonomiska politiken [1], särskilt artikel 9.3,
med beaktande av kommissionens rekommendation, och
efter att ha hört Ekonomiska och finansiella kommittén.
HÄRIGENOM FRAMFÖRS FÖLJANDE.
(1) Den 8 mars 2005 granskade rådet Sloveniens uppdaterade konvergensprogram, som omfattar perioden 2004–2007. Programmet uppfyller delvis uppgiftskraven i "uppförandekoden för stabilitets- och konvergensprogrammens innehåll och utformning". Den offentliga sektorns redovisning följer inte helt ENS 95, vilket framgår av den stora andelen "övriga" intäkter och utgifter som andel av BNP. Slovenien anmodas därför se till att uppgiftskraven följs.
(2) Enligt tillgängliga uppgifter verkar programmets bakomliggande makroekonomiska scenario bygga på rimliga tillväxtantaganden. År 2004 beräknas den reala BNP-tillväxten bli 4,0 % och förväntas ligga kvar på ungefär samma nivå under resten av programperioden. Inflationsprognosen förefaller realistisk, men risker kvarstår.
(3) Programmets bakomliggande budgetstrategi syftar till sunda offentliga finanser i form av ett saldo nära balans, dock inte under programperioden. I programmet planeras en gradvis minskning av det offentliga underskottet under perioden, i form av en konsekvent sänkning av utgifternas procentandel av BNP. Inkomstkvoten skall successivt sjunka till och med 2006 men åter stiga mot slutet av programperioden, till följd av EU-medlemskapets positiva nettoeffekter på budgeten. Enligt anpassningsbanan skall underskottet halveras under de fyra följande åren och uppgå till drygt 1 % år 2007. Den aktuella uppdateringen bekräftar huvudsakligen det föregående programmets planerade korrigeringar med ett något gynnsammare makroekonomiskt scenario.
(4) De risker som omgärdar programmets budgetprognoser verkar i stort sett uppväga varandra. Å ena sidan understöds underskottsmålen av ett rimligt makroekonomiskt scenario. Vidare ankommer det på regeringen att avvisa krav på ytterligare utgifter om underskottsmålet hotas av ogynnsamma omständigheter, vilket också skedde 2004. Dessutom kan den årliga förlusten av momsintäkter på 0,3 % av BNP i budgeten 2005–2007 vara för högt beräknad, vilket gör att skatteintäktsprognoserna är överdrivet försiktiga. Å andra sidan kan nivån på skatteintäkterna vara osäker efter skattereformen. Samtidigt beror utfallet 2007 delvis på EU:s nya budgetplan för 2007–2013 och förutsätter en betydande ökning av budgetens nettointäkter från EU-budgeten Det finns dessutom en risk för att utgiftsmålen överskrids, vilket särskilt kan gälla pensionsutgifterna om översynen år 2006 av nuvarande pensionsindex leder till mindre strikta parametrar.
(5) Mot bakgrund av denna riskbedömning är det inte uppenbart att programmets finanspolitiska inriktning ger en tillräcklig säkerhetsmarginal för att hålla underskottet inom referensvärdet på 3 % av BNP, vid normala konjunktursvängningar utom under programmets sista år. Den räcker heller inte till för att till 2007 uppnå stabilitets- och tillväxtpaktens medelfristiga mål på offentliga finanser nära balans.
(6) Offentliga sektorns bruttoskuld är relativt låg: skuldkvoten beräknas ha uppgått till 30,2 % av BNP 2004, betydligt lägre än fördragets referensvärde på 60 % av BNP, och beräknas uppgå till 29,7 % år 2007.
(7) Slovenien är i farozonen när det gäller de offentliga finansernas hållbarhet på lång sikt, där en viktig aspekt är den förväntade budgetkostnaden för en åldrande befolkning. Den pågående pensionsreformen har påverkat budgeten positivt, men pensionsutgifternas beräknade ökning efter 2020 är fortfarande mycket stor. Trots vissa rationaliseringsåtgärder inom hälso- och sjukvårdssystemet under 2004 skulle även en mer genomgripande reform av hälso- och sjukvårdssystemet bidra till att förbättra de offentliga finansernas hållbarhet på lång sikt.
Mot bakgrund av denna bedömning anser rådet att Slovenien bör
i) utnyttja alla möjligheter att snabbare minska underskottet i de offentliga finanserna, och
ii) ytterligare reformera pensionssystemet samt hälso- och sjukvårdssystemet för att förbättra de offentliga finansernas hållbarhet på lång sikt.
Jämförelse av nyckeltal i makroekonomiska prognoser och budgetprognoser
Konvergensprogram (KP) och kommissionens höstprognos för 2004 (KOM).
| 2004 | 2005 | 2006 | 2007 |
Real BNP-tillväxt(i %) | KP januari 2005 | 4,0 | 3,8 | 3,9 | 4,0 |
KOM oktober 2004 | 4,0 | 3,6 | 3,8 | — |
KP maj 2004 | 3,6 | 3,7 | 3,8 | 3,9 |
HIKP-inflation(i %) | KP januari 2005 | 3,6 | 3,0 | 2,7 | 2,6 |
KOM oktober 2004 | 3,9 | 3,4 | 3,0 | — |
KP maj 2004 | 3,3 | 3,0 | 2,7 | 2,6 |
Saldo i de offentliga finanserna(i % av BNP) | KP januari 2005 | – 2,1 | – 2,1 | – 1,8 | – 1,1 |
KOM oktober 2004 | – 2,3 | – 2,2 | – 1,9 | — |
KP maj 2004 | – 1,9 | – 1,8 | – 1,5 | – 0,9 |
Primärt saldo(i % av BNP) | KP januari 2005 | – 0,3 | – 0,4 | – 0,2 | 0,4 |
KOM oktober 2004 | – 0,3 | – 0,2 | – 0,1 | — |
KP maj 2004 | – 0,3 | – 0,4 | – 0,2 | 0,4 |
Offentliga sektorns bruttoskuld (i % av BNP) | KP januari 2005 | 30,2 | 30,7 | 30,9 | 29,7 |
KOM oktober 2004 | 30,9 | 30,8 | 30,6 | — |
KP maj 2004 | 29,1 | 29,5 | 29,4 | 28,4 |
[1] EGT L 209, 2.8.1997, s. 1. De dokument som denna text hänvisar till återfinns på följande webbplats:http://europa.eu.int/comm/economy_finance/about/activities/sgp/main_en.htm.
--------------------------------------------------
Kommissionens beslut
av den 14 mars 2005
om ändring av beslut 2003/526/EG när det gäller skyddsåtgärder mot klassisk svinpest i Tyskland, Frankrike, Luxemburg och Slovakien
[delgivet med nr K(2005) 600]
(Text av betydelse för EES)
(2005/225/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättande av Europeiska gemenskapen,
med beaktande av rådets direktiv 90/425/EEG av den 26 juni 1990 om veterinära och avelstekniska kontroller i handeln med vissa levande djur och varor inom gemenskapen med sikte på att förverkliga den inre marknaden [1], särskilt artikel 10.4 i detta, och
av följande skäl:
(1) Till följd av utbrotten av klassisk svinpest i vissa medlemsstater antog kommissionen beslut 2003/526/EG av den 18 juli 2003 om skyddsåtgärder mot klassisk svinpest i Belgien, Frankrike, Tyskland och Luxemburg [2]. I det beslutet föreskrivs det vissa ytterligare åtgärder för bekämpning av klassisk svinpest.
(2) Situationen när det gäller klassisk svinpest i vissa delar av Rheinland-Pfalz i Tyskland, i departementet Moselle i Frankrike samt i Luxemburg har förbättrats avsevärt. Detta gäller också i Veterinärdistriktet och livsmedelsförvaltningsområdet Levice, Nitra, Topoľčany, Nové Mesto nad Váhom och distriktet Púchov i Slovakien. De åtgärder som antogs genom beslut 2003/526/EG rörande dessa områden bör därför inte längre tillämpas.
(3) Med tanke på det allmänna sjukdomsläget när det gäller klassisk svinpest i andra områden i Tyskland, Frankrike och Slovakien bör giltighetstiden för beslut 2003/526/EG förlängas.
(4) Beslut 2003/526/EG bör därför ändras i enlighet med detta.
(5) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Beslut 2003/526/EG ändras enligt följande:
1. I artikel 11 skall "den 30 april 2005" ersättas med "den 30 april 2006".
2. Bilagan skall ersättas med bilagan till detta beslut.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 14 mars 2005
om ändring av beslut 2005/59/EG beträffande de områden där planerna för utrotning av klassisk svinpest bland viltlevande svin och nödvaccinering av viltlevande svin mot klassisk svinpest skall genomföras i Slovakien
[delgivet med nr K(2005) 601]
(Endast den slovakiska texten är giltig)
(Text av betydelse för EES)
(2005/226/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 2001/89/EG av den 23 oktober 2001 om gemenskapsåtgärder för bekämpning av klassisk svinpest [1], särskilt artiklarna 16.1 och 20.2 i detta, och
av följande skäl:
(1) Kommissionen antog sitt beslut 2005/59/EG av den 26 januari 2005 om att godkänna planerna för utrotning av klassisk svinpest hos vildlevande svin och nödvaccinering av sådana svin i Slovakien [2] som en av flera åtgärder för bekämpning av klassisk svinpest.
(2) De slovakiska myndigheterna har informerat kommissionen om hur denna sjukdom har utvecklats under den senaste tiden bland viltlevande svin. Av denna information framgår att klassisk svinpest bland viltlevande svin har utrotats i Veterinärdistriktet och livsmedelsförvaltningsområdet Levice, Nitra, Topoľčany, Nové Mesto nad Váhom och distriktet Púchov och att den godkända planen för utrotning inte längre behöver tillämpas i dessa områden. Mot bakgrund av den epidemiologiska informationen bör planen för vaccinering utvidgas så att viltlevande svin även i distrikten Ilava, Žiar nad Hronom, Žarnovica and Banská Štiavnica vaccineras mot klassisk svinpest.
(3) Beslut 2005/59/EG bör därför ändras i enlighet med detta.
(4) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till beslut 2005/59/EG skall ersättas med bilagan till det här beslutet.
Artikel 2
Detta beslut riktar sig till Republiken Slovakien.
Kommissionens beslut
av den 29 april 2005
om undantag från vissa bestämmelser i rådets direktiv 2000/29/EG beträffande obarkade stockar av ek (Quercus L.) med ursprung i Amerikas förenta stater
[delgivet med nr K(2005) 1298]
(2005/359/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 2000/29/EG av den 8 maj 2000 om skyddsåtgärder mot att skadegörare på växter eller växtprodukter förs in till gemenskapen och mot att de sprids inom gemenskapen [1], särskilt artikel 15.1 i detta, och
av följande skäl:
(1) Enligt direktiv 2000/29/EG får obarkade stockar av ek (Quercus L.) med ursprung i Amerikas förenta stater i princip inte föras in i gemenskapen på grund av risken för införsel av Ceratocystis fagacearum (Bretz) Hunt, som orsakar ekvissnesjuka.
(2) Erfarenheten har visat att med avseende på Amerikas förenta stater kan risken att Ceratocystis fagacearum (Bretz) Hunt sprids elimineras genom tillämpning av vissa åtgärder.
(3) En sådan åtgärd är gasning. Vissa medlemsstater har begärt att införsel av gasade ekstockar bara skall äga rum i angivna hamnar där nödvändiga hanterings- och inspektionsfaciliteter finns tillgängliga.
(4) Det är också möjligt att avstå från gasning när det gäller ekvirke som tillhör viteksgruppen, om vissa tekniska villkor föreligger. Vissa medlemsstater har dessutom begärt undantag för att tillåta införsel av vitek under vissa månader på året. Detta senare undantag bör begränsas till de delar av gemenskapen där potentiella vektorer för Ceratocystis fagacearum (Bretz) Hunt har liten eller ingen aktivitet under vintern, dvs. områden norr om 45° nordlig bredd.
(5) Kommissionen kommer att se till att Amerikas förenta stater tillhandahåller all teknisk information som krävs för att övervaka tillämpningen av de nödvändiga skyddsåtgärderna.
(6) Medlemsstaterna bör därför bemyndigas att tillämpa ett tidsbegränsat undantag för införsel av obarkade stockar av ek (Quercus L.) från Amerikas förenta stater.
(7) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för växtskydd.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Genom undantag från artikel 5.1 i direktiv 2000/29/EG och från artikel 13.1 i tredje strecksatsen i det direktivet med avseende på bilaga IV A I 3 i det direktivet bemyndigas medlemsstaterna att med verkan från och med den 1 januari 2005 tillåta införsel på sitt territorium av obarkade stockar av ek (Quercus L.) med ursprung i Amerikas förenta stater (nedan kallade "stockarna"), förutsatt att villkoren i artiklarna 2–7 uppfylls.
Artikel 2
1. För att detta undantag skall kunna tillämpas måste stockarna ha gasats och identifierats i enlighet med bilaga I.
2. Medlemsstaterna får undanta gasade stockar från de krav som anges i artikel 5.1 med avseende på våtlagring, artiklarna 5.2 och 6.2.
Artikel 3
1. Stockarna får endast lossas i de hamnar som förtecknas i bilaga II.
2. På begäran av den berörda medlemsstaten får förteckningen över lossningshamnar i bilaga II ändras av kommissionen efter samråd med övriga medlemsstater.
Artikel 4
1. De inspektioner som krävs i enlighet med artikel 13 i direktiv 2000/29/EG skall utföras av tjänstemän som har fått särskild instruktion eller utbildning angående detta beslut, med bistånd av sådana experter som avses i artikel 21 i direktiv 2000/29/EG på det sätt som anges där, antingen i de hamnar som förtecknas i bilaga II eller på den första lagerplatsen i enlighet med artikel 5.
Om lossningshamnen och den första lagerplatsen är belägna i olika medlemsstater skall de medlemsstaterna träffa överenskommelser om var inspektionerna skall utföras och utbyta information om ankomst och lagring av sändningarna.
2. Inspektionerna skall omfatta följande:
a) En granskning av varje sundhetscertifikat.
b) En identitetskontroll som innebär att märkningen på varje stock och antalet stockar jämförs med uppgifterna i det tillhörande sundhetscertifikatet.
c) Ett färgreaktionstest för påvisande av gasning, enligt bilaga III, av ett lämpligt antal slumpvis utvalda stockar från varje sändning.
3. Om inspektionerna inte visar att sändningen fullständigt uppfyller villkoren i artikel 2.1 skall hela sändningen avvisas och avlägsnas från gemenskapen.
Kommissionen och de behöriga officiella organen i alla medlemsstater skall omedelbart underrättas om uppgifterna om den berörda sändningen.
Artikel 5
1. Stockarna skall endast lagras på platser som har anmälts till och godkänts av behörigt officiellt organ i den berörda medlemsstaten och som har lämpliga anordningar för våtlagring som är tillgängliga under den tid som anges i punkt 2.
2. Stockarna skall hållas under ständig våtlagring, med början senast vid lövsprickningen i närliggande ekbestånd.
3. Närliggande ekbestånd skall av de behöriga officiella organen regelbundet inspekteras för symtom på Ceratocystis fagacearum (Bretz) Hunt med lämpliga intervall.
Om symtom som kan ha orsakats av Ceratocystis fagacearum (Bretz) Hunt upptäcks skall ytterligare officiella tester utföras på lämpligt sätt för att avgöra huruvida svampen förekommer.
Om förekomst av Ceratocystis fagacearum (Bretz) Hunt bekräftas skall kommissionen omedelbart underrättas om detta.
Artikel 6
1. Stockarna får bearbetas endast vid anläggningar som har anmälts till och godkänts av behörigt officiellt organ.
2. Bark och annat avfall från bearbetningen skall omedelbart destrueras på den plats där bearbetningen sker.
Artikel 7
1. Före införsel skall importören anmäla varje sändning i tillräckligt god tid till behörigt officiellt organ i den medlemsstat där den första lagerplatsen ligger, och lämna följande uppgifter:
a) Mängd stockar.
b) Ursprungsland.
c) Utskeppningshamn.
d) Lossningshamn(ar).
e) Lagerplats(er).
f) Plats(er) där bearbetning kommer att äga rum.
2. När en importör anmäler avsikt att föra in en sändning enligt punkt 1 skall han eller hon före införseln underrättas av det behöriga officiella organet om de villkor som anges i detta beslut.
3. Kopior av de uppgifter som avses i punkterna 1 och 2 skall lämnas av det behöriga officiella organet i den berörda medlemsstaten till den myndighet som svarar för tillsyn över lossningshamnen.
Artikel 8
1. Medlemsstaterna får undanta stockar av arten Quercus L. tillhörande viteksgruppen från den gasning som avses i artikel 2.1, förutsatt att följande villkor är uppfyllda:
a) Stockarna skall ingå i sändningar som består endast av stockar från viteksgruppen.
b) Stockarna skall vara identifierade enligt bilaga IV.
c) Stockarna skall skickas från utskeppningshamnen tidigast den 15 oktober och nå lagerplatsen senast den 30 april nästföljande år.
d) Stockarna skall våtlagras.
e) Stockarna får inte föras in i eller genom områden som ligger söder om 45° nordlig bredd; Marseille får dock användas som lossningshamn förutsatt att det tillses att sändningen omedelbart forslas till områden som ligger norr om 45° nordlig bredd.
f) De inspektioner som avses i artikel 4 skall i stället för färgreaktionstestet för påvisande av gasning omfatta ett färgtest för identifiering av vitekstockar enligt bilaga IV, vilket skall utföras på minst 10 % av stockarna från varje sändning efter ett slumpvis urval.
Med avvikelse från punkt c får växtskyddsorganisationen i den medlemsstat där stockarna lagras tillåta att sändningar lossas och förs till våtlager efter den 30 april nästföljande år i enlighet med den punkten, om deras ankomst till lossningshamnen försenats på grund av oförutsedda omständigheter.
2. Punkt 1 skall inte tillämpas på Grekland, Spanien, Italien, Cypern, Malta och Portugal.
Artikel 9
Medlemsstaterna skall till kommissionen och de andra medlemsstaterna överlämna texten till de bestämmelser som de antar i kraft av bemyndigandet i artikel 1.
Artikel 10
De medlemsstater som har utnyttjat det undantag som anges i detta beslut skall rapportera om dess tillämpning senast den 30 juni 2007. Rapporten skall innehålla uppgifter om införd mängd.
I förekommande fall skall en liknande rapport lämnas senast den 30 juni 2009.
Artikel 11
Detta beslut skall upphöra att gälla den 31 december 2010.
Artikel 12
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 18 maj 2005
om ändring för femte gången av beslut 2004/122/EG beträffande vissa skyddsåtgärder mot aviär influensa i Nordkorea
[delgivet med nr K(2005) 1451]
(Text av betydelse för EES)
(2005/390/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/496/EEG av den 15 juli 1991 om fastställande av regler för hur veterinärkontroller skall organiseras för djur som importeras till gemenskapen från tredje land och om ändring av direktiven 89/662/EEG, 90/425/EEG och 90/675/EEG [1], särskilt artikel 18.7 i detta,
med beaktande av rådets direktiv 97/78/EG av den 18 december 1997 om principerna för organisering av veterinärkontroller av produkter från tredje land som förs in i gemenskapen [2], särskilt artikel 22.6 i detta, och
av följande skäl:
(1) I kommissionens beslut 2000/666/EG av den 16 oktober 2000 om djurhälsokrav och utfärdande av veterinärintyg vid import av fåglar utom fjäderfä samt villkor för karantän [3] föreskrivs att medlemsstaterna skall tillåta import av fåglar från tredjeländer som är medlemmar i Internationella byrån för epizootiska sjukdomar (OIE) samt att fåglarna efter införseln till gemenskapen skall placeras i karantän och genomgå provtagning.
(2) Demokratiska folkrepubliken Korea (Nordkorea) har bekräftat ett utbrott av aviär influensa i landet. Eftersom landet är medlem i OIE skall medlemsstaterna enligt beslut 2000/666/EG tillåta import från Nordkorea av ovan nämnda fåglar. Som en försiktighetsåtgärd och med hänsyn till den risk för allvarliga konsekvenser som föreligger i samband med den särskilda stam av aviärt influensavirus som förekommer i övriga Asien bör importen från Nordkorea av dessa fåglar avbrytas.
(3) Enligt Europaparlamentets och rådets förordning (EG) nr 1774/2002 av den 3 oktober 2002 om hälsobestämmelser för animaliska biprodukter som inte är avsedda att användas som livsmedel [4] är import av obearbetade fjädrar och delar av fjädrar med ursprung i Nordkorea tillåten. Med beaktande av det rådande sjukdomsläget i Nordkorea bör dock importen av sådana produkter avbrytas.
(4) Kommissionens beslut 2004/122/EG av den 6 februari 2004 om vissa skyddsåtgärder mot aviär influensa i flera asiatiska länder [5] antogs som en följd av utbrotten av denna sjukdom i ett antal asiatiska länder. I artikel 4 i det beslutet föreskrivs att medlemsstaterna skall avbryta import från vissa tredjeländer av obearbetade fjädrar och delar av fjädrar samt levande fåglar utom fjäderfä enligt definitionen i beslut 2000/666/EG. Med hänsyn till djurs och människors hälsa bör Nordkorea läggas till i uppräkningen av de tredjeländer som avses i artikel 4 i beslut 2004/122/EG.
(5) Beslut 2004/122/EG bör ändras i enlighet med detta.
(6) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 4.1 i beslut 2004/122/EG skall ersättas med följande:
"1. Medlemsstaterna skall avbryta import från Kambodja, Kina inklusive Hongkong, Indonesien, Laos, Malaysia, Nordkorea, Pakistan, Thailand och Vietnam av
- obearbetade fjädrar och delar av fjädrar, och
- "levande fåglar utom fjäderfä" enligt definitionen i beslut 2000/666/EG, inklusive fåglar som åtföljer sin ägare (sällskapsdjur)."
Artikel 2
Medlemsstaterna skall ändra de åtgärder som de tillämpar för import så att dessa överensstämmer med detta beslut och skall omedelbart på lämpligt sätt offentliggöra de åtgärder som har antagits. De skall utan dröjsmål informera kommissionen om dessa.
Artikel 3
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 9 juni 2005
om ändring av beslut 2005/393/EG avseende undantag från utförselförbudet för inhemska förflyttningar av djur från restriktionszonerna
[delgivet med nr K(2005) 1689]
(Text av betydelse för EES)
(2005/434/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 2000/75/EG av den 20 november 2000 om fastställande av särskilda bestämmelser om åtgärder för bekämpning och utrotning av bluetongue [1], särskilt artikel 9.1 c och artikel 19 tredje stycket i detta, och
av följande skäl:
(1) I direktiv 2000/75/EG fastställs kontrollregler och åtgärder för bekämpning av bluetongue i gemenskapen, däribland inrättande av skydds- och övervakningszoner och förbud mot förflyttning av djur från dessa zoner.
(2) I kommissionens beslut 2005/393/EG [2] avgränsas geografiska områden inom vilka medlemsstaterna skall upprätta skydds- och övervakningszoner (restriktionszoner) när det gäller bluetongue. I beslutet fastställs även villkoren för att vissa förflyttningar av djur, sperma, ägg och embryon från dessa djur kan undantas från utförselförbudet i direktiv 2000/75/EG (utförselförbudet).
(3) När en hjord har vaccinerats i enlighet med ett vaccinationsprogram har virusspridningen minskats så mycket att förflyttningar av ungdjur från restriktionszonen till anläggningar utanför zonen, där vektorerna är under kontroll, bör anses utgöra en acceptabel risk.
(4) Den 14 mars 2005 lämnade kommissionens arbetsgrupp om OIE:s Terrestrial Animal Health Code en rapport om olika aspekter av de bestämmelser som bör tillämpas på förflyttningar av djur när det gäller bluetongue.
(5) Arbetsgruppen kom fram till att viremi som förekommer mer än 60 dagar inte bör anses utgöra en avsevärd risk i samband med förflyttningar av levande djur och därför bör djur som har skyddats mot attacker av vektorer i mer än 60 dagar anses säkra.
(6) Arbetsgruppen kom därutöver fram till att eftersom 28 dagar är den maximala perioden för serokonversion efter en infektion, är ett djur säkert när det har skyddats mot attacker av vektorer under en period på mer än 28 dagar och det har testats serologiskt med negativt resultat vid endast ett tillfälle efter denna 28-dagarsperiod.
(7) Arbetsgruppen kom slutligen fram till att eftersom ett virologiskt test alltid är positivt sju dagar efter infektionen är ett djur säkert när det har skyddats mot attacker av vektorer i mer än sju dagar och det har testats virologiskt med negativt resultat vid ett tillfälle efter denna sjudagarsperiod.
(8) Beslut 2005/393/EG bör därför ändras i enlighet med detta.
(9) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Ändringar i beslut 2005/393/EG
Direktiv 2005/393/EG ändras på följande sätt:
1. Artikel 3.2 skall ersättas med följande:
"2. De behöriga myndigheterna skall undanta inhemska förflyttningar enligt punkt 1 från utförselförbudet om
a) djuren härstammar från en hjord som vaccinerats i enlighet med ett vaccinationsprogram som antagits av den behöriga myndigheten, och
b) djuren
i) har vaccinerats mot den eller de serotyper som förekommer eller eventuellt förekommer i det epidemiologiskt relevanta ursprungsområdet mer än 30 dagar men mindre än tolv månader före dagen för förflyttningen, eller
ii) är mindre än två månader gamla dagen för förflyttningen och skall sändas till en anläggning för uppfödning; en sådan anläggning skall vara skyddad mot attacker av vektorer och registrerad hos den behöriga myndigheten som uppfödningsanläggning."
2. I bilaga II skall del A ersättas med följande:
"A. Levande djur skall ha skyddats från attacker av Culicoides
1. under minst 60 dagar före dagen för förflyttningen, eller
2. under minst 28 dagar före dagen för förflyttning och under den perioden med negativt resultat ha genomgått ett serologiskt test för påvisande av antikroppar mot bluetongue-virus, som ett kompetitivt ELISA-test för påvisande av antikroppar mot bluetongue eller ett AGID-test, varvid testet utfördes på prov som tagits minst 28 dagar efter dagen då perioden för skyddet mot attacker från vektorer började, eller
3. under minst sju dagar före dagen för förflyttning och skall under den perioden med negativt resultat ha genomgått test för isolering av bluetongue-virus eller polymeraskedjereaktionstest, varvid testet utfördes på blodprov som tagits minst sju dagar efter dagen då perioden för skyddet mot attacker från vektorer började, och
4. under transporten till avsändningsplatsen."
Artikel 2
Tillämpning
Detta beslut skall tillämpas från och med den 4 juli 2005.
Artikel 3
Adressater
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 16 september 2005
om ändring av tillägget till bilaga XIV till 2003 års anslutningsakt beträffande vissa anläggningar inom köttsektorn i Slovakien
[delgivet med nr K(2005) 3451]
(Text av betydelse för EES)
(2005/661/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Anslutningsakten för Tjeckien, Estland, Cypern, Lettland, Litauen, Ungern, Malta, Polen, Slovenien och Slovakien [1], särskilt kapitel 5 avsnitt B led d i bilaga XIV till denna, och
av följande skäl:
(1) I kapitel 5 avsnitt B led a i bilaga XIV till 2003 års anslutningsakt fastställs att de strukturella kraven i bilaga I till rådets direktiv 64/433/EEG av den 26 juni 1964 om hygienproblem som påverkar handeln med färskt kött inom gemenskapen [2] samt i bilagorna A och B till rådets direktiv 77/99/EEG av den 21 december 1976 om hygienproblem som påverkar handeln med köttprodukter inom gemenskapen [3], fram till och med den 31 december 2006 inte skall gälla för de anläggningar i Slovakien som förtecknas i tillägget [4] till bilaga XIV till anslutningsakten, med förbehåll för vissa villkor.
(2) Tillägget till bilaga XIV till 2003 års anslutningsakt har ändrats genom kommissionens beslut 2004/463/EG [5] och 2005/189/EG [6].
(3) Enligt ett officiell uttalande från den behöriga slovakiska myndigheten har tre köttanläggningar slutfört sin uppgradering och uppfyller nu kraven enligt gemenskapslagstiftningen. Dessa anläggningar bör därför utgå från förteckningen över anläggningar med övergångsbestämmelser.
(4) En köttanläggning i förteckningen över anläggningar med övergångsbestämmelser har gjort avsevärda ansträngningar för att uppfylla de strukturella krav som fastställs i gemenskapslagstiftningen. Denna anläggning kan emellertid på grund av exceptionella tekniska problem inte avsluta sin uppgradering inom den föreskrivna tidsfristen. Anläggningen bör därför få mer tid på sig för att avsluta uppgraderingen.
(5) Tillägget till bilaga XIV till 2003 års anslutningsakt bör därför ändras i enlighet med detta. För tydlighetens skull bör förteckningen ersättas.
(6) Ständiga kommittén för livsmedelskedjan och djurhälsa har informerats om de åtgärder som föreskrivs i detta beslut.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Tillägget till bilaga XIV till 2003 års anslutningsakt skall ersättas med bilagan till detta beslut.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 20 oktober 2005
om ändring av beslut 2005/693/EG om vissa skyddsåtgärder i samband med aviär influensa i Ryssland
[delgivet med nr K(2005) 4176]
(Text av betydelse för EES)
(2005/740/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA BESLUT
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/496/EEG av den 15 juli 1991 om fastställande av regler för hur veterinärkontroller skall organiseras för djur som importeras till gemenskapen från tredje land och om ändring av direktiven 89/662/EEG, 90/425/EEG och 90/675/EEG [1], särskilt artikel 18.1 och 18.6,
med beaktande av rådets direktiv 97/78/EG av den 18 december 1997 om principerna för organisering av veterinärkontroller av produkter från tredje land som förs in i gemenskapen [2], särskilt artikel 22.1 och 22.5, och
av följande skäl:
(1) Aviär influensa är en smittsam virussjukdom hos fjäderfä och fåglar, som orsakar dödlighet och störningar som snabbt kan nå epizootiska proportioner, vilket i sin tur kan utgöra ett allvarligt hot mot djur- och folkhälsan och starkt minska lönsamheten i uppfödningen av fjäderfä.
(2) Kommissionens beslut 2005/693/EG av den 6 oktober 2005 om vissa skyddsåtgärder i samband med aviär influensa i Ryssland [3] antogs efter utbrott av aviär influensa i Ryssland. Genom det beslutet hävs tills vidare importen från Ryssland av fåglar utom fjäderfä.
(3) Genom beslut 2005/693/EG hävs dessutom tills vidare importen av obearbetade fjädrar och obearbetade delar av fjädrar från de regioner i Ryssland som förtecknas i bilaga I till det beslutet. Importen av obearbetade fjädrar och delar av obearbetade fjädrar tillåts dock fortfarande på vissa villkor från de områden i Ryssland som inte förtecknas i bilaga I till det beslutet, även de områden som ligger väster om Uralbergen, där utbrott ännu inte hade förekommit den dag då beslut 2005/693/EG antogs.
(4) Den 19 oktober 2005 underrättade Ryssland kommissionen om ett utbrott av aviär influensa i Tula i det centrala federala distriktet i Ryssland, varifrån inga utbrott tidigare hade rapporterats och från vilket obearbetade fjädrar och delar av obearbetade fjädrar fortfarande får importeras enligt beslut 2005/693/EG.
(5) När det gäller den senaste tidens utbrott av högpatogen aviär influensa orsakad av influensavirus A av subtyp H5N1 i Turkiet, Rumänien och Ryssland, tyder indicier och molekylärepidemiologiska uppgifter starkt på att det aviära influensaviruset spridits till dessa tredjeländer från Centralasien via flyttfåglar. Detta framgår också av den rapport som offentliggjordes den 14 oktober 2005 från ett besök nyligen i Ryssland som genomfördes av Världsorganisationen för djurens hälsa (OIE).
(6) Importen till gemenskapen av obearbetade fjädrar och delar av obearbetade fjädrar bör därför förbjudas från de områden i Ryssland där utbrott av aviär influensa nyligen har förekommit eller där det föreligger en särskild risk, enligt nuvarande kännedom om flyttvägarna för flyttfåglar som kommer från de områden i Centralasien och Sibirien där sjukdomen har konstaterats.
(7) Bilaga I till kommissionens beslut 2005/693/EG bör därför ändras i enlighet med detta.
(8) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I bilaga I till beslut 2005/693/EG skall följande punkter 4, 5, 6 och 7 läggas till:
"4. Centrala federala distriktet
Omfattar följande federationssubjekt: länet Belgorod, länet Bryansk, länet Ivanovo, länet Kaluga, länet Kostroma, länet Kursk, länet Lipetsk, den federala staden Moskva, länet Moskva, länet Oryol, länet Ryazan, länet Smolensk, länet Tambov, länet Tver, länet Tula, länet Vladimir, länet Voronezh, länet Yaroslavl.
5. Södra federala distriktet
Omfattar följande federationssubjekt: Delrepubliken Adygeya, Astrakhan, delrepubliken Chechnya, delrepubliken Dagestan, delrepubliken Ingushetia, delrepubliken Kabardino-Balkaria, delrepubliken Kalmykia, delrepubliken Karachay-Cherkessia, Krasnodar Krai, delrepubliken Nordossetien, Stavropol Krai, länet Rostov, länet Volgograd.
6. Nordvästra federala distriktet
Omfattar följande federationssubjekt: länet Arkhangelsk, delrepubliken Komi, länet Novgorod, länet Pskov, länet Vologda.
7. Federala distriktet Privolzhsky (Volga)
Omfattar följande federationssubjekt: delrepubliken Bashkortostan, delrepubliken Chuvashia, länet Kirov, delrepubliken Mari El, delrepubliken Mordovia, länet Nizhny Novgorod, länet Orenburg, länet Penza, länet Perm, autonoma området Permyakia, länet Samara, länet Saratov, delrepubliken Tatarstan, delrepubliken Udmurtia, länet Ulyanovsk."
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 19 oktober 2005
om tillstånd för medlemsstaterna att förlänga provisoriska tillstånd för de nya verksamma ämnena boscalid, indoxacarb, spinosad och Spodoptera exigua nuclear polyhedrosis virus
[delgivet med nr K(2005) 4002]
(Text av betydelse för EES)
(2005/743/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/414/EEG av den 15 juli 1991 om utsläppande av växtskyddsmedel på marknaden [1], särskilt artikel 8.1 fjärde stycket i detta, och
av följande skäl:
(1) I enlighet med artikel 6.2 i direktiv 91/414/EEG mottog Tyskland i april 2001 en ansökan från BASF AG om införande av det verksamma ämnet boscalid (tidigare kallat nicobifen) i bilaga I till direktiv 91/414/EEG. Genom kommissionens beslut 2002/268/EG [2] bekräftades att dokumentationen var fullständig och i princip kunde anses uppfylla uppgiftskraven i bilagorna II och III till det direktivet.
(2) I oktober 1997 mottog Nederländerna en ansökan från DuPont de Nemours rörande indoxacarb (tidigare kallat DPX-KN128). Genom kommissionens beslut 98/398/EG [3] bekräftades att dokumentationen var fullständig och i princip kunde anses uppfylla uppgiftskraven i bilagorna II och III till direktivet.
(3) I juli 1999 mottog Nederländerna en ansökan från Dow Agrosciences rörande spinosad. Genom kommissionens beslut 2000/210/EG [4] bekräftades att dokumentationen var fullständig och i princip kunde anses uppfylla uppgiftskraven i bilagorna II och III till direktivet.
(4) I juli 1996 mottog Nederländerna en ansökan från Biosys rörande Spodoptera exigua nuclear polyhedrosis virus. Genom kommissionens beslut 97/865/EG [5] bekräftades att dokumentationen var fullständig och i princip kunde anses uppfylla uppgiftskraven i bilagorna II och III till direktivet.
(5) Bekräftelsen av att dokumentationen var fullständig var nödvändig för att en detaljerad granskning av ärendena skulle kunna äga rum, och för att medlemsstaterna skulle kunna utfärda provisoriska tillstånd för högst tre år för de växtskyddsmedel som innehåller de verksamma ämnena i fråga samtidigt som villkoren i artikel 8.1 i direktiv 91/414/EEG uppfylls, särskilt kravet på att en detaljerad utvärdering av det verksamma ämnet och av växtskyddsmedlet skall göras i enlighet med direktivets bestämmelser.
(6) Effekterna av dessa verksamma ämnen på människors hälsa och på miljön har bedömts i enlighet med artikel 6.2 och 6.4 i direktiv 91/414/EEG för de användningsområden som har föreslagits av de respektive sökande företagen. De medlemsstater som handlägger ärendena lade fram sina utkast till utvärderingsrapporter för kommissionen den 22 november 2002 (boscalid), den 7 februari 2000 (indoxacarb), den 5 mars 2001 (spinosad) respektive den 19 november 1999 (Spodoptera exigua nuclear polyhedrosis virus).
(7) Sedan de föredragande medlemsstaterna lämnade in utkasten till utvärderingsrapporter har det blivit nödvändigt att begära ytterligare upplysningar från de sökande och att låta de föredragande medlemsstaterna granska uppgifterna och lämna in en bedömning av ärendet. Granskningen av ärendena pågår därför fortfarande och kommer inte att kunna avslutas inom den tid som anges i direktiv 91/414/EEG.
(8) Eftersom utvärderingen hittills inte har gett någon anledning till oro bör medlemsstaterna få möjlighet att förlänga provisoriska tillstånd för de växtskyddsmedel som innehåller dessa verksamma ämnen med 24 månader i enlighet med artikel 8 i direktiv 91/414/EEG, så att granskningen av ärendena kan fortsätta. Utvärderingen och beslutet om att eventuellt införa de verksamma ämnena i fråga i bilaga I kommer att ha avslutats inom 24 månader.
(9) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från Ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Medlemsstaterna får förlänga provisoriska tillstånd för de växtskyddsmedel som innehåller boscalid, indoxacarb, spinosad eller Spodoptera exigua nuclear polyhedrosis virus med högst 24 månader från och med den dag detta beslut antas.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 8 december 2005
om beviljande av ett undantag på begäran av Nederländerna i enlighet med rådets direktiv 91/676/EEG om skydd mot att vatten förorenas av nitrater från jordbruket
[delgivet med nr K(2005) 4778]
(Endast den nederländska texten är giltig)
(2005/880/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR FATTAT DETTA BESLUT
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/676/EEG av den 12 december 1991 om skydd mot att vatten förorenas av nitrater från jordbruket [1], särskilt bilaga III, stycke 2 b, och
av följande skäl:
(1) Om mängden gödsel som en medlemsstat avser att sprida per hektar och år skiljer sig från den mängd som anges i de inledande meningarna i punkt 2 samt i punkt 2 a i bilaga 3 till direktiv 91/676/EEG, skall den fastställas så att den inte inverkar på möjligheten att uppnå de mål som anges i artikel 1 i det direktivet och skall bestämmas på grundval av objektiva kriterier, exempelvis lång växtperiod och grödor med stor kväveupptagningsförmåga.
(2) Den 8 april 2005 lämnade Nederländerna till kommissionen in en begäran om undantag enligt punkt 2 b i bilaga III till direktiv 91/676/EEG.
(3) Undantaget rör Nederländernas planer på att tillåta användning av 250 kg kväve per hektar och år från stallgödsel i lantbruk med minst 70 % vall- och betesmark. Undantaget berör cirka 25000 gårdar och cirka 900000 hektar i Nederländerna.
(4) Nederländerna har antagit den lagstiftning som genomför direktiv 91/676/EEG och som även gäller det begärda undantaget.
(5) Den nederländska lagstiftning som genomför direktiv 91/676/EEG omfattar tillämpningsstandarder för både kväve och fosfat. Tillämpningsnormer för fosfat har som mål att det senast 2015 skall uppnås jämvikt i fråga om tillförsel och upptagning av kväve vid gödsling.
(6) Nederländerna behandlade frågan om näringsämnesöverskott från gödsel och mineraliska gödselmedel med hjälp av flera politiska instrument och under perioden 1992–2002 minskade man antalet nötkreatur med 17 %, grisar med 14 % och får och getter med 21 %. Kväve och fosfor i gödsel minskade med 29 respektive 34 % under perioden 1985–2002. Kväve- och fosforöverskotten minskade med 25 respektive 37 % under perioden 1992–2002.
(7) Enligt uppgifter om vattenkvaliteten sjunker nitrathalten i grundvatten och i ytvatten. I ytvatten sjunker även fosforhalten.
(8) Av de tekniska och vetenskapliga dokument som åtföljer den nederländska begäran framgår att den föreslagna mängden på 250 kg kväve per hektar och år från gödsel från nötkreatur på lantbruk med minst 70 % är förenlig med nivån på 11,3 mg/l N (vilket motsvarar 50 mg/l NO3) i vatten i alla marktyper och med ett uppskattningsvis obefintligt fosforöverskott, vid optimala förvaltningsvillkor.
(9) De tekniska och vetenskapliga dokumenten visar vidare att den föreslagna mängden 250 kg kväve per hektar och år från stallgödsel på lantbruk med minst 70 % vall- och betesmark kan motiveras med hjälp av objektiva kriterier som lång växtsäsong och grödor med högt kväveupptag.
(10) Kommissionen anser därför att den mängd gödsel som Nederländerna begärt undantag för inte påverkar uppfyllandet av målen enligt direktiv 91/676/EEG under förutsättning att vissa stränga villkor uppfylls.
(11) Det rör sig bland annat om följande mål: fastställandet av gödselplaner för varje jordbruk, dokumentation om gödslingsmetoder i form av gödslingsplaner, periodiska markanalyser, täckgröda på vintern för fodermajs, särskilda bestämmelser om gräsbrytning, förbud mot gödsling för gräsbrytning och justering av gödselmängderna för att ta hänsyn till påverkan från baljväxter. Syftet är att se till att gödslingen sker med växternas behov som grundval och att kväveförlusterna till vatten minskas eller hindras.
(12) För att undvika att det begärda undantaget leder till ökad tillförsel bör de behöriga myndigheterna se till att de mängder kväve och fosfor som uppstår vid gödselproduktionen inte överstiger nivån för år 2002 i enlighet med det handlingsprogram Nederländerna skall genomföra.
(13) Det begärda undantaget bör följaktligen beviljas.
(14) Detta beslut bör tillämpas i samband med Nederländernas handlingsprogram för 2006 till 2009.
(15) Åtgärderna i detta beslut är förenliga med yttrandet från den kvävekommitté som har inrättats i enlighet med artikel 9 i direktiv 91/676/EEG.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Det undantag som Nederländerna begärde i en skrivelse av den 8 april 2005 för att tillåta en högre nivå stallgödsel än vad som fastställs i de inledande meningarna i punkt 2 och i punkt 2 a i bilaga III till direktiv 91/676/EEG beviljas under förutsättning att de villkor som anges i det här beslutet uppfylls.
Artikel 2
Definitioner
I detta beslut används följande beteckningar med de betydelser som här anges:
jordbruksföretag med betesdrift : gård där minst 70 % av den areal som är tillgänglig för gödselspridning utgörs av gräs.
betesdjur : nötkreatur (med undantag av gödkalvar), får, getter, hästar, åsnor, hjort och rådjur samt vattenbuffel.
jordbruksmark : den areal som ägs, arrenderas eller förvaltas av lantbrukaren genom ett skriftligt kontrakt och för vilken han/hon har ett direkt förvaltningsansvar.
gräs : permanent eller tillfälligt gräsbevuxen mark (tillfälligt innebär i regel mindre än fyra år).
Artikel 3
Tillämpningsområde
Det här beslutet gäller på individuell basis och på de villkor som anges i artiklarna 4, 5 och 6 för jordbruksföretag med betesdrift.
Artikel 4
Årligt godkännande och åtagande
1. Lantbrukare som vill utnyttja ett undantag skall en gång per år lämna in en ansökan till behörig myndighet.
2. Tillsammans med denna årliga ansökan skall de skriftligen åta sig att uppfylla villkoren i artiklarna 5 och 6.
3. De behöriga myndigheterna skall se till att ansökningarna om undantag och redovisningar av gödselmedel granskas. Om den myndighetskontroll av de ansökningar som avses i punkt 1 avslöjar att villkoren i artiklarna 5 och 6 inte är uppfyllda, skall den sökande informeras om detta. I sådana fall skall ansökan inte godkännas.
Artikel 5
Spridning av stallgödsel och annan gödsel
1. Den mängd gödsel från betesdjur, inklusive från djuren själva, som varje år sprids på jordbruksföretag med betesdrift skall inte överstiga den mängd gödsel som innehåller 250 kg kväve per år, i enlighet med villkoren i punkterna 2–7.
2. Den totala kvävetillförseln skall motsvara näringsbehovet hos den berörda grödan och kvävetillförseln från marken.
3. För varje jordbruksföretag skall det finnas en gödslingsplan som beskriver växtföljden och den planerade spridningen av gödsel, kväve- och fosfathaltigt gödsel. Planen skall finnas på jordbruksföretaget senast den 1 februari och omfatta följande:
a) Antalet kreatur, en beskrivning av lagringslokalerna, inklusive volymen på lagringskapaciteten för gödsel.
b) En beräkning av kväve- och fosforhalten i det stallgödsel (med avdrag för förluster vid lagring) som produceras vid jordbruksföretaget.
c) Växtföljden och arealen för varje gröda, inklusive en skiss över de enskilda åkrarnas placering.
d) Grödornas förväntade kväve- och fosforbehov.
e) Mängd och typ av gödsel som levererats till underleverantörer och som inte används på jordbruksföretaget.
f) Mängd inköpt gödsel som används på jordbruksföretaget.
g) En beräkning av bidraget från mineralisering av organiskt material, baljväxter och atmosfäriskt nedfall samt den mängd kväve som finns i marken vid den tidpunkt då grödan börjar använda den i nämnvärd utsträckning.
h) Tillförsel av kväve och fosfor från gödsling på varje åker (jordlotter som är likartade i fråga om grödor och jordtyp).
i) Tillförsel av kväve och fosfor från konstgödsel och andra gödselmedel på varje åker.
j) Kalkyler för bedömning av överensstämmelse med normerna för användning av kväve och fosfor.
Planerna skall ses över senast sju dagar efter det att ändringar i jordbruksmetoderna företagits, för att garantera att de överensstämmer med de använda jordbruksmetoderna.
4. Gödselredogörelser skall finnas på varje jordbruksföretag. De skall skickas till den behöriga myndigheten för varje kalenderår och skall innehålla följande:
a) Grödarealen.
b) Antal och typ av kreatur.
c) Gödselproduktion per djur.
d) Mängd gödsel som jordbruksföretaget köper in.
e) Mängd gödsel som levereras från jordbruksföretaget och vem mottagaren är.
5. De jordbruksföretag med betesdrift som utnyttjar ett enskilt undantag skall godta att ansökan och gödselredogörelser kan komma att kontrolleras.
6. Periodiska analyser av kväve- och fosfalthalten i jorden skall ske på de jordbruksföretag som gynnas av ett enskilt undantag minst vart fjärde år för varje likartat område på jordbruksföretaget, i fråga om växtföljden och jordegenskaperna.
Kväveanalyser i fråga om mineraliskt kväve och parametrar för att bedöma kvävetillförseln från mineralisering av organiskt material skall ske efter gräsbrytning för varje likartat område på jordbruksföretaget.
Minimikravet för analyserna i första och andra stycket är en analys per fem hektar mark.
7. Gödselspridning får inte ske under hösten före odling av gräs.
Artikel 6
Marktäcke
1. 70 % eller mer av de arealer som är disponibla för gödselspridning på jordbruksföretagen skall odlas med gräs. Jordbrukare som omfattas av ett individuellt undantag skall vidta följande åtgärder:
a) Efter majs skall sand- och lössjordar odlas med gräs eller andra grödor som garanterar marktäckning under vintern, i syfte att väsentligt minska läckagepotentialen.
b) Fånggrödor skall inte brytas före den 1 februari så att jordbruksmarken garanteras ett växttäcke som återför höstens nitratförluster från de lägre markskikten och begränsar vinterförlusterna.
c) Gräs på sand- och lössjordar skall brytas på våren.
d) Gräs som brutits skall på alla jordarter omedelbart följas av en gröda med högt nitratbehov och gödslingen skall baseras på jordanalys avseende mineraliskt kväve och andra parametrar som erbjuder referenser för uppskattning av mängden kväve som avges från mineralisering av organiskt material i jorden.
e) Om växtföljden omfattar baljväxter eller andra växter som fixerar atmosfäriskt kväve skall gödselspridningen minskas i motsvarande grad.
2. Genom undantag från punkt c skall gräsbrytning vara tillåtet under hösten för plantering av blomsterlökar.
Artikel 7
Åtgärder mot gödselproduktion
De nationella myndigheterna skall se till att gödselproduktionen varken när det gäller kväve eller fosfor överstiger produktionsnivån för 2002.
Artikel 8
Övervakning
1. Varje år skall den behöriga myndigheten framställa kartor som visar andelen jordbruksföretag med betesdrift, andelen djur och andelen jordbruksmark (uttryckt i procent) som omfattas av det individuella undantaget i varje kommun, och kartorna skall uppdateras varje år.
Kartorna skall skickas in till kommissionen en gång om året från och med andra kvartalet 2006.
2. Ett övervakningsnät av provtagningpunkter i markvatten, vattendrag och ytnära grundvatten skall upprättas och användas för övervakning av undantagen.
Övervakningsnätet, i vilket minst 300 jordbruksföretag som omfattas av individuellt undantag skall ingå, skall vara representativt för alla jordarter (ler-, torv-, sand- och sandiga lössjordar) samt för gödslingsmetoder och växtföljd. Övervakningsnätets sammansättning får inte ändras under tillämpningsperioden för det här beslutet.
3. Undersökningar och löpande näringsämnesanalyser skall tillhandahålla uppgifter om lokal markanvändning, växtföljd och jordbruksmetoder på jordbruksföretag som omfattas av individuella undantag. Dessa uppgifter kan användas för modellbaserade beräkningar av omfattningen av nitratläckaget och fosforförlusterna från åkrar där upp till 250 kg kväve i stallgödsel sprids per hektar och år.
4. Ytnära grundvatten, markvatten, dräneringsvatten och vattendrag på jordbruksföretag som ingår i övervakningsnätet skall tillhandahålla uppgifter om koncentrationen av nitrat och fosfor i vatten som lämnar rotzonen och tränger ut i grundvatten- och ytvattensystemet.
5. En stärkt övervakning skall riktas mot områden med avrinning från jordbruket i sandjordar.
Artikel 9
Kontroller
1. Den behöriga nationella myndigheten skall göra administrativa kontroller av alla jordbruksföretag som omfattas av ett individuellt undantag, i syfte att bedöma om den maximala mängden på 250 kg kväve per hektar och år från betesgödsel har efterlevts och att normerna för spridning av kväve och fosfat och villkoren för markanvändning har iakttagits.
2. Det skall upprättas ett inspektionsprogram grundat på riskanalys samt på resultaten av kontrollerna från tidigare år och resultaten av allmänna stickprovskontroller av tillämpningen av den lagstiftning genom vilken direktiv 91/676/EEG genomförs.
Minst 5 % av de jordbruksföretag som omfattas av individuellt undantag skall kontrolleras med avseende på markanvändning, antal djur och gödselproduktion.
Minst 3 % av jordbruksföretagen skall omfattas av åkerinspektioner för kontroll av om villkoren enligt artiklarna 5 och 6 iakttas.
Artikel 10
Rapportering
1. Den behöriga myndigheten skall överlämna övervakningsresultaten till kommissionen varje år, och i dessa skall ingå en konkret rapport om utvärderingsrutiner (kontroller på jordbruksföretagen, inklusive uppgifter om jordbruksföretag som inte uppfyller kraven baserat på resultaten från de administrativa åkerinspektionerna) och vattenkvalitetens utveckling (baserat på övervakning av läckage från rotzonen, yt/grundvattenkvaliteten och modellbaserade beräkningar).
Den första rapporten skall skickas in senast i mars 2007 och efter det varje år senast i mars 2008, 2009 och 2010.
2. Förutom uppgifterna enligt punkt 1 skall rapporten innehålla följande:
a) Uppgifter rörande gödsling för alla jordbruksföretag som omfattas av undantaget,
b) utvecklingen i fråga om antalet djur per kategori i Nederländerna och på de jordbruksföretag som omfattas av undantaget,
c) utvecklingen inom den nationella gödselproduktionen när det gäller kväve och fosfater i gödsel,
d) en sammanfattning av resultaten av kontrollerna knutna till utsöndringskoefficienten för gris- och fjäderfägödsel på nationell nivå.
3. De erhållna resultaten kommer att beaktas av kommissionen vid en eventuell ny begäran om undantag från de holländska myndigheterna.
4. Den behöriga myndigheten skall utarbeta en årlig rapport om gödsling och avkastning för olika jordarter och grödor och skicka in den till kommissionen, så att denna får uppgifter om förvaltningen på de jordbruksföretag med betesdrift som omfattas av undantag och om i vilken mån förvaltningen är optimal.
Artikel 11
Tillämpning
Detta beslut skall tillämpas från och med den 1 januari 2006.
Det skall löpa ut den 31 december 2009.
Artikel 12
Detta beslut riktar sig till Konungariket Nederländerna.
Kommissionens Direktiv 2005/30/EG
av den 22 april 2005
om ändring, för att anpassa dem till den tekniska utvecklingen, av Europarlamentets och rådets direktiv 97/24/EG och 2002/24/EG avseende typgodkännande av två- och trehjuliga motorfordon
(Text av betydelse för EES)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA DIREKTIV
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av Europaparlamentets och rådets direktiv 97/24/EG av den 17 juni 1997 om vissa komponenter och karakteristiska egenskaper hos två- eller trehjuliga motorfordon [1], särskilt artikel 7 i detta,
med beaktande av Europaparlamentets och rådets direktiv 2002/24/EG av den 18 mars 2002 om typgodkännande av två- och trehjuliga motorfordon och om upphävande av rådets direktiv 92/61/EEG [2], särskilt artikel 17 i detta, och
av följande skäl:
(1) Direktiv 97/24/EG är ett av särdirektiven inom ramen för det förfarande för EG typgodkännande som fastställs i direktiv 2002/24/EG.
(2) Tekniska regler för typgodkännande av ersättningskatalysatorer som separata tekniska enheter bör införas för att säkerställa att utsläppen håller en lämplig nivå. Regler bör införas för att främja tillämpningen i medlemsstaterna genom krav på märkning av ersättningskatalysatorer och deras förpackningar.
(3) Typgodkännandekoden för medlemsstaterna Malta och Cypern i bilaga V till direktiv 2002/24/EG bör uppdateras.
(4) Direktiven 97/24/EG och 2002/24/EG bör därför ändras i enlighet med detta.
(5) Bestämmelserna i detta direktiv är förenliga med yttrandet från Kommittén för anpassning till den tekniska utvecklingen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE:
Artikel 1
Texten som bifogas direktiv 97/24/EG skall ändras i enlighet med bilaga I till det här direktivet.
Artikel 2
Bilagorna II och V till direktiv 2002/24/EG skall ändras i enlighet med bilaga II till det här direktivet.
Artikel 3
1. När det gäller nya ersättningskatalysatorer som är avsedda att monteras på fordon som har erhållit typgodkännande i enlighet med direktiv 97/24/EG, får medlemsstaterna från och med den 18 maj 2006 inte längre
a) vägra att bevilja EG-typgodkännande i enlighet med artikel 4.1 i direktiv 2002/24/EG, eller
b) förbjuda försäljning eller installation i fordon.
2. Från och med den 18 maj 2006 får medlemsstaterna inte längre, av skäl som hänför sig till åtgärder mot luftföroreningar, tillåten ljudnivå eller åtgärder för att förhindra otillåtna förändringar, bevilja EG-typgodkännande enligt artikel 4.1 i direktiv 2002/24/EG för en ny ersättningskatalysator om den inte uppfyller bestämmelserna i direktiv 97/24/EG, ändrat genom det här direktivet.
Artikel 4
1. Medlemsstaterna skall anta och offentliggöra de lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 17 maj 2006. De skall genast överlämna texten till dessa bestämmelser till kommissionen tillsammans med en jämförelsetabell för dessa bestämmelser och bestämmelserna i detta direktiv.
De skall tillämpa dessa bestämmelser från och med den 18 maj 2006.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texterna till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av det här direktivet.
Artikel 5
Detta direktiv träder i kraft den tjugonde dagen efter det att det har offentliggjorts i Europeiska unionens officiella tidning.
Artikel 6
Detta direktiv riktar sig till medlemsstaterna.
Europaparlamentets och rådets direktiv 2005/65/EG
av den 26 oktober 2005
om ökat hamnskydd
(Text av betydelse för EES)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 80.2,
med beaktande av kommissionens förslag,
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande [1],
med beaktande av Regionkommitténs yttrande [2],
i enlighet med förfarandet i artikel 251 i fördraget [3], och
av följande skäl:
(1) Säkerhetstillbud till följd av terrorism hör till de allvarligaste hoten mot de ideal i fråga om demokrati, frihet och fred som utgör själva grunden för Europeiska unionen.
(2) Människor, infrastruktur och utrustning i hamnar bör skyddas mot säkerhetstillbud och de förödande effekter sådana kan få. Ett sådant skydd gagnar både dem som använder transporterna och ekonomin och samhället som helhet.
(3) Den 31 mars 2004 antog Europaparlamentet och Europeiska unionens råd förordning (EG) nr 725/2004 om förbättrat sjöfartsskydd på fartyg och i hamnanläggningar [4]. Åtgärderna för ökat sjöfartsskydd enligt den förordningen är bara ett led i de åtgärder som krävs för att man skall uppnå tillräckligt hög skyddsnivå i hela transportkedjan med koppling till sjöfarten. Den förordningens räckvidd är begränsad till skyddsåtgärder ombord på fartyg och till samverkan mellan fartyg och hamn.
(4) För säkerställande av bästa möjliga skydd för sjöfarts- och hamnverksamhet bör det införas hamnskyddsåtgärder som omfattar varje hamn inom de gränser som den berörda medlemsstaten har fastställt så att de skyddsåtgärder som vidtagits med tillämpning av förordning (EG) nr 725/2004 förbättras genom ökat skydd i områden med hamnverksamhet. Åtgärderna bör gälla alla hamnar med en eller flera av de hamnanläggningar som omfattas av förordning (EG) nr 725/2004.
(5) Skyddsmålet i detta direktiv bör kunna uppnås genom att lämpliga åtgärder antas utan att det påverkar medlemsstaternas bestämmelser inom området nationell säkerhet och de åtgärder som kan vidtas enligt avdelning VI i fördraget om Europeiska unionen.
(6) Medlemsstaterna bör ta ingående skyddsutredningar till hjälp när de fastställer de exakta gränserna för det skyddsvärda hamnområdet och fattar beslut om vilka åtgärder som krävs för att säkerställa tillräckligt hamnskydd. Beroende på gällande skyddsnivå och skillnaderna mellan olika hamnområdens riskprofiler bör olika åtgärder vidtas.
(7) Medlemsstaterna bör godkänna sådana hamnskyddsplaner som omsätter hamnskyddsutredningens resultat i praktiken. För att skyddsåtgärderna verkligen skall fungera krävs det dessutom regelbundna övningar och en tydlig uppgiftsdelning mellan de berörda parterna. En hamnskyddsplan som innehåller bestämmelser om uppgiftsdelning och övningar anses avsevärt öka effektiviteten av både förebyggande och korrigerande hamnskyddsåtgärder.
(8) Ro-ro-fartyg är särskilt sårbara för säkerhetstillbud, i synnerhet om fartygen medför både passagerare och gods. Lämpliga åtgärder grundade på riskanalyser bör vidtas för att säkerställa att bil- och godsfordon som transporteras på ett ro-ro-fartyg på nationella och internationella rutter inte utgör någon risk för fartyg, passagerare, fartygsbesättning eller gods. Åtgärderna bör genomföras på ett sådant sätt att verksamhetsflödet hämmas i så liten omfattning som möjligt.
(9) Medlemsstaterna bör kunna inrätta hamnskyddskommittéer som har till uppgift att komma med praktiska råd i de hamnar som omfattas av detta direktiv.
(10) Medlemsstaterna bör se till att alla berörda parter är helt införstådda med ansvarsfördelningen i fråga om hamnskyddet. Medlemsstaterna bör övervaka skyddsbestämmelsernas efterlevnad, inrätta en myndighet med tydligt ansvar för landets samtliga hamnar, ansvara för godkännandet av alla skyddsutredningar och skyddsplaner för sina hamnar, fastställa och meddela skyddsnivåer på lämpligt sätt samt se till att åtgärderna meddelas, genomförs och samordnas väl.
(11) Medlemsstaterna bör godkänna utredningar och planer och övervaka genomförandet i sina hamnar. För att minimera störningarna av hamnverksamheten och den administrativa bördan för övervakningsorganen, bör kommissionens övervakning av genomförandet av detta direktiv göras samtidigt som de inspektioner som föreskrivs i artikel 9.4 i förordning (EG) nr 725/2004.
(12) Medlemsstaterna bör se till att en sambandspunkt för hamnskydd sköter förbindelserna mellan kommissionen och medlemsstaterna. De bör informera kommissionen om vilka hamnar som omfattas av detta direktiv på grundval av de skyddsutredningar som gjorts.
(13) Ett effektivt och enhetligt genomförande av åtgärderna inom ramen för en denna skyddspolitik väcker viktiga frågor om finansieringsaspekten. Finansieringen av extra skyddsåtgärder bör inte leda till att konkurrensen snedvrids. Senast den 30 juni 2006 bör kommissionen för Europaparlamentet och rådet lägga fram resultaten av en undersökning om kostnaderna för de åtgärder som vidtas enligt detta direktiv, och särskilt behandla frågan om hur kostnaderna fördelas mellan de offentliga myndigheterna, hamnmyndigheterna och operatörerna.
(14) Detta direktiv respekterar de grundläggande rättigheter och principer som erkänns framför allt i Europeiska unionens stadga om de grundläggande rättigheterna.
(15) De åtgärder som är nödvändiga för att genomföra detta direktiv bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter [5].
(16) Det bör fastställas ett förfarande för anpassning av detta direktiv med hänsyn till den utveckling som internationella instrument genomgår och, mot bakgrund av gjorda erfarenheter, för anpassning och komplettering av de enskilda bestämmelserna i bilagorna till detta direktiv, utan att direktivets räckvidd utvidgas.
(17) Eftersom målet för detta direktiv, nämligen väl avvägt införande av lämpliga åtgärder på det sjöfarts- och hamnpolitiska området, inte i tillräcklig utsträckning kan uppnås av medlemsstaterna och det därför, på grund av detta direktivs europeiska dimension, bättre kan uppnås på gemenskapsnivå, kan gemenskapen vidta åtgärder i enlighet med subsidiaritetsprincipen i artikel 5 i fördraget. I enlighet med proportionalitetsprincipen i samma artikel går detta direktiv inte utöver vad som är nödvändigt för att uppnå detta mål.
(18) Eftersom detta direktiv gäller kusthamnar bör de skyldigheter som anges i direktivet ej vara tillämpliga för Luxemburg, Slovakien, Tjeckien, Ungern och Österrike.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Syfte
1. Huvudsyftet med detta direktiv är att införa gemenskapsåtgärder för att förbättra hamnskyddet inför hot om säkerhetstillbud.
Detta direktiv skall även säkerställa att sådana skyddsåtgärder som vidtas med tillämpning av förordning (EG) nr 725/2004 drar fördel av ett ökat skydd i hamnar.
2. Åtgärderna enligt punkt 1 skall bestå av följande:
a) Gemensamma grundregler för hamnskyddsåtgärder.
b) En mekanism för genomförande av dessa regler.
c) Lämpliga mekanismer för övervakning av att reglerna följs.
Artikel 2
Räckvidd
1. Detta direktiv fastställer skyddsåtgärder som skall beaktas i hamnar. Medlemsstaterna får tillämpa detta direktiv på områden som har anknytning till hamnarna.
2. De åtgärder som fastställs i detta direktiv skall tillämpas på alla hamnar i en medlemsstat där det finns en eller flera av de hamnanläggningar som omfattas av en godkänd skyddsplan för hamnanläggningar i enlighet med förordning (EG) nr 725/2004. Detta direktiv skall inte tillämpas på militära anläggningar i hamnar.
3. Medlemsstaterna skall för varje hamn fastställa de gränser inom vilka detta direktiv skall vara tillämpligt, med vederbörlig hänsyn tagen till hamnskyddsutredningens resultat.
4. Om en medlemsstat har fastställt gränserna för en hamnanläggning i den betydelse som avses i förordning (EG) nr 725/2004 på ett sådant sätt att den i praktiken omfattar en hamn, skall de relevanta bestämmelserna i förordning (EG) nr 725/2004 ha företräde framför bestämmelserna i detta direktiv.
Artikel 3
Definitioner
I detta direktiv används följande beteckningar med de betydelser som här anges:
1) hamn: ett specificerat land- och vattenområde, med gränser som fastställts av den medlemsstat i vilken hamnen befinner sig, vilket består av sådana anläggningar och sådan utrustning som underlättar kommersiella sjöfartstransporter.
2) samverkan mellan fartyg och hamn: det samspel som sker när ett fartyg direkt och omedelbart berörs av åtgärder som innebär förflyttning av personer eller gods eller tillhandahållande av hamntjänster till eller från fartyget.
3) hamnanläggning: en plats där samverkan mellan fartyg och hamn äger rum. Detta inkluderar, i tillämpliga fall, områden såsom ankarplatser, väntekajer och insegling från sjösidan.
4) sambandspunkt för hamnskydd: det organ som utsetts av varje medlemsstat och som skall utgöra en kontaktpunkt för kommissionen och andra medlemsstater och underlätta, följa upp och informera om genomförandet av de hamnskyddsåtgärder som anges i detta direktiv.
5) hamnskyddsmyndighet: myndighet med ansvar för skyddsfrågor i en viss hamn.
Artikel 4
Samordning med åtgärder enligt förordning (EG) nr 725/2004
Medlemsstaterna skall se till att hamnskyddsåtgärderna enligt detta direktiv noga samordnas med de åtgärder som vidtas med tillämpning av förordning (EG) nr 725/2004.
Artikel 5
Hamnskyddsmyndighet
1. Medlemsstaterna skall för varje hamn som omfattas av detta direktiv utse en hamnskyddsmyndighet. En hamnskyddsmyndighet får utses för flera hamnar.
2. Hamnskyddsmyndigheten skall ansvara för upprättande och genomförande av hamnskyddsplaner som grundar sig på resultatet av hamnskyddsutredningar.
3. Medlemsstaterna får som hamnskyddsmyndighet utse en behörig sjöfartsskyddsmyndighet enligt förordning (EG) nr 725/2004.
Artikel 6
Hamnskyddsutredning
1. Medlemsstaterna skall se till att det för de hamnar som omfattas av detta direktiv görs hamnskyddsutredningar. I samband med utredningarna skall vederbörlig hänsyn tas till de olika hamndelarnas särart och, i de fall där berörda myndigheter i medlemsstaten anser det tillämpligt, även till närliggande områden, om dessa påverkar säkerheten i hamnen, samt till de utredningar för det berörda områdets hamnanläggningar som har gjorts med tillämpning av förordning (EG) nr 725/2004.
2. Varje hamnskyddsutredning skall genomföras med beaktande av de specifika kraven i bilaga I som ett minimum.
3. Hamnskyddsutredningarna kan göras av en erkänd skyddsorganisation som avses i artikel 11.
4. Hamnskyddsutredningarna skall godkännas av den berörda medlemsstaten.
Artikel 7
Hamnskyddsplan
1. Medlemsstaterna skall se till att hamnskyddsplaner utarbetas, upprätthålls och uppdateras mot bakgrund av resultatet av hamnskyddsutredningarna. I planerna skall dels vederbörlig hänsyn tas till de olika hamndelarnas särart, dels de skyddsplaner integreras som har tagits fram för det berörda områdets hamnanläggningar med tillämpning av förordning (EG) nr 725/2004.
2. För var och en av de skyddsnivåer som avses i artikel 8 skall det i hamnskyddsplanerna fastställas
a) vilka förfaranden som skall tillämpas,
b) vilka åtgärder som skall vidtas,
c) vilka insatser som krävs.
3. Varje hamnskyddsplan skall utarbetas med beaktande av de specifika kraven i bilaga II som ett minimum. Hamnskyddsplanen skall vid behov särskilt innehålla skyddsåtgärder som skall tillämpas på passagerare och fordon innan de embarkerar havsgående fartyg som medför passagerare och fordon. När det gäller internationella sjötransporttjänster skall de berörda medlemsstaterna delta i utredningen av skyddet i hamnen.
4. Hamnskyddsplanerna får utarbetas av en erkänd skyddsorganisation som avses i artikel 11.
5. Hamnskyddsplanerna skall godkännas av den berörda medlemsstaten innan de genomförs.
6. Medlemsstaterna skall se till att hamnskyddsplanernas genomförande övervakas. Övervakningen skall samordnas med annan kontrollverksamhet i hamnen.
7. Medlemsstaterna skall sörja för lämpliga övningar med hänsyn till de grundläggande kraven på skyddsutbildningsövningar i bilaga III.
Artikel 8
Skyddsnivåer
1. Medlemsstaterna skall införa ett system med skyddsnivåer för hamnar eller delar av hamnar.
2. Det skall finnas tre skyddsnivåer enligt definitionen i förordning (EG) nr 725/2004:
- Skyddsnivå 1: den nivå på vilken de minst omfattande skyddsåtgärderna alltid skall upprätthållas.
- Skyddsnivå 2: den nivå på vilken tillämpliga ytterligare skyddsåtgärder skall upprätthållas under en viss tidsperiod på grund av en förhöjd risk för säkerhetstillbud.
- Skyddsnivå 3: den nivå på vilken ytterligare specifika skyddsåtgärder skall upprätthållas under en begränsad tidsperiod i samband med att säkerhetstillbud kan förväntas eller är överhängande, även om det kanske inte är möjligt att identifiera något specifikt mål.
3. Medlemsstaterna skall bestämma vilken skyddsnivå som skall gälla för varje hamn eller del av hamn. En medlemsstat får på varje skyddsnivå fastställa att olika skyddsåtgärder skall vidtas i olika delar av hamnen beroende på hamnskyddsutredningens resultat.
4. Medlemsstaterna skall för varje hamn eller del av hamn meddela gällande skyddsnivå och eventuella ändringar av denna till lämplig person eller lämpliga personer.
Artikel 9
Hamnskyddschef
1. En hamnskyddschef skall godkännas av den berörda medlemsstaten för varje hamn. Varje hamn skall om möjligt ha en egen hamnskyddschef, men får, om det är lämpligt, dela skyddschef med andra hamnar.
2. Hamnskyddscheferna skall fungera som kontaktpunkter i hamnskyddsfrågor.
3. Om hamnskyddschefen inte är samma person som hamnanläggningens/hamnanläggningarnas skyddschefer enligt förordning (EG) nr 725/2004, skall ett nära samarbete mellan dem säkerställas.
Artikel 10
Översyn
1. Medlemsstaterna skall se till att hamnskyddsutredningarna och hamnskyddsplanerna ses över vid behov. Översynen skall göras åtminstone en gång vart femte år.
2. Översynsförfarandet skall omfatta artikel 6 eller artikel 7, beroende på omständigheterna.
Artikel 11
Erkänd skyddsorganisation
Medlemsstaterna får utse erkända skyddsorganisationer inom ramen för detta direktiv. Erkända skyddsorganisationer skall uppfylla villkoren i bilaga IV.
Artikel 12
Sambandspunkt för hamnskydd
Medlemsstaterna skall utse en sambandspunkt för hamnskydd. Medlemsstaterna får utse den sambandspunkt för sjöfartsskydd som har utsetts enligt förordning (EG) nr 725/2004. Sambandspunkten för hamnskydd skall till kommissionen överlämna en förteckning över de hamnar som berörs av detta direktiv och informera kommissionen om varje ändring av förteckningen.
Artikel 13
Genomförande och kontroll av efterlevnaden
1. Medlemsstaterna skall införa ett system för att säkerställa adekvat och regelbunden övervakning av hamnskyddsplanerna och deras genomförande.
2. Kommissionen skall, i samarbete med de sambandspunkter som avses i artikel 12, övervaka medlemsstaternas genomförande av detta direktiv.
3. Denna övervakning skall genomföras samtidigt med de inspektioner som föreskrivs i artikel 9.4 i förordning (EG) nr 725/2004.
Artikel 14
Ändringar
Bilagorna I–IV får ändras i enlighet med förfarandet i artikel 15.2, utan att detta direktivs räckvidd utvidgas.
Artikel 15
Kommittéförfarande
1. Kommissionen skall biträdas av den kommitté som inrättats enligt förordning (EG) nr 725/2004.
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i beslut 1999/468/EG tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Den tid som avses i artikel 5.6 i beslut 1999/468/EG skall vara en månad.
3. Kommittén skall själv anta sin arbetsordning.
Artikel 16
Sekretess och spridning av information
1. Vid tillämpningen av detta direktiv skall kommissionen, i enlighet med beslut 2001/844/EG, EKSG, Euratom [6], vidta lämpliga åtgärder för att skydda den sekretessbelagda information som den har tillgång till eller som medlemsstaterna har lämnat till kommissionen.
Medlemsstaterna skall vidta likvärdiga åtgärder i enlighet med gällande nationell lagstiftning.
2. Personal som genomför skyddsinspektioner eller handhar sekretessbelagd information inom ramen för detta direktiv skall genomgå lämplig säkerhetsprövning, som skall utföras av den medlemsstat där den berörda personen är medborgare.
Artikel 17
Sanktioner
Medlemsstaterna skall se till att det finns effektiva, proportionerliga och avskräckande sanktioner för överträdelser av de nationella bestämmelser som antas i enlighet med detta direktiv.
Artikel 18
Genomförande
1. Medlemsstaterna skall sätta i kraft de bestämmelser i lagar och andra författningar som är nödvändiga för att följa detta direktiv senast den 15 juni 2007. De skall genast underrätta kommissionen om detta.
När en medlemsstat antar dessa bestämmelser skall de innehålla en hänvisning till detta direktiv eller åtföljas av en sådan hänvisning när de offentliggörs. Närmare föreskrifter om hur hänvisningen skall göras skall varje medlemsstat själv utfärda.
2. Medlemsstaterna skall till kommissionen överlämna texten till de centrala bestämmelser i nationell lagstiftning som de antar inom det område som omfattas av detta direktiv.
Artikel 19
Utvärderingsrapport
Senast den 15 december 2008 och därefter vart femte år skall kommissionen för Europaparlamentet och rådet lägga fram en utvärderingsrapport som bland annat skall grunda sig på de uppgifter som erhålls enligt artikel 13. Kommissionen skall i rapporten analysera om medlemsstaterna efterlever detta direktiv och hur effektiva de vidtagna åtgärderna är. Vid behov skall kommissionen lägga fram förslag till nya åtgärder.
Artikel 20
Ikraftträdande
Detta direktiv träder i kraft den tjugonde dagen efter det att det har offentliggjorts i Europeiska unionens officiella tidning.
Artikel 21
Adressater
Detta direktiv riktar sig till de medlemsstater som har sådana hamnar som avses i artikel 2.2.
Europaparlamentets och rådets direktiv 2005/82/EG
av den 14 december 2005
om upphävande av rådets direktiv 90/544/EEG om frekvensband för det samordnade införandet av alleuropeisk, landbaserad, allmänt tillgänglig, radiobaserad personsökning i gemenskapen
(Text av betydelse för EES)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DETTA DIREKTIV
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 95,
med beaktande av kommissionens förslag,
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande [1],
med beaktande av Regionkommitténs yttrande [2],
i enlighet med förfarandet i artikel 251 i fördraget [3], och
av följande skäl:
(1) Enligt direktiv 90/544/EEG [4] skulle medlemsstaterna senast den 31 december 1992 ange fyra kanaler på frekvensbandet 169,4–169,8 MHz för den alleuropeiska, landbaserade, allmänt tillgängliga, radiobaserade personsökningstjänsten (nedan kallad "ERMES") samt så snabbt som möjligt utarbeta planer så att den alleuropeiska, allmänt tillgängliga, radiobaserade personsökningstjänsten kan uppta hela bandet 169,4–169,8 MHz i takt med den kommersiella efterfrågan.
(2) Användningen av spektrumbandet 169,4–169,8 MHz för ERMES i gemenskapen har minskat eller till och med upphört, vilket innebär att detta band för närvarande inte utnyttjas effektivt av ERMES och skulle kunna utnyttjas bättre för att tillgodose andra gemenskapspolitiska behov.
(3) Genom Europaparlamentets och rådets beslut nr 676/2002/EG av den 7 mars 2002 om ett regelverk för radiospektrumpolitiken i Europeiska gemenskapen (radiospektrumbeslut) [5] inrättades politiska och rättsliga ramar inom gemenskapen för att säkerställa samordning av policystrategier och i förekommande fall harmoniserade villkor när det gäller tillgång till och effektiv användning av det radiospektrum som krävs för att upprätta en välfungerande inre marknad. Det beslutet gör det möjligt för kommissionen att anta tekniska genomförandeåtgärder för att säkerställa harmoniserade villkor för tillgång till och effektiv användning av spektrumbandet.
(4) Eftersom frekvensbandet 169,4–169,8 MHz är lämpligt för tillämpningar som är till nytta för personer med funktionshinder eller handikapp, och med tanke på att främjande av sådana tillämpningar utgör ett gemenskapspolitiskt mål tillsammans med det generella målet att säkerställa en välfungerande inre marknad, har kommissionen i enlighet med artikel 4.2 i radiospektrumbeslutet gett Europeiska post- och telesammanslutningen (nedan kallad "CEPT") i uppdrag att bland annat undersöka tillämpningar som kan utgöra stöd till personer med funktionshinder.
(5) I enlighet med uppdraget har CEPT utarbetat en ny frekvensplan och en kanalfördelning som gör det möjligt att låta sex typer av utvalda tillämpningar dela på bandet i syfte att tillgodose flera gemenskapspolitiska behov.
(6) Av dessa skäl och i enlighet med målen i radiospektrumbeslutet bör direktiv 90/544/EEG upphöra att gälla.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Direktiv 90/544/EEG skall upphöra att gälla med verkan från och med den 27 december 2005.
Artikel 2
Detta direktiv träder i kraft samma dag som det offentliggörs i Europeiska unionens officiella tidning.
Artikel 3
Detta direktiv riktar sig till medlemsstaterna.
Kommissionens förordning (EG) nr 295/2005
av den 22 februari 2005
om ändring för tredje gången av rådets förordning (EG) nr 1763/2004 om införande av vissa restriktiva åtgärder till stöd för ett effektivt genomförande av Internationella krigsförbrytartribunalens för f.d. Jugoslavien (ICTY) uppgift
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1763/2004 om införande av vissa restriktiva åtgärder till stöd för ett effektivt genomförande av Internationella krigsförbrytartribunalens för f.d. Jugoslavien (ICTY) uppgift [1], särskilt artikel 10 a i denna, och
av följande skäl:
(1) Bilaga I till förordning (EG) nr 1763/2004 innehåller en förteckning över personer vars penningmedel och ekonomiska resurser har spärrats enligt den förordningen.
(2) Kommissionen är bemyndigad att ändra den bilagan med beaktande av rådets beslut om genomförande av gemensam ståndpunkt 2004/694/GUSP om ytterligare åtgärder till stöd för ett effektivt genomförande av Internationella tribunalen för f.d. Jugoslaviens (ICTY) uppgift [2]. Den gemensamma ståndpunkten genomförs genom rådets beslut 2005/148/GUSP [3] Bilaga I till förordning (EG) nr 1763/2004 bör därför ändras i enlighet med detta.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga I till förordning (EG) nr 1763/2004 skall ändras i enlighet med bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 619/2005
av den 21 april 2005
om fastställande av den största sänkningen av importtullar för majs inom ramen för den anbudsinfordran som avses i förordning (EG) nr 2277/2004
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1784/2003 av den 29 september 2003 om den gemensamma organisationen av marknaden för spannmål [1], särskilt artikel 12.1 i denna, och
av följande skäl:
(1) En anbudsinfordran om den största sänkningen av importtullar för majs till Spanien från tredjeland har inletts genom kommissionens förordning (EG) nr 2277/2004 [2].
(2) I enlighet med artikel 7 i kommissionens förordning (EG) nr 1839/95 [3] kan kommissionen, enligt förfarandet som föreskrivs i artikel 25 i förordning (EG) nr 1784/2003, besluta att fastställa den största sänkningen av importtullar. Vid fastställande av denna måste särskild hänsyn tas till kriterierna i artiklarna 6 och 7 i förordning (EG) nr 1839/95. Kontrakt tilldelas alla anbudsgivare vars anbud ligger på samma nivå som den största sänkningen av importtullar eller på en lägre nivå.
(3) Tillämpningen av ovannämnda kriterier på det nuvarande marknadsläget för ifrågavarande spannmålsslag medför att den största sänkningen av importtullar fastställs till det belopp som anges i artikel 1.
(4) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för spannmål.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
För de anbud som meddelats från och med den 15 till den 21 april 2005, inom ramen för den anbudsinfordran som avses i förordning (EG) nr 2277/2004, är den största sänkningen av importtullar för majs fastställd till 28,49 EUR/t för en maximal mängd av totalt 141000 t.
Artikel 2
Denna förordning träder i kraft den 22 april 2005.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 702/2005
av den 3 maj 2005
om fastställande av enhetsvärdena för tullvärdesbestämmelse när det gäller vissa lättfördärvliga varor
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2913/92 av den 12 oktober 1992 om upprättandet av en tullkodex för gemenskapen [1],
med beaktande av kommissionens förordning (EEG) nr 2454/93 [2] om fastställande av tillämpningsföreskrifter till förordning (EEG) nr 2913/92, särskilt artikel 173.1 i denna, och
av följande skäl:
(1) I artiklarna 173–177 i förordning (EEG) nr 2454/93 fastställer kommissionens kriterier för bestämmande av de periodiska enhetsvärdena för de produkter som avses i klassificeringen i bilaga 26 i den förordningen.
(2) Genom tillämpningen av de regler och kriterier som fastställs i ovannämnda artiklar på de uppgifter som meddelats kommissionen i enlighet med bestämmelserna i artikel 173.2 i den förordningen kan enhetsvärdena för de avsedda produkterna fastställas i enlighet med vad som föreskrivs i bilagan till den här förordningen.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De enhetsvärden som avses i artikel 173.1 i förordning (EEG) nr 2454/93 skall fastställas i enlighet med vad som anges i tabellen i bilagan.
Artikel 2
Denna förordning träder i kraft den 6 maj 2005.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 810/2005
av den 26 maj 2005
om fastställande av den största sänkningen av importtullar för majs inom ramen för den anbudsinfordran som avses i förordning (EG) nr 641/2005
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1784/2003 av den 29 september 2003 om den gemensamma organisationen av marknaden för spannmål [1], särskilt artikel 12.1 i denna, och
av följande skäl:
(1) En anbudsinfordran om den största sänkningen av importtullar för majs till Spanien från tredjeland har inletts genom kommissionens förordning (EG) nr 641/2005 [2].
(2) I enlighet med artikel 7 i kommissionens förordning (EG) nr 1839/95 [3] kan kommissionen, enligt förfarandet som föreskrivs i artikel 25 i förordning (EG) nr 1784/2003, besluta att fastställa den största sänkningen av importtullar. Vid fastställande av denna måste särskild hänsyn tas till kriterierna i artiklarna 6 och 7 i förordning (EG) nr 1839/95. Kontrakt tilldelas alla anbudsgivare vars anbud ligger på samma nivå som den största sänkningen av importtullar eller på en lägre nivå.
(3) Tillämpningen av ovannämnda kriterier på det nuvarande marknadsläget för ifrågavarande spannmålsslag medför att den största sänkningen av importtullar fastställs till det belopp som anges i artikel 1.
(4) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för spannmål.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
För de anbud som meddelats från och med den 20 till den 26 maj 2005, inom ramen för den anbudsinfordran som avses i förordning (EG) nr 641/20054, är den största sänkningen av importtullar för majs fastställd till 29,99 EUR/t för en maximal mängd av totalt 50900 t.
Artikel 2
Denna förordning träder i kraft den 27 maj 2005.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 925/2005
av den 17 juni 2005
om fastställande av det lägsta försäljningspriset för skummjölkspulver för den 20:e enskilda anbudsinfordran inom ramen för den stående anbudsinfordran som avses i förordning (EG) nr 214/2001
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1255/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter [1], särskilt artikel 10 c i denna, och
av följande skäl:
(1) I enlighet med artikel 21 i kommissionens förordning (EG) nr 214/2001 av den 12 januari 2001 om tillämpningsföreskrifter till rådets förordning (EG) nr 1255/1999 beträffande interventionsåtgärder på marknaden för skummjölkspulver [2] har interventionsorganen genom stående anbudsinfordran bjudit ut vissa kvantiteter skummjölkspulver som de innehar till försäljning.
(2) På grundval av de anbud som mottas för varje enskild anbudsinfordran skall det, i enlighet med artikel 24a i förordning (EG) nr 214/2001, fastställas ett lägsta försäljningspris eller beslutas att inget anbud skall antas.
(3) På grundval av de anbud som mottagits bör det fastställas ett lägsta försäljningspris.
(4) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för mjölk och mjölkprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
För den 20:e enskilda anbudsinfordran i enlighet med förordning (EG) nr 214/2001, för vilken tidsfristen för inlämnande av anbud löpte ut den 14 juni 2005, fastställs det lägsta försäljningspriset för skummjölkspulver härmed till 198,24 EUR/100 kg.
Artikel 2
Denna förordning träder i kraft den 18 juni 2005.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1263/2005
av den 28 juli 2005
om ändring för femte gången av rådets förordning (EG) nr 798/2004 om förlängning av de restriktiva åtgärderna mot Burma/Myanmar och om upphävande av förordning (EG) nr 1081/2000
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 798/2004 av den 26 april 2004 om förlängning av de restriktiva åtgärderna mot Burma/Myanmar och om upphävande av förordning (EG) nr 1081/2000 [1], särskilt artikel 12 i denna, och
av följande skäl:
(1) I bilaga II till förordning (EG) nr 798/2004 anges de behöriga myndigheter vilka det åligger att utföra särskilda arbetsuppgifter med anknytning till genomförandet av den förordningen.
(2) Belgien, Italien, Nederländerna och Förenade kungariket har begärt att adressuppgifterna avseende deras behöriga myndigheter skall ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilaga II till förordning (EG) nr 798/2004 skall ändras i enlighet med bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Förordningen är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1571/2005
av den 28 september 2005
om fastställande av schablonvärden vid import för bestämning av ingångspriset för vissa frukter och grönsaker
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av kommissionens förordning (EG) nr 3223/94 av den 21 december 1994 om tillämpningsföreskrifter för importordningen för frukt och grönsaker [1], särskilt artikel 4.1 i denna, och
av följande skäl:
(1) I förordning (EG) nr 3223/94 anges som tillämpning av resultaten av de multilaterala förhandlingarna i Uruguayrundan kriterierna för kommissionens fastställande av schablonvärdena vid import från tredje land för de produkter och de perioder som anges i bilagan till den förordningen.
(2) Vid tillämpningen av dessa kriterier bör schablonvärdena vid import fastställas till de nivåer som anges i bilagan till denna förordning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De schablonvärden vid import som avses i artikel 4 i förordning (EG) nr 3223/94 skall fastställas enligt tabellen i bilagan.
Artikel 2
Denna förordning träder i kraft den 29 september 2005.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1599/2005
av den 29 september 2005
om de anbud som meddelats för export av havre inom ramen för den anbudsinfordran som avses i förordning (EG) nr 1438/2005
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1784/2003 av den 29 september 2003 om den gemensamma organisationen av marknaden för spannmål [1] särskilt artikel 7 i denna,
med beaktande av kommissionens förordning (EG) nr 1501/95 av den 29 juni 1995 om vissa tillämpningsföreskrifter för rådets förordning (EEG) nr 1766/92 vad avser beviljande av exportbidrag och de åtgärder som skall vidtas vid störningar inom spannmålssektorn [2], särskilt artikel 7 i denna,
med beaktande av kommissionens förordning (EG) nr 1438/2005 av den 2 september 2005 om en särskild interventionsåtgärd för havre i Finland och Sverige för regletringsåret 2005/06 [3], och
av följande skäl:
(1) En anbudsinfordran för bidrag för export av havre som producerats i Finland och Sverige för export från Finland eller Sverige till alla tredjeländer utom Bulgarien, Norge, Rumänien och Schweiz har inletts genom förordning (EG) nr 1438/2005.
(2) Särskilt med hänsyn till de kriterier som avses i artikel 1 i förordning (EG) nr 1501/95 är det inte uppenbart att ett högsta exportbidrag skall fastställas.
(3) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för spannmål.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De anbud som meddelats från den 23 till den 29 september 2005 inom ramen för den anbudsinfordran för exportbidrag för havre som avses i förordning (EG) nr 1438/2005 skall inte fullföljas.
Artikel 2
Denna förordning träder i kraft den 30 september 2005.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1962/2005
av den 30 november 2005
om undantag från förordning (EG) nr 800/1999 när det gäller fastställandet av bidragssatsen för mjölk och mjölkprodukter vid leveranser, enligt artiklarna 36 och 44 i den förordningen, under perioden 1– 16 juni 2005
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1255/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter [1], särskilt artikel 31.14, och
av följande skäl:
(1) Från och med den 17 juni 2005 ges enligt kommissionens förordning (EG) nr 909/2005 av den 16 juni 2005 om fastställande av exportbidragen för mjölk och mjölkprodukter [2] inte längre exportbidrag för sådana leveranser som avses i artiklarna 36 och 44 i kommissionens förordning (EG) nr 800/1999 av den 15 april 1999 om gemensamma tillämpningsföreskrifter för systemet med exportbidrag för jordbruksprodukter [3].
(2) I enlighet med artikel 37 i förordning (EG) nr 800/1999 får medlemsstaterna tillåta exportörer att följa ett förfarande som innebär att den sista dagen i månaden är den avgörande dagen för bestämning av bidragssatsen för sådana leveranser som avses i artiklarna 36 och 44 i den förordningen och som lastas varje månad. Därmed är det inte möjligt att bestämma vilken bidragssats som skall tillämpas på sådana leveranser av mjölk och mjölkprodukter som genomförs i enlighet med det förfarandet under perioden 1– 16 juni 2005.
(3) Detta bör dock inte påverka rätten till bidrag för leveranser som har utförts enligt förfarandet i artikel 37 i förordning (EG) nr 800/1999 innan förordning (EG) nr 909/2005 trädde i kraft. För att kunna fastställa den bidragssatsen är det därför nödvändigt att, genom undantag från artikel 37.2 i förordning (EG) nr 800/1999, ange det datum som skall användas för detta syfte.
(4) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för mjölk och mjölkprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Genom undantag från artikel 37.2 i förordning (EG) nr 800/1999 skall den 16 juni 2005 användas för att fastställa bidragssatsen för mjölk och mjölkprodukter vid sådana leveranser som avses i artiklarna 36.1 a och c och 44.1 a och b i den förordningen och som sker under perioden 1– 16 juni 2005 i enlighet med förfarandet i artikel 37 i den förordningen.
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Den skall tillämpas från och med den 1 juni 2005.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 2134/2005
av den 22 december 2005
om fastställande av exportbidragen för bearbetade produkter av spannmål och ris
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1784/2003 av den 29 september 2003 om den gemensamma organisationen av marknaden för spannmål [1], särskilt artikel 13.3 i denna,
med beaktande av rådets förordning (EG) nr 1785/2003 av den 29 september 2003 om den gemensamma organisationen av marknaden för ris [2], särskilt artikel 14.3 i denna, och
av följande skäl:
(1) Artikel 13 i förordning (EG) nr 1784/2003 och artikel 14 i förordning (EG) nr 1785/2003 fastställer att skillnaden mellan noteringarna eller priserna på världsmarknaden för de produkter som anges i artikel 1 i de förordningarna och priserna för de produkterna inom gemenskapen kan täckas av ett exportbidrag.
(2) Artikel 14 i förordning (EG) nr 1785/2003 föreskriver att då exportbidragen fastställs måste hänsyn tas till den rådande situationen och den förväntade utvecklingen vad avser priser för och tillgängliga kvantiteter av spannmål, ris, brutet ris och spannmålsprodukter på gemenskapens marknad å ena sidan och priser för spannmål, ris, brutet ris och spannmålsprodukter på världsmarknaden å andra sidan. Samma artiklar föreskriver att det också är viktigt att säkerställa jämvikten hos och den naturliga utvecklingen av priserna och handeln på marknaderna för spannmål och ris och dessutom att ta hänsyn till den planerade exportens ekonomiska aspekt, och behovet av att undvika störningar på gemenskapens marknad.
(3) Artikel 4 i kommissionens förordning (EG) nr 1518/95 [3], om import- och exportsystemet för bearbetade produkter baserade på spannmål respektive ris definierar de särskilda kriterier som det bör tas hänsyn till då exportbidraget för dessa produkter beräknas.
(4) Det exportbidrag som beviljas för vissa bearbetade produkter bör graderas på grundval av innehållet av aska, råfibrer, skal, proteiner, fett och stärkelse i varje enskild berörd produkt, eftersom detta innehåll är en särskilt god indikator på den kvantitet basprodukter som faktiskt ingår i den bearbetade produkten.
(5) Det finns för närvarande inget behov av att, på grundval av den ekonomiska aspekten av en eventuell export och särskilt produkternas natur och ursprung, fastställa ett exportbidrag för maniok, andra tropiska rötter och knölar eller finmalet mjöl erhållna av dessa. För vissa bearbetade produkter av spannmål är det, på grund av gemenskapens obetydliga deltagande i världshandeln, för närvarande onödigt att fastställa ett exportbidrag.
(6) Förhållandena på världsmarknaden, eller de särskilda krav som vissa marknader ställer, kan göra det nödvändigt att variera exportbidraget för vissa produkter i enlighet med destination.
(7) Exportbidraget måste fastställas en gång per månad. Det kan ändras under den mellanliggande perioden.
(8) Vissa bearbetade produkter av majs får undergå en värmebehandling efter vilken ett exportbidrag som inte motsvarar produktens kvalitet kanske betalas ut. Det bör därför specificeras att för dessa produkter, som innehåller förgelatinerad stärkelse, bör inget exportbidrag betalas ut.
(9) Förvaltningskommittén för spannmål har inte yttrat sig inom den tid som ordföranden har bestämt.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Exportbidragen för de produkter som anges i artikel 1 i förordning (EG) nr 1518/95 fastställs så som det anges i bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft den 23 december 2005.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 2183/2005
av den 22 december 2005
om ändring av rådets förordning (EG) nr 1782/2003 om upprättande av gemensamma bestämmelser för system för direktstöd inom den gemensamma jordbrukspolitiken och om upprättande av vissa stödsystem för jordbrukare och om ändring av förordning (EG) nr 795/2004 om tillämpningsföreskrifter för det system med samlat gårdsstöd som föreskrivs i rådets förordning (EG) nr 1782/2003
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1782/2003 av den 29 september 2003 om upprättande av gemensamma bestämmelser för system för direktstöd inom den gemensamma jordbrukspolitiken och om upprättande av vissa stödsystem för jordbrukare och om ändring av förordningarna (EEG) nr 2019/93, (EG) nr 1452/2001, (EG) nr 1453/2001, (EG) nr 1454/2001, (EG) nr 1868/94, (EG) nr 1251/1999, (EG) nr 1254/1999, (EG) nr 1673/2000, (EEG) nr 2358/71 och (EG) nr 2529/2001 [1], särskilt artikel 145 c, h, i, s och artikel 155, och
av följande skäl:
(1) Genom kommissionens förordning (EG) nr 795/2004 [2] införs tillämpningsföreskrifter för det system med samlat gårdsstöd som gäller från och med 2005.
(2) I förordning (EG) nr 1782/2003, ändrad genom förordning (EG) nr 864/2004 [3], fastställs reglerna för kopplat stöd för bomull, olivolja, råtobak och humle samt det frikopplade stödet och integrationen av dessa sektorer i systemet med samlat gårdsstöd.
(3) För att fastställa summan och stödrättigheterna inom ramen för integrationen av stödet för tobak, olivolja, bomull och humle i systemet med samlat gårdsstöd, bör särskilda regler fastställas för dels de nationella tak som anges i artikel 41 i förordning (EG) nr 1782/2003, dels de olika aspekter på den nationella reserv som anges i artikel 42.1 och 42.8 i den förordningen.
(4) I de medlemsstater där systemet med samlat gårdsstöd tillämpades under 2005 bör man, som följd av referensbeloppen och hektar från integrationen av stödet för tobak, olivolja och bomull, räkna om värdet på och antalet stödrättigheter för de jordbrukare som tilldelades, köpte eller mottog stödrättigheter vid det senaste ansökningsdatumet för fastställande av sådana rättigheter för 2006. Arealuttagsrättigheter bör inte tas med i den här beräkningen.
(5) Man bör tillåta att det privata kontrakt som det hänvisas till i artikel 27 i förordning (EG) nr 795/2004 kan infogas eller ändras i ett arrendekontrakt till sista dagen för inlämnande av ansökan om samlat gårdsstöd under 2006.
(6) För de medlemsstater som tillämpar den regionala modell som fastställs i artikel 59.1 och 59.3 i förordning (EG) nr 1782/2003, bör samtliga stödrättigheter ökas med ett kompletterande belopp som är en följd av referensbeloppen från integrationen av stödet för tobak, olivolja, bomull och humle.
(7) Genom tillämpning av artikel 71.1 i förordning (EG) nr 1782/2003 har Malta och Slovenien beslutat tillämpa systemet med samlat gårdsstöd år 2007. I artikel 71.1 tredje stycket i den förordningen fastställs att övergångsperioden inte skall gälla för bomull, olivolja, bordsoliver samt tobak och endast fram till och med den 31 december 2005 för humle. Malta och Slovenien skulle följaktligen vara tvungna att tillämpa systemet med samlat gårdsstöd enbart för de sektorerna och integrera övriga sektorer under 2007. För att underlätta övergången till systemet med samlat gårdsstöd bör man därför tillåta övergångsregler så att man under 2006 kan tillämpa dagens system för olivodlingar i Malta och Slovenien och för humle i Slovenien, som är de enda sektorer i de länderna som berörs. Malta och Slovenien skulle därmed kunna införa systemet med samlat gårdsstöd år 2007 för samtliga sektorer.
(8) I artikel 37 i förordning (EG) nr 1782/2003, ändrad genom förordning (EG) nr 864/2004, sägs att för olivoljesektorn skall referensbeloppet för enskilda jordbrukare vara genomsnittet under fyra år av de sammanlagda belopp som beviljats en jordbrukare inom produktionsstödet för olivolja, beräknat och justerat i enlighet med bilaga VII till den förordningen, under regleringsåren 1999/2000, 2000/01, 2001/02 och 2002/03. När förordning (EG) nr 864/2004 antogs hade kommissionen ännu inte fastställt det slutliga stödbeloppet för regleringsåret 2002/03. Det är lämpligt att ändra punkt H i bilaga VII till förordning (EG) nr 1782/2003 i syfte att ta hänsyn till enhetsbeloppet för produktionsstödet för olivolja för regleringsåret 2002/03 som fastställts i kommissionens förordning (EG) nr 1299/2004 [4].
(9) I artikel 43 i förordning (EG) nr 1782/2003 fastställs att det totala antalet stödrättigheter skall vara detsamma som det genomsnittliga antalet hektar för vilket direktstöd har beviljats under referensperioden. I fråga om olivoljesektorn skall antalet hektar beräknas med den gemensamma metod som det hänvisas till i punkt H i bilaga VII till den förordningen som underlag. Det är nödvändigt att definiera den gemensamma metoden för att fastställa antalet hektar samt stödrättigheterna och användningen av stödrättigheterna i olivoljesektorn.
(10) Enligt artiklarna 44 och 51 i förordning (EG) nr 1782/2003 är områden med olivträd planterade efter den 1 maj 1998 inom godkända planteringsplaner bidragsberättigande inom systemet med samlat gårdsstöd. Sådana plantor kan likställas med investeringar inom ramen för artikel 21 i förordning (EG) nr 795/2004. Slutdatumet för godkända plantor enligt de planerna har fastställts till den 31 december 2006. Det är nödvändigt att fastställa ett senare datum för investeringar för olivträdsplanteringar.
(11) Förordningarna (EG) nr 1782/2003 och (EG) nr 795/2004 bör därför ändras i enlighet med detta.
(12) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från förvaltningskommittén för direktstöd.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 1782/2003 skall ändras på följande sätt:
1. Bilaga I ändras på följande sätt:
a) Kolumnen för "olivolja" skall ersättas med följande:
Sektor | Rättslig grund | Anmärkningar |
"Olivolja | Avdelning IV kapitel 10b i denna förordning | Arealstöd |
Artikel 48a 10 i kommissionens förordning (EG) nr 795/2004 | För Malta och Slovenien under 2006 |
b) Kolumnen för "humle" skall ersättas med följande:
Sektor | Rättslig grund | Anmärkningar |
"Humle | Avdelning IV kapitel 10d i denna förordning (***) (*****) | Arealstöd |
Artikel 48a 11 i förordning (EG) nr 795/2004 | För Slovenien under 2006" |
2. I bilaga VII skall första meningen i punkt H "(EG) nr 1794/2003" och motsvarande fotnot ersättas med följande:
"(EG) nr 1299/2004 [6]
Artikel 2
Förordning (EG) nr 795/2004 skall ändras på följande sätt:
1. I artikel 21.1 skall följande stycke läggas till:
"I fråga om investeringar för plantering av olivträd inom ramen för program som kommissionen godkänt, skall det datum som fastställs i första stycket vara den 31 december 2006."
2. I artikel 21.2 skall följande stycke läggas till:
"I fråga om de investeringar som omnämns i andra stycket i punkt 1 skall planen eller programmet vara genomfört senast den 31 december 2006."
3. Följande artikel 31b skall läggas till kapitel 4:
"Artikel 31b
Fastställande och användande av stödrättigheter i olivoljesektorn
1. Medlemsstaterna skall beräkna det antal hektar som skall beaktas när man fastställer de stödrättigheter som det hänvisas till i artikel 43 och i punkt H i bilaga VII till förordning (EG) nr 1782/2003 i GIS-olivhektar i enlighet med den gemensamma metod som anges i bilaga XXIV till förordning (EG) nr 1973/2004.
2. I fråga om jordbruksskiften som upptas av dels olivträd, dels andra grödor som omfattas av systemet med gårdsstöd, inklusive arealuttag, skall den areal som upptas av olivträd beräknas med hjälp av den metod som anges i punkt 1. Den del av det jordbruksskifte som upptas av andra grödor som omfattas av systemet med gårdsstöd skall beräknas med hjälp av det integrerade system som anges i kapitel 4 i avdelning II i förordning (EG) nr 1782/2003.
Dessa två beräkningsmetoder får inte leda till en areal som överstiger jordbruksarealen för jordbruksskiftet.
3. Trots vad som sägs i punkt 1, skall den gemensamma metod som anges i bilaga XXIV inte tillämpas i följande fall:
a) Jorbruksskiftet med olivodling är av minimal storlek, som skall fastställas av medlemsstaten och som högst får vara 0,1 hektar.
b) Jordbruksskiftet befinner sig i en administrativ enhet för vilken medlemsstaten upprättat ett alternativt system för GIS-olivsystemet.
I dessa fall skall medlemsstaten fastställa den stödberättigande arealen med objektiva kriterier som underlag och på ett sätt som garanterar likabehandling av jordbrukarna.
4. Den areal som skall beaktas vid användningen av stödrättigheter i enlighet med artikel 44 i förordning (EG) nr 1782/2003 skall beräknas i enlighet med punkterna 1–3 i den här artikeln."
4. I artikel 48a skall följande punkter läggas till:
"10. Malta och Slovenien får bevilja stöd för olivodlingar per GIS-olivhektar under 2006 för högst fem kategorier olivodlingar i enlighet med definitionen i artikel 110i.2 i förordning (EG) nr 1782/2003 och inom det maximibelopp som fastställs i punkt 3 i den artikeln, i enlighet med objektiva kriterier och på ett sätt som garanterar likabehandling av jordbrukarna.
11. För Sloveniens del skall artiklarna 12 och 13 i rådets förordning (EEG) nr 1696/71 [7] och rådets förordning (EG) nr 1098/98 [8] fortsätta att gälla för 2006 års skörd och till den 31 december 2006.
5. Följande kapitel skall föras in:
"KAPITEL 6b
INTEGRATION AV STÖDET FÖR TOBAK, OLIVOLJA, BOMULL OCH HUMLE I SYSTEMET MED SAMLAT GÅRDSSTÖD
Artikel 48c
Allmänna regler
1. Om en medlemsstat har använt sig av möjligheten i artikel 71 i förordning (EG) nr 1782/2003 och beslutat att använda systemet med samlat gårdsstöd under 2006, skall reglerna i avdelning III i förordning (EG) nr 1782/2003 och i kapitel 1–6 i den här förordningen gälla.
2. Om en medlemsstat har tillämpat systemet med samlat gårdsstöd under 2005, utan att det påverkat tillämpningen av tredje stycket i artikel 71.1 i förordning (EG) nr 1782/2003, för att fastställa summan och stödrättigheterna för 2006 inom ramen för integrationen av stödet för tobak, olivolja och bomull i systemet med samlat gårdsstöd skall artiklarna 37 och 43 i den förordningen gälla i enlighet med reglerna i artikel 48d i den här förordningen och, om medlemsstaten har använt sig av möjligheten i artikel 59 i förordning (EG) nr 1782/2003, i artikel 48e i den här förordningen.
3. Om en medlemsstat har tillämpat systemet med samlat gårdsstöd under 2005 ansvarar den för att det nationella tak som fastställs i bilaga VIII till förordning (EG) nr 1782/2003 respekteras.
4. I givna fall skall artikel 41.2 i förordning (EG) nr 1782/2003 gälla i fråga om värdet på samtliga befintliga stödrättigheter under 2006, före integrationen av stödet för tobak, olivolja, bomull och/eller mjölk, och för referensbeloppen för stödet för tobak, olivolja, bomull och/eller mjölk.
5. Om en medlemsstat har tillämpat systemet med samlat gårdsstöd under 2005, skall den procentuella minskning medlemsstaterna fastställt i enlighet med artikel 42.1 i förordning (EG) nr 1782/2003 gälla under 2006 för de referensbelopp för tobak, olivolja och bomull som skall integreras i systemet med samlat gårdsstöd.
6. Den femårsperiod som anges i artikel 42.8 i förordning (EG) nr 1782/2003 skall inte starta på nytt för de stödrättigheter som kommer från den nationella reserven och som räknats om eller ökats i enlighet med artiklarna 48d och 48e i den förordningen.
7. Första tillämpningsåret för det system med samlat gårdsstöd som det hänvisas till i artiklarna 7.1, 12–17 och 20 skall vara 2006 när det gäller att fastställa stödrättigheterna för bomull, tobak och olivolja.
Artikel 48d
Särskilda regler
1. Den jordbrukare som inte tilldelats eller som inte köpt stödrättigheter före sista ansökningsdagen för fastställandet av stödrättigheter för 2006, skall få stödrättigheter för tobak, olivolja och bomull som beräknats i enlighet med artiklarna 37 och 43 i förordning (EG) nr 1782/2003.
Det första stycket skall också gälla om jordbrukaren har arrenderat stödrättigheter för 2005 eller 2006.
2. Om jordbrukaren tilldelats, köpt eller mottagit stödrättigheter före sista ansökningsdagen för fastställandet av stödrättigheter för 2006, skall värdet på och antalet stödrättigheter räknas om enligt följande metod:
a) Antalet stödrättigheter skall vara samma som det antal jordbrukaren äger, plus det antal hektar som det i enlighet med artikel 43 i förordning (EG) nr 1782/2003 beviljades tobaks-, olivolje- och bomullsstöd för under referensperioden.
b) Värdet skall räknas fram genom att man dividerar summan av värdet på de stödrättigheter jordbrukaren äger och den referenssumma som beräknats i enlighet med artikel 37 i förordning (EG) nr 1782/2003 för de arealer som det under referensperioden beviljades tobaks-, olivolje- och bomullsstöd för, med det antal som fastställts i enlighet med punkt a i det här stycket.
Arealuttagsrättigheter skall inte ingå i beräkningen i punkt a.
3. Genom undantag från artikel 27 kan den kontraktsklausul som det hänvisas till i den artikeln infogas i eller ändras genom ett arrendekontrakt senast den sista ansökningsdagen för samlat gårdsstöd 2006.
4. Stödrättigheter som arrenderats ut före sista dagen för inlämnande av ansökan om samlat gårdsstöd under 2006 skall tas med i den beräkning som avses i punkt 2. Stödrättigheter som före den 15 maj 2004 arrenderas ut via en kontraktsklausul i enlighet med artikel 27 skall tas med i den beräkning som avses i punkt 2 i den här artikeln endast om arrendevillkoren kan ändras.
Artikel 48e
Regionalt genomförande
1. Om en medlemsstat har använt sig av möjligheten i artikel 59.1 i förordning (EG) nr 1782/2003, skall samtliga stödrättigheter ökas med ett kompletterande belopp motsvarande ökningen av det regionala taket under 2006, dividerad med det totala antalet stödrättigheter som tilldelades under 2005.
2. Om en medlemsstat har använt sig av möjligheten i artikel 59.1 och 59.3 i förordning (EG) nr 1782/2003, och utan att det påverkar tillämpningen av artikel 48 i den förordningen, skall jordbrukaren erhålla ett kompletterande belopp per stödrättighet.
Detta belopp skall bestå av summan av följande:
a) Motsvarande del av ökningen av det regionala taket dividerad med det totala antalet stödrättigheter som tilldelades under 2005.
b) Referenssumman för varje jordbrukare, som motsvarar den återstående delen av ökningen av det regionala taket dividerat med det antal stödrättigheter den jordbrukaren äger den sista ansökningsdagen för samlat gårdsstöd 2006.
I fråga om arealuttagsrättigheter skall jordbrukaren dock endast erhålla det kompletterande belopp som för varje arealuttagsrättighet beräknats i enlighet med stycke a."
6. Följande artikel skall införas som artikel 49a:
"Artikel 49a
Integration av tobak, bomull, olivolja och humle
1. Om en medlemsstat har använt sig av möjligheten i artikel 59.1 och 59.3 i förordning (EG) nr 1782/2003, skall den senast den 1 oktober 2005 meddela kommissionen vilket skäl som fanns för den partiella uppdelningen av ökningen av taket.
2. Senast den 1 oktober 2005 skall medlemsstaterna meddela kommissionen vilket beslut medlemsstaten fattat före den 1 augusti i fråga om de möjligheter som anges i artikel 68a i förordning (EG) nr 1782/2003, i punkterna H och I i bilaga VII i den förordningen och i artikel 69 i den förordningen i fråga om bomull, tobak, olivolja och humle."
Artikel 3
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska unionens officiella tidning.
Den skall tillämpas från och med den 1 januari 2006.
Artikel 2.6 i den här förordningen och stycke 7 i artikel 48c i förordning (EG) nr 795/2004, som lagts till genom artikel 2.5 i den här förordningen, skall gälla från och med den 1 oktober 2005.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Rådets yttrande
av den 24 januari 2006
om Tjeckiens uppdaterade konvergensprogram för 2005–2008
(2006/C 55/02)
EUROPEISKA UNIONENS RÅD HAR AVGIVIT FÖLJANDE YTTRANDE
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1466/97 av den 7 juli 1997 om förstärkning av övervakningen av de offentliga finanserna samt övervakningen och samordningen av den ekonomiska politiken [1], särskilt artikel 9.3,
med beaktande av kommissionens rekommendation, och
efter att ha hört Ekonomiska och finansiella kommittén.
HÄRIGENOM FRAMFÖRS FÖLJANDE.
(1) Den 24 januari 2006 behandlade rådet Tjeckiens uppdaterade konvergensprogram, som omfattar perioden 2005–2008.
(2) Efter en period av framgång i fråga om ekonomiska reformer och stabilisering under mitten av nittiotalet drabbades Tjeckien av makroekonomiska obalanser som i maj 1997 ledde till en valutakris och ekonomisk nedgång 1997-1999. Omfattande strukturreformer inom finans- och företagssektorerna möjliggjorde en återhämtning av ekonomin från och med 2000. Sedan dess har den genomsnittliga reala BNP-tillväxten legat på cirka 3 % per år, jämfört med en genomsnittlig årlig tillväxt på 1,7 % inom EU. Programmet innehåller tre olika scenarier för de makroekonomiska prognoserna och budgetprognoserna: ett "optimistiskt scenario", ett "huvudscenario" och ett "pessimistiskt scenario". "Huvudscenariot" betraktas som referensscenario vid bedömningen av budgetprognoserna, eftersom det enligt tillgängliga uppgifter tycks utgå från rimliga tillväxtantaganden som dock närmast är optimistiska för slutåret. I detta antas den reala BNP-tillväxten sjunka något, från 4,8 % 2005 till i genomsnitt 4,3 % under resten av programperioden. Konjunkturkomponenten i tillväxten är sannolikt högre än i programmets beräkningar. Inflationsberäkningarna i programmet förefaller vara tilltagna i underkant.
(3) Den 5 juli 2004 bedömde rådet att Tjeckiens underskott var alltför stort. Enligt rådets rekommendation av den 5 juli 2004 enligt artikel 104.7 skulle det alltför stora underskottet korrigeras till 2008. I sitt yttrande av den 18 januari 2005 om den föregående uppdateringen av Tjeckiens konvergensprogram för 2004–2007 rekommenderade rådet Tjeckien "att utnyttja eventuella inkomster utöver vad som planerats i budgeten till att minska underskottet samt att strikt iaktta de utgiftstak på medellång sikt för den centrala myndigheten vilka blir rättsligt bindande från och med 2006." Tjeckien uppmanades vidare att "påskynda pensionsreformen och genomföra reformen av vårdsystemet för att förbättra de offentliga finansernas långsiktiga hållbarhet."
(4) Programmet motsvarar i stora drag den modell och de krav beträffande inlämning av uppgifter för stabilitets- och konvergensprogram som anges i den nya uppförandekoden [2].
(5) Enligt kommissionens höstprognos 2005 beräknas underskottet i den offentliga sektorns finanser för 2005 till 3,2 % av BNP, vilket kan jämföras med ett planerat underskott på 4,7 % i den föregående uppdateringen och en mycket försiktig uppskattning på 4,8 % av BNP i den aktuella uppdateringen. Kommissionens uppskattning av underskottet avspeglar nyare information om utfallet för den centrala myndigheten, särskilt statsbudgeten, som kunnat registrera skatteintäkter utöver de planerade och underutnyttjande av anslag på cirka 1,5 % av BNP.
(6) Det uppdaterade programmet syftar till att senast 2008 få ned det offentliga underskottet under referensvärdet på 3 % av BNP, i linje med rådets rekommendation enligt artikel 104.7. Särskilt beräknas underskottet minskas med drygt 2 procentenheter av BNP mellan 2005 och 2008 och det primära underskottet med 2,3 procentenheter. Om man utesluter effekterna av två engångsutgifter under 2005, stannar dock minskningen av det nominella underskottet vid cirka 1 procentenhet av BNP. Minskningen av underskottet är främst ett resultat av att utgiftskvoten minskas under programperioden (med 2,3 procentenheter av BNP), medan intäkterna i stort sett är oförändrade (-0,2 procentenheter). Offentlig konsumtion och sociala överföringar är de utgiftsslag vars procentuella andel av BNP väntas sjunka mest. De offentliga investeringarna väntas öka kraftigt, från 5 % av BNP 2004 till över 6 % 2008, dvs. betydligt högre än EU-genomsnittet (2,5 % av BNP 2005). Jämfört med det föregående programmet är uppdateringen från november 2005 i stort sett en bekräftelse på den planerade anpassningen, även om det bakomliggande makroekonomiska scenariot är avsevärt starkare.
(7) Enligt beräkningar med den allmänt vedertagna metoden väntas det strukturella saldot (dvs. det konjunkturrensade saldot netto efter engångsåtgärder och andra tillfälliga åtgärder) förbättras med 12 % av BNP under programperioden. Programmets mål för de offentliga finanserna på medellång sikt är ett strukturellt underskott på "cirka" 1 % av BNP, men detta mål skall inte nås under programperioden. Eftersom programmets mål på medellång sikt är mer ambitiöst än det lägsta riktmärket (ett beräknat underskott på cirka 112 % av BNP), bör dess slutliga uppfyllande motsvara målet med en säkerhetsmarginal mot ett alltför stort underskott. Programmets mål på medellång sikt ligger enligt den aktuella bedömningen på en rimlig nivå, eftersom det i tillräcklig grad tar hänsyn till skuldkvoten och den genomsnittliga potentiella produktionstillväxten på lång sikt.
(8) De risker som omgärdar programmets prognoser för de offentliga finanserna verkar i stort sett uppväga varandra. Å ena sidan tyder tidigare erfarenheter av försiktig budgetplanering på att resultaten kan överträffa målen (vilket var fallet 2004 och vilket kommissionen också förutspår för 2005). De grundläggande tillväxtantagandena om de offentliga finanserna har vanligtvis varit realistiska och antagandena om skatteelasticiteten försiktiga. Dessutom har budgeterade utgifter inte alltid verkställts, främst för att outnyttjade medel från tidigare budgetår kan föras över. Å andra sidan hänvisar programmet till olika (föreslagna) åtgärder på det sociala utgiftsområdet som skulle öka motsvarande utgifter i stället för att enligt programmets beräkningar minska dem. Dessutom har outnyttjade medel på drygt 1 % av BNP ackumulerats under 2004 och kommissionen väntar att de skall öka ytterligare 2005. Dessa outnyttjade medel från tidigare budgetår är betydande och skulle de och de budgeterade utgifterna tas i anspråk – vilket inte kan uteslutas särskilt under valåret 2006 – kan budgetutfallet bli sämre än planerat, särskilt 2006. Dessutom framstår tillväxtantagandet för programmets slutår som optimistiskt.
(9) Med hänsyn till dessa risker förefaller programmets finanspolitiska inriktning vara förenlig med den korrigering av det alltför stora underskottet senast 2008 som rådet rekommenderat. Emellertid skulle den planerade strukturella anpassningsvägen kunna stärkas, särskilt med hänsyn till att ett mycket bättre resultat eventuellt kan uppnås 2005 och till uppjusteringen av tillväxtantagandena.
(10) Skuldkvoten beräknas 2005 uppgå till 37,4 % av BNP, vilket är betydligt lägre än fördragets referensvärde 60 %. I programmet väntas skuldkvoten öka med 12 procentenhet under programperioden.
(11) När det gäller de offentliga finansernas hållbarhet förefaller Tjeckien löpa stora risker, till följd av de beräknade budgetkostnaderna för en åldrande befolkning. Jämfört med EU i stort är den nuvarande skuldkvoten relativt låg, men det stora underskottet bidrar till att skuldkvoten ökar i långtidsprognoserna fram till 2050, vilket innebär ökade risker för en hållbar skuld. Att pensionsutgifterna beräknas öka kraftigt under prognosperioden väntas samtidigt anstränga de offentliga finanserna. För att minska riskerna för de offentliga finansernas hållbarhet [3] är det ytterst viktigt att strikt genomföra den planerade konsolideringen av de offentliga finanserna på medellång sikt och fortsätta stärka dessa, samtidigt som ytterligare strukturreformer för att styra ökningen av åldersrelaterade utgifter särskilt för pensioner, hälso- och sjukvård, genomförs.
(12) De planerade åtgärderna för de offentliga finanserna överensstämmer i huvudsak med de allmänna riktlinjerna för den ekonomiska politiken, som ingår i de integrerade riktlinjerna för perioden 2005–2008. I programmet planeras särskilt en korrigering av det alltför stora underskottet enligt rådets rekommendationer. Det innehåller också åtgärder för tillväxt- och sysselsättningsfrämjande resursfördelning, särskilt genom att minska den offentliga sektorns betydelse för ekonomin och genom en övergång från direkt till indirekt beskattning. Även om regeringen är medveten om problemet med långsiktig hållbarhet, innehåller programmet inga konkreta insatser för att åtgärda det.
(13) Tjeckien lade den 14 oktober 2005 fram ett nationellt reformprogram i samband med den förnyade Lissabonstrategin för tillväxt och sysselsättning. I detta anges långsiktig hållbarhet som det största problemet för de offentliga finanserna. Budgetkonsekvenserna av det begränsade antal konkreta reformåtgärder som anges i det nationella reformprogrammet återspeglas i konvergensprogrammets budgetprognoser. Konvergensprogrammets åtgärder för de offentliga finanserna ligger i linje med de insatser som anges i det nationella reformprogrammet. Mer specifikt anges i konvergensprogrammet åtgärder för sysselsättning och tillväxt genom förändrad inkomst- och utgiftsstruktur (särskilt genom en övergång från direkt till indirekt beskattning och minskning av offentlig konsumtion och offentliga överföringar) samt genom en prioritering av offentliga investeringar. Emellertid anges, såsom nämns ovan, inga konkreta reforminsatser för att åtgärda problemet med långsiktig hållbarhet. I programmet planeras vidare en stärkning på medellång sikt av utgiftstakens roll genom att bindande principer tillämpas på statsbudgetens och de statliga medlens olika rubriker och genom att lokala myndigheter engageras i budgetplaneringen.
Utifrån denna bedömning noterar rådet att programmet följer den väg för underskottsanpassning som fastställts i rådets rekommendationer enligt artikel 104.7. Mot bakgrund av dessa rekommendationer anser rådet att Tjeckien bör
i) med hänsyn till möjligheten till ett bättre budgetresultat 2005, samt utsikterna till fortsatt stark tillväxt, öka ansträngningarna att anpassa budgeten strukturellt med tanke på den lilla marginal under referensvärdet som planeras för 2008 (tidsfristen för korrigering av det alltför stora underskottet) och för att se till att målen på medellång sikt uppnås snabbare,
ii) höja budgetplaneringens kvalitet, särskilt genom att analysera orsakerna till de betydande outnyttjade medlen från tidigare budgetår och genom på medellång sikt stärka utgiftstakens roll,
iii) förbättra de offentliga finansernas hållbarhet på lång sikt, särskilt genom att påskynda pensionsreformen och genomföra reformen av vårdsystemet.
Jämförelse av centrala makroekonomiska och finansiella prognoser
Anmärkningar:
Källor:
Konvergensprogram (KP); kommissionens höstprognos 2005 (KOM); samt kommissionens beräkningar
| 2004 | 2005 | 2006 | 2007 | 2008 |
Real BNP (förändring i %) | KP nov. 2005 | 4,4 | 4,8 | 4,4 | 4,2 | 4,3 |
KOM nov. 2005 | 4,4 | 4,8 | 4,4 | 4,3 | — |
KP dec. 2004 | 3,8 | 3,6 | 3,7 | 3,8 | — |
Inflation (HIKP, i %) | KP nov. 2005 | 2,6 | 1,5 | 2,2 | 2,0 | 2,1 |
KOM nov. 2005 | 2,6 | 1,7 | 2,9 | 2,6 | — |
KP dec. 2004 | 2,7 | 3,2 | 2,6 | 2,2 | — |
BNP-gap (i % av potentiell BNP) | KP nov. 2005 [4] | – 1,9 | – 0,8 | – 0,1 | 0,3 | 0,8 |
KOM nov. 2005 [8] | – 1,4 | – 0,2 | 0,6 | 1,2 | — |
KP dec. 2004 [4] | – 1,3 | – 0,9 | – 0,4 | 0,3 | — |
Saldot för de offentliga finanserna (i % av BNP) | KP nov. 2005 | – 3,0 | – 4,8 | – 3,8 | – 3,3 | – 2,7 |
KOM nov. 2005 | – 3,0 | – 3,2 | – 3,7 | – 3,3 | — |
KP dec. 2004 | – 5,2 | – 4,7 | – 3,8 | – 3,3 | — |
Primärt saldo (i % av BNP) | KP nov. 2005 | – 1,8 | – 3,5 | – 2,5 | – 2,0 | – 1,2 |
KOM nov. 2005 | – 1,8 | – 1,9 | – 2,3 | – 1,9 | — |
KP dec. 2004 | – 4,0 | – 3,4 | – 2,4 | – 1,7 | — |
Konjunkturrensat saldo (i % av BNP) | KP nov. 2005 [4] | – 2,4 | – 4,5 | – 3,8 | – 3,4 | – 3,0 |
KOM nov. 2005 | – 2,5 | – 3,1 | – 3,9 | – 3,8 | — |
KP dec. 2004 [4] | — | — | — | — | — |
Strukturellt saldo [5] (i % av BNP) | KP nov. 2005 [6] | – 1,9 | – 3,4 | – 3,8 | – 3,4 | – 3,0 |
KOM nov. 2005 [7] | – 2,0 | – 2,0 | – 3,9 | – 3,8 | — |
KP dec. 2004 | — | — | — | — | — |
Offentliga sektorns bruttoskuld (i % av BNP) | KP nov. 2005 | 36,8 | 37,4 | 37,1 | 37,9 | 37,8 |
KOM nov. 2005 | 36,8 | 36,2 | 36,6 | 36,9 | — |
KP dec. 2004 | 38,6 | 38,3 | 39,2 | 40,0 | — |
[1] EGT L 209, 2.8.1997, s. 1. Förordningen ändrad genom förordning (EG) nr 1055/2005 (EUT L 174, 7.7.2005, s. 1). De dokument som det hänvisas till i texten återfinns på följande webbplats:http://europa.eu.int/comm/economy_finance/about/activities/sgp/main_en.htm
[2] I programmet redovisas alla obligatoriska och flertalet av de frivilliga uppgifter som föreskrivs i den nya uppförandekoden.
[3] Närmare uppgifter om hållbarhet på lång sikt finns i kommissionens tekniska bedömning av programmet, som kommer att offentliggöras på följande webbplats:http://europa.eu.int/comm/economy_finance/about/activities/sgp/main_en.htm
[4] Kommissionens beräkningar på grundval av uppgifterna i programmet.
[5] Konjunkturrensat saldo (se föregående rad), utan beaktande av engångsåtgärder och andra tillfälliga åtgärder.
[6] Engångsåtgärder och andra tillfälliga åtgärder enligt rapporten om de offentliga finanserna (0,5 % 2004) och enligt programmet (1,1 % 2005). Bägge ökar underskottet.
[7] Engångsåtgärder och andra tillfälliga åtgärder enligt kommissionens höstprognos 2005 (0,5 % av BNP 2004, 1,1 % av BNP 2005. Bägge ökar underskottet).
[8] Baseras på en beräknad potentiell tillväxt på 3,5 %, 3,5 %, 3,6 % och 3,7 % per år under perioden 2004-2007.
--------------------------------------------------
Sammanställning över inkomster och utgifter för Europeiska arbetsmiljöbyrån för budgetåret 2006 – ändringsbudget 1
(2006/341/EG)
REDOGÖRELSE FÖR INKOMSTER
Avdelning Kapitel | Rubrik | Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
1
BIDRAG FRÅN EUROPEISKA GEMENSKAPERNA
1 0 | BIDRAG FRÅN EUROPEISKA GEMENSKAPERNA | 13342216 | 489142 | 13831358 |
| Avdelning 1 – Totalt | 13342216 | 489142 | 13831358 |
| TOTALSUMMA | 13522519 | 489142 | 14011661 |
AVDELNING 1
BIDRAG FRÅN EUROPEISKA GEMENSKAPERNA
KAPITEL 1 0 — BIDRAG FRÅN EUROPEISKA GEMENSKAPERNA
Artikel Punkt | Rubrik | Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
KAPITEL 1 0
1 0 0 | Bidrag från Europeiska gemenskapen | 13200000 | — | 13200000 |
1 0 1 | Phareprogram III (öronmärkt) | 142216 | 187222 | 329438 |
1 0 2 | Phareprogram IV (öronmärkt) | 142216 | 159704 | 301920 |
| KAPITEL 1 0 TOTALT | 13342216 | 489142 | 13831358 |
| Avdelning 1 – Totalt | 13342216 | 489142 | 13831358 |
| TOTALSUMMA | 13522519 | 489142 | 14011661 |
Anmärkningar
Bidrag från Europeiska gemenskapen, totalt.
KAPITEL 1 0 —BIDRAG FRÅN EUROPEISKA GEMENSKAPERNA
1 0 0Bidrag från Europeiska gemenskapen
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
13200000 | — | 13200000 |
Anmärkningar
Rådets förordning (EG) nr 2062/94 av den 18 juli 1994 om upprättande av en europeisk arbetsmiljöbyrå (EGT L 216, 20.8.1994, s. 1), ändrad genom förordning (EG) nr 1643/95 (EGT L 156, 7.7.1995, s. 1). Enligt artikel 12.3 i denna förordning förs ett bidrag till arbetsmiljöbyrån in i avsnittet "Kommissionen" i den allmänna budgeten.
1 0 1Phareprogram III (öronmärkt)
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
142216 | 187222 | 329438 |
Anmärkningar
Detta kapitel motsvarar öronmärkta inkomster för Phare och innefattar finansiering av ett Phare III-program som undertecknats tillsammans med gemenskapen och kommer att omfatta perioden 2005–2006 till ett totalt belopp av 500000 euro. Verksamheten inom ramen för Phare III är knuten till det godkända arbetsprogrammet med öronmärkta inkomster och utgifter. Siffran för 2005 motsvarar det faktiska genomförandet för detta år. Saldot avseende det totala beloppet på 500000 euro framgår av budgeten för 2006.
1 0 2Phareprogram IV (öronmärkt)
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
142216 | 159704 | 301920 |
Anmärkningar
Detta kapitel motsvarar öronmärkta inkomster för Phare och innefattar finansiering av ett Phare IV-program som godkänts av gemenskapen och kommer att omfatta perioden 2006–2007 till ett totalt belopp av 450000 euro. Verksamheten inom ramen för Phare III är knuten till det godkända arbetsprogrammet med öronmärkta inkomster och utgifter.
REDOGÖRELSE FÖR UTGIFTER
Avdelning Kapitel | Rubrik | Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
3
DRIFTSUTGIFTER
3 0 | ALLMÄNNA DRIFTSUTGIFTER | 5750000 | — | 5750000 |
3 1 | SMÅ OCH MEDELSTORA FÖRETAG | | | |
3 2 | PHAREPROGRAM | 142216 | 187222 | 329438 |
3 3 | HANDLINGSPLAN FÖR UTVIDGNINGEN | 1550000 | — | 1550000 |
3 4 | PHAREPROGRAM IV (ÖRONMÄRKT) | | 301920 | 301920 |
| Avdelning 3 – Totalt | 7442216 | 489142 | 7931358 |
| TOTALSUMMA | 13522519 | 489142 | 14011661 |
AVDELNING 3
DRIFTSUTGIFTER
KAPITEL 3 0 — ALLMÄNNA DRIFTSUTGIFTER
KAPITEL 3 1 — SMÅ OCH MEDELSTORA FÖRETAG
KAPITEL 3 2 — PHAREPROGRAM
KAPITEL 3 3 — HANDLINGSPLAN FÖR UTVIDGNINGEN
KAPITEL 3 4 — PHAREPROGRAM IV (ÖRONMÄRKT)
Artikel Punkt | Rubrik | Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
KAPITEL 3 0
3 0 0
Kontaktpunkternas verksamhet inklusive expertgruppsverksamhet, kostnader för möten och tolkning
3 0 0 0 | Begäran om information och övriga kostnader | p.m. | p.m. | p.m. |
3 0 0 1 | Bidrag till kontaktpunkterna | 940000 | — | 940000 |
3 0 0 2 | Kontaktpunkternas möten | 88500 | — | 88500 |
3 0 0 3 | Extern utvärdering av arbetsmiljöbyrån och kontaktpunkternas nätverk | 150000 | — | 150000 |
| Artikel 3 0 0 – Totalt | 1178500 | — | 1178500 |
3 0 1
Upprättande och administration av informationsnätverket på Internet
3 0 1 0 | Upprättande och administration av informationsnätverket på Internet | 180000 | — | 180000 |
| Artikel 3 0 1 – Totalt | 180000 | — | 180000 |
3 0 2
Informationsprojekt och Informationssystem/ämnescentrum och externa uppdragstagare
3 0 2 0 | Riskcentrum | 628500 | — | 628500 |
3 0 2 1 | God arbetsmiljöpraxis (ämnescentrum) | | | |
3 0 2 2 | Forskning om arbetsmiljö (ämnescentrum) | | | |
3 0 2 3 | God arbetsmiljöpraxis (ämnescentrum) – nya medlemsstater | | | |
3 0 2 4 | Arbetsmiljö | 1100000 | — | 1100000 |
| Artikel 3 0 2 – Totalt | 1728500 | | 1728500 |
3 0 3
Konferenser, seminarier, workshopar och offentliga evenemang, reklamverksamhet, osv.
3 0 3 0 | Konferenser, seminarier, workshopar och offentliga evenemang, reklamverksamhet, osv. | 480000 | — | 480000 |
3 0 3 2 | Övriga möten | 66690 | — | 66690 |
| Artikel 3 0 3 – Totalt | 546690 | — | 546690 |
3 0 4
Redigering, publicering och distribution av information, samt övrig verksamhet
3 0 4 0 | Publicering och distribution av undersökningsresultat samt övrig informationsverksamhet och gemensamma produkter | 380000 | — | 380000 |
3 0 4 4 | Redigering | 51250 | — | 51250 |
| Artikel 3 0 4 – Totalt | 431250 | — | 431250 |
3 0 6
Översättning och tolkning
3 0 6 0 | Översättning av undersökningar, rapporter och arbetsdokument | 705811 | — | 705811 |
3 0 6 1 | Tolkning | p.m. | p.m. | p.m. |
| Artikel 3 0 6 – Totalt | 705811 | — | 705811 |
3 0 7
Förberedelser, anordnande och administration av Europeiska arbetsmiljöveckan
3 0 7 2 | Förberedelser, anordnande och administration av Europeiska arbetsmiljöveckan | 480000 | — | 480000 |
| Artikel 3 0 7 – Totalt | 480000 | — | 480000 |
3 0 8
Styrelsens och presidiets möten
3 0 8 0 | Styrelsens och presidiets möten | 271202 | — | 271202 |
| Artikel 3 0 8 – Totalt | 271202 | — | 271202 |
3 0 9
Utgifter för tjänsteresor, mottagningar och representation
3 0 9 1 | Utgifter för tjänsteresor, resekostnader och andra tillhörande utgifter | 219351 | — | 219351 |
3 0 9 2 | Mottagnings- och representationskostnader | 8696 | — | 8696 |
| Artikel 3 0 9 – Totalt | 228047 | — | 228047 |
| KAPITEL 3 0 TOTALT | 5750000 | — | 5750000 |
KAPITEL 3 1
3 1 1
Projektstöd
3 1 1 0 | Stöd till projekt | | | |
| Artikel 3 1 1 – Totalt | | | |
3 1 2
Arbetsmiljöbyråns informationsverksamhet
3 1 2 0 | Arbetsmiljöbyråns informationsverksamhet | | | |
| Artikel 3 1 2 – Totalt | | | |
3 1 4
Utvärdering SMF
3 1 4 0 | Utvärdering SMF | | | |
| Artikel 3 1 4 – Totalt | | | |
| KAPITEL 3 1 TOTALT | | | |
KAPITEL 3 2
3 2 0
PHAREPROGRAM III (öronmärkt)
3 2 0 0 | Löner för utlandsstationerad/internationell personal | 53240 | 27627 | 80867 |
3 2 1 0 | Resekostnader (internationella) | 31757 | 44400 | 76157 |
3 2 1 1 | Utgifter för tjänsteresor för projektpersonal utomlands | 2170 | 1629 | 3799 |
3 2 1 2 | Utgifter för tjänsteresor för deltagande i seminarier/konferenser | 2700 | 6797 | 9497 |
3 2 2 0 | Översättning/tolkar | 17600 | — | 17600 |
3 2 3 0 | Workshop i samband med Europaveckan | — | 14376 | 14376 |
3 2 4 0 | Webbansvariga | 13336 | 6564 | 19900 |
3 2 4 1 | Teknisk utrustning | | 10000 | 10000 |
3 2 5 0 | Ämnescentrum för god praxis | | — | — |
3 2 6 0 | Förvaltningskostnader | 1413 | 2057 | 3470 |
3 2 7 0 | Tryckning av informationsmaterial | 20000 | 7772 | 27772 |
3 2 8 0 | Seminarier och konferenser inom ramen för Healthy workplace initiative (initiativet för hälsosamma arbetsplatser) | | 48000 | 48000 |
3 2 8 1 | Mediatjänster | | 10000 | 10000 |
3 2 8 2 | Hantering och distribution av listor | | 8000 | 8000 |
| Artikel 3 2 0 – Totalt | 142216 | 187222 | 329438 |
| KAPITEL 3 2 TOTALT | 142216 | 187222 | 329438 |
KAPITEL 3 3
3 3 0 | Handlingsplan för utvidgningen | 1550000 | — | 1550000 |
| KAPITEL 3 3 TOTALT | 1550000 | — | 1550000 |
KAPITEL 3 4
3 4 0
PHAREPROGRAM IV (öronmärkt)
3 4 0 0 | Löner för utlandsstationerad/internationell personal | | 67500 | 67500 |
3 4 1 0 | Resekostnader (internationella) | | 45000 | 45000 |
3 4 1 1 | Utgifter för tjänsteresor för projektpersonal utomlands | | 3110 | 3110 |
3 4 1 2 | Utgifter för tjänsteresor för seminarie-/konferensdeltagare | | 6000 | 6000 |
3 4 2 0 | Översättning/tolkar | | 27840 | 27840 |
3 4 3 0 | Workshop i samband med Europaveckan | | 44000 | 44000 |
3 4 4 0 | Webbansvariga, stöd till kontaktpunkterna | | 75600 | 75600 |
3 4 4 1 | Datautrustning | | 4800 | 4800 |
3 4 5 0 | Inventarier | | 4000 | 4000 |
3 4 6 0 | Tryckning av informationsmaterial | | 24070 | 24070 |
| Artikel 3 4 0 – Totalt | | 301920 | 301920 |
| KAPITEL 3 4 TOTALT | | 301920 | 301920 |
| Avdelning 3 – Totalt | 7442216 | 489142 | 7931358 |
| TOTALSUMMA | 13522519 | 489142 | 14011661 |
Anmärkningar
Totalt anslag för driftsutgifter.
KAPITEL 3 0 —ALLMÄNNA DRIFTSUTGIFTER
3 0 0Kontaktpunkternas verksamhet inklusive expertgruppsverksamhet, kostnader för möten och tolkning
3 0 0 0Begäran om information och övriga kostnader
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
p.m. | p.m. | p.m. |
Anmärkningar
Detta anslag är avsett att täcka kostnader för besvarande av begäran om information (som skall besvaras av kontaktpunkterna) och upprättandet av små rapporter som bygger på resultaten, samt täcka övriga kostnader som rör förvaltningen av kontaktpunktssystemet).
3 0 0 1Bidrag till kontaktpunkterna
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
940000 | — | 940000 |
Anmärkningar
Detta anslag är avsett att täcka utgifter till förmån för verksamheterna inom ramen för arbetsmiljöbyråns nätverk av kontaktpunkter för att säkerställa att byråns information och kampanjbudskap sprids på medlemsstatsnivå. Detta genomförs genom bidragsavtal mellan arbetsmiljöbyrån och kontaktpunkterna om samfinansiering av lämpliga verksamheter, som till exempel för att stimulera verksamheter inom ramen för Europaveckan och andra åtgärder för spridning.
3 0 0 2Kontaktpunkternas möten
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
88500 | — | 88500 |
Anmärkningar
Detta anslag är avsett att täcka driftskostnaderna för kontaktpunktsnätverket, däribland kostnader för resor och traktamenten, kostnader för tolkning och eventuell hyra av rum.
3 0 0 3Extern utvärdering av arbetsmiljöbyrån och kontaktpunkternas nätverk
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
150000 | — | 150000 |
Anmärkningar
Detta anslag är avsett att täcka kontraktskostnaderna för en utvärdering av arbetsmiljöbyråns arbete och dess nätverk av kontaktpunkter.
3 0 1Upprättande och administration av informationsnätverket på Internet
3 0 1 0Upprättande och administration av informationsnätverket på Internet
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
180000 | — | 180000 |
Anmärkningar
Detta anslag är avsett att täcka administration och utveckling av arbetsmiljöbyråns elektroniska kommunikationer. Detta omfattar "tredje generationens" webbplatser inklusive flerspråkiga webbplatser med upp till 20 språk, byråns extranät och intranät.
3 0 2Informationsprojekt och Informationssystem/ämnescentrum och externa uppdragstagare
Anmärkningar
Detta anslag är avsett att täcka det arbete som utförs av de ämnescentrum som utsetts av styrelsen som en del av byråns arbetsprogram, eller särskilda projekt och rapporter som bidrar till genomförandet av de viktigaste verksamhetsområdena i byråns arbetsprogram.
3 0 2 0Riskcentrum
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
628500 | — | 628500 |
Anmärkningar
Detta anslag täcker inrättandet och utvecklingen av riskcentrumet. Det innefattar särskilt insamling, analys och konsolidering av befintlig statistik; förutseende av nya och framväxande risker; skapande av en webbplats för riskcentrumet; utformning av och testfas för en företagspanel/företagsundersökning för hela EU; fastställande av prioriteringar för arbetsmiljöforskning och främjande av projekt för arbetsmiljöforskning på EU-nivå.
3 0 2 1God arbetsmiljöpraxis (ämnescentrum)
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| | |
Anmärkningar
Detta anslag har för 2005 förts upp under posterna 3 0 2 0 och 3 0 2 4.
3 0 2 2Forskning om arbetsmiljö (ämnescentrum)
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| | |
Anmärkningar
Detta anslag har för 2005 förts upp under punkterna 3 0 2 0 och 3 0 2 4.
3 0 2 3God arbetsmiljöpraxis (ämnescentrum) – nya medlemsstater
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| | |
Anmärkningar
Detta anslag har för 2005 förts upp under punkt 3 0 2 4.
3 0 2 4Arbetsmiljö
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
1100000 | — | 1100000 |
Anmärkningar
Detta anslag avser utveckling av en rad ämnen som genom att kombinera granskning och analys av befintlig forskning med insamling och tillhandahållande av exempel på policy och god praxis. Det avser särskilt bidrag till Europaveckan om unga arbetstagare, en sektorgranskning (hotell och restauranger), förberedelse av Europaveckan 2007 om muskuloskeletala sjukdomar och fortsatt förbättring av webbresurserna.
3 0 3Konferenser, seminarier, workshopar och offentliga evenemang, reklamverksamhet, osv.
3 0 3 0Konferenser, seminarier, workshopar och offentliga evenemang, reklamverksamhet, osv.
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
480000 | — | 480000 |
Anmärkningar
Detta anslag är avsett att täcka kostnaderna för marknadsföring och kommunikationsaktiviteter för arbetsmiljöbyråns informationsprodukter och informationstjänster, vilket skall bidra till genomförandet av arbetsprogrammet. Dessa aktiviteter kan omfatta anordnandet av marknadsförings-, marknadsundersöknings-, press- och reklamverksamhet beträffande arbetsmiljöbyråns arbete (undersökningar, broschyrer, videor, affischer, offentliga evenemang, möten, seminarier, utställningar, kampanjer osv.) samt bidrag till liknande aktiviteter som anordnas av andra, vilket medverkar till genomförandet och utvecklingen av arbetsprogrammet.
3 0 3 2Övriga möten
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
66690 | — | 66690 |
Anmärkningar
Detta anslag är avsett att täcka driftskostnader för andra möten som ad hoc-gruppmöten eller andra expertmöten (inklusive reskostnader och traktamenten, eventuella tolkningskostnader och hyra av rum).
3 0 4Redigering, publicering och distribution av information, samt övrig verksamhet
3 0 4 0Publicering och distribution av undersökningsresultat samt övrig informationsverksamhet och gemensamma produkter
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
380000 | — | 380000 |
Anmärkningar
Detta anslag är avsett att täcka publicerings- och distributionskostnader (inklusive databaser och utskick) för undersökningsresultat, övrig informationsverksamhet och gemensamma publikationer (årsrapporter, tidskrifter, byråns budget osv.), som bidrar till genomförandet av arbetsmiljöbyråns arbetsprogram.
3 0 4 4Redigering
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
51250 | — | 51250 |
Anmärkningar
Detta anslag är avsett att täcka redigeringskostnader.
3 0 6Översättning och tolkning
3 0 6 0Översättning av undersökningar, rapporter och arbetsdokument
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
705811 | — | 705811 |
Anmärkningar
Detta anslag är avsett att täcka utgifter för översättningen av undersökningar, rapporter och arbetsdokument för styrelsen och presidiet samt för kongresser, seminarier osv. till de olika gemenskapsspråken. Översättningsarbetet kommer i huvudsak att utföras av Översättningscentrum för Europeiska unionens organ i Luxemburg.
3 0 6 1Tolkning
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
p.m. | p.m. | p.m. |
Anmärkningar
Detta anslag är avsett att täcka utgifter för den tolkning som faktureras byrån av institutionerna, särskilt kommissionen. Det är också avsett att täcka betalning till frilanstolkar som anlitats för att arbetsmiljöbyrån skall kunna stå för tolkning vid enstaka konferenser, om kommissionen inte kan ställa tolkningsresurser till förfogande. Ersättningen innefattar, förutom arbetsersättning, avgifter till livförsäkring, sjuk- och olycksfallsförsäkring och ersättning vid dödsfall, ersättning för reseutlägg samt schablonersättning för resor för de frilanstolkar vars yrkesmässiga hemort inte sammanfaller med tjänsteorten.
3 0 7Förberedelser, anordnande och administration av Europeiska arbetsmiljöveckan
3 0 7 2Förberedelser, anordnande och administration av Europeiska arbetsmiljöveckan
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
480000 | — | 480000 |
Anmärkningar
Detta anslag skall täcka kostnaderna för produktion och distribution av kampanjmaterial, anordnande och administration av konferenser (avslutningsevenemang och program för utdelande av pris för god praxis), seminarier, utställningar, offentliga evenemang, pr-verksamhet och utvärderingar inom ramen för Europeiska arbetsmiljöveckan.
3 0 8Styrelsens och presidiets möten
3 0 8 0Styrelsens och presidiets möten
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
271202 | — | 271202 |
Anmärkningar
Detta anslag skall täcka styrelsens och presidiets driftsutgifter inklusive utgifter för resor och traktamenten, kostnader för tolkning, och eventuell hyra av rum.
3 0 9Utgifter för tjänsteresor, mottagningar och representation
3 0 9 1Utgifter för tjänsteresor, resekostnader och andra tillhörande utgifter
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
219351 | — | 219351 |
Anmärkningar
Detta anslag skall täcka utgifter för transport, betalning av dagtraktamenten och tillkommande eller särskilda utgifter som etablerad personal haft i tjänstens intresse, i enlighet med tjänsteföreskrifterna för tjänstemännen i Europeiska gemenskaperna.
3 0 9 2Mottagnings- och representationskostnader
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
8696 | — | 8696 |
Anmärkningar
Detta anslag skall täcka underhållnings- och representationsutgifter.
KAPITEL 3 1 —SMÅ OCH MEDELSTORA FÖRETAG
3 1 1Projektstöd
3 1 1 0Stöd till projekt
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| | |
Anmärkningar
Detta anslag är avsett att täcka finansieringsåtgärder för små och medelstora företag för utveckling och utbyte av effektiva goda exempel som minskar arbetsmiljöriskerna.
3 1 2Arbetsmiljöbyråns informationsverksamhet
3 1 2 0Arbetsmiljöbyråns informationsverksamhet
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| | |
Anmärkningar
Detta anslag är avsett att täcka arbetsmiljöbyråns informationsverksamhet, särskilt för att främja de belönade projektresultaten.
3 1 4Utvärdering SMF
3 1 4 0Utvärdering SMF
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| | |
Anmärkningar
Detta anslag skall täcka en extern uppdragstagares utvärdering och rapportering av SMF-finansieringsprogrammen.
KAPITEL 3 2 —PHAREPROGRAM
3 2 0PHAREPROGRAM III (öronmärkt)
Anmärkningar
Detta kapitel innefattar förberedelser för Rumäniens och Bulgariens kommande deltagande i arbetsmiljöbyrån. Ett Phare III-program till ett totalt belopp av 500000 euro har undertecknats tillsammans med gemenskapen och kommer att omfatta perioden 2005–2006. Verksamheten inom ramen för Phare III är knuten till det godkända arbetsprogrammet med öronmärkta inkomster och utgifter. Siffrorna för 2005 motsvarar det faktiska genomförandet för detta år. Saldot avseende det totala beloppet på 500000 euro framgår av budgeten för 2006.
3 2 0 0Löner för utlandsstationerad/internationell personal
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
53240 | 27627 | 80867 |
3 2 1 0Resekostnader (internationella)
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
31757 | 44400 | 76157 |
3 2 1 1Utgifter för tjänsteresor för projektpersonal utomlands
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
2170 | 1629 | 3799 |
3 2 1 2Utgifter för tjänsteresor för deltagande i seminarier/konferenser
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
2700 | 6797 | 9497 |
3 2 2 0Översättning/tolkar
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
17600 | — | 17600 |
3 2 3 0Workshop i samband med Europaveckan
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
— | 14376 | 14376 |
3 2 4 0Webbansvariga
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
13336 | 6564 | 19900 |
3 2 4 1Teknisk utrustning
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 10000 | 10000 |
3 2 5 0Ämnescentrum för god praxis
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| — | — |
3 2 6 0Förvaltningskostnader
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
1413 | 2057 | 3470 |
3 2 7 0Tryckning av informationsmaterial
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
20000 | 7772 | 27772 |
3 2 8 0Seminarier och konferenser inom ramen för Healthy workplace initiative (initiativet för hälsosamma arbetsplatser)
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 48000 | 48000 |
3 2 8 1Mediatjänster
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 10000 | 10000 |
3 2 8 2Hantering och distribution av listor
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 8000 | 8000 |
KAPITEL 3 3 —HANDLINGSPLAN FÖR UTVIDGNINGEN
3 3 0Handlingsplan för utvidgningen
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
1550000 | — | 1550000 |
Anmärkningar
Detta anslag är avsett att täcka genomförandet av handlingsplanen för utvidgningen för att förbättra arbetsmiljönivån i de tio nya medlemsstaterna. Aktiviteterna omfattar i synnerhet åtgärder för att höja medvetenheten och kunskapsöverföring till små och medelstora företag.
KAPITEL 3 4 —PHAREPROGRAM IV (ÖRONMÄRKT)
3 4 0PHAREPROGRAM IV (öronmärkt)
Anmärkningar
Detta kapitel innefattar förberedande åtgärder för Kroatiens och Turkiets framtida deltagande i arbetsmiljöbyrån. Ett Phare IV-program till ett totalt belopp av 450000 euro har godkänts av gemenskapen och kommer att omfatta perioden 2006–2007. Verksamheten inom ramen för Phare IV är knuten till det godkända arbetsprogrammet med öronmärkta inkomster och utgifter. Siffrorna visar verksamhetsnivåer 2006 och 2007. Saldon för vilka inga åtaganden gjorts kommer att överföras till 2007.
3 4 0 0Löner för utlandsstationerad/internationell personal
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 67500 | 67500 |
3 4 1 0Resekostnader (internationella)
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 45000 | 45000 |
3 4 1 1Utgifter för tjänsteresor för projektpersonal utomlands
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 3110 | 3110 |
3 4 1 2Utgifter för tjänsteresor för seminarie-/konferensdeltagare
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 6000 | 6000 |
3 4 2 0Översättning/tolkar
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 27840 | 27840 |
3 4 3 0Workshop i samband med Europaveckan
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 44000 | 44000 |
3 4 4 0Webbansvariga, stöd till kontaktpunkterna
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 75600 | 75600 |
3 4 4 1Datautrustning
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 4800 | 4800 |
3 4 5 0Inventarier
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 4000 | 4000 |
3 4 6 0Tryckning av informationsmaterial
Budgetår 2006 | ÄB 1/2006 | Totalt 2006 |
| 24070 | 24070 |
--------------------------------------------------
Kommissionens beslut
av den 17 februari 2006
om vissa skyddsåtgärder i samband med högpatogen aviär influensa hos vilda fåglar i gemenskapen och om upphävande av besluten 2006/86/EG, 2006/90/EG, 2006/91/EG, 2006/94/EG, 2006/104/EG och 2006/105/EG
[delgivet med nr K(2006) 554]
(Text av betydelse för EES)
(2006/115/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA BESLUT
med beaktande av rådets direktiv 89/662/EEG av den 11 december 1989 om veterinära kontroller vid handeln inom gemenskapen i syfte att fullborda den inre marknaden [1], särskilt artikel 9.4,
med beaktande av rådets direktiv 90/425/EEG av den 26 juni 1990 om veterinära och avelstekniska kontroller i handeln med vissa levande djur och varor inom gemenskapen med sikte på att förverkliga den inre marknaden [2], särskilt artikel 10.4,
med beaktande av Europaparlamentets och rådets förordning (EG) nr 998/2003 av den 26 maj 2003 om djurhälsovillkor som skall tillämpas vid transporter av sällskapsdjur utan kommersiellt syfte och om ändring av rådets direktiv 92/65/EEG [3], särskilt artikel 18, och
av följande skäl:
(1) Aviär influensa är en smittsam virussjukdom hos fjäderfä och fåglar, som orsakar dödlighet och störningar som snabbt kan anta epizootiska proportioner, vilket i sin tur kan utgöra ett allvarligt hot mot djur- och folkhälsan och starkt minska lönsamheten inom fjäderfäuppfödningen. Det finns en risk för att sjukdomsagenset sprids från vilda fåglar till tamfåglar, framför allt fjäderfä, och från en medlemsstat till andra medlemsstater och tredjeländer via internationell handel med levande fåglar eller produkter från dem.
(2) Fall av högpatogen aviär influensa av subtyp H5N1 misstänks eller har bekräftats i flera medlemsstater. Kommissionen har redan antagit tillfälliga skyddsåtgärder. Med hänsyn till den epidemiologiska situationen bör de skyddsåtgärder som är nödvändiga vidtas på gemenskapsnivå i syfte att förhindra att sjukdomen sprids från vilda fåglar till fjäderfä.
(3) Om ett aviärt influensavirus av subtyp H5 har isolerats i ett kliniskt fall hos vilda fåglar inom en medlemsstats territorium och om, i avvaktan på att neuraminidastyp (N) och patogenitetsindex bestäms, den kliniska bilden och de epidemiologiska omständigheterna ger anledning att misstänka att det rör sig om högpatogen aviär influensa orsakad av influensavirus A av subtyp H5N1 eller förekomsten av denna subtyp har bekräftats, skall den berörda medlemsstaten tillämpa vissa skyddsåtgärder för att minimera risken för fjäderfä.
(4) De särskilda åtgärder som föreskrivs i detta beslut skall tillämpas utan att det påverkar de åtgärder som medlemsstaterna skall vidta enligt rådets direktiv 92/40/EEG av den 19 maj 1992 om införande av gemenskapsåtgärder för bekämpning av aviär influensa [4].
(5) För konsekvensens skull bör vissa definitioner som fastställs i rådets direktiv 2005/94/EG av den 20 december 2005 om gemenskapsåtgärder för bekämpning av aviär influensa och om upphävande av direktiv 92/40/EEG [5], rådets direktiv 90/539/EEG av den 15 oktober 1990 om djurhälsovillkor för handel inom gemenskapen med och för import från tredje land av fjäderfä och kläckningsägg [6], Europaparlamentets och rådets förordning (EG) nr 853/2004 av den 29 april 2004 om fastställande av särskilda hygienregler för livsmedel av animaliskt ursprung [7] och i Europaparlamentets och rådets förordning (EG) nr 998/2003 av den 26 maj 2003 om djurhälsovillkor som skall tillämpas vid transporter av sällskapsdjur utan kommersiellt syfte och om ändring av rådets direktiv 92/65/EEG [8] tillämpas på det här beslutet.
(6) Skydds- och övervakningsområden bör upprättas runt den plats där sjukdomen påvisats hos vilda fåglar. Dessa områden bör begränsas till det nödvändiga för att förhindra att viruset införs i kommersiella och icke kommersiella fjäderfäflockar.
(7) Förflyttning av främst levande fåglar och kläckägg bör kontrolleras och begränsas medan kontrollerad sändning av dessa fåglar och fågelprodukter bör tillåtas på vissa villkor.
(8) De åtgärder som fastställs i kommissionens beslut 2005/734/EG av den 19 oktober 2005 om fastställande av åtgärder för biosäkerhet för att minska risken för överföring av högpatogen aviär influensa orsakad av influensavirus A av subtyp H5N1 från viltlevande fåglar till fjäderfä och andra fåglar i fångenskap och om ett system för tidig upptäckt i särskilt riskutsatta områden [9] bör tillämpas i skydds- och övervakningsområden, oberoende av den riskstatus som fastställts för det område där högpatogen aviär influensa misstänks eller har bekräftats hos vilda fåglar.
(9) I rådets direktiv 92/65/EEG av den 13 juli 1992 om fastställande av djurhälsokrav i handeln inom och importen till gemenskapen av djur, sperma, ägg (ova) och embryon som inte faller under de krav som fastställs i de specifika gemenskapsregler som avses i bilaga A.I till direktiv 90/425/EEG [10] fastställs godkända organ, institut och center samt en förlaga till hälsointyg som skall åtfölja djuren eller deras könsceller mellan sådana godkända anläggningar i olika medlemsstater. Ett undantag från transportrestriktioner bör göras för fåglar från och på väg till organ, institut och center som godkänts enligt det direktivet.
(10) Transport av kläckägg från skyddszonerna bör tillåtas på vissa villkor. Sändning av kläckägg till andra länder får tillåtas framför allt om de uppfyller villkoren i direktiv 2005/94/EG. I sådana fall bör det djurhälsointyg som utfärdas i enlighet med direktiv 90/529/EEG innehålla en hänvisning till det här beslutet.
(11) Sändning av kött, malet kött, köttberedningar och köttprodukter från skyddsområdena bör tillåtas under förutsättning att vissa villkor, främst vissa krav i förordning (EG) nr 853/2004 och i Europaparlamentets och rådets förordning (EG) nr 854/2004 av den 29 april 2004 om fastställande av särskilda bestämmelser för genomförandet av offentlig kontroll av produkter av animaliskt ursprung avsedda att användas som livsmedel [11] uppfylls.
(12) I rådets direktiv 2002/99/EG av den 16 december 2002 om fastställande av djurhälsoregler för produktion, bearbetning, distribution och införsel av produkter av animaliskt ursprung avsedda att användas som livsmedel [12] upprättas en förteckning över behandlingar som gör kött från områden där restriktioner gäller säkra samt fastställs möjligheten att inrätta ett särskilt kontrollmärke och den identifieringsmärkning som krävs för kött som av djurhälsoskäl inte får släppas ut på marknaden. Det bör vara tillåtet att från skyddsområdena sända kött som är märkt med det kontrollmärke som fastställs i det direktivet och köttprodukter som genomgått den behandling som avses i det direktivet.
(13) Enligt Europaparlamentets och rådets förordning (EG) nr 1774/2002 av den 3 oktober 2002 om hälsobestämmelser för animaliska biprodukter som inte är avsedda att användas som livsmedel [13] är det tillåtet att släppa ut en rad animaliska biprodukter på marknaden, t.ex. gelatin för teknisk användning, material för farmaceutiska ändamål och annat, med ursprung i områden i gemenskapen som omfattas av restriktioner av djurhälsoskäl, eftersom dessa produkter anses säkra på grund av de särskilda villkoren för produktion, bearbetning och användning som effektivt inaktiverar eventuella patogener eller förhindrar kontakt med mottagliga djur.
(14) Detta beslut bör ses över mot bakgrund av genomförandet av direktiv 2005/94/EG i medlemsstaterna.
(15) Efter anmälan av fall av högpatogen aviär influensa orsakad av influensavirus A av subtyp H5N1 hos vilda fåglar i Grekland, Italien och Slovenien antog kommissionen i samarbete med de berörda medlemsstaterna besluten 2006/86/EG [14], 2006/90/EG [15], 2006/91/EG [16], 2006/94/EG [17], 2006/104/EG [18] och 2006/105/EG [19] om vissa tillfälliga skyddsåtgärder i samband med misstänkta fall av högpatogen aviär influensa hos vilda fåglar i respektive medlemsstat. Dessa beslut bör upphöra att gälla.
(16) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Syfte, tillämpningsområde och definitioner
1. I detta beslut fastställs vissa skyddsåtgärder som skall tillämpas när högpatogen aviär influensa orsakad av influensavirus A av subtyp H5 har isolerats hos vilda fåglar inom en medlemsstats territorium (nedan kallad %quot%berörd medlemsstat%quot%) och som misstänks eller har bekräftats vara av neuraminidastyp N1, för att förhindra spridning av aviär influensa från vilda fåglar till fjäderfä eller andra fåglar i fångenskap liksom kontaminering av produkter av dessa fåglar.
2. Om inte annat fastställs skall definitionerna i direktiv 2005/95/EG gälla. Därutöver skall följande definitioner gälla:
kläckägg : ägg enligt definitionen i artikel 2.2 i direktiv 90/539/EEG.
viltlevande fågelvilt : vilt enligt definitionen i punkt 1.5 andra strecksatsen och punkt 1.7 i bilaga I till förordning (EG) nr 853/2004.
andra fåglar i fångenskap i) sällskapsdjur av de fågelarter som avses i artikel 3 a i förordning (EG) nr 998/2003 samt
ii) fåglar för djurparker, cirkusar, nöjesparker och försökslaboratorier.
Artikel 2
Upprättande av skydds- och övervakningsområden
1. Den berörda medlemsstaten skall runt det område där högpatogen aviär influensa orsakad av influensavirus A av subtyp H5 har bekräftats hos vilda fåglar och neuraminidastyp N1 antingen misstänks eller har bekräftats upprätta
a) ett skyddsområde med en radie på minst 3 km och
b) ett övervakningsområde med en radie på minst 10 km innefattande skyddsområdet.
2. De skydds- och övervakningsområden som avses i punkt 1 skall upprättas med hänsyn till geografiska, administrativa, ekologiska och epizootologiska faktorer i samband med aviär influensa och med hänsyn till kontrollmöjligheterna.
3. Om skydds- eller övervakningsområdena omfattar andra medlemsstaters territorium skall den berörda medlemsstaten samarbeta med myndigheterna i dessa medlemsstater för att upprätta områdena.
4. Den berörda medlemsstaten skall till kommissionen och de övriga medlemsstaterna överlämna närmare uppgifter om eventuella skydds- och övervakningsområden som upprättas enligt denna artikel samt på lämpligt sätt informera allmänheten om de åtgärder som vidtagits.
Artikel 3
Åtgärder i skyddsområdet
1. Den berörda medlemsstaten skall se till att minst följande åtgärder vidtas i skyddsområdet:
a) Kartläggning av samtliga anläggningar inom området.
b) Regelbundna och dokumenterade besök i alla kommersiella anläggningar med en klinisk undersökning av fjäderfän och, vid behov, provtagning för laboratorieundersökning.
c) Genomförande av lämpliga åtgärder för biosäkerhet på jordbruksföretaget, inklusive användning av lämpliga desinfektionsmedel vid anläggningens in- och utgångar, inhysning eller instängning av fjäderfä i byggnader där direkt eller indirekt kontakt med annat fjäderfä eller andra fåglar i fångenskap kan förhindras.
d) Genomförande av de åtgärder för biosäkerhet som fastställs i beslut 2005/734/EG.
e) Kontroll av förflyttningar av fjäderfäprodukter i enlighet med artikel 9.
f) Aktiv sjukdomsövervakning bland vildfågelpopulationen, främst bland sjöfåglar, vid behov i samarbete med jägare och fågelskådare, som har fått särskilda instruktioner om hur de skall skydda sig själva mot infektion av viruset och hur man kan förhindra att viruset sprids till mottagliga djur.
g) Kampanjer för att informera allmänheten och för att öka medvetenheten om sjukdomen bland fågelägare, jägare och fågelskådare.
2. Den berörda medlemsstaten skall se till att följande förbjuds i skyddsområdet:
a) Avlägsnande av fjäderfä och andra fåglar i fångenskap från den anläggning där de hålls.
b) Sammanförande av fjäderfä och andra fåglar i fångenskap vid mässor, marknader, uppvisningar och övriga sammankomster.
c) Transport av fjäderfä och andra fåglar i fångenskap genom området, utom transitering på huvudleder eller järnväg samt transport till ett slakteri för direkt slakt.
d) Sändning av kläckägg från området.
e) Sändning av färskt kött, malet kött, köttberedningar och köttprodukter från fjäderfä, andra fåglar i fångenskap och viltlevande fågelvilt från området.
f) Transport eller spridning av obearbetat använt strö eller fjäderfägödsel utanför området från anläggningar inom området, utom transport för behandling i enlighet med förordning (EG) nr 1774/2002.
g) Jakt på vilda fåglar.
Artikel 4
Åtgärder i övervakningsområdet
1. Den berörda medlemsstaten skall se till att minst följande åtgärder vidtas i övervakningsområdet:
a) Kartläggning av samtliga anläggningar inom området.
b) Genomförande av lämpliga åtgärder för biosäkerhet på jordbruksföretaget, inklusive användning av lämpliga desinfektionsmedel vid anläggningens in- och utgångar.
c) Genomförande av de åtgärder för biosäkerhet som fastställs i beslut 2005/734/EG.
d) Kontroll av förflyttningar av fjäderfä, andra fåglar i fångenskap och kläckägg inom området.
2. Den berörda medlemsstaten skall se till att följande förbjuds i övervakningsområdet:
a) Förflyttning av fjäderfä och andra fåglar i fångenskap ut ur området under de första 15 dagarna efter det att området har upprättats.
b) Sammanförande av fjäderfä och andra fåglar vid mässor, marknader, uppvisningar och övriga sammankomster.
c) Jakt på vilda fåglar.
Artikel 5
Åtgärdernas varaktighet
Om neuraminidastypen bekräftas vara en annan än N1 eller om viruset har låg patogenitet skall åtgärderna i artiklarna 3 och 4 upphävas.
Om förekomst av ett högpatogent influensavirus A, särskilt av subtyp H5N1, bekräftas hos vilda fåglar skall åtgärderna i artiklarna 3 och 4 vidtas så länge det är nödvändigt med hänsyn till de geografiska, administrativa, ekologiska och epizootologiska faktorerna i samband med aviär influensa och i minst 21 dagar inom skyddsområdet och i minst 30 dagar inom övervakningsområdet efter den dag då ett aviärt influensavirus av subtyp H5 isolerades i ett kliniskt fall hos vilda fåglar.
Artikel 6
Undantag för levande fåglar och dagsgamla kycklingar
1. Genom undantag från artikel 3.2 a får den berörda medlemsstaten tillåta transport av värpfärdiga unghöns, slaktkalkoner och annat fjäderfä och fågelvilt i hägn till anläggningar under officiell översyn i antingen skydds- eller övervakningsområdet.
2. Genom undantag från artiklarna 3.2 a och 4.2 a får den berörda medlemsstaten tillåta transport av
a) fjäderfä, inklusive uttjänta värphöns, för omedelbar slakt till ett slakteri i skydds- eller övervakningsområdet eller, om detta inte är möjligt, till ett slakteri som den behöriga myndigheten anvisat utanför områdena,
b) dagsgamla kycklingar från skyddsområdet till anläggningar som står under officiell översyn inom den berörda medlemsstatens territorium, under förutsättning att det på den mottagande anläggningen inte finns några andra fjäderfän eller fåglar i fångenskap, bortsett från sällskapsfåglar enligt artikel 1.2 c i som hålls avskilda från fjäderfä, eller att transporten sker enligt de villkor som beskrivs i artikel 24.1 a och 24.1 b i direktiv 2005/94/EG och fjäderfäna stannar kvar på den mottagande anläggningen under 21 dagar,
c) dagsgamla kycklingar från övervakningsområdet till anläggningar som står under officiell översyn på den berörda medlemsstatens territorium,
d) värpfärdiga unghöns, slaktkalkoner och annat fjäderfä och fågelvilt i hägn från övervakningsområdet till anläggningar under officiell översyn på den berörda medlemsstatens territorium,
e) sällskapsfåglar enligt artikel 1.2 c i till anläggningar på den berörda medlemstatens territorium där inget fjäderfä hålls, om sändningen består av högst fem burfåglar, trots nationella regler enligt artikel 1 tredje stycket i direktiv 92/65/EEG,
f) fåglar enligt artikel 1.2 c ii från organ, institut och center och på väg mot andra sådana organ, institut och center som godkänts i enlighet med artikel 13 i direktiv 92/65/EEG.
Artikel 7
Undantag för kläckägg
1. Genom undantag från artikel 3.2 d får den berörda medlemsstaten tillåta
a) transport av kläckägg från skyddsområdet till ett anvisat kläckeri inom den berörda medlemsstatens territorium,
b) sändning av kläckägg från skyddsområdet till kläckerier utanför den berörda medlemsstatens territorium, under förutsättning att
i) kläckäggen har samlats in från flockar som
- inte misstänks vara smittade med aviär influensa och
- med negativt resultat har genomgått en serologisk undersökning för aviär influensa som kan påvisa en prevalens på 5 % med ett konfidensintervall på minst 95 % och
ii) villkoren i artikel 26.1 b, 26.1 c och 26.1 d i direktiv 2005/94/EG har uppfyllts.
2. Djurhälsointygen i enlighet med förlaga 1 i bilaga IV till rådets direktiv 90/539/EEG som åtföljer sändningar av de kläckägg som avses i punkt 1 b till andra medlemsstater skall innehålla följande fras:
%quot%Denna sändning uppfyller djurhälsovillkoren i kommissionens beslut 2006/115/EG.%quot%
Artikel 8
Undantag för kött, malet kött, köttberedningar, maskinurbenat kött och köttprodukter
1. Genom undantag från artikel 3.2 e får den berörda medlemsstaten tillåta sändning av följande från skyddsområdet:
a) Färskt fjäderfäkött, inklusive kött från ratiter, med ursprung i eller utanför området som har producerats i enlighet med bilaga II och avsnitten II och III i bilaga III till förordning (EG) nr 853/2004 och kontrollerats i enlighet med avsnitten I, II och III samt avsnitt IV kapitlen V och VII i bilaga I till förordning (EG) nr 854/2004.
b) Malet kött, köttberedningar, maskinurbenat kött och köttprodukter som innehåller kött som avses i punkt a och som producerats i enlighet med avsnitten V och VI i bilaga III till förordning (EG) nr 853/2004.
c) Färskt kött av viltlevande fågelvilt med ursprung i området, om köttet är märkt med det kontrollmärke som fastställs i bilaga II till direktiv 2002/99/EG och är avsett för transport till en anläggning för den behandling som krävs för aviär influensa i enlighet med bilaga III till det direktivet.
d) Köttprodukter av kött från viltlevande fågelvilt som har genomgått en behandling som krävs för aviär influensa i enlighet med bilaga III till direktiv 2002/99/EG.
e) Färskt kött av viltlevande fågelvilt med ursprung utanför skyddsområdet som producerats på anläggningar inom skyddsområdet i enlighet med avsnitt IV i bilaga III till förordning (EG) nr 853/2004 och kontrollerats i enlighet med avsnitt IV kapitel VIII i bilaga I till förordning (EG) nr 854/2004.
f) Malet kött, köttberedningar, maskinurbenat kött och köttprodukter som innehåller kött som avses i punkt e och som producerats på anläggningar inom skyddsområdet i enlighet med avsnitten V och VI i bilaga III till förordning (EG) nr 853/2004.
2. Den berörda medlemsstaten skall se till att de produkter som avses i punkt 1 e och 1 f åtföljs av ett handelsdokument där följande anges:
%quot%Denna sändning uppfyller djurhälsovillkoren i kommissionens beslut 2006/115/EG.%quot%
Artikel 9
Villkor för animaliska biprodukter
1. I enlighet med artikel 3.1 e får den berörda medlemsstaten tillåta sändning av följande:
a) Animaliska biprodukter som uppfyller villkoren i kapitlen II.A, III.B, IV.A, VI.A, VI.B, VII.A, VIII.A, IX.A och X.A i bilaga VII, och kapitlen II.B och III.II.A i bilaga VIII till förordning (EG) nr 1774/2002.
b) Obearbetade fjädrar och delar av fjädrar enligt kapitel VIII.A.1 a i bilaga VIII till förordning (EG) nr 1774/2002 från fjäderfä som kommer från utanför skyddsområdet.
c) Bearbetade fjädrar från fjäderfä eller delar av fjädrar från fjäderfä som har behandlats med ånga eller med någon annan metod som säkerställer att inga patogener återstår.
d) Produkter som härrör från fjäderfä eller andra fåglar i fångenskap som i enlighet med gemenskapslagstiftningen inte omfattas av några djurhälsokrav eller som inte omfattas av några förbud eller restriktioner av djurhälsoskäl, inklusive de produkter som avses i kapitel VII.A.1 a i bilaga VIII till förordning (EG) nr 1774/2002.
2. Den berörda medlemsstaten skall se till att de produkter som anges i punkt 1 b och 1 c i denna artikel åtföljs av ett handelsdokument i enlighet med kapitel X i bilaga II till förordning (EG) nr 1774/2002 och i punkt 6.1 i det dokumentet, för de produkter som avses i punkt 1 c i denna artikel, ange att dessa produkter har behandlats med ånga eller med någon annan metod som säkerställer att inga patogener återstår.
Handelsdokumentet skall dock inte krävas för bearbetade dekorationsfjädrar, bearbetade fjädrar som medförs av resande för privat bruk eller sändningar av bearbetade fjädrar som sänts till privatpersoner för icke-industriellt syfte.
Artikel 10
Villkor för förflyttning
1. Om förflyttning av djur eller produkter från dessa som omfattas av detta beslut tillåts enligt artikel 6, 7, 8 eller 9, skall tillståndet grundas på ett positivt resultat av en riskbedömning som gjorts av den behöriga myndigheten och alla åtgärder vidtas som ur biosäkerhetssynpunkt är nödvändiga för att förhindra spridning av aviär influensa.
2. Om sändning, förflyttning eller transport av produkter som avses i punkt 1 tillåts enligt artikel 7, 8 eller 9, enligt motiverade villkor eller restriktioner, skall de produceras, hanteras, behandlas, lagras och transporteras på ett sådant sätt att de inte äventyrar djurhälsosituationen för andra produkter som uppfyller samtliga djurhälsokrav för handel, utsläppande på marknaden eller export till tredjeländer.
Artikel 11
Efterlevnad av bestämmelserna
Alla medlemsstater skall genast anta och offentliggöra de åtgärder som är nödvändiga för att följa detta beslut. De skall genast underrätta kommissionen om detta.
Den berörda medlemsstaten skall tillämpa dessa åtgärder så snart den rimligen misstänker förekomst av virus av högpatogen aviär influensa, särskilt av subtyp H5N1.
Den berörda medlemsstaten skall till kommissionen och de övriga medlemsstaterna regelbundet överlämna nödvändig information om sjukdomsepidemiologin, i lämpliga fall om ytterligare kontroll- och övervakningsåtgärder och upplysningskampanjer, och alltid förhandsinformation om planerat upphävande av åtgärder i enlighet med artikel 5.
Artikel 12
Upphävande
Kommissionens beslut 2006/86/EG, 2006/90/EG, 2006/91/EG, 2006/94/EG, 2006/104/EG och 2006/105/EG skall upphöra att gälla.
Artikel 13
Adressat
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 12 april 2006
om ändring av beslut 2003/526/EG när det gäller skyddsåtgärder mot klassisk svinpest i Tyskland
[delgivet med nr K(2006) 1521]
(Text av betydelse för EES)
(2006/284/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA BESLUT
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 90/425/EEG av den 26 juni 1990 om veterinära och avelstekniska kontroller i handeln med vissa levande djur och varor inom gemenskapen med sikte på att förverkliga den inre marknaden [1], särskilt artikel 10.4, och
av följande skäl:
(1) Till följd av utbrotten av klassisk svinpest i vissa medlemsstater antogs kommissionens beslut 2003/526/EG av den 18 juli 2003 om skyddsåtgärder mot klassisk svinpest i vissa medlemsstater [2]. I det beslutet fastställs vissa ytterligare åtgärder för bekämpning av klassisk svinpest.
(2) Tyskland har informerat kommissionen om den senaste utvecklingen av sjukdomen bland viltlevande svin i delstaten Nordrhein-Westfalen. Mot bakgrund av tillgängliga epidemiologiska uppgifter bör de områden i Tyskland där det vidtas åtgärder för att bekämpa sjukdomen utvidgas till att omfatta vissa områden i Nordrhein-Westfalen och angränsande områden i Rheinland-Pfalz.
(3) Situationen i andra områden av delstaten Rheinland-Pfalz har förbättrats markant. De åtgärder som föreskrivs i beslut 2003/526/EG angående dessa områden bör därför inte längre tillämpas.
(4) Beslut 2003/526/EG bör därför ändras i enlighet med detta.
(5) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Bilagan till beslut 2003/526/EG skall ersättas med bilagan till det här beslutet.
Artikel 2
Detta beslut riktar sig till medlemsstaterna.
Kommissionens beslut
av den 19 april 2006
om tillsättande av en expertgrupp som skall ge kommissionen råd i policyfrågor i kampen mot radikalisering med ökat våld
(2006/299/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR BESLUTAT FÖLJANDE
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, och
av följande skäl:
(1) Enligt artikel 2 i fördraget om Europeiska unionen skall unionen bevara och utveckla unionen som ett område med frihet, säkerhet och rättvisa.
(2) Europeiska unionen skall ge medborgarna en hög säkerhetsnivå inom området med frihet, säkerhet och rättvisa. Detta mål skall nås genom bekämpande av terrorism, även den yttre dimensionen av detta hot, och genom att vidta åtgärder mot de faktorer som bidrar till radikalisering med ökat våld.
(3) I sitt meddelande Terroristattacker: förebyggande, beredskap och insatser [1] fastslog kommissionen att kampen mot extremistiskt våld i samhället och försvårandet av rekryteringen av terrorister måste vara grundläggande prioriteringar i en strategi för att förebygga terrorism.
(4) I sitt meddelande Rekrytering till terrorism: faktorer som bidrar till radikalisering med ökat våld [2] erkände kommissionen behovet av att anlita sakkunskapen hos specialister för att vidareutveckla sin politik på detta område.
(5) Gruppen skall bestå av specialister från olika vetenskapsgrenar med erfarenhet av att analysera och forska i radikalisering med ökat våld eller på områden med direkt anknytning till detta.
(6) En expertgrupp om radikalisering med ökat våld bör därför tillsättas och dess behörighet och struktur fastställas närmare.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Härmed tillsätter kommissionen en expertgrupp som skall ge råd i policyfrågor, expertgruppen om radikalisering med ökat våld (nedan kallad "gruppen").
2. Expertgruppen skall bestå av kvalificerade personer med tillräcklig kompetens att kunna bedöma frågor som gäller radikalisering med ökat våld och terrorism.
Artikel 2
Uppgifter
Kommissionen kan rådfråga gruppen i alla frågor som gäller radikalisering med ökat våld och terrorism.
Gruppen skall ha följande uppgifter:
- Samla ledamöternas sakkunskap för att ge kommissionen råd i policyfrågor. Sådan rådgivning kan ske antingen på gruppens eget initiativ eller på kommissionens uttryckliga begäran.
- Hjälpa kommissionen att identifiera nya områden för nödvändig forskning i fenomenet radikalisering med ökat våld och terrorism.
- Utbyta sakkunskap med nätverk, institut eller andra EU-organ, i medlemsstaterna, tredjeland eller med internationella organisationer som är verksamma på samma område.
- Särskilt utarbeta en sammanfattande rapport senast i juni 2006 om forskningsläget på området radikalisering med ökat våld.
Gruppens ordförande kan meddela kommissionen om att det vore lämpligt att höra gruppen i en viss fråga.
Artikel 3
Sammansättning och utnämning av gruppens ledamöter
1. Gruppens ledamöter skall utses av generaldirektören för Europeiska kommissionens generaldirektorat för rättvisa, frihet och säkerhet bland specialister med kompetens på områdena radikalisering med ökat våld och terrorism. En sådan kompetens måste omfatta erfarenhet förvärvad genom akademisk forskning och publicerade arbeten.
2. Gruppen skall bestå av högst 20 ledamöter.
3. Följande skall gälla:
- Ledamöterna skall utnämnas personligen och ha i uppgift att ge råd till kommissionen oberoende av påverkan utifrån.
- Gruppens ledamöter skall utnämnas för en mandatperiod på ett år, som kan förlängas av kommissionen. De skall ha kvar sitt uppdrag till dess att de avgår, ersätts eller deras mandat upphör.
- De ledamöter som inte längre på ett effektivt sätt kan medverka i gruppens arbete, som avgår eller som bryter mot de bestämmelser som fastställs i den första eller andra strecksatsen i denna artikel eller i artikel 287 i fördraget om upprättandet av Europeiska gemenskapen får ersättas under resten av sitt mandat.
- Medlemmarna skall varje år avge en skriftlig försäkran om att de förbinder sig att agera i allmänhetens intresse och en försäkran om avsaknaden eller förekomsten av intressekonflikter som skulle kunna påverka deras oberoende ställning.
Artikel 4
Verksamhet
1. Generaldirektören för generaldirektoratet för rättvisa, frihet och säkerhet utnämner gruppens ordförande.
Gruppen skall lägga fram yttranden och rapporter för kommissionen. Innehållet i sådana rapporter och yttranden är inte bindande för kommissionen eller någon annan EU-institution. Kommissionen får fastställa en tidsfrist inom vilken ett yttrande eller en rapport skall läggas fram.
Om gruppen är enig om ett yttrande eller en rapport skall den utarbeta gemensamma slutsatser som skall bifogas mötesprotokollen. Om gruppen inte kan enas om ett yttrande eller en rapport, skall den underrätta kommissionen om de skiljaktiga ståndpunkterna.
2. Med kommissionens samtycke får undergrupper inrättas för att undersöka särskilda frågor inom ramen för ett mandat som fastställs av gruppen; dessa undergrupper skall upplösas när uppdraget har slutförts. Rapporter som sammanställts av sådana undergrupper måste godkännas av gruppen, och samma bestämmelser i stycket ovan gäller i fall där enighet inte nås.
3. Företrädaren för kommissionen har rätt att be andra experter eller observatörer med särskild kompetens i ett ämne på dagordningen att medverka i gruppens eller undergruppens överläggningar om detta är nyttigt och/eller nödvändigt.
4. Information som erhålls genom deltagande i gruppens eller undergruppernas överläggningar måste betraktas som konfidentiell och får endast röjas om kommissionen uttryckligen säger att detta får göras. Varje ledamot av gruppen och/eller dess undergrupper förblir bunden av sekretessreglerna efter det att deras mandat löpt ut.
5. Gruppen och dess undergrupper skall normalt sammanträda i kommissionens lokaler i enlighet med de förfaranden och tidsplaner som kommissionen fastställer. Kommissionen tillhandahåller sekreterartjänster. Berörda tjänstemän från kommissionen får delta i sammanträdena.
6. Gruppen skall anta sin arbetsordning på grundval av den standardiserade arbetsordning som antagits av kommissionen.
7. Kommissionen får offentliggöra på Internet alla sammanfattningar, slutsatser, delar av slutsatser eller arbetsdokument från gruppen på det aktuella dokumentets originalspråk som inte är konfidentiella. De dokument som gruppen lägger fram omfattas av bestämmelserna i Europaparlamentets och rådets förordning (EG) nr 1049/2001 [3].
Artikel 5
Sammanträdesutgifter
Kommissionen skall ersätta utgifter för resor och, om det anses lämpligt, uppehälle för ledamöter, andra experter och observatörer i samband med gruppens verksamhet i enlighet med kommissionens interna regler om ersättning av externa experters utgifter.
Ledamöterna, eller andra experter och observatörer som kan bjudas in ibland, skall inte få ersättning för sin verksamhet och sina funktioner.
Artikel 6
Ikraftträdande
Detta beslut börjar gälla samma dag som det offentliggörs i Europeiska unionens officiella tidning. Det gäller till den 19 mars 2007. Före detta datum skall kommissionen bestämma om eventuell förlängning.
Rådets beslut
av den 14 februari 2006
om ingående av Europa–Medelhavsavtalet om upprättande av en associering mellan Europeiska gemenskapen och dess medlemsstater, å ena sidan, och Republiken Libanon, å andra sidan
(2006/356/EG)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 310 jämförd med artikel 300.2 första stycket andra meningen och artikel 300.3 andra stycket,
med beaktande av kommissionens förslag,
med beaktande av Europaparlamentets samtycke, och
av följande skäl:
(1) Europa–Medelhavsavtalet om upprättande av en associering mellan Europeiska gemenskapen och dess medlemsstater, å ena sidan, och Republiken Libanon, å andra sidan, undertecknades på Europeiska gemenskapens vägnar i Luxemburg den 17 juni 2002, med förbehåll för dess ingående.
(2) Avtalet bör godkännas.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Europa–Medelhavsavtalet om upprättande av en associering mellan Europeiska gemenskapen och dess medlemsstater, å ena sidan, och Republiken Libanon, å andra sidan, bilagorna och protokollen till avtalet samt de gemensamma förklaringar och förklaringar från Europeiska gemenskapen som åtföljer slutakten godkänns härmed på Europeiska gemenskapens vägnar.
2. De texter som nämns i punkt 1 åtföljer detta beslut.
Artikel 2
1. Den ståndpunkt som gemenskapen skall inta i associeringsrådet och associeringskommittén skall fastställas av rådet på förslag av kommissionen eller, i förekommande fall, av kommissionen i enlighet med de relevanta bestämmelserna i fördragen.
2. Rådets ordförande skall i enlighet med artikel 75 i Europa–Medelhavsavtalet utöva ordförandeskapet i associeringsrådet. En företrädare för kommissionen skall utöva ordförandeskapet i associeringskommittén i enlighet med de överenskomna förfarandereglerna.
3. Beslut om att offentliggöra associeringsrådets och associeringskommitténs beslut i Europeiska unionens officiella tidning skall fattas från fall till fall av rådet respektive av kommissionen.
Artikel 3
Rådets ordförande bemyndigas härmed att utse den eller de personer som på Europeiska gemenskapens vägnar har rätt att deponera den anmälan som avses i artikel 91 i avtalet.
Rådets beslut
av den 29 april 2004
om undertecknande och provisorisk tillämpning av ett protokoll till avtalet om partnerskap och samarbete om upprättande av ett partnerskap mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Republiken Uzbekistan, å andra sidan, för att beakta Republiken Tjeckiens, Republiken Estlands, Republiken Cyperns, Republiken Lettlands, Republiken Litauens, Republiken Ungerns, Republiken Maltas, Republiken Polens, Republiken Sloveniens och Republiken Slovakiens anslutning till Europeiska unionen
(2006/458/EG)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artiklarna 44.2, 47.2 sista meningen, artikel 55, artikel 57.2, artikel 71, artikel 80.2, artiklarna 93, 94, 133 och 181a jämförda med artikel 300.2 första stycket första meningen,
med beaktande av anslutningsfördraget av den 16 april 2003, särskilt artikel 2.3,
med beaktande av den akt, som är bifogad anslutningsfördraget, särskilt artikel 6.2,
med beaktande av kommissionens förslag, och
av följande skäl:
(1) Den 8 december 2003 bemyndigade rådet kommissionen att, på gemenskapens och dess medlemsstaters vägnar, med Republiken Uzbekistan förhandla fram ett protokoll till avtalet om partnerskap och samarbete i syfte att beakta Republiken Tjeckiens, Republiken Estlands, Republiken Cyperns, Republiken Lettlands, Republiken Litauens, Republiken Ungerns, Republiken Maltas, Republiken Polens, Republiken Sloveniens och Republiken Slovakiens anslutning till Europeiska unionen samt att föreskriva vissa tekniska anpassningar som sammanhänger med den institutionella och rättsliga utvecklingen inom Europeiska unionen.
(2) Protokollet har förhandlats fram mellan parterna och bör nu undertecknas på Europeiska gemenskapens och dess medlemsstaters vägnar, med förbehåll för att det senare ingås.
(3) Protokollet bör tillämpas provisoriskt från och med dagen för anslutningen till dess att de relevanta förfarandena för det formella ingåendet har slutförts.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Rådets ordförande bemyndigas att utse den eller de personer som, på Europeiska gemenskapens och dess medlemsstaters vägnar, skall ha rätt att underteckna protokollet till avtalet om partnerskap och samarbete om upprättande av ett partnerskap mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Republiken Uzbekistan, å andra sidan, i syfte att beakta Republiken Tjeckiens, Republiken Estlands, Republiken Cyperns, Republiken Lettlands, Republiken Litauens, Republiken Ungerns, Republiken Maltas, Republiken Polens, Republiken Sloveniens och Republiken Slovakiens anslutning till Europeiska unionen, med förbehåll för att protokollet ingås i ett senare skede.
Texten till protokollet åtföljer detta beslut [1].
Artikel 2
I avvaktan på att det skall träda i kraft skall protokollet tillämpas provisoriskt från och med dagen för anslutningen.
Kommissionens beslut
av den 28 juli 2006
om vissa tillfälliga skyddsåtgärder i samband med högpatogen aviär influensa i Sydafrika
[delgivet med nr K(2006) 3350]
(Text av betydelse för EES)
(2006/532/EG)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DETTA BESLUT
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets direktiv 91/496/EEG av den 15 juli 1991 om fastställande av regler för hur veterinärkontroller skall organiseras för djur som importeras till gemenskapen från tredje land och om ändring av direktiven 89/662/EEG, 90/425/EEG och 90/675/EEG [1], särskilt artikel 18.1 och 18.6,
med beaktande av rådets direktiv 97/78/EG av den 18 december 1997 om principerna för organisering av veterinärkontroller av produkter från tredje land som förs in i gemenskapen [2], särskilt artikel 22.1 och 22.5, och
av följande skäl:
(1) Aviär influensa är en smittsam virussjukdom hos fjäderfä och andra fåglar, som orsakar dödlighet och störningar som snabbt kan nå epizootiska proportioner, vilket i sin tur kan utgöra ett allvarligt hot mot djur- och folkhälsan och starkt minska lönsamheten inom fjäderfäuppfödningen. Det finns risk för att sjukdomsagenset sprids via internationell handel med levande fjäderfä och andra fåglar eller produkter av dessa.
(2) Den 29 juni 2006 bekräftade Sydafrika att högpatogen aviär influensa hade brutit ut på en strutsfarm i Västra Kapprovinsen.
(3) Den virusstam av aviär influensa som upptäcktes under detta utbrott är av subtyp H5N2 och skiljer sig därför från den stam som orsakar den nuvarande epidemin i Asien, Nordafrika och Europa. Enligt aktuell kunskap utgör denna subtyp en mindre risk för folkhälsan än den virusstam som för närvarande är i omlopp i Asien, nämligen subtypen H5N1.
(4) Enligt nuvarande gemenskapslagstiftning har Sydafrika endast tillstånd att exportera till gemenskapen levande ratiter och kläckägg från dessa liksom färskt kött, köttberedningar och köttprodukter innehållande kött av dessa arter.
(5) Med hänsyn till den risk för djurhälsan som det skulle innebära om högpatogen aviär influensa kom in i gemenskapen bör som en omedelbar åtgärd all import från Sydafrika av levande ratiter och kläckägg från dessa arter tillfälligt upphävas.
(6) Dessutom är det lämpligt att tillfälligt upphäva import till gemenskapen från Sydafrika av färskt kött av ratiter och av köttberedningar och köttprodukter som består av eller innehåller kött av dessa arter. Med hänsyn till att sjukdomen kom in på de drabbade farmerna i mitten på juni är det dock lämpligt att besluta om ett undantag för färskt kött och köttberedningar som består av eller innehåller kött från sådana arter om fågeln slaktades före den 1 maj 2006, vilket bör vara underställt vissa villkor.
(7) Sydafrika har tillämpat stränga åtgärder för sjukdomsbekämpning och har sänt uppgifter om sjukdomssituationen till kommissionen, vilket motiverar en begränsning av importförbudet till den drabbade delen av Sydafrikas territorium.
(8) Kommissionens beslut 2005/432/EG av den 3 juni 2005 om djur- och folkhälsovillkor och förlagor till hälsointyg för import från tredjeländer av köttprodukter avsedda att användas som livsmedel och om upphävande av besluten 97/41/EG, 97/221/EG och 97/222/EG [3] innehåller en förteckning över de tredjeländer från vilka medlemsstaterna får tillåta import av köttprodukter och fastställer behandlingar som anses effektiva när det gäller att göra patogener för vissa djursjukdomar inaktiva. För att man skall förhindra risk för sjukdomsspridning via sådana produkter måste produkterna genomgå lämplig behandling beroende på hälsoläget i ursprungslandet och beroende på vilken art produkten härrör från. Import av köttprodukter och köttberedningar som består av eller innehåller kött av ratiter med ursprung i Sydafrika vilka genomgått lämplig behandling enligt det beslutet bör därför även fortsättningsvis vara tillåten.
(9) Så snart Sydafrika har inkommit med ytterligare information om sjukdomssituationen i fråga om högpatogen aviär influensa och de bekämpningsåtgärder som vidtagits mot sjukdomen, bör de åtgärder som vidtagits på gemenskapsnivå till följd av det nyligen inträffade utbrottet i Sydafrika ses över. Detta beslut bör därför endast gälla till och med den 31 oktober 2006.
(10) De åtgärder som föreskrivs i detta beslut är förenliga med yttrandet från ständiga kommittén för livsmedelskedjan och djurhälsa.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Medlemsstaterna skall tillfälligt upphäva importen från den del av Sydafrikas territorium som anges i bilagan till detta beslut av följande:
a) levande ratiter och kläckägg från ratiter,
b) färskt kött av ratiter, och
c) köttberedningar och köttprodukter som består av eller innehåller kött av ratiter.
Artikel 2
1. Genom undantag från artikel 1.b och 1.c skall medlemsstaterna tillåta import av färskt kött, köttprodukter och köttberedningar som avses i dessa punkter om de härrör från fåglar som har slaktats före den 1 maj 2006.
2. I de veterinärintyg som åtföljer sändningar av det kött och de köttprodukter och köttberedningar som avses i punkt 1 skall följande omnämnande ingå:
%quot%Färskt kött av ratiter/köttprodukter som består av eller innehåller kött av ratiter/köttberedningar som består av eller innehåller kött av ratiter [4] från fåglar som slaktats före den 1 maj 2006 i enlighet med artikel 2.1 i kommissionens beslut 2006/532/EC.
3. Genom undantag från artikel 1 c skall medlemsstaterna tillåta import av köttprodukter och köttberedningar som består av eller innehåller kött av ratiter förutsatt att köttet har genomgått minst en av de särskilda behandlingar som fastställs i B, C eller D i del 4 i bilaga II till beslut 2005/432/EG.
Artikel 3
Medlemsstaterna skall genast vidta de åtgärder som är nödvändiga för att följa detta beslut och offentliggöra dessa åtgärder. De skall genast underrätta kommissionen om detta.
Artikel 4
Detta beslut skall tillämpas till och med den 31 oktober 2006.
Artikel 5
Detta beslut riktar sig till medlemsstaterna.
Rådets beslut
av den 24 juli 2006
om fastställande av datum för tillämpningen av artikel 1.4 och 1.5 i förordning (EG) nr 871/2004 om införande av ett antal nya funktioner för Schengens informationssystem bland annat i kampen mot terrorism
(2006/628/EG)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av rådets förordning (EG) nr 871/2004 av den 29 april 2004 om införande av ett antal nya funktioner för Schengens informationssystem bland annat i kampen mot terrorism [1], särskilt artikel 2.2, och
av följande skäl:
(1) I artikel 2.2 i förordning (EG) nr 871/2004 anges det att förordningen skall tillämpas från och med ett datum som rådet skall fastställa så snart de nödvändiga förutsättningarna har uppfyllts och att rådet får besluta att fastställa olika tidpunkter för tillämpningen av olika bestämmelser.
(2) De förutsättningar som avses i artikel 2.2 i förordning (EG) nr 871/2004 har uppfyllts i fråga om artikel 1.4 och 1.5.
(3) När det gäller Schweiz utgör detta beslut, i enlighet med avtalet mellan Europeiska unionen, Europeiska gemenskapen och Schweiziska edsförbundet om Schweiziska edsförbundets associering till genomförandet, tillämpningen och utvecklingen av Schengenregelverket, en utveckling av de bestämmelser i Schengenregelverket vilka omfattas av det område som avses i artikel 1 G i rådets beslut 1999/437/EG av den 17 maj 1999 om vissa tillämpningsföreskrifter för det avtal som har ingåtts mellan Europeiska unionens råd och Republiken Island och Konungariket Norge om dessa båda staters associering till genomförandet, tillämpningen och utvecklingen a
Kommissionens förordning (EG) nr 94/2006
av den 19 januari 2006
om fastställande av exportbidrag för sirap och vissa andra sockerprodukter i obearbetat skick
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1260/2001 av den 19 juni 2001 om den gemensamma organisationen av marknaden för socker [1], särskilt artikel 27.5 andra stycket i denna, och
av följande skäl:
(1) I enlighet med artikel 27 i förordning (EG) nr 1260/2001 kan skillnaderna mellan kurserna eller priserna på världsmarknaden för de produkter som avses i artikel 1.1 d i nämnda förordning och priserna på dessa produkter inom gemenskapen, täckas av ett exportbidrag.
(2) I enlighet med artikel 3 i kommissionens förordning (EG) nr 2135/95 av den 7 september 1995 om tillämpningsföreskrifter för beviljande av exportbidrag vid sockerexport [2], skall bidraget för 100 kg av de produkter som avses i artikel 1.1 d i förordning (EG) nr 1260/2001 i samband med export vara lika med basbeloppet multiplicerat med sackarosinnehållet, i tillämpliga fall inklusive halten av andra sockerarter omräknade till sackaros. Den sackaroshalt som konstateras för produkten i fråga fastställs i enlighet med bestämmelserna i artikel 3 i kommissionens förordning (EG) nr 2135/95.
(3) I enlighet med artikel 30.3 i förordning (EG) nr 1260/2001 skall basbeloppet för bidrag för sorbos i obearbetat skick vara lika med basbeloppet för bidraget minskat med en hundradel av produktionsbidraget i enlighet med kommissionens förordning (EG) nr 1265/2001 av den 27 juni 2001 om tillämpningsföreskrifter för rådets förordning (EG) nr 1260/2001 när det gäller beviljande av produktionsbidrag för vissa sockerprodukter som används inom den kemiska industrin [3], när det gäller de produkter som avses i bilagan till den sistnämnda förordningen.
(4) I enlighet med artikel 30.1 i förordning (EG) nr 1260/2001 skall basbeloppet för bidraget för de övriga produkter som avses i artikel 1.1 d i denna förordning vid export i obearbetat skick vara lika med hundradelen av ett belopp som fastställs med hänsyn till skillnaden mellan interventionspriset för vitsocker inom områden inom gemenskapen utan underskott, under den månad för vilken basbeloppet fastställs och de kurser eller priser på vitsocker som noteras på världsmarknaden och behovet av att åstadkomma en balans mellan användningen av gemenskapens basprodukter vid export till tredje land av förädlingsprodukter och användningen av produkter importerade från dessa länder i förädlingssyfte.
(5) I enlighet med artikel 30.4 i förordning (EG) nr 1260/2001 kan tillämpningen av basbeloppet begränsas till vissa av de produkter som avses i artikel 1.1 d i denna förordning.
(6) I enlighet med artikel 27 i förordning (EG) nr 1260/2001 får exportbidrag ges för de produkter som avses i artikel 1.1 f, 1.1 g och 1.1 h i den förordningen. Bidragets storlek skall fastställas per 100 kg torrvara med beaktande, framför allt, av de bidrag som gäller vid export av de produkter som omfattas av KN-nummer 17023091, det bidrag som är tillämpligt vid export av de produkter som avses i artikel 1.1 d i förordning (EG) nr 1260/2001 och de ekonomiska aspekter som gäller för denna export. För de produkter som avses i artikel 1.1 f och 1.1 g skall bidrag beviljas endast för de produkter som uppfyller de villkor som fastställs i artikel 5 i förordning (EG) nr 2135/95. För de produkter som avses i 1.1 h skall bidrag beviljas endast för de produkter som uppfyller villkoren i artikel 6 i förordning (EG) nr 2135/95.
(7) De exportbidrag som avses ovan måste fastställas varje månad. De kan ändras däremellan.
(8) Enligt artikel 27.5 första stycket i förordning (EG) nr 1260/2001 kan världsmarknadssituationen eller särskilda krav på vissa marknader göra det nödvändigt att differentiera bidraget för de produkter som avses i artikel 1 i den förordningen, beroende på produkternas destination.
(9) Den avsevärda och snabba ökningen av å ena sidan förmånsimport av socker från länderna på västra Balkan sedan början av år 2001 och å andra sidan av sockerexporten från gemenskapen till dessa länder tycks vara synnerligen konstlad.
(10) För att undvika missbruk i form av återimport till Europeiska unionen av sockerprodukter för vilka det beviljats exportbidrag bör det inte finnas något bidrag för de produkter som avses i den här förordningen när det gäller länderna på västra Balkan.
(11) Med hänsyn till detta bör exportbidragen för de ifrågavarande produkterna uppgå till de belopp som anses lämpliga.
(12) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för socker.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De exportbidrag som skall beviljas vid export i oarbetat skick av de produkter som avses i artikel 1.1 d, 1.1 f, 1.1 g och 1.1 h i förordning (EG) nr 1260/2001 skall fastställas i enlighet med bilagan til den här förordning.
Artikel 2
Denna förordning träder i kraft den 20 januari 2006.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 412/2006
av den 9 mars 2006
om de anbud som meddelats för export av vanligt vete inom ramen för den anbudsinfordran som avses i förordning (EG) nr 1059/2005
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1784/2003 av den 29 september 2003 om den gemensamma organisationen av marknaden för spannmål [1], särskilt artikel 13.3 första stycket i denna, och
av följande skäl:
(1) En anbudsinfordran för bidrag för export av vanligt vete till vissa tredjeländer har inletts genom kommissionens förordning (EG) nr 1059/2005 [2].
(2) I enlighet med artikel 7 i kommissionens förordning (EG) nr 1501/95 av den 29 juni 1995 om vissa tillämpningsföreskrifter för rådets förordning (EEG) nr 1766/92 vad avser beviljande av exportbidrag och de åtgärder som skall vidtas vid störningar inom spannmålssektorn [3] kan kommissionen besluta att inte fullfölja anbudsinfordran.
(3) Särskilt med hänsyn till de kriterier som avses i artikel 1 i förordning (EG) nr 1501/95 är det inte uppenbart att ett högsta exportbidrag skall fastställas.
(4) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från Förvaltningskommittén för spannmål.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De anbud som meddelats från den 3 till den 9 mars 2006 inom ramen för den anbudsinfordran för exportbidrag för vanligt vete som avses i förordning (EG) nr 1059/2005 skall inte fullföljas.
Artikel 2
Denna förordning träder i kraft den 10 mars 2006.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 691/2006
av den 4 maj 2006
om de anbud som meddelats för export av korn inom ramen för den anbudsinfordran som avses i förordning (EG) nr 1058/2005
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1784/2003 av den 29 september 2003 om den gemensamma organisationen av marknaden för spannmål [1], särskilt artikel 13.3 första stycket, och
av följande skäl:
(1) En anbudsinfordran för bidrag för export av korn till vissa tredje länder har inletts genom kommissionens förordning (EG) nr 1058/2005 [2].
(2) I enlighet med artikel 7 i kommissionens förordning (EG) nr 1501/95 [3] av den 29 juni 1995 om vissa tillämpningsföreskrifter för rådets förordning (EEG) nr 1766/92 vad avser beviljande av exportbidrag och de åtgärder som skall vidtas vid störningar inom spannmålssektorn kan kommissionen besluta att inte fullfölja anbudsinfordran.
(3) Särskilt med hänsyn till de kriterier som avses i artikel 1 i förordning (EG) nr 1501/95 är det inte uppenbart att ett högsta exportbidrag skall fastställas.
(4) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från förvaltningskommittén för spannmål.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De anbud som meddelats från den 28 april– 4 maj 2006 inom ramen för den anbudsinfordran för exportbidrag för korn som avses i förordning (EG) nr 1058/2005 skall inte fullföljas.
Artikel 2
Denna förordning träder i kraft den 5 maj 2006.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 800/2006
av den 30 maj 2006
om öppnande och förvaltning av en tullkvot för import av unga handjur av nötkreatur avsedda för gödning ( 1 juli 2006– 30 juni 2007)
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1254/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för nötkött [1], särskilt artikel 32.1, och
av följande skäl:
(1) Enligt Världshandelsorganisationens lista CXL skall gemenskapen öppna en årlig tullkvot för import av 169000 unga handjur av nötkreatur avsedda för gödning. Till följd av de förhandlingar som ledde till avtalet i form av skriftväxling mellan Europeiska gemenskapen och Amerikas Förenta stater i enlighet med artikel XXIV:6 och artikel XXVIII i Allmänna tull- och handelsavtalet (GATT) 1994 [2], godkänt genom rådets beslut 2006/333/EG [3], åtog sig dock gemenskapen att i sin bindningslista för samtliga medlemsstater justera den importtullkvoten.
(2) I bestämmelserna för förvaltningen av denna tullkvot bör det för perioden 1 juli 2006– 30 juni 2007 fastställas att den tillgängliga kvoten bör fördelas över året på ett lämpligt sätt i den mening som avses i artikel 32.4 i förordning (EG) nr 1254/1999.
(3) Mot bakgrund av att fördraget om Bulgariens och Rumäniens anslutning till Europeiska unionen kommer att träda i kraft, och utan att det påverkar tillämpningen av artikel 39 i det fördraget, bör kvotperioden delas in i två delperioder och den kvantitet som finns tillgänglig inom kvoten fördelas mellan dessa perioder med hänsyn till den traditionella handeln mellan gemenskapen och leverantörsländerna inom ramen för den här kvoten. Syftet med detta är att se till att aktörer från dessa länder kan utnyttja kvoten från och med anslutningsdagen.
(4) För att man skall kunna sörja både för en jämnare fördelning av kvoten och ett ekonomiskt lönsamt antal djur per ansökan, bör en nedre och en övre gräns för antalet djur gälla för varje ansökan om importlicenser.
(5) För att undvika spekulation bör de tillgängliga kvantiteterna inom kvoten ställas till sådana aktörers förfogande som kan visa att de bedriver en seriös importverksamhet av betydande omfattning med tredjeländer. Med tanke på detta och för att säkerställa en effektiv förvaltning bör det krävas av de berörda aktörerna att de importerat minst 50 djur under perioden 1 maj 2005– 30 april 2006, eftersom ett parti på 50 djur kan betraktas som en ekonomiskt lönsam sändning.
(6) För att dessa kriterier skall kunna kontrolleras krävs att ansökan lämnas in i den medlemsstat där importören är upptagen i ett register för mervärdesskatt.
(7) För att undvika spekulation bör importörer som den 1 januari 2006 inte längre bedrev handel med levande nötkreatur nekas tillgång till kvoten, och licenserna bör inte kunna överlåtas.
(8) De kvantiteter för vilka ansökan om importlicens kan lämnas in bör tilldelas efter en viss betänketid och eventuellt med tillämpning av en enhetlig tilldelningskoefficient.
(9) Det bör föreskrivas att systemet skall förvaltas med hjälp av importlicenser. Det bör för detta ändamål införas närmare bestämmelser om inlämnande av ansökningar och om de uppgifter som skall lämnas i ansökningar och licenser, i förekommande fall genom tillägg till eller undantag från relevanta bestämmelser i kommissionens förordning (EG) nr 1445/95 av den 26 juni 1995 om tillämpningsföreskrifter för ordningen med import- och exportlicenser inom nötköttssektorn och om upphävande av förordning (EEG) nr 2377/80 [4] och i kommissionens förordning (EG) nr 1291/2000 av den 9 juni 2000 om gemensamma tillämpningsföreskrifter för systemet med import- och exportlicenser samt förutfastställelselicenser för jordbruksprodukter [5].
(10) Erfarenheten har visat att det för en korrekt förvaltning av kvoten också krävs att licensinnehavaren verkligen är importör. En importör bör därför aktivt delta i uppköp, transport och import av djuren i fråga. Uppvisande av handlingar som styrker sådan verksamhet bör därför också vara ett primärt krav när det gäller den säkerhet som skall ställas för licensen i den mening som avses i kommissionens förordning (EEG) nr 2220/85 av den 22 juli 1985 om gemensamma tillämpningsföreskrifter för systemet med säkerheter för jordbruksprodukter [6].
(11) För att garantera en strikt statistisk kontroll av de djur som importeras inom kvoten bör den tolerans som avses i artikel 8.4 i förordning (EG) nr 1291/2000 inte tillämpas.
(12) För tillämpningen av denna tullkvot krävs effektiva kontroller beträffande bestämmelseorten för de importerade djuren i varje enskilt fall. Gödningen bör därför ske i den medlemsstat som har utfärdat importlicensen.
(13) En säkerhet bör ställas som garanti för att djuren göds under minst 120 dagar på de anläggningar som utsetts. Säkerheten bör täcka skillnaden mellan tullarna i Gemensamma tulltaxan och de lägre tullar som tas ut den dag då djuren i fråga övergår till fri omsättning.
(14) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från förvaltningskommittén för nötkött.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. En tullkvot omfattande 24070 unga handjur av nötkreatur med KN-nummer 01029005, 01029029 eller 01029049 avsedda för gödning inom gemenskapen, öppnas härmed för perioden 1 juli 2006– 30 juni 2007.
Löpnumret för denna kvot skall vara 09.4005.
2. För den kvot som avses i punkt 1 skall importtullen uppgå till en värdetull på 16 % plus 582 euro per ton netto.
Tillämpningen av den tullsats som föreskrivs i första stycket förutsätter att gödningen av de importerade djuren har ägt rum under minst 120 dagar i den medlemsstat som utfärdat importlicensen.
3. De kvantiteter som avses i punkt 1 skall fördelas enligt följande:
a) 12035 levande nötkreatur under perioden 1 juli 2006– 31 december 2006.
b) 12035 levande nötkreatur under perioden 1 januari 2007– 30 juni 2007.
4. Om den kvantitet som omfattas av licensansökningar under den period som nämns i punkt 3 a är mindre än den kvantitet som finns tillgänglig för den perioden skall den återstående kvantiteten för den perioden läggas till den tillgängliga kvantiteten för den period som nämns i punkt 3 b.
Artikel 2
1. För att få ta del av den kvot som avses i artikel 1 krävs det att de sökande är fysiska eller juridiska personer som vid ansökningstillfället på ett för de behöriga myndigheterna i den berörda medlemsstaten tillfredsställande sätt kan styrka att de under perioden 1 maj 2005– 30 april 2006 har importerat minst 50 djur med KN-nummer 010290.
Förutsatt att fördraget om Bulgariens och Rumäniens anslutning till Europeiska unionen träder i kraft den 1 januari 2007 får aktörerna i dessa länder ansöka om importlicenser inom ramen för den kvantitet som finns tillgänglig för den andra delperioden för den här kvoten enligt artikel 1.3 b, om de har importerat minst 50 djur med KN-nummer 010290 under perioden 1 maj 2005– 30 april 2006.
De sökande skall vara införda i ett nationellt register för mervärdesskatt.
2. Import skall styrkas uteslutande med hjälp av ett tulldokument om övergång till fri omsättning, som attesterats av tullmyndigheterna och i vilket sökanden i fråga uppges som mottagare.
Medlemsstaterna får godta kopior av det dokument som avses i första stycket, om dessa styrkts av den behöriga myndigheten. Om en sådan kopia godtas, skall medlemsstaten för varje berörd sökande anmäla detta i det meddelande som avses i artikel 3.5.
3. Aktörer som den 1 januari 2006 hade upphört med sin handelsverksamhet med tredjeländer inom nötköttssektorn får inte ansöka om licens.
4. Ett företag som bildats genom fusion av företag som vart för sig hade en referensimport på minst den mängd som anges i punkt 1 får lägga dessa referensimporter till grund för sin ansökan.
Artikel 3
1. Ansökan om importlicenser får endast lämnas in i den medlemsstat där den sökande är upptagen i ett nationellt register för mervärdesskatt.
2. Ansökan om importlicens för var och en av perioderna enligt artikel 1.3
a) skall avse minst 50 djur,
b) får avse högst 5 % av den tillgängliga kvantiteten.
Om ansökan avser en större kvantitet än den som anges i första stycket led b, skall den överskjutande kvantiteten inte beaktas.
3. Ansökningar om importlicenser för den period som avses i artikel 1.3 a skall lämnas in under de tio arbetsdagarna efter offentliggörandet av denna förordning i Europeiska unionens officiella tidning.
Ansökningar om importlicenser för den period som avses i artikel 1.3 b skall lämnas in under de första tio arbetsdagarna i den perioden.
4. En sökande får endast lämna in en ansökan för var och en av de perioder som nämns i artikel 1.3. Om samma sökande lämnar in fler än en ansökan, skall ingen av dessa ansökningar behandlas.
5. Efter en kontroll av dokumenten skall medlemsstaterna, senast den femte arbetsdagen efter det att perioden för inlämnande av ansökningar löpt ut, till kommissionen lämna en förteckning över de sökande med adressuppgifter samt uppgift om de kvantiteter som de ansökt om.
Alla meddelanden, även om att ingen ansökan har lämnats in, skall skickas per fax eller e-post, i förekommande fall med användning av förlagan i bilaga I.
Artikel 4
1. Efter anmälan enligt artikel 3.5 skall kommissionen snarast möjligt besluta i vilken utsträckning ansökningarna kan tillgodoses.
2. Om kvantiteten i licensansökningarna enligt artikel 3 överstiger de kvantiteter som finns tillgängliga för perioden i fråga, skall kommissionen fastställa en enhetlig koefficient för tilldelning som skall tillämpas på de begärda kvantiteterna.
Om den tilldelningskoefficient som avses i första stycket resulterar i en kvantitet på mindre än 50 djur per ansökan, skall importrättigheter för partier på 50 djur fördelas av de berörda medlemsstaterna genom lottdragning. Om den återstående kvantiteten är mindre än 50 djur, skall den anses utgöra ett enda parti.
3. Om kommissionen beslutar att ansökningarna kan godtas, skall licenserna utfärdas så snart som möjligt.
Artikel 5
1. Importlicenserna skall utfärdas i den ansökande aktörens namn.
2. Licensansökan och licensen skall innehålla följande uppgifter:
a) I fält 8, ursprungslandet.
b) I fält 16, ett eller flera av följande KN-nummer: 01029005, 01029029 eller 01029049;
c) I fält 20, kvotens löpnummer (09.4005) och en av de uppgifter som anges i bilaga II.
Artikel 6
1. Genom avvikelse från artikel 9.1 i förordning (EG) nr 1291/2000 får importlicenser som har utfärdats i enlighet med den här förordningen inte överlåtas, och de skall ge tillgång till tullkvoten endast om de är utfärdade med samma namn- och adressuppgifter som dem som uppges för mottagaren i de tulldeklarationer om övergång till fri omsättning som åtföljer dem.
2. Genom avvikelse från artikel 3 i förordning (EG) nr 1445/95 skall importlicenser gälla under 180 dagar från och med utfärdandet i enlighet med artikel 4.3 i föreliggande förordning. Inga licenser skall gälla efter den 30 juni 2007.
3. Säkerheten för importlicensen skall vara 15 euro per djur och skall ställas av den sökande tillsammans med licensansökan.
4. De utfärdade licenserna skall vara giltiga i hela gemenskapen.
5. Enligt artikel 50.1 i förordning (EG) nr 1291/2000 skall hela den tull enligt Gemensamma tulltaxan som tillämpas den dag då tulldeklarationen om övergång till fri omsättning godkänns tas ut på alla kvantiteter som importeras utöver de kvantiteter som anges i importlicensen.
6. Genom avvikelse från bestämmelserna i avdelning III avsnitt 4 i förordning (EG) nr 1291/2000 får säkerheten inte frisläppas förrän handlingar har uppvisats som styrker att licensinnehavaren har varit kommersiellt och logistiskt ansvarig för inköp, transport och klarering för fri omsättning av de berörda djuren. Dessa handlingar skall minst omfatta följande:
a) Handelsfakturan i original eller en bestyrkt kopia utfärdad i licensinnehavarens namn av säljaren eller dennes företrädare, vilka båda skall vara etablerade i det exporterande tredjelandet, samt licensinnehavarens betalningsbevis eller bevis för att licensinnehavaren har öppnat en ouppsägbar remburs till förmån för säljaren.
b) Konossement eller i tillämpliga fall väg- eller lufttransportdokument, utfärdat i licensinnehavarens namn för de berörda djuren.
c) Handling som styrker att varorna har deklarerats för övergång till fri omsättning med uppgift om licensinnehavarens namn och adress och att denna är mottagare.
Artikel 7
1. Vid importtillfället skall importören styrka
a) att han har undertecknat ett skriftligt åtagande att inom en månad underrätta den behöriga myndigheten i medlemsstaten om vid vilken eller vilka anläggningar de unga nötkreaturen skall gödas,
b) att han har ställt en säkerhet på det belopp som fastställs för varje godkänt KN-nummer i bilaga III hos den behöriga myndigheten i medlemsstaten. Det skall vara ett primärt krav i den mening som avses i artikel 20.2 i förordning (EEG) nr 2220/85 att gödningen av de importerade djuren sker i den medlemsstaten under minst 120 dagar räknat från och med den dag då tulldeklarationen om övergång till fri omsättning godkändes.
2. Utom vid force majeure skall den säkerhet som avses i punkt 1 b inte frisläppas förrän de behöriga myndigheterna i medlemsstaten har erhållit handlingar som styrker att djuren
a) har götts i den anläggning eller de anläggningar som anges i punkt 1,
b) inte har slaktats inom 120 dagar räknat från importdagen, eller
c) före utgången av denna tid har slaktats av hälsoskäl, eller har dött till följd av sjukdom eller olyckshändelse.
Säkerheten skall frisläppas omedelbart efter det att sådana handlingar har framlagts.
Om tidsfristen enligt punkt 1 a inte har iakttagits, skall emellertid det säkerhetsbelopp som skall frisläppas minskas med
- 15 %, och med
- 2 % av det återstående beloppet för varje dags överskridande.
De belopp som inte frisläpps skall anses vara förverkade och skall behållas som tull.
3. Om de handlingar som avses i punkt 2 inte framläggs inom 180 dagar från importdagen, skall säkerheten anses vara förverkad och behållas som tull.
Om sådana handlingar inte har framlagts inom den period på 180 dagar som föreskrivs i första stycket men framläggs inom sex månader efter dessa 180 dagar, skall det förverkade beloppet återbetalas, minskat med 15 % av säkerheten.
Artikel 8
Förordningarna (EG) nr 1291/2000 och (EG) nr 1445/95 skall tillämpas, om inte annat följer av den här förordningen.
Artikel 9
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 832/2006
av den 2 juni 2006
om fördelningen mellan %quot%leveranser%quot% och %quot%direktförsäljning%quot% av de nationella referenskvantiteter som fastställts för 2005/2006 i bilaga I till rådets förordning (EG) nr 1788/2003
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1788/2003 av den 29 september 2003 om införande av en avgift inom sektorn för mjölk och mjölkprodukter [1], särskilt artikel 6.4 och artikel 8, och
av följande skäl:
(1) I artikel 6 i förordning (EG) nr 1788/2003 föreskrivs att medlemsstaterna skall fastställa individuella referenskvantiteter för producenterna. En producent kan ha antingen en eller två individuella referenskvantiteter, en för leverans och en för direktförsäljning, och omställningen mellan en producents referenskvantiteter kan göras på vederbörligen motiverad begäran från producenten.
(2) I kommissionens förordning (EG) nr 490/2005 av den 29 mars 2005 om fördelningen mellan %quot%leveranser%quot% och %quot%direktförsäljning%quot% av de nationella referenskvantiteter som fastställts för 2004/2005 i bilaga I till rådets förordning (EG) nr 1788/2003 [2] fastställs fördelningen mellan %quot%leveranser%quot% och %quot%direktförsäljning%quot% för perioden 1 april 2004– 31 mars 2005 för Belgien, Tjeckien, Danmark, Tyskland, Estland, Grekland, Spanien, Frankrike, Irland, Italien, Cypern, Lettland, Litauen, Luxemburg, Ungern, Malta, Nederländerna, Österrike, Portugal, Slovakien, Finland, Sverige och Förenade kungariket.
(3) För Polen och Slovenien fastställs grunden för de individuella referenskvantiteterna i tabell f i bilaga I till förordning (EG) nr 1788/2003.
(4) I enlighet med artikel 25.2 i kommissionens förordning (EG) nr 595/2004 av den 30 mars 2004 om tillämpningsföreskrifter för rådets förordning (EG) nr 1788/2003 om införande av en avgift inom sektorn för mjölk och mjölkprodukter [3] har Belgien, Tjeckien, Danmark, Tyskland, Estland, Grekland, Spanien, Frankrike, Irland, Italien, Cypern, Lettland, Litauen, Ungern, Nederländerna, Österrike, Polen, Portugal, Slovenien, Slovakien, Finland och Förenade kungariket anmält hur stora kvantiteter som på producenternas begäran har ställts om definitivt mellan individuella referenskvantiteter för leveranser och direktförsäljning.
(5) I artikel 6.4 i förordning (EG) nr 1788/2003 fastställs att den del av den finländska nationella referenskvantitet som är avdelad för sådana leveranser som avses i artikel 1 i den förordningen kan ökas upp till högst 200000 ton som kompensation till de finländska Slom-producenterna. I enlighet med artikel 6 i kommissionens förordning (EG) nr 671/95 av den 29 mars 1995 om tilldelning av en särskild referenskvantitet till vissa producenter av mjölk och mjölkprodukter i Österrike och Finland [4], har Finland meddelat kvantiteterna för regleringsåret 2005/2006.
(6) Det är därför lämpligt att fastställa fördelningen mellan %quot%leveranser%quot% och %quot%direktförsäljning%quot% av de nationella referenskvantiteterna för perioden 1 april 2005– 31 mars 2006 som fastställts i bilaga I till förordning (EG) nr 1788/2003.
(7) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från förvaltningskommittén för mjölk och mjölkprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Fördelningen mellan %quot%leveranser%quot% och %quot%direktförsäljning%quot% av de nationella referenskvantiteter för perioden 1 april 2005– 31 mars 2006 som fastställts i bilaga I till förordning (EG) nr 1788/2003 anges i bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 877/2006
av den 15 juni 2006
om fastställande av det högsta exportbidraget för smör inom ramen för den stående anbudsinfordran som fastställs i förordning (EG) nr 581/2004
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1255/1999 av den 17 maj 1999 om den gemensamma organisationen av marknaden för mjölk och mjölkprodukter [1], särskilt artikel 31.3 tredje stycket och
av följande skäl:
(1) I kommissionens förordning (EG) nr 581/2004 av den 26 mars 2004 om inledande av en stående anbudsinfordran för exportbidrag för vissa typer av smör [2] fastställs bestämmelser för en stående anbudsinfordran.
(2) Enligt artikel 5 i kommissionens förordning (EG) nr 580/2004 av den 26 mars 2004 om fastställande av ett anbudsförfarande för exportbidrag för vissa mjölkprodukter [3] och en granskning av de anbud som inlämnats inom ramen för anbudsförfarandet är det lämpligt att fastställa ett högsta exportbidrag för den anbudsperiod som löper ut den 13 juni 2006.
(3) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från förvaltningskommittén för mjölk och mjölkprodukter.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
För den stående anbudsinfordran som inleddes genom förordning (EG) nr 581/2004 för den anbudsperiod som löper ut den 13 juni 2006 skall det högsta bidragsbeloppet för de produkter som avses i artikel 1.1 i den förordningen vara det som anges i bilagan till den här förordningen.
Artikel 2
Denna förordning träder i kraft den 16 juni 2006.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1108/2006
av den 19 juli 2006
om fastställande av schablonvärden vid import för bestämning av ingångspriset för vissa frukter och grönsaker
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av kommissionens förordning (EG) nr 3223/94 av den 21 december 1994 om tillämpningsföreskrifter för importordningen för frukt och grönsaker [1], särskilt artikel 4.1, och
av följande skäl:
(1) I förordning (EG) nr 3223/94 anges som tillämpning av resultaten av de multilaterala förhandlingarna i Uruguayrundan kriterierna för kommissionens fastställande av schablonvärdena vid import från tredje land för de produkter och de perioder som anges i bilagan till den förordningen.
(2) Vid tillämpningen av dessa kriterier bör schablonvärdena vid import fastställas till de nivåer som anges i bilagan till denna förordning.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
De schablonvärden vid import som avses i artikel 4 i förordning (EG) nr 3223/94 skall fastställas enligt tabellen i bilagan.
Artikel 2
Denna förordning träder i kraft den 20 juli 2006.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1191/2006
av den 4 augusti 2006
om ändring av förordning (EG) nr 1458/2003 om öppnande och förvaltning av tullkvoter för griskött
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EEG) nr 2759/75 av den 29 oktober 1975 om den gemensamma organisationen av marknaden för griskött [1], särskilt artiklarna 8.2 och 11.1, och
av följande skäl:
(1) Förordning (EG) nr 1458/2003 [2] avser öppnande och förvaltning av tullkvoter för griskött.
(2) I det avtal genom skriftväxling mellan Europeiska gemenskapen och Amerikas förenta stater enligt artikel XXIV:6 och artikel XXVIII i Allmänna tull- och handelsavtalet (GATT) 1994 [3], som godkänns genom rådets beslut 2006/333/EG [4], föreskrivs en ökning av den årliga importtullkvoten för griskött med 1430 ton griskött.
(3) Den hänvisning som måste göras i ansökningar om importlicens bör göras på gemenskapens samtliga officiella språk.
(4) Med tanken på Bulgariens och Rumäniens eventuella anslutning till Europeiska unionen den 1 januari 2007 bör det föreskrivas en särskild ansökningsperiod för importlicenser under första kvartalet 2007.
(5) Förordning (EG) nr 1458/2003 bör ändras i enlighet med detta.
(6) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från förvaltningskommittén för griskött.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EG) nr 1458/2003 skall ändras på följande sätt:
1. I artikel 4 skall leden d och e ersättas med följande:
%quot%d) I fält 20 i ansökningarna och i licenserna skall en av de texter som förtecknas i bilaga Ia anges.
e) I fält 24 i licenserna skall en av de texter som förtecknas i bilaga Ib anges.%quot%
2. I artikel 5.1 skall följande stycke läggas till:
%quot%Avseende perioden 1 januari– 31 mars 2007 får licensansökningarna emellertid lämnas in under de första femton dagarna i januari 2007.%quot%
3. Bilagorna I–IV skall ersättas med bilagorna till denna förordning.
Artikel 2
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska unionens officiella tidning.
Den skall tillämpas från och med den 1 juli 2006.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1238/2006
av den 16 augusti 2006
om fastställande av en enhetlig tilldelningskoefficient som skall tillämpas på tullkvoten för vete i enlighet med förordning (EG) nr 573/2003
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1784/2003 av den 29 september 2003 om den gemensamma organisationen av marknaden för spannmål [1],
med beaktande av kommissionens förordning (EG) nr 573/2003 av den 28 mars 2003 om tillämpningsföreskrifter för rådets beslut 2003/18/EG beträffande medgivanden i form av gemenskapstullkvoter för vissa spannmålsprodukter med ursprung i Rumänien och om ändring av förordning (EG) nr 2809/2000 [2], särskilt artikel 2.3, och
av följande skäl:
(1) Genom förordning (EG) nr 573/2003 öppnas en årlig tullkvot på 230000 ton vete (löpnummer 09.4766) för regleringsåret 2006/2007.
(2) De kvantiteter som begärdes måndagen den 14 augusti 2006, i enlighet med artikel 2.1 i förordning (EG) nr 573/2003, överskrider de kvantiteter som finns tillgängliga. Det bör därför beslutas i vilken omfattning licenser skall utfärdas. Det bör ske genom fastställande av en enhetlig tilldelningskoefficient som skall tillämpas på de begärda kvantiteterna.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Samtliga ansökningar om importlicens för tullkvoten för vete från Rumänien som, i enlighet med artikel 2.1 och 2.2 i förordning (EG) nr 573/2003, lämnades in och vidarebefordrades till kommissionen måndagen den 14 augusti 2006, skall godkännas för 1,744760634 % av de begärda kvantiteterna.
Artikel 2
Denna förordning träder i kraft den 17 augusti 2006.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1601/2006
av den 26 oktober 2006
om utfärdande av importlicenser för ris avseende de ansökningar som lämnats in under de tio första arbetsdagarna i oktober 2006 i enlighet med förordning (EG) nr 327/98
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1785/2003 av den 29 september 2003 om den gemensamma organisationen av marknaden för ris [1],
med beaktande av kommissionens förordning (EG) nr 327/98 av den 10 februari 1998 om öppnande och förvaltning av vissa tullkvoter för import av ris och brutet ris [2], särskilt artikel 5.2, och
av följande skäl:
Vid en genomgång av de kvantiteter för vilka ansökningar om importlicenser för ris lämnades in under ansökningsomgången för oktober 2006 framgick det dels att licenser bör utfärdas för de kvantiteter som ansökningarna gäller och som i tillämpliga fall omfattas av en nedsättningsprocentsats, dels att den slutliga utnyttjandeprocenten under 2006 bör meddelas för varje tullkvot.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. De ansökningar om importlicenser för de tullkvoter för ris som öppnas genom förordning (EG) nr 327/98, som lämnats in under de tio första arbetsdagarna i oktober 2006 och som meddelats kommissionen, skall omfattas av nedsättningskoefficienter i enlighet med bilagan till denna förordning.
2. I bilagan anges slutlig procentsats som gäller för 2006 för varje berörd kvot.
Artikel 2
Denna förordning träder i kraft den 27 oktober 2006.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1659/2006
av den 9 november 2006
om fastställande av exportbidrag för sirap och vissa andra sockerprodukter som exporteras i obearbetat skick
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 318/2006 av den 20 februari 2006 om den gemensamma organisationen av marknaden för socker [1], särskilt artikel 33.2 andra stycket, och
av följande skäl:
(1) I artikel 32 i förordning (EG) nr 318/2006 fastställs att skillnaden mellan priserna på världsmarknaden för de produkter som förtecknas i artikel 1.1 c, d och g i den förordningen och priserna för dessa produkter inom gemenskapen får täckas av ett exportbidrag.
(2) Med hänsyn till den situation som för närvarande råder på sockermarknaden bör exportbidrag fastställas i enlighet med bestämmelserna och vissa kriterier i artiklarna 32 och 33 i förordning (EG) nr 318/2006.
(3) Enligt artikel 33.2 första stycket i förordning (EG) nr 318/2006 kan världsmarknadssituationen eller de särskilda behoven på vissa marknader vara sådana att bidraget måste varieras beroende på destination.
(4) Bidrag bör endast beviljas för produkter som omfattas av den fria rörligheten för varor inom gemenskapen och som uppfyller kraven i kommissionens förordning (EG) nr 951/2006 av den 30 juni 2006 om tillämpningsföreskrifter till förordning (EG) nr 318/2006 för handel med tredjeländer i sockersektorn [2].
(5) Förhandlingarna inom ramen för Europaavtalen mellan Europeiska gemenskapen och Rumänien och Bulgarien syftar främst till att avreglera handeln med de produkter som omfattas av den gemensamma organisationen av den berörda marknaden. Exportbidragen för Rumänien och Bulgarien bör därför avskaffas.
(6) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från förvaltningskommittén för socker.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Exportbidrag enligt artikel 32 i förordning (EG) nr 318/2006 skall beviljas för de produkter och med de belopp som anges i bilagan till den här förordningen om inte annat följer av villkoren i punkt 2 i den här artikeln.
2. För att berättiga till bidrag enligt punkt 1 skall produkterna uppfylla tillämpliga krav i artiklarna 3 och 4 i förordning (EG) nr 951/2006.
Artikel 2
Denna förordning träder i kraft den 10 november 2006.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Kommissionens förordning (EG) nr 1850/2006
av den 14 december 2006
om närmare bestämmelser om certifiering av humle och humleprodukter
EUROPEISKA GEMENSKAPERNAS KOMMISSION HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen,
med beaktande av rådets förordning (EG) nr 1952/2005 av den 23 november 2005 om den gemensamma organisationen av marknaden för humle och om upphävande av förordningarna (EEG) nr 1696/71, (EEG) nr 1037/72, (EEG) nr 879/73 och (EEG) nr 1981/82 [1], särskilt artikel 17, och
av följande skäl:
(1) I artikel 4.1 i förordning (EG) nr 1952/2005 anges det att reglerna för certifiering skall tillämpas för de produkter som avses i artikel 1 i den förordningen och som skördats eller framställts inom gemenskapen.
(2) Närmare bestämmelser om certifiering av humle fastställs i rådets förordning (EEG) nr 1784/77 av den 19 juli 1977 om certifiering av humle [2] och kommissionens förordning (EEG) nr 890/78 av den 28 april 1978 om närmare bestämmelser om certifiering av humle [3]. Eftersom ytterligare ändringar skall göras är det för tydlighetens skull lämpligt att upphäva förordningarna (EEG) nr 1784/77 och (EEG) nr 890/78 och ersätta dem med en enda förordning.
(3) För att skapa ett i huvudsak enhetligt certifieringsförfarande i medlemsstaterna är det nödvändigt att precisera vilka produkter som kommer i fråga, hur hanteringen skall gå till och vilken information som skall ges i de dokument som åtföljer produkterna.
(4) Vissa produkter bör på grund av sin särskilda karaktär och användning undantas från certifieringsförfarandet.
(5) För att humlekottar skall kunna kontrolleras bör en beskrivning som undertecknats av producenten åtfölja humlekottar som görs tillgängliga för certifiering. Denna beskrivning bör innehålla upplysningar som gör det möjligt att identifiera humlet från den tidpunkt då det görs tillgängligt för certifiering till dess att certifikatet är utfärdat.
(6) Enligt artikel 4.2 i förordning (EG) nr 1952/2005 får certifikat utfärdas endast för produkter med de kvalitetsegenskaper som anges som minimikrav. Det bör därför fastställas att sådana minimikrav för avsättning skall gälla för humlekottar från det första handelsledet.
(7) När de kvalitetsegenskaper skall fastställas som humlet måste ha, bör vattenhalten och halten främmande beståndsdelar medräknas. Eftersom humle från gemenskapen är känt för att vara av hög kvalitet, bör nuvarande praxis inom handeln användas som utgångspunkt.
(8) Det bör överlåtas åt medlemsstaterna att besluta vilken metod som skall användas för att fastställa vattenhalten, förutsatt att de metoder som används leder till jämförbara resultat. Vid eventuella tvister bör en gemenskapsmetod användas.
(9) Det bör fastställas strikta regler för blandningar. Därför bör blandningar av humlekottar bara tillåtas om de består av certifierade produkter av samma sort, från samma skörd och från samma produktionsområde. Det bör också fastställas att blandningar skall göras under tillsyn och underkastas samma certifieringsförfarande som de produkter som ingår i blandningen.
(10) När det gäller tillverkning av pulver och extrakt är det, med hänsyn till användarnas krav, lämpligt att på vissa villkor tillåta blandningar av certifierat humle som inte är av samma sort och som kommer från olika produktionsområden.
(11) Humle som framställs av obehandlat certifierat humle får certifieras endast om framställningen sker i en sluten tillverkningsprocess.
(12) För att säkerställa att certifieringsreglerna följs när det gäller humleprodukter bör lämpliga bestämmelser om tillsyn fastställas.
(13) Om en humleprodukt omförpackas under officiell tillsyn utan bearbetning bör det efterföljande certifieringsförfarandet också förenklas.
(14) För att säkerställa att certifierade produkter kan identifieras, bör det fastställas att förpackningarna skall förses med de uppgifter som krävs för den officiella tillsynen och som information till köparna.
(15) För att användarna skall få exakta upplysningar om ursprung och egenskaper hos de produkter som avsätts, bör gemensamma bestämmelser fastställas om märkning av förpackningar och referensnummer på certifikaten.
(16) Med hänsyn till nuvarande handelspraxis inom vissa områden i gemenskapen bör det anges om humlet avsätts på marknaden med eller utan frö och det bör fastställas att detta skall framgå av certifikatet.
(17) Humle från försökssorter under utveckling kan identifieras genom en namn- eller nummeruppgift.
(18) Det bör ställas särskilda krav på produkter som undantas från certifieringsförfarandet så att det säkerställs dels att dessa produkter inte kan störa den normala avsättningen av certifierade produkter, dels att de är lämpliga för den avsedda användningen och bara används av avsedda mottagare.
(19) Medlemsstaterna bör certifiera produkter i enlighet med denna förordning genom behöriga organ som särskilt utsetts för detta. Förteckningarna över dessa organ bör sändas till kommissionen.
(20) Medlemsstaterna bör fastställa vilka områden som skall betraktas som produktionsområden för humle och sända denna förteckning till kommissionen.
(21) De åtgärder som föreskrivs i denna förordning är förenliga med yttrandet från förvaltningskommittén för humle.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
KAPITEL 1
ALLMÄNNA BESTÄMMELSER
Artikel 1
Syfte och tillämpningsområde
1. I denna förordning fastställs närmare bestämmelser om certifiering av humle och humleprodukter.
2. Denna förordning skall tillämpas på
a) produkter som avses i artikel 1 i förordning (EG) nr 1952/2005 och som har skördats inom gemenskapen,
b) produkter framställda av sådana produkter som avses i artikel 1 i nämnda förordning vilka antingen har skördats inom gemenskapen eller importerats från tredjeland i enlighet med artikel 9 i den förordningen.
3. Denna förordning skall inte tillämpas på
a) humle som skördats på arealer som tillhör ett bryggeri och som används av bryggeriet i obearbetat eller bearbetat skick,
b) produkter som härrör från humle och under avtal bearbetats för ett bryggeris räkning, under förutsättning att produkterna används av samma bryggeri,
c) humle och produkter som härrör från humle, i små förpackningar avsedda för försäljning till privatpersoner för eget bruk,
d) produkter som tillverkats av isomeriserade humleprodukter.
Artikel 20 skall dock tillämpas på de produkter som avses i a, b och c i den här punkten.
4. Utan att det påverkar tillämpningen av punkt 3 a får bara certifierat humle, certifierade humleprodukter som framställts av certifierat humle och humle som importerats från tredjeländer i enlighet med artikel 9 i förordning (EG) nr 1952/2005 användas vid tillverkning av produkter som framställs av humle.
Artikel 2
Definitioner
I denna förordning gäller följande definitioner:
a) obehandlat humle : humle som bara preliminärt har torkats och förpackats.
b) behandlat humle : humle som slutgiltigt har torkats och slutgiltigt förpackats.
c) humle med frö : humle som avsätts med ett fröinnehåll på mer än 2 % av vikten.
d) humle utan frö : humle som avsätts med ett fröinnehåll på högst 2 % av vikten.
e) försegling : förslutning av förpackningar under officiell tillsyn och på ett sådant sätt att förslutningen går sönder när den öppnas.
f) sluten tillverkningsprocess : process för behandling eller bearbetning av humle vilken genomförs under officiell tillsyn och på ett sådant sätt att varken humle eller bearbetade produkter kan tillsättas eller avlägsnas under processen. Den slutna tillverkningsprocessen inleds med öppnandet av den förseglade förpackningen med det humle eller de humleprodukter som skall behandlas eller bearbetas och avslutas med förseglingen av den förpackning som innehåller det bearbetade humlet eller humleprodukterna.
g) parti : ett antal förpackningar med humle eller humleprodukter som har samma egenskaper och som görs tillgängliga för certifiering samtidigt av en och samma enskilde producent eller producent i en sammanslutning eller av samma bearbetningsanläggning.
h) produktionsområden för humle : de områden för produktion som anges i den förteckning som upprättas av berörda medlemsstater.
i) koncentrerat humlepulver : produkt som erhålls genom lösningsmedels inverkan på den produkt som erhålls genom malning av humlet, innehållande alla naturliga beståndsdelar av humle.
j) behörig certifieringsmyndighet : myndighet eller organ som medlemsstaten har utsett för att genomföra certifieringen och godkänna och kontrollera certifieringscentraler.
k) märkning : etikettering och identifiering.
l) certifieringscentral : plats där certifieringen sker.
m) företrädare för en behörig certifieringsmyndighet : person som är anställd hos den behöriga certifieringsmyndigheten eller hos en tredje part och som har den behöriga certifieringsmyndighetens tillstånd att genomföra certifiering.
n) officiell tillsyn : den behöriga certifieringsmyndighetens eller dess företrädares övervakning av certifieringsverksamheten.
o) isomeriserad humleprodukt : humleprodukt i vilken alfasyrorna så gott som fullständigt isomeriserats.
KAPITEL 2
HUMLE
Artikel 3
Humle som görs tillgängligt för certifiering
1. Varje parti humle som görs tillgängligt för certifiering skall åtföljas av en beskrivning som undertecknats av producenten och innehåller följande uppgifter:
a) Producentens namn och adress.
b) Skördeår.
c) Sort.
d) Produktionsplats.
e) Skiftesbeteckningen i det integrerade administrations- och kontrollsystemet enligt artikel 17 i rådets förordning (EG) nr 1782/2003 [4] eller utdrag ur fastighetsregistret eller en officiell motsvarighet till detta.
f) Antalet förpackningar i partiet.
2. Beskrivningen enligt punkt 1 skall åtfölja humlepartiet under all bearbetning eller blandning och i varje fall till dess att certifikatet är utfärdat.
Artikel 4
Krav för avsättning
1. Humle skall för att kunna certifieras uppfylla villkoren i artikel 2 a i förordning (EG) nr 1952/2005 och de minimikrav för avsättning som anges i bilaga I till den här förordningen.
2. Företrädare för den behöriga certifieringsmyndigheten skall med tillämpning av någon av metoderna i bilaga II B kontrollera att de minimikrav för avsättning som gäller humlets vattenhalt uppfylls.
Den metod som anges i bilaga II B 2 skall godkännas av den behöriga certifieringsmyndigheten och måste ge resultat med en standardavvikelse på högst 2,0. Om det uppstår en tvist skall kontrollen göras enligt den metod som anges i bilaga II B 1.
3. Kontrollen av att minimikraven för avsättning uppfylls förutom vad gäller vattenhalten skall göras i enlighet med normal handelspraxis.
Om det uppstår en tvist skall kontrollen göras enligt den metod som anges i bilaga II C.
Artikel 5
Provtagning
För genomförandet av de kontroller som avses i artikel 4.2 och 4.3 skall prover tas och behandlas i enlighet med den metod som anges i bilaga II A.
I varje parti skall prover tas från minst en förpackning av tio och i varje fall från minst två förpackningar i ett parti.
Artikel 6
Certifieringsförfarande
1. Certifieringsförfarandet skall omfatta utfärdande av certifikaten samt märkning och försegling av förpackningarna.
2. Certifieringen skall genomföras innan produkten bjuds ut till försäljning och alltid före bearbetning.
Den skall ske senast den 31 mars året efter skördeåret. Medlemsstaterna får fastställa ett tidigare datum.
3. Märkningen skall göras enligt anvisningarna i bilaga III, under officiell tillsyn och efter försegling, på varje förpackning i vilken produkten skall avsättas.
4. Certifieringsförfarandet skall äga rum på odlingen eller i certifieringscentraler.
5. Om humlet byter emballage efter certifieringen, eventuellt i samband med bearbetning, skall humlet genomgå ett nytt certifieringsförfarande.
Artikel 7
Blandningar
1. Humle som certifierats i enlighet med denna förordning får blandas endast under officiell tillsyn i certifieringscentraler.
2. Humle som skall blandas måste komma från samma produktionsområde för humle, samma skörd och vara av samma sort.
3. Genom avvikelse från punkt 2 får dock certifierat humle av gemenskapsursprung som kommer från samma skörd men är av olika sorter och från olika produktionsområden för humle blandas vid tillverkning av pulver och extrakt, under förutsättning att det certifikat som åtföljer produkten anger
a) vilka sorter som använts, humlets produktionsområden och skördeår,
b) procentuell vikt för varje sort som ingår i blandningen; om humleprodukter har använts i kombination med humlekottar vid tillverkningen av humleprodukter, eller om olika humleprodukter har använts, skall den procentuella vikten för varje sort anges baserat på den kvantitet humlekottar som användes vid framställningen av de använda produkterna,
c) referensnummer på de certifikat som utfärdats för det humle och de humleprodukter som ingår.
Artikel 8
Återförsäljning
Humle som återförsäljes inom gemenskapen efter det att ett certifierat parti har delats upp, skall åtföljas av en faktura eller annat dokument upprättat av säljaren som anger certifikatets referensnummer.
Följande upplysningar från certifikatet skall också anges på fakturan eller i dokumentet:
a) Produktens beteckning.
b) Bruttovikt och/eller nettovikt.
c) Produktionsplats.
d) Skördeår.
e) Sort.
KAPITEL 3
HUMLEPRODUKTER
Artikel 9
Certifieringsförfarande
1. Certifieringsförfarandet skall omfatta utfärdande av certifikaten samt märkning och försegling av förpackningarna.
2. Certifieringen skall genomföras innan produkten bjuds ut till försäljning.
3. Märkningen skall göras enligt anvisningarna i bilaga III, under officiell tillsyn och efter försegling, på varje förpackning i vilken produkten skall avsättas.
4. Certfieringsförfarandet skall äga rum i certifieringscentraler.
5. Om humleprodukterna byter emballage efter certifieringen, eventuellt i samband med vidare bearbetning, skall produkten genomgå ett nytt certifieringsförfarande.
Artikel 10
Behandling i en sluten tillverkningsprocess
1. Behandlat humle, framställt av humle som certifierats i obehandlat skick, får certifieras endast om behandlingen ägt rum i en sluten tillverkningsprocess.
Första stycket gäller även produkter som framställs av humle som avses i artikel 1.4.
2. Om humlet behandlas i en certifieringscentral gäller följande:
a) Certifikatet skall inte utfärdas förrän efter behandlingen.
b) Det ursprungliga obehandlade humlet skall åtföljas av den beskrivning som avses i artikel 3.1.
3. Före behandlingen skall det ursprungliga obehandlade humlepartiet tilldelas ett identifieringsnummer. Detta nummer måste anges på det certifikat som utfärdas för det behandlade humlet.
4. Med undantag av de substanser som anges i bilaga IV får endast certifierat humle och certifierade humleprodukter som avses i artikel 1.4 i denna förordning tillsättas den slutna tillverkningsprocessen. De får endast tillsättas i samma skick som då de certifierades.
5. Om bearbetningen i den slutna tillverkningsprocessen vid produktion av extrakt, som framställs med användning av koldioxid, måste avbrytas av tekniska skäl, skall företrädarna för den behöriga certifieringsmyndigheten säkerställa att den förpackning som innehåller mellanprodukten förseglas i det ögonblick då processen avbryts. Förseglingen får endast brytas av företrädare för den behöriga certifieringsmyndigheten när processen sätts igång på nytt.
Artikel 11
Officiell tillsyn vid framställning av humleprodukter
1. Vid framställningen av humleprodukter skall företrädare för den behöriga certifieringsmyndigheten vara närvarande under hela den tid då bearbetningen sker. De skall på lämpligt sätt övervaka alla skeden i framställningen, från det att den förseglade förpackning öppnas som innehåller det humle eller de humleprodukter som skall bearbetas, till dess att förpackning, försegling och märkning av humleprodukten har avslutats. Företrädare för den behöriga certifieringsmyndigheten får vara frånvarande om det genom tekniska åtgärder, som den behöriga certifieringsmyndigheten har godkänt, kan garanteras att bestämmelserna i denna förordning ändå iakttas.
2. Före byte till en annan sats i tillverkningssystemet skall företrädarna för den behöriga certifieringsmyndigheten genom officiell tillsyn försäkra sig om att tillverkningssystemet är tomt, åtminstone i den utsträckning som krävs för att kunna konstatera att innehållet i två olika satser inte kan blandas.
Om humle, humleprodukter, humlerester eller någon annan produkt som härrör från humle finns kvar i tillverkningssystemet, exempelvis i blandnings- eller påfyllningsbehållarna, medan humle från en annan sats bearbetas, måste dessa delar kopplas ifrån genom lämpliga tekniska åtgärder och under officiell tillsyn. De får kopplas tillbaka till tillverkningssystemet endast under officiell tillsyn.
Det får inte finnas någon fysisk förbindelse mellan tillverkningslinjerna för koncentrerat humlepulver och icke-koncentrerat humlepulver när någon av dem är i drift.
Artikel 12
Information och uppgiftsregistrering
1. Driftsledningen på bearbetningsanläggningen skall förse företrädarna för den behöriga certifieringsmyndigheten med all information som rör de tekniska funktionerna i anläggningen.
2. Driftsledningen skall göra exakta noteringar om de bearbetade humlemängderna. För varje sats humle som skall bearbetas skall det upprättas en redogörelse med uppgifter om den ingående och den bearbetade produktens vikt.
Vad beträffar den ingående produkten skall certifikatets referensnummer anges för alla berörda humlepartier och humlesorter. Om mer än en sort används i samma sats skall deras respektive andel av vikten anges i noteringarna.
Vad beträffar den bearbetade produkten skall sorten också framgå av noteringarna eller, om produkten är en blandning, sortsammansättningen anges.
Alla viktangivelser får avrundas till närmaste kilogram.
3. Så snart bearbetningen av en sats har avslutats skall en förteckning över de producerade mängderna upprättas under officiell tillsyn och undertecknas av företrädare för den behöriga certifieringsmyndigheten.
Handlingarna skall förvaras av anläggningens driftsledning under minst tre år.
Artikel 13
Ompackning
1. När humlepulver och humleextrakt fortfarande är i omlopp får ompackning med eller utan vidare bearbetning ske bara under officiell tillsyn.
2. Om ompackning sker utan bearbetning av produkten skall det nya certifieringsförfarandet bara omfatta
a) märkning av den nya förpackningen,
b) angivande av denna märkning och av ompackningen på det ursprungliga certifikatet.
Artikel 14
Blandningar
1. Humleprodukter som certifierats i enlighet med denna förordning får blandas endast under officiell tillsyn i certifieringscentraler.
2. Certifierade humleprodukter som framställts av certifierat humle av gemenskapsursprung som kommer från samma skörd men är av olika sorter och från olika produktionsområden för humle får dock blandas vid tillverkning av pulver och extrakt, under förutsättning att det certifikat som åtföljer produkten anger
a) vilka sorter som använts, humlets produktionsområden och skördeår,
b) procentuell vikt för varje sort som ingår i blandningen; om humleprodukter har använts i kombination med humlekottar vid tillverkningen av humleprodukter, eller om olika humleprodukter har använts, skall den procentuella vikten för varje sort anges baserad på den kvantitet humlekottar som användes vid framställningen av de använda produkterna,
c) referensnummer på de certifikat som utfärdats för det humle och de humleprodukter som ingår.
Artikel 15
Återförsäljning
Humleprodukter som återförsäljes inom gemenskapen efter det att ett certifierat parti har delats upp, skall åtföljas av en faktura eller annat dokument upprättat av säljaren som anger certifikatets referensnummer. Följande upplysningar från certifikatet skall också anges på fakturan eller i dokumentet:
a) Produktens beteckning.
b) Bruttovikt och/eller nettovikt.
c) Produktionsplats.
d) Skördeår.
e) Sort.
f) Plats och datum för bearbetningen.
KAPITEL 4
CERTIFIERING OCH MÄRKNING
Artikel 16
Certifikat
1. Certifikatet skall utfärdas i det handelsled för vilket minimikraven för avsättning gäller.
2. När det gäller humlekottar skall certifikatet innehålla minst följande uppgifter:
a) En beskrivning av produkten.
b) Certifikatets referensnummer.
c) Nettovikt och/eller bruttovikt.
d) Humlets produktionsområde eller produktionsplatsen enligt artikel 4.3 a i förordning (EG) nr 1952/2005.
e) Skördeår.
f) Sort.
g) Uppgiften "humle med frö" eller "humle utan frö".
h) Åtminstone en av de uppgifter som anges i bilaga V och som används av den behöriga certifieringsmyndigheten.
3. När det gäller produkter som framställts av humle skall certifikatet, utöver de uppgifter som anges i punkt 2, innehålla uppgift om plats och datum för bearbetningen.
4. Det referensnummer på certifikatet som avses i punkt 2 b skall bestå av koder som i enlighet med bilaga VI anger certifieringscentral, medlemsstat, skördeår och parti.
Referensnumret skall vara detsamma på alla förpackningar som ingår i ett parti.
Artikel 17
Information på förpackningen
På varje förpackning skall minst följande uppgifter lämnas på ett av gemenskapens språk:
a) En beskrivning av produkten samt uppgiften "humle med frö" respektive "humle utan frö" och "behandlat humle" respektive "obehandlat humle", allt efter omständigheterna.
b) Sort eller sorter.
c) Certifikatets referensnummer.
Uppgifterna skall anges med lättläsliga bokstäver av enhetlig storlek med outplånligt tryck.
Artikel 18
Humle från försökssorter
När det gäller humle från försökssorter under utveckling, producerat av ett forskningsinstitut på dess egna odlingar eller av en producent för ett sådant instituts räkning, får de uppgifter som avses i artikel 16.2 f och artikel 17 b ersättas av ett namn eller nummer som identifikation av sorten i fråga.
Artikel 19
Bevis på certifiering
Uppgifterna på varje förpackning och certifikatet som åtföljer produkten skall utgöra bevis om att certifiering har skett.
KAPITEL 5
UNDANTAG
Artikel 20
Särskilda krav
1. I det fall som avses i artikel 1.3 a skall bryggeriet, för varje skörd, senast den 15 november varje år till den behöriga certifieringsmyndigheten sända upplysningar om vilka sorter som odlats, vilka kvantiteter som skördats, produktionsplatser och planterade arealer, samt skiftesbeteckningen i det integrerade administrations- och kontrollsystemet eller utdrag ur fastighetsregister eller en motsvarande officiell beteckning.
Punkt 2 a–d och 2 f skall dessutom gälla i tillämpliga delar, utom när humlet bearbetas eller används i obearbetat skick av bryggeriet självt.
2. I det fall som avses i artikel 1.3 b skall den behöriga certifieringsmyndigheten på bryggeriets begäran, när humlet levererats till den anläggning där det skall bearbetas, upprätta ett dokument där minst följande uppgifter skall införas under bearbetningens gång:
a) Avtalets referensnummer.
b) Det bryggeri som produkterna är avsedda för.
c) Bearbetningsanläggningen.
d) En beskrivning av den bearbetade produkten.
e) Referensnumret på certifikatet eller det likvärdiga intyget för det ursprungliga humlet.
f) Den bearbetade produktens vikt.
Det dokument som avses i första stycket skall förses med ett referensnummer som också skall anges på förpackningen.
När det gäller blandningar av humle skall dessutom följande anges i dokumentet och på förpackningen:
"Blandning av humle för eget bruk. Får inte säljas."
3. I det fall som avses i artikel 1.3 c får förpackningens vikt inte överstiga
a) 1 kg för humlekottar eller humlepulver,
b) 300 g för extrakt, pulver och nya isomeriserade produkter.
En beskrivning av produkten samt vikten måste anges på förpackningen.
KAPITEL 6
CERTIFIERINGSORGAN
Artikel 21
Behörig certifieringsmyndighet
1. Medlemsstaterna skall utse en behörig certifieringsmyndighet och se till att nödvändiga kontroller och förfaranden genomförs för att garantera att humlet och humleprodukterna håller minimikvalitet och kan spåras.
2. Den behöriga certifieringsmyndigheten eller dess företrädare skall genomföra certifieringen. Den skall ha de resurser som krävs för att kunna utföra sina arbetsuppgifter.
3. Den behöriga certifieringsmyndigheten ansvarar för kontrollen av att bestämmelserna i denna förordning efterlevs. Regelbundenheten eller frekvensen för dessa kontroller skall bestämmas av medlemsstaten på grundval av en riskanalys, men minst en kontroll per månad skall genomföras. Varje år skall det göras en utvärdering av hur effektiva parametrarna i tidigare års riskanalyser har varit.
Artikel 22
Godkännande av certifieringscentraler
1. Den behöriga certifieringsmyndigheten skall godkänna certifieringscentraler som är juridiska personer eller som har tillräcklig rättskapacitet för att enligt den nationella lagstiftningen kunna inneha rättigheter och skyldigheter, och den skall se till att dessa har tillräckliga resurser för att kunna utföra de arbetsuppgifter som krävs för provtagning, analyser, statistikföring och registrering.
Den behöriga certifieringsmyndigheten skall på grundval av en riskanalys, men minst två gånger per kalenderår, genomföra stickprovskontroller på plats i certifieringscentralerna för att kontrollera att bestämmelserna i föregående stycke efterlevs. Varje år skall det göras en utvärdering av hur effektiva parametrarna i tidigare års riskanalyser har varit.
2. Om det konstateras att beståndsdelar som inte är tillåtna har använts vid framställningen av humleprodukter, eller om de beståndsdelar som använts inte motsvarar uppgifterna i certifikatet enligt artikel 16, och om detta kan tillskrivas certifieringscentralen som en medveten handling eller allvarligt fel, skall den behöriga certifieringsmyndigheten återkalla godkännandet av certifieringscentralen.
Ett nytt godkännande får inte beviljas inom de första tolv månaderna efter återkallandet. På anhållan av den certifieringscentral vars godkännande har återkallats skall ett nytt godkännande utfärdas efter två år, eller i allvarliga fall efter tre år, efter det att godkännandet återkallades.
KAPITEL 7
MEDDELANDEN OCH OFFENTLIGGÖRANDE AV FÖRTECKNINGARNA
Artikel 23
Meddelanden
1. Medlemsstaterna skall senast den 30 juni 2007 till kommissionen lämna uppgifter om
a) den behöriga certifieringsmyndighetens namn och adress,
b) de åtgärder som vidtagits för att genomföra denna förordning.
2. Medlemsstaterna skall senast den 30 juni varje år till kommissionen överlämna
a) en förteckning över produktionsområden för humle,
b) en förteckning över certifieringscentralerna och den kod som varje central har tilldelats,
c) uppgifter om ändringar som skett av den behöriga certifieringsmyndighetens namn och adress under det föregående året.
Artikel 24
Offentliggörande av förteckningarna
Kommissionen skall se till att förteckningen över produktionsområdena för humle och förteckningen över certifieringscentralerna och deras koder uppdateras varje år och finns tillgänglig på kommissionens webbplats [5].
KAPITEL 8
SLUTBESTÄMMELSER
Artikel 25
Upphävande
Förordning (EEG) nr 1784/77 och förordning (EEG) nr 890/78 skall upphöra att gälla.
Hänvisningar till de upphävda förordningarna skall anses som hänvisningar till denna förordning och skall läsas i enlighet med jämförelsetabellen i bilaga VII.
Artikel 26
Ikraftträdande
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Den skall tillämpas från och med den 1 april 2007.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
BESLUT FATTAT AV DE I RÅDET FÖRSAMLADE FÖRETRÄDARNA FÖR MEDLEMSSTATERNAS REGERINGAR av den 18 december 1987 om nomenklaturen och konventionella tullsatser för vissa produkter och om allmänna regler för tolkning och tillämpning av nämnda nomenklatur och tullar (87/597/EKSG)
DE I RÅDET FÖRSAMLADE FÖRETRÄDARNA FÖR REGERINGARNA I EUROPEISKA KOL- OCH STÅLGEMENSKAPENS MEDLEMSSTATER HAR BESLUTAT FÖLJANDE
Artikel 1
Från och med den 1 januari 1988 skall medlemsstaternas gemensamma tullnomenklatur samt de konventionella tullar som tillämpas på produkter som omfattas a
VERKSTÄLLANDE KOMMITTÉNS BESLUT
av den 14 december 1993
om ministrarnas och statssekreterarnas förklaringar
(SCH/Com-ex (93) 10)
VERKSTÄLLANDE KOMMITTÉN HAR FATTAT DETTA BESLUT
med beaktande av artikel 132 i konventionen om tillämpning av Schengenavtalet.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Ministrarnas och statssekreterarnas förklaringar av den 19 juni 1992(1) och den 30 juni 1993 om genomförandet av Schengenavtalets tillämpningskonvention och om uppfyllande av villkoren bekräftas härmed.
Paris den 14 december 1993.
Alain Lamassoure
Ordförande
(1) Förklaringarna av den 19 juni 1992 har inte överförts till regelverket.
MINISTRARNAS OCH STATSSEKRETERARNAS FÖRKLARINGAR
Madrid den 30 juni 1993.
SCH/M (93) 14
1. Ministrarna och statssekreterarna är härmed eniga om att fastställa det politiska målet om tillämpning av 1990 års konvention till den 1 december 1993.
2. Ministrarna och statssekreterarna noterar att följande villkor har uppfyllts:
- den gemensamma handboken,
- bestämmelserna om utfärdande av enhetliga viseringar och gemensamma konsulära anvisningar,
- handläggning av asylansökningar,
- flygplatserna, enligt överenskommelse i ministrarnas och statssekreterarnas förklaring av den 19 juni 1992.
Stora framsteg har gjorts beträffande de andra villkoren, som redan har uppfyllts i sådan utsträckning att ovannämnda tillämpning bör vara möjlig från och med den 1 december 1993. Därför, och i överensstämmelse med 1990 års Schengenkonvention, behövs det ytterligare insatser för att genomföra de bestämmelser som redan har fastställts beträffande kontroll av de yttre gränserna och av narkotika.
Ministrarna och statssekreterarna bekräftar att ett operationellt SIS är en ovillkorlig förutsättning för avskaffandet av kontrollerna vid de inre gränserna. Betydande framsteg har gjorts inom detta område. De är eniga om att öka tempot i arbetet för att möjliggöra att SIS gradvis blir operationellt, allteftersom staterna genomför framgångsrika test och de nationella delarna av SIS blir operationella.
3. Vid mötet i oktober kommer Verkställande kommittén att slutligen ta ställning till genomförandet av de övriga insatser som nämns ovan.
4. 1990 års Schengenkonvention kommer att gälla i alla de medlemsstater som har uppfyllt villkoren och som har ett operationellt nationellt SIS.
För att kunna åstadkomma detta åtar sig alla medlemsstater att genomföra alla nödvändiga åtgärder för att fullfölja de nationella förfaranden som krävs för att ratificera konventionen och anslutningsavtalen.
5. Ministrarna och statssekreterarna är eniga om att de stater som ursprungligen undertecknade 1990 års konvention snarast möjligt måste deponera sina ratifikationsinstrument, om de inte redan har gjort detta, och senast vid en tidpunkt som möjliggör att det datum som anges i punkt 1 iakttas. Medlemsstaterna samtycker även till att, om det inte redan har gjorts, snarast möjligt och senast vid en tidpunkt som möjliggör att datumet i punkt 1 iakttas, deponera sina ratificeringsinstrument för de stater vars nationella SIS skall integreras i systemet. Detta åtagande skall även gälla allteftersom de andra medlemsstaterna uppnår en likvärdig nivå i sitt nationella SIS.
Ministrarna och statssekreterarna är eniga om att förklaringen till artikel 139 i slutakten till konventionen innebär att konventionen kan börja tillämpas när Verkställande kommittén fattat beslut om detta vilket skall ske så snart som villkoren är uppfyllda.
till konventionen om tillämpning av Schengenavtalet av den 14 juni 1985 mellan regeringarna i Beneluxstaterna, Förbundsrepubliken Tyskland och Franska republiken om gradvis avskaffande av kontroller vid de gemensamma gränserna, undertecknad i Schengen den 19 juni 1990, till vilken Italienska republiken anslutit sig genom avtal undertecknat i Paris den 27 november 1990 KONUNGARIKET BELGIEN, FÖRBUNDSREPUBLIKEN TYSKLAND, FRANSKA REPUBLIKEN, STORHERTIGDÖMET LUXEMBURG och KONUNGARIKET NEDERLÄNDERNA, som är parter i konventionen om tillämpning av Schengenavtalet av den 14 juni 1985 mellan regeringarna i Beneluxstaterna, Förbundsrepubliken Tyskland och Franska republiken om gradvis avskaffande av kontroller vid de gemensamma gränserna, undertecknad i Schengen den 19 juni 1990, nedan kallad %quot%1990 års konvention%quot%, och Italienska republiken, som anslutit sig till 1990 års konvention genom avtal undertecknat i Paris den 27 november 1990, å ena sidan,
som beaktar undertecknandet i Bonn den 25 juni 1991 av protokollet om Portugisiska republikens regerings anslutning till Schengenavtalet av den 14 juni 1985 mellan regeringarna i Beneluxstaterna, Förbundsrepubliken Tyskland och Franska republiken, om gradvis avskaffande av kontroller vid de gemensamma gränserna, ändrat genom Italienska republikens regerings anslutningsprotokoll, undertecknat i Paris den 27 november 1990, och som stöder sig på artikel 140 i 1990 års konvention,
1. De polismän som avses i artikel 40.4 i 1990 års konvention är, när det gäller Portugisiska republiken, polismän i Policía Judiciária samt tulltjänstemän när de biträder åklagarmyndigheten, på de villkor som fastställs i de lämpliga bilaterala avtal som avses i artikel 40.6 i 1990 års konvention, när det gäller deras åligganden i fråga om olaglig handel med narkotika och psykotropa ämnen, olaglig handel med vapen och sprängämnen samt olaglig transport av giftigt och farligt avfall. 2. Den myndighet som avses i artikel 40.5 i 1990 års konvention är, när det gäller Portugisiska republiken, Direccão geral de la Policía Judiciária.
Artikel 3
1. De polismän som avses i artikel 41.7 i 1990 års konvention är, när gäller Portugisiska republiken, polismän i Policía Judiciária (kriminalpolisen) samt tulltjänstemän när de biträder åklagarmyndigheten, på de villkor som fastställs i de lämpliga bilaterala avtal som avses i artikel 41.10 i 1990 års konvention, när det gäller deras åligganden i fråga om olaglig handel med narkotika och psykotropa ämnen, olaglig handel med vapen och sprängämnen samt olaglig transport av giftigt och farligt avfall. 2. Vid undertecknandet av detta avtal skall Portugisiska republikens regering avge en förklaring, när det gäller Konungariket Spaniens regering, i vilken det fastställs, på grundval av artikel 41.2, 41.3 och 41.4 i 1990 års konvention, vilka förfaranden som skall gälla för förföljande över gränserna in på dess territorium.
Artikel 4 Det behöriga ministerium som avses i artikel 65.2 i 1990 års konvention är, när det gäller Portugisiska republiken, justitieministeriet.
När det gäller utlämning mellan de avtalsslutande parterna i 1990 års konvention skall stycket under c i Portugisiska republikens förklaring om artikel 1 i den europeiska utlämningskonventionen av den 13 december 1957, lyda på följande sätt: Portugisiska republiken kommer inte att medge utlämning av personer vars utlämning begärs för ett brott som kan bestraffas med fängelsestraff på livstid. Likväl kan utlämning medges om den ansökande staten försäkrar att den i enlighet med sin lagstiftning och sin praxis för verkställande av straff kommer att förespråka anpassningsåtgärder som den person vars utlämning begärs skulle kunna komma i åtnjutande av.
1. Detta avtal skall ratificeras, godkännas eller godtas. Ratifikations-, godkännande- eller godtagandeinstrumenten skall deponeras hos Storhertigdömet Luxemburgs regering, som skall underrätta samtliga avtalsslutande parter om deponeringen. 2. Detta avtal träder i kraft den första dagen i den andra månaden efter det att de fem signatärstaterna till 1990 års konvention och Portugisiska republiken har deponerat sina ratifikations-, godkännande- eller godtagandeinstrument, och tidigast den dag då 1990 års konvention träder i kraft. I förhållande till Italienska republiken träder avtalet i kraft den första dagen i den andra månaden efter det att den staten har deponerat sina ratifikations-, godkännande- eller godtagandeinstrument, och tidigast den dag då avtalet träder i kraft mellan de övriga avtalsslutande parterna.
3. Storhertigdömet Luxemburgs regering skall underrätta samtliga avtalsslutande parter om datum för ikraftträdandet. Artikel 8
1. Storhertigdömet Luxemburgs regering skall till Portugisiska republikens regering överlämna en bestyrkt kopia av 1990 års konvention på tyska, franska, italienska och nederländska. 2. Texten till 1990 års konvention, upprättad på portugisiska, bifogas detta avtal och gäller på samma villkor som de texter till 1990 års konvention som är upprättade på tyska, franska, italienska och nederländska.
Till bevis härför har undertecknade befullmäktigade undertecknat detta avtal. Upprättat i Bonn den tjugofemte juni nittonhundranittioett i ett enda original på tyska, franska, italienska, nederländska och portugisiska, vilka samtliga fem texter är lika giltiga, som skall deponeras i arkiven hos Storhertigdömet Luxemburgs regering, som skall överlämna en bestyrkt kopia därav till varje avtalsslutande part.
%gt%PIC FILE= %quot%L_2000239SV.007701.TIF%quot%%gt% För Förbundsrepubliken Tysklands regering
%gt%PIC FILE= %quot%L_2000239SV.007803.TIF%quot%%gt% För Konungariket Nederländernas regering
SLUTAKT I. Vid undertecknandet av avtalet om Portugisiska republikens anslutning till konventionen om tillämpning av Schengenavtalet av den 14 juni 1985 om gradvis avskaffande av kontroller vid de gemensamma gränserna, undertecknad i Schengen den 19 juni 1990 mellan regeringarna i Beneluxstaterna, Förbundsrepubliken Tyskland och Franska republiken, till vilket Italienska republiken anslutit sig genom avtal undertecknat i Paris den 27 november 1990, ansluter sig Portugisiska republikens regering till slutakten, protokollet och ministrarnas och statssekreterarnas gemensamma förklaring, som undertecknades i samband med undertecknandet av 1990 års konvention.
Portugisiska republikens regering ansluter sig till de gemensamma förklaringarna och noterar de ensidiga förklaringarna i dessa. Storhertigdömet Luxemburgs regering skall till Portugisiska republikens regering överlämna en bestyrkt kopia av slutakten, protokollet och ministrarnas och statssekreterarnas gemensamma förklaring, som undertecknades i samband med undertecknandet av 1990 års konvention på tyska, franska, italienska och nederländska.
Texterna till slutakten, protokollet och ministrarnas och statssekreterarnas gemensamma förklaring, som undertecknades i samband med undertecknandet av 1990 års konvention, upprättade på portugisiska, bifogas denna slutakt och är giltiga på samma villkor som de texter som är upprättade på tyska, franska, italienska och nederländska. II. Vid undertecknandet av avtalet om Portugisiska republikens anslutning till konventionen om tillämpning av Schengenavtalet av den 14 juni 1985 mellan regeringarna i Beneluxstaterna, Förbundsrepubliken Tyskland och Franska republiken om gradvis avskaffande av kontroller vid de gemensamma gränserna, undertecknad i Schengen den 19 juni 1990, till vilken Italienska republiken anslutit sig genom avtal undertecknat i Paris den 27 november 1990, har de avtalsslutande parterna antagit följande förklaringar:
1) Gemensam förklaring om artikel 7 i anslutningsavtalet Signatärstaterna skall redan innan anslutningsavtalet träder i kraft underrätta varandra om alla omständigheter av betydelse för de frågor som avses i 1990 års konvention och för genomförandet av anslutningsavtalet.
Detta anslutningsavtal skall inte genomföras mellan de fem signatärstaterna till 1990 års konvention och Portugisiska republiken förrän villkoren för tillämpning av 1990 års konvention har uppfyllts i dessa sex stater och bevakningen av de yttre gränserna blivit genomförd. I förhållande till Italienska republiken skall detta anslutningsavtal inte genomföras förrän villkoren för tillämpning av 1990 års konvention har uppfyllts i signatärstaterna till det avtalet och bevakningen av de yttre gränserna blivit genomförd. 2) Gemensam förklaring om artikel 9.2 i 1990 års konvention
De avtalsslutande parterna slår fast att vid tiden för undertecknandet av avtalet om Italienska republikens anslutning till 1990 års konvention är de gemensamma viseringsregler som avses i artikel 9.2 i 1990 års konvention de gemensamma regler som från och med den 19 juni 1990 tillämpas mellan signatärstaterna till den konventionen. 3) Gemensam förklaring om skydd av personuppgifter
De avtalsslutande parterna noterar att Portugisiska republiken den 29 april 1991 offentliggjorde en lag om skydd av personuppgifter vid automatisk databehandling. De avtalsslutande parterna noterar att Portugisiska republikens regering åtar sig att före ratifikationen av avtalet om anslutning till 1990 års konvention ta alla nödvändiga initiativ för att komplettera den portugisiska lagstiftningen så att samtliga bestämmelser i 1990 års konvention som rör skyddet av personuppgifter kan tillämpas fullt ut.
1) Förklaring om brasilianska medborgare som reser in i Portugal enligt avtalet om avskaffande av visering mellan Portugal och Brasilien av den 9 augusti 1960 Portugisiska republikens regering åtar sig att på sitt territorium tillåta återinresa av brasilianska medborgare vilka, efter att ha rest in på de avtalsslutande parternas territorium via Portugal i enlighet med avtalet om avskaffande av visering mellan Portugal och Brasilien, återfinns på de avtalsslutande parternas territorium efter den tidsperiod som avses i artikel 20.1 i 1990 års konvention.
Portugisiska republikens regering åtar sig att tillåta inresa av brasilianska medborgare endast om de uppfyller de villkor som anges i artikel 5 i 1990 års konvention och vidta alla åtgärder för att se till att deras resehandlingar stämplas när de passerar de yttre gränserna. 2) Förklaring om den europeiska konventionen om inbördes rättshjälp i brottmål
Portugisiska republikens regering åtar sig att ratificera den europeiska konventionen om inbördes rättshjälp i brottmål av den 20 april 1959 och dess tilläggsprotokoll innan 1990 års konvention träder i kraft för Portugal. 3) Förklaring om överenskommelsen om exportrestriktioner för missilteknik och -utrustning (MTCR)
För tillämpningen av artikel 123 i 1990 års konvention åtar sig Portugisiska republikens regering att snarast möjligt, och senast när 1990 års konvention träder i kraft för Portugal, ansluta sig till överenskommelsen om exportrestriktioner för missilteknik och -utrustning (MTCR), i dess lydelse av den 16 april 1987. 4) Förklaring om artikel 121 i 1990 års konvention
Portugisiska republikens regering förklarar att den, utom när det gäller färska frukter av citrus, skall tillämpa den förenkling av växtskyddskontroller som avses i artikel 121 i 1990 års konvention från tidpunkten för undertecknandet av avtalet om anslutning till 1990 års konvention. Portugisiska republiken förklarar att den före den 1 januari 1992 skall utföra en bedömning av risken för skadliga organismer (pest risk assessment) på färska frukter av citrus, vilken, om den visar att det finns risk för att skadliga organismer förs in eller sprids, i förekommande fall kan motivera undantaget enligt artikel 121.2 i 1990 års konvention efter det att avtalet om Konungariket Spaniens anslutning har trätt i kraft.
5) Förklaring om avtalet om Konungariket Spaniens anslutning till 1990 års konvention
Vid undertecknandet av detta avtal noterar Portugisiska republiken innehållet i avtalet om Konungariket Spaniens anslutning till 1990 års konvention liksom i den till det avtalet fogade slutakten och förklaringen. Upprättad i Bonn den tjugofemte juni nittonhundranittioett i ett enda original på spanska, tyska, franska, italienska och nederländska, vilka samtliga fem texter är lika giltiga, som skall deponeras i arkiven hos Storhertigdömet Luxemburgs regering, som skall överlämna en bestyrkt kopia till varje avtalsslutande part.
%gt%PIC FILE= %quot%L_2000239SV.008101.TIF%quot%%gt% För Förbundsrepubliken Tysklands regering
FÖRKLARING AV MINISTRARNA OCH STATSSEKRETERARNA Den 25 juni 1991 undertecknade företrädare för regeringarna i Konungariket Belgien, Förbundsrepubliken Tyskland, Franska republiken, Italienska republiken, Storhertigdömet Luxemburg, Konungariket Nederländerna och Portugisiska republiken i Bonn avtalet om Portugisiska republikens anslutning till konventionen om tillämpning a
Beslut av företrädarna för medlemsstaternas regeringar
av den 6 april 2006
om utnämning av domare och generaladvokater vid Europeiska gemenskapernas domstol
(2006/281/EG, Euratom)
FÖRETRÄDARNA FÖR REGERINGARNA I EUROPEISKA GEMENSKAPERNAS MEDLEMSSTATER HAR BESLUTAT FÖLJANDE
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 223,
med beaktande av fördraget om upprättandet av Europeiska atomenergigemenskapen, särskilt artikel 139, och
av följande skäl:
(1) Mandattiden för domarna Peter JANN, Christiaan TIMMERMANS, Konrad SCHIEMANN, Jiří MALENOVSKÝ, Jean-Pierre PUISSOCHET, Ninon COLNERIC och Stig VON BAHR, Antonio TIZZANO, José Narciso DA CUNHA RODRIGUES, Pranas KŪRIS, George ARESTIS, Anthony BORG BARTHET, Egils LEVITS och för generaladvokaterna Christine STIX-HACKL, Philippe LÉGER, Leendert GEELHOED och Paolo MENGOZZI, vid Europeiska gemenskapernas domstol, löper ut den 6 oktober 2006.
(2) Sammansättningen av Europeiska gemenskapernas domstol behöver delvis förnyas för tiden från och med den 7 oktober 2006 till och med den 6 oktober 2012. En domare kan dock inte utses förrän vid ett senare tillfälle, eftersom det saknas förslag.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Följande personer utnämns härmed till domare vid Europeiska gemenskapernas domstol för tiden från och med den 7 oktober 2006 till och med den 6 oktober 2012:
George ARESTIS
Jean-Claude BONICHOT
Anthony BORG BARTHET
José Narciso DA CUNHA RODRIGUES
Peter JANN
Pranas KŪRIS
Egils LEVITS
Pernilla LINDH
Jiří MALENOVSKÝ
Christiaan TIMMERMANS
Antonio TIZZANO
Konrad SCHIEMANN
2. Följande personer utnämns härmed till generaladvokater vid Europeiska gemenskapernas domstol för tiden från och med den 7 oktober 2006 till och med den 6 oktober 2012:
Yves BOT
Ján MAZÁK
Paolo MENGOZZI
Verica TRSTENJAK
Artikel 2
Detta beslut skall offentliggöras i Europeiska unionens officiella tidning.
P6_TA(2004)0073
Säkerhetsdetaljer och biometriska kännetecken i EU-medborgarnas pass * Europaparlamentets lagstiftningsresolution om komissionens förslag till rådets förordning om standarder för säkerhetsdetaljer och biometriska kännetecken i EU-medborgarnas pass (KOM(2004)0116 - C5-0101/2004 - 2004/0039(CNS))
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
- med beaktande av kommissionens förslag (KOM(2004)0116) [1],
- med beaktande av rådets riktlinjer enligt dokument 15139/2004 som överlämnades till parlamentet den 24 november 2004,
- med beaktande av artikel 62.2 a i EG-fördraget,
- med beaktande av artikel 67 i EG-fördraget, i enlighet med vilken rådet har hört parlamentet (C5-0101/2004),
- med beaktande av protokollet om införlivande av Schengenregelverket inom Europeiska unionens ramar, i enlighet med vilket rådet har hört parlamentet,
- med beaktande av artikel 51 i arbetsordningen,
- med beaktande av betänkandet från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor (A6-0028/2004).
1. Europaparlamentet godkänner kommissionens förslag såsom ändrat av parlamentet.
2. Kommissionen uppmanas att ändra sitt förslag i överensstämmelse härmed i enlighet med artikel 250.2 i EG-fördraget.
3. Rådet uppmanas att underrätta Europaparlamentet om rådet har för avsikt att avvika från den text som parlamentet har godkänt.
4. Europaparlamentet begär att medlingsförfarandet enligt den gemensamma förklaringen av den 4 mars 1975 inleds om rådet har för avsikt att avvika från den text som parlamentet har godkänt.
5. Rådet uppmanas att höra Europaparlamentet om rådet har för avsikt att avvika från kommissionens förslag.
6. Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
KOMMISSIONENS FÖRSLAG | PARLAMENTETS ÄNDRINGAR |
Ändring 1
Skäl 2
(2) Minimisäkerhetsstandarder för pass infördes genom en resolution antagen av företrädarna för medlemsstaternas regeringar, församlade i rådet, av den 17 oktober 2000. Denna resolution bör nu ersättas och uppdateras genom en gemenskapsåtgärd i syfte att skapa mer harmoniserade säkerhetsstandarder för pass som ger ett bättre skydd mot förfalskning. Samtidigt bör biometriska kännetecken integreras i passet för att skapa en tillförlitlig koppling mellan den egentliga innehavaren och handlingen. | (2) Minimisäkerhetsstandarder för pass infördes genom en resolution antagen av företrädarna för medlemsstaternas regeringar, församlade i rådet, av den 17 oktober 2000. Europeiska rådet har beslutat att denna resolution nu bör ersättas och uppdateras genom en gemenskapsåtgärd i syfte att skapa mer harmoniserade säkerhetsstandarder för pass som ger ett bättre skydd mot förfalskning. Samtidigt bör biometriska kännetecken integreras i passet för att skapa en tillförlitlig koppling mellan den egentliga innehavaren och handlingen. |
Ändring 2
Skäl 2a (nytt)
| (2a) Biometriska uppgifter i pass bör användas endast för att kontrollera dokumentets äkthet och innehavarens identitet genom direkt tillgängliga jämförbara uppgifter när pass skall framläggas enligt lag. |
Ändring 3
Skäl 3
(3) Harmoniseringen av säkerhetsdetaljer och införandet av biometriska kännetecken är ett viktigt steg i användningen av nya element mot bakgrund av utvecklingen på EU-nivå för att göra resehandlingar säkrare och skapa en mer tillförlitlig koppling mellan innehavaren och passet, och därigenom hindra att passet används i bedrägligt syfte. Specifikationerna i Internationella civila luftfartsorganisationens (ICAO) dokument nr 9303 om maskinläsbara resehandlingar bör beaktas. | (3) Harmoniseringen av säkerhetsdetaljer och införandet av biometriska kännetecken är ett viktigt steg i användningen av nya element mot bakgrund av utvecklingen på EU-nivå för att göra resehandlingar säkrare och skapa en mer tillförlitlig koppling mellan innehavaren och passet, och därigenom hindra att passet används i bedrägligt syfte. |
Ändring 4
Skäl 7
(7) Beträffande vilka personuppgifter som kommer att användas för passändamål gäller Europaparlamentets och rådets direktiv 95/46/EG av den 24 oktober 1995 om skydd för enskilda personer med avseende på behandling av personuppgifter och om det fria flödet av sådana uppgifter. Det måste säkerställas att inga andra uppgifter lagras i passet om det inte föreskrivs i förordningen eller dess bilagor eller anges i den aktuella resehandlingen. | (7) Beträffande vilka personuppgifter som kommer att användas för passändamål gäller Europaparlamentets och rådets direktiv 95/46/EG av den 24 oktober 1995 om skydd för enskilda personer med avseende på behandling av personuppgifter och om det fria flödet av sådana uppgifter. Inga andra uppgifter bör lagras i passet. |
Ändring 5
Artikel 1, punkt 2
2. Passet skall vara försett med ett väl skyddat lagringsmedium som har tillräcklig kapacitet och som innehåller en ansiktsbild. Medlemsstaterna får även inkludera fingeravtryck i driftskompatibla format. | 2. Passet skall vara försett med ett väl skyddat lagringsmedium som har tillräcklig kapacitet och som kan säkra de lagrade uppgifternas integritet, äkthet och konfidentialitet. Det skall innehålla en ansiktsbild. Medlemsstaterna får även inkludera fingeravtryck i driftskompatibla format. Ingen central databas för Europeiska unionens pass och resehandlingar får upprättas som innehåller biometriska och andra uppgifter om samtliga innehavare av EU-pass. |
Ändring 6
Artikel 2, punkt 1, inledningen
1. Kompletterande tekniska specifikationer för passet som rör följande skall fastställas i enlighet med det förfarande som anges i artikel 5.2: | 1. Kompletterande tekniska specifikationer för passet som rör följande skall fastställas i enlighet med det förfarande som anges i artikel 5: |
Ändring 7
Artikel 2, punkt 1, led b
b)Tekniska specifikationer för lagringsmediet för de biometriska uppgifterna och skyddet av dessa. | b)Tekniska specifikationer för lagringsmediet för de biometriska uppgifterna och skyddet av dessa, i synnerhet för att säkra uppgifternas integritet, äkthet och konfidentialitet och för att garantera att de utnyttjas i enlighet med de ändamål som fastställs i denna förordning. |
Ändring 8
Artikel 2, punkt 1a (ny)
| 1a. Lagringsmediet får endast användas av a)de myndigheter i medlemsstaterna som är behöriga att ta del av, lagra, ändra och stryka uppgifter, ochb)godkända organ som enligt lag har rätt att ta del av uppgifterna, i syfte att ta del av uppgifterna. |
Ändring 9
Artikel 3, punkt 2a (ny)
| 2a. Varje medlemsstat skall upprätta en förteckning över behöriga myndigheter samt över godkända organ enligt artikel 2.1 a. Medlemsstaten skall översända denna förteckning med, om så behövs, regelbundna uppdateringar till kommissionen som skall upprätthålla en aktuell sammanställning online av de nationella förteckningarna. Kommissionen skall årligen offentliggöra denna sammanställning. |
Ändring 10
Artikel 4, punkt 1
1. Utan att det påverkar bestämmelserna om skydd av personuppgifter, har personer till vilka pass utfärdas rätt att kontrollera personuppgifterna i passet och begära att få uppgifter rättade eller strukna. | 1. Utan att det påverkar bestämmelserna om skydd av personuppgifter, har personer till vilka pass utfärdas rätt att kontrollera personuppgifterna i passet och begära att få uppgifter rättade eller strukna. Varje kontroll, rättelse eller strykning skall utföras kostnadsfritt av den utsedda nationella myndigheten. |
Ändring 11
Artikel 4, punkt 2
2. Uppgifter i maskinläsbar form får inte finnas i passet, om inte annat följer av förordningen eller bilagan till denna eller anges i passet. | 2. Uppgifter i maskinläsbar form får inte finnas i passet, om inte annat följer av förordningen eller bilagan till denna eller anges i passet. Inga andra uppgifter skall finnas i passet. |
Ändring 12
Artikel 4, punkt 2a (ny)
| 2a. De biometriska uppgifterna i pass skall endast utnyttjas för att kontrollera a)dokumentets äkthet,b)innehavarens identitet genom direkt tillgängliga jämförbara uppgifter när pass skall framläggas enligt lag. |
Ändring 13
Artikel 4, punkt 2b (ny)
| 2b. Medlemsstaterna skall regelbundet översända granskningsrapporter om genomförandet av denna förordning till kommissionen, på grundval av gemensamt överenskomna standarder, särskilt vad gäller syftet och reglerna om tillgångsbegränsningar. De skall även informera kommissionen om alla problem som uppkommer vid tillämpningen av denna förordning samt utbyta goda metoder med kommissionen och med varandra. |
Ändring 14
Artikel 5, punkt 3a (ny)
| 3a. Kommittén skall bistås av experter som utses av den arbetsgrupp som instiftats genom artikel 29 i direktiv 95/46/EG. |
Ändring 15
Artikel 5, punkt 3b (ny)
| 3b. När kommittén har slutfört de kompletterande tekniska specifikationer som avses i artikel 2.1 skall den arbetsgrupp som instiftats genom artikel 29 i direktiv 95/46/EG avge ett yttrande om dessa specifikationers överensstämmelse med standarder för uppgiftsskydd, vilket skall översändas till Europaparlamentet, rådet och kommissionen. |
Ändring 16
Artikel 5, punkt 3c (ny)
| 3c. Kommissionen skall översända sitt förslag till beslut om de kompletterande tekniska specifikationerna som avses i artikel 2.1 till Europaparlamentet, som inom tre månader kan anta en resolution genom vilken det motsätter sig detta förslag. |
Ändring 17
Artikel 5, punkt 3d (ny)
| 3d. Kommissionen skall informera Europaparlamentet om hur den avser att rätta sig efter Europaparlamentets resolution samt om skälen för detta. |
Ändring 18
Artikel 5, punkt 3e (ny)
| 3e. De kompletterande tekniska specifikationer som avses i artikel 2.1 skall hållas konfidentiella. |
Ändring 19
Artikel 6, punkt 2
2. Medlemsstaterna skall börja tillämpa denna förordning senast ett år efter antagandet av de åtgärder som avses i artikel 2. Detta påverkar dock inte giltigheten av redan utfärdade pass. | 2. För att denna förordning skall kunna tillämpas måste de nationella dataskyddsmyndigheterna intyga att de har de undersökande befogenheter och de resurser som krävs för att genomföra direktiv 95/46/EG när det gäller uppgifter som inhämtats i enlighet med detta. Medlemsstaterna skall börja tillämpa denna förordning senast 18 månader efter antagandet av de åtgärder som avses i artikel 2. Detta påverkar dock inte giltigheten av redan utfärdade pass. |
[1] Ännu ej offentliggjort i EUT.
--------------------------------------------------
Rådets yttrande
av den 7 juli 1997
om Polens konvergensprogram, 2004–2007
(2004/C 320/08)
EUROPEISKA UNIONENS RÅD HAR AVGETT FÖLJANDE YTTRANDE
med beaktande a
Yttrande från Europeiska ekonomiska och sociala kommittén om "XXXIII:e rapporten om konkurrenspolitiken – 2003"
(SEK(2004) 658 slutlig)
(2005/C 221/01)
Den 4 juni 2004 beslutade kommissionen att i enlighet med artikel 262 i EG-fördraget rådfråga Europeiska ekonomiska och sociala kommittén om "XXXIII:e rapporten om konkurrenspolitiken – 2003"
Facksektionen för inre marknaden, produktion och konsumtion, som svarat för kommitténs beredning av ärendet, antog sitt yttrande den 11 januari 2005. Föredragande var Franco Chiriaco.
Vid sin 414:e plenarsession den 9– 10 februari 2005 (sammanträdet den 9 februari) antog Europeiska ekonomiska och sociala kommittén följande yttrande med 75 röster för och 1 nedlagd röst:
1. Inledning
1.1 Syftet med 2003 års rapport om konkurrenspolitiken är att återspegla de viktiga förändringarna i kommissionens interna organisation och arbetsmetoder och att visa hur kommissionen bidrar till att samordna behovet av kontinuitet och behovet av nya grepp inom den ekonomiska styrningen i Europa.
1.2 EU:s konkurrenspolitik spelar en viktig roll för att nå de mål för konkurrenskraften som fastställts i Lissabonstrategin. Denna politik omfattar inte endast antitrust- och koncentrationsregler, utan även tillämpningen av en effektiv och strikt disciplin för statligt stöd.
1.3 För att möjliggöra en anslutning utan negativa återverkningar för de tio nya medlemsländerna har kommissionen utarbetat ett regelsystem på konkurrensområdet som är gemensamt för alla medlemsstater så att reglerna om statligt stöd tillämpas lika inom hela EU. Med detta vill man understryka att det är lika viktigt att ta itu med statliga ingripanden som snedvrider konkurrensen som att tillämpa konkurrensbestämmelser för företagen.
1.4 Under 2003 registrerades 815 nya fall av överträdelser mot konkurrenslagstiftningen. Dessutom inrättades en ny post: "Kontaktperson för konsumentfrågor". Posten inrättades för att garantera att en ständig dialog förs med Europas konsumenter. konsumenternas väl är konkurrenspolitikens huvuduppgift, men konsumenterna kommer inte till tals i tillräcklig utsträckning då enskilda ärenden behandlas eller policyfrågor diskuteras. Kontaktpersonen för konsumentfrågor har en roll som inte är begränsad till kontroll av koncentrationer, utan som även omfattar antitrustområdet – karteller och missbruk av dominerande ställning – liksom andra ärenden och policyfrågor på konkurrensområdet.
1.5 I oktober 2003 offentliggjorde kommissionen ett utkast till regler och riktlinjer för licensieringsavtal om tekniköverföring som EESK redan har avgivit ett yttrande om [1]. Mot bakgrund av den utveckling som har ägt rum under de senaste åren när det gäller denna typ av avtal har förslaget som mål att förenkla gemenskapens undantagsbestämmelser och bredda tillämpningsområdet. De nya bestämmelserna har följande fördelar:
- Gruppundantagsförordningen kommer endast att ha en svart lista: allt som inte uttryckligen utesluts från gruppundantaget är nu undantaget.
- Det görs en klar skillnad mellan licensiering mellan konkurrenter och licensiering mellan icke-konkurrenter.
- Man har redan planerat att anta ett "moderniseringspaket".
1.6 Kommissionen har för övrigt redan utnämnt en chefsekonom för konkurrensområdet, vars mandat inleddes den 1 september 2003, och samtidigt har man på ett positivt sätt stärkt förhörsombudets roll. Chefsekonomen för konkurrensområdet har tre huvuduppgifter:
- Rådgivning i ekonomiska och ekonometriska frågor vid tillämpningen av EU:s konkurrensregler. Detta kan även innefatta hjälp vid utvecklandet av allmänna policyinstrument.
- Allmän rådgivning redan på ett tidigt stadium i enskilda konkurrensärenden.
- Detaljerad rådgivning i de viktigaste konkurrensärendena som berör komplicerade ekonomiska frågor, särskilt sådana som kräver avancerade kvantitativa analyser.
1.7 Förhörsombudet får större befogenheter och oberoende att säkerställa rätten till försvar i vissa konkurrensförfaranden. Förhörsombudet är direkt knutet till kommissionsledamoten med ansvar för konkurrens och tar inte emot några instruktioner från GD Konkurrens. Ombudet kan alltid ingripa om det föreskrivna förfarandet står på spel. Han eller hon organiserar och genomför muntliga förhör objektivt och beslutar om tredje part skall höras. Dessutom kan nya handlingar endast läggas fram med tillstånd av förhörsombudet. Förhörsombudet har hela tiden kontakt med ansvarig kommissionsledamot.
2. Tillämpningen av reglerna om konkurrensbegränsande samverkan (antitrustbestämmelserna) – artiklarna 81 och 82 i fördraget 2.1 I oktober 2003 inledde kommissionen slutfasen i reformeringen av tillämpningen av antitrustreglerna (det så kallade moderniseringspaket), som syftar till att underlätta konkurrensmyndigheternas myndighetsutövande och att skapa de mekanismer för samarbete med nationella konkurrensmyndigheter och nationella domstolar som föreskrivs i förordning 1/2003.
2.2 I synnerhet innehåller moderniseringspaketet en ny tillämpningsförordning som behandlar formerna för att höra de berörda parterna samt en rad andra förfarandefrågor, t.ex. tillgång till handlingarna och behandling av sekretessbelagda uppgifter. De sex utkasten till tillkännagivanden behandlar bl.a. formerna för samarbetet inom det europeiska konkurrensnätverket och mellan kommissionen och de nationella domstolarna, effekterna på handeln mellan medlemsstaterna, behandlingen av klagomål och de riktlinjer som kommissionen tänker utfärda för att hjälpa företagen att bedöma nya eller olösta frågor. Hela detta moderniseringspaket behandlas i EESK:s yttrande om "Kommissionens förordning om kommissionens förfaranden enligt artiklarna 81 och 82 i EG-fördraget samt utkasten till kommissionens tillkännagivanden" [1].
2.3 Under 2003 har kommissionen utfärdat fem beslut riktade mot olagliga horisontella avtal: Det har gällt franskt nötkött, sorbater, elektriska och mekaniska kol- och grafitprodukter, organiska peroxider och industrirör av koppar. De böter som utdömdes uppgick till 400 miljoner euro, en summa som borde säkerställa en avskräckande verkan. I undersökningarna ingår inspektioner på företaget. Fullständig immunitet mot böter ges till det företag som först träder fram och som tillhandahåller tillräckliga bevis för att föranleda en undersökning. Däremot föreskrivs endast ett godkännande från kommissionen när avtalen mellan företagen inte begränsar konkurrensen på de berörda marknaderna och konsumenterna gynnas av samarbetet. Under 2003 uttalade sig också kommissionen om tre fall av överträdelser mot artikel 82, nämligen om
- de avgifter som Deutsche Telekom AG tog ut av konkurrerande företag för tillgången till den lokala infrastrukturen i det egna telekommunikationsnätet,
- Wanadoos prisstrategi för sina ADSL-tjänster,
- Ferrovie dello Stato S.p.A (FS), för missbruk av företagets dominerande ställning i fråga om tillgången till järnvägsinfrastrukturen för dragning och passagerartrafik.
3. Konkurrensutvecklingen i olika sektorer
3.1 Under 2003 gjordes stora framsteg (som dock kunde ha varit ännu större) i avregleringen av energisektorn (el och gas), och i juni antogs ett lagstiftningspaket som innebär att alla användare av el och gas i Europa fritt kan välja leverantör senast den 1 juli 2007. Genom dessa bestämmelser har man försökt balansera behovet av incitament till ny infrastruktur mot skapandet av en gemensam marknad.
3.2 Bland konsumenterna och företagen i olika EU-länder finns emellertid fortfarande en viss otillfredsställelse med prisnivån, som upplevs vara alltför hög, och tjänsternas effektivitet. Arbetsmarknadsparterna och konsumentorganisationerna, särskilt i de nya medlemsstaterna, framhåller i synnerhet kravet på att oberoendet för de nationella konkurrensmyndigheterna och för tillsynsmyndigheterna för offentliga tjänster skall respekteras i full omfattning.
3.2.1 När en adekvat och fullständig konkurrenslagstiftning väl har införts händer det ibland, särskilt i de nya medlemsstaterna, att myndigheterna för kontroll och reglering stöter på motstånd när de vill fullgöra sina uppdrag på ett självständigt sätt. Lagstiftningen på detta område har därför ibland inte kunnat försvara vare sig konsumenternas eller marknadernas intressen. Kommittén förordar ett mer funktionellt förhållande mellan konkurrenspolitiken och konsumentskyddspolitiken. En bättre organiserad och aktivare konsumentrörelse kommer också att kunna bidra till beslutsfattandet och tillhandahålla information om marknader och snedvridning av konkurrensen.
3.3 I fråga om posttjänster är det nya postdirektivet, som antogs 2002, ett led i fullbordandet av en inre marknad, framför allt genom en gradvis minskning av det monopoliserade området och genom avreglering av utgående gränsöverskridande post. Kommissionen skall för övrigt på grundval av en överenskommelse inom Europeiska rådet under 2006 genomföra en studie som underlag för en bedömning av konsekvenserna av de samhällsomfattande tjänsterna i de olika medlemsstaterna. På grundval av resultatet av denna studie antar sedan kommissionen ett förslag om ett fullständigt öppnande av marknaden för posttjänster från och med 2009 eller motsvarande åtgärd för att garantera de samhällsomfattande tjänsterna.
3.4 När det gäller elektronisk kommunikation löpte tidsfristen för att införliva den nya lagstiftningen om elektronisk kommunikation ut i juli 2004. I sin rapport i frågan har kommissionen i synnerhet framhållit följande principer: marknaderna bör analyseras mot bakgrund av principerna för konkurrens; bindande krav kan endast ställas på företag som har en dominerande marknadsställning; alla elektroniska kommunikationstjänster och kommunikationsnät behandlas på samma sätt ("teknisk neutralitet"). Utvecklingen av elektronisk kommunikation och den allmänna tillgången till sådan räcker inte för att säkerställa en återhämtning i den ekonomiska tillväxten. För en sådan återhämtning krävs ökad kunskap och kompetens hos alla dem som skall utnyttja informations- och kommunikationstekniken.
3.5 För lufttrafiksektorn beslutade kommissionen 2003 att inleda en omfattande branschdialog med berörda parter inom luftfartsnäringen, oberoende av enskilda ärenden. Syftet är att utarbeta en öppen policyvägledning för konkurrensfrågor i samband med allianser och koncentrationer mellan flygbolag.
3.5.1 Framsteg har gjorts när det gäller att fastställa och genomföra gemensamma riktlinjer för tillämpningen av antitrustreglerna i järnvägssektorn, i fråga om både godstransporter och persontrafik.
3.5.2 Branschdialogen har också utvecklats inom sektorerna för sjöfart, återförsäljning av bilar samt försäkringar, i syfte att se över eller anta lämpliga bestämmelser om gruppundantag.
3.5.3 Denna dialog bör också ta hänsyn till jämförbarheten i beskattningsformerna.
3.6 Media: Kommissionen anser att mångfalden i media är av grundläggande betydelse för utvecklingen av både Europeiska unionen och medlemsstaternas kulturella identitet, men att kontrollen av koncentrationer i mediebranschen i huvudsak skall utövas av medlemsstaterna. I mediebranschen tillämpas konkurrenspolitiska instrument endast på den underliggande marknaden och de ekonomiska effekterna av medieföretagens agerande och på kontroll av statligt stöd. Dessa instrument kan inte ersätta nationella kontroller av koncentrationer i mediebranschen eller åtgärder för att säkra mångfald inom media. Konkurrensreglerna tillämpas endast för att lösa problem till följd av att en dominerande ställning skapas eller förstärks på en viss marknad och för att kontrollera att konkurrenter inte utestängs från denna marknad.
3.6.1 Vi kan konstatera att kommissionens hållning här visserligen är formellt korrekt men att man inte har kunnat hindra eller upphäva dominerande marknadspositioner och därmed sammanhängande konkurrenshämmande metoder, framför allt i vissa länder. De berörda marknaderna är olika, och bland dem har TV-reklammarknaden en allt större betydelse när det gäller att bevara mångfalden, och den har hittills inte utretts på ett tillfredsställande sätt.
3.6.2 Kontrollerna har för övrigt förbisett de metoder som används av vissa företagskoncerner inom mediaområdet för att stärka den dominerande ställningen, framför allt defensiva åtgärder som syftar till att avvärja fientliga övertaganden genom skuldsättning av målbolaget eller genom införande av aktier med olika röststyrka som gör det lättare för aktieägare med minoritetsinnehav att kontrollera företaget.
3.6.3 Kommissionen bör således vara mycket vaksam i fråga om tillämpningen av normer och konkurrensmetoder.
3.7 Fria yrken: Kommissionen har offentliggjort en studie genomförd av Institut für Höhere Studien (IHS) i Wien. Studien visade att regleringen av de tjänster som erbjuds av de fria yrkena skiljer sig mycket mellan medlemsstaterna och även mellan olika yrken. I studien drogs slutsatsen att det fanns möjligheter att skapa ökat totalt välstånd i de länder där regleringen var mindre och friheten i yrkesutövningen var större.
3.7.1 Vid den konferens om regleringen av fria yrken som hölls i oktober 2003 i Bryssel samlades 260 företrädare för de berörda aktörerna för att diskutera regleringens och bestämmelsernas effekter på marknadsstrukturen och konsumentskyddet.
3.7.2 Vid samma tillfälle tillkännagav kommissionsledamot Mario Monti att han hade för avsikt att i början av 2004 offentliggöra en kommissionsrapport om konkurrensen i de fria yrkena. Denna rapport, som innehåller mycket viktiga riktlinjer och vägledande anvisningar, offentliggjordes den 9 februari 2004.
4. Reform av koncentrationskontrollen
4.1 Den 27 november 2003 uppnådde rådet politisk enighet om en omarbetad koncentrationsförordning, som i huvudsak införlivar de reformer som kommissionen föreslog i december 2002. Ändringarna innehåller andra åtgärder än lagstiftning, i syfte att effektivisera beslutsprocessen, förstärka den ekonomiska analysen och på ett effektivare sätt respektera företagens rätt till försvar. Bland annat har man utnämnt en chefsekonom för konkurrensområdet och inrättat en panel för att säkerställa helt oberoende slutsatser. EESK:s bedömning av företagsfusioner återfinns i kommitténs yttrande om "Förslag till Europaparlamentets och rådets direktiv om gränsöverskridande fusioner av aktiebolag och andra bolag med begränsat ansvar" [2].
4.2 Syftet med kommissionen reformförslag var att se till att substanstestet (dominanstestet) i koncentrationsförordningen faktiskt skulle täcka alla konkurrensbegränsande koncentrationer och samtidigt garantera fortsatt rättssäkerhet. Substanstestet jämfördes med testet "märkbar begränsning av konkurrensen", och slutligen enades man om följande nya lydelse för kriteriet: "En koncentration som påtagligt skulle hämma den effektiva konkurrensen inom den gemensamma marknaden eller en väsentlig del av den, i synnerhet till följd av att en dominerande ställning skapas eller förstärks, skall förklaras oförenlig med den gemensamma marknaden".
4.2.1 De nya bestämmelsernas formulering "i synnerhet till följd av att en dominerande ställning skapas eller förstärks" öppnar för en eventuell utvidgning av tillämpningsområdet för förbudet som inte är strikt kopplat till dominanskravet. Denna bestämmelse bör dock tolkas och tillämpas med beaktande av rådets och kommissionens gemensamma uttalande om artikel 2, där man hänvisar till skäl 25 i förordningen [3], enligt vilket begreppet "påtagligt hinder för effektiv konkurrens" bör "tolkas så att det, utöver begreppet 'dominerande ställning', endast sträcker sig till en koncentrations konkurrenshämmande effekter till följd av ett icke-samordnat beteende hos företag som inte skulle få någon dominerande ställning på den berörda marknaden". Därav följer att tillämpningsområdet även fortsättningsvis kommer att definieras i förhållande till dominansbegreppet.
4.3 Riktlinjer för bedömning av horisontella koncentrationer – sammanslagningar av faktiskt eller potentiellt konkurrerande företag. Sådana koncentrationer är endast olagliga om de förstärker företags marknadsinflytande på ett sätt som sannolikt får negativa konsekvenser för konsumenterna, särskilt i form av högre priser, produkter av sämre kvalitet eller minskad valfrihet. Detta gäller oavsett om de konkurrenshämmande effekterna följer av att en enda dominerande marknadsaktör skapas eller stärks eller av en oligopolsituation. Effekterna av en koncentration skall dessutom bedömas i reaktion till vad som annars skulle ha hänt på marknaden. Det innebär, t.ex. att ett uppköp av ett konkurshotat företag inte skulle motivera något ingripande från kommissionen.
4.4 Nya riktlinjer för bästa praxis: Som en del av reformpaketet 2002 genomfördes ett offentligt samråd som avslutades i februari 2003. Syftet var att ge berörda parter vägledning om det dagliga arbetet i EU:s förfaranden för kontroll av företagskoncentrationer.
5. Internationellt samarbete
5.1 Kommissionen har aktivt deltagit i det internationella konkurrensnätverkets (ICN) arbetsgrupp om kontroll av företagskoncentrationer som omfattar flera jurisdiktioner. Arbetsgruppen har bedrivit sin verksamhet i tre olika undergrupper:
- Anmälningar och förfaranden.
- Utredningstekniker.
- Analysramar.
5.1.1 Kommissionen deltar i alla tre undergrupperna. Det grundläggande målet är att främja ömsesidig förståelse mellan olika jurisdiktioner för att effektivisera koncentrationskontrollen.
5.1.2 ICN inrättades som ett virtuellt nätverk av olika konkurrensmyndigheter för att underlätta internationellt samarbete och utarbeta förslag för att sänka tillsynskostnaderna och harmonisera förfarandena och innehållet i regelverken.
5.1.3 Vid ICN:s andra konferens, som hölls i Merida, Mexiko, i juni 2003, framhölls särskilt behovet av att i konkurrensfrågor använda ett tydligt och lättillgängligt språk. Man underströk också den strategiska betydelse som främjandet av konkurrensen i de reglerade sektorerna har för att sänka tillsynskostnaderna och övervinna hinder för förståelsen mellan olika jurisdiktioner i frågan om koncentrationspolitiken.
6. Statligt stöd
6.1 Kontrollen av statligt stöd inriktar sig på de konkurrenseffekter som uppstår när medlemsstaterna beviljar stöd till företag. Målet är att se till att statliga ingripanden inte inverkar negativt på den inre marknadens funktion, liksom att främja konkurrens och konkurrenskraftiga marknader samt strukturella reformer. Man försöker särskilt se till att bevisligen gynnsamma effekter från avregleringen inte undergrävs av statliga stödåtgärder. Europeiska rådet i Stockholm: Medlemsstaterna måste generellt minska stödnivåerna samtidigt som stödet omdirigeras mot övergripande mål av gemenskapsintresse, till exempel en förstärkning av den ekonomiska och sociala sammanhållningen, sysselsättning, miljöskydd, främjande av forskning och utveckling av små och medelstora företag. Kommissionen har fastslagit att återkrav av stöd som olagligen beviljats av medlemsstaterna skall vara en prioritet.
6.1.1 I detta sammanhang finns det skäl att beklaga den bristande öppenheten i en rad medlemsstater gentemot anbudsgivare från andra medlemsstater när det gäller offentlig upphandling. Inom EU har den offentliga upphandlingen en årlig omsättning på mer än 1500 miljarder euro, och den praxis som finns i några medlemsstater att gynna de inhemska företagen hämmar konkurrensen och ökar beskattningen av konsumenterna.
6.2 Stöd till undsättning och omstrukturering av företag i svårigheter. Enligt de riktlinjer som löpte ut i oktober 2004 kunde stödet anses vara legitimt endast om det uppfyller stränga villkor. Dessa riktlinjer har setts över, och översynen har särskilt inriktats på följande:
- Att se till att undsättningsstöd begränsas till återbetalningsbart, tillfälligt och kortsiktigt finansiellt stöd som bara beviljas så länge det är nödvändigt för att genomföra en genomgripande omstruktureringsplan.
- Att koncentrera kontrollen av statligt stöd till stora företag som handlar inom hela EU.
- Att, särskilt för stora företag, förstärka principen att mottagaren av statligt stöd skall finansiera en stor del av omstruktureringskostnaderna utan något statligt stöd.
- Att principen om att stöd endast får beviljas en gång skall tillämpas.
6.3 Sektorsövergripande rambestämmelser för stora investeringsprojekt: Strikta regler för sektorer med strukturproblem. En förteckning över sådana sektorer skulle ha upprättats i slutet av 2003. På grund av de praktiska och tekniska svårigheterna med att sammanställa den har kommissionen beslutat att skjuta antagandet av förteckningen på framtiden. De befintliga övergångsreglerna för stora investeringsprojekt inom "känsliga" sektorer förlängs t.o.m. december 2006.
6.4 Stöd till forskning och utveckling i små och medelstora företag kan bidra till ekonomisk tillväxt, stärkt konkurrenskraft och ökad sysselsättning. För de små och medelstora företagen är stöden särskilt viktiga.
6.5 Miljöstöd, FoU-stöd, utbildningsstöd och skattestöd: I fråga om skattestöd granskades särskilt alternativa beskattningsmetoder, såsom kostnadsplusmetoden (den beskattningsbara inkomsten bestäms schablonmässigt och motsvarar en procentandel av summan av utgifter och driftskostnader). När det gäller sektorsstöd (jfr särskilt tillämpningen av tillfälliga skyddsordningar) behandlades följande sektorer: stålindustrin, telekommunikationer, kol, järnvägstransporter, kombinerade transporter, vägtransporter, lufttransporter och sjötransporter.
6.6 Jordbruk: Den 23 december antog kommissionen en ny förordning som innebär undantag för vissa typer av statligt stöd som medlemsstaterna inte längre behöver förhandsanmäla till kommissionen för godkännande. Den nya förordningen, som träder i kraft i slutet av 2006, gäller statligt stöd som beviljats små och medelstora företag inom jordbrukssektorn. Mot bakgrund av definitionen av små och medelstora företag (högst 250 anställda, 40 miljoner euro i omsättning eller 27 miljoner euro som tillgångar i balansräkningen) uppfyller nästan alla rörelser och företag inom jordbrukssektorn dessa krav. Kommissionen inför också en ny norm för öppenhet och insyn: en sammanställning över allt statligt stöd som beviljats av medlemsstaterna skall publiceras på Internet senast fem dagar innan utbetalningen av stöden påbörjas, för att säkerställa att alla berörda parter har tillgång till informationen.
7. Allmänna kommentarer
7.1 Efter att ha sammanfattat och delvis kommenterat kommissionens XXXIII:e rapport om konkurrenspolitiken (2003) finns det nu skäl att formulera några bedömningar av rapporten som helhet och vissa av de viktigaste aspekterna samt av framtidsutsikterna.
7.2 Förhållandet mellan konkurrenspolitiken och politiken för ekonomisk utveckling
7.2.1 EU:s konkurrenspolitik har blivit mer effektiv och öppen för ett positivt förhållande mellan företagen och konsumenterna tack vare införandet av nya tillämpningsförfaranden för antitrustbestämmelserna, översynen av koncentrationsförordningen och förändringar i kommissionens interna organisationsstruktur.
7.2.2 Tack vare konkurrenspolitiken har EU gjort avsevärda framsteg när det gäller avreglering, och återfört hela ekonomiska sektorer till marknadens funktion och dynamik samtidigt som man har arbetat konkret med inrättandet av en europeisk inre marknad. Konkurrenspolitiken är således central, och dess oberoende måste alltid bevaras.
7.2.3 Konkurrenspolitiken kan emellertid inte själv tillfredställa det för närvarande i hela EU djupt kända behovet av en ordentlig tillväxtåterhämtning och en långsiktig ekonomisk politik grundad på innovation och social dialog. De strukturella förändringar som har ägt rum inom produktion och handel i hela världen, med början i de förändringar som orsakats av ny teknik, ställer krav på kommissionen att initiera och samordna andra instrument inom ramen för den ekonomiska politiken för att kunna säkerställa och ge ny kraft åt den europeiska ekonomins konkurrenskraft och för att kunna stärka den ekonomiska och sociala sammanhållningen, öka sysselsättningen och miljöskyddet samt främja omfattande och krävande forsknings- och utvecklingsprogram. Kommissionens ståndpunkt i meddelandet "Att stödja strukturomvandlingarna: En industripolitik för ett utvidgat EU" och EESK:s yttrande i ärendet [4] ligger i linje med detta. Lissabondagordningen stakar ut den väg som måste följas. Genomförandet av den måste emellertid möjliggöras och påskyndas, såväl generellt som sektorsvis.
7.2.3.1 På sektorsnivå framhåller EESK behovet av att föra fram det nya helt integrerade arbetssätt som rådet (konkurrensfrågor) fastställde i november 2003 för att stärka den industriella konkurrenskraften och inom alla sektorer uppmuntra forskning, utveckling och innovation. Kommittén bekräftar därmed de ståndpunkter som framfördes i yttrandet av den 30 juni 2004 om "LeaderSHIP 2015 – Framtiden för varvs- och reparationsvarvsindustrin inom EU – Konkurrenskraft genom spetskompetens" [5].
7.3 Statsstöd till tjänster av allmänt intresse
7.3.1 Den reformprocess som syftar till att rationalisera och förenkla förfarandena för kontroll av statligt stöd har gjort stora framsteg i den riktning som utstakades av Europeiska rådet i Stockholm när det gäller att minska stödnivåerna samtidigt som stödet omdirigeras mot övergripande mål av gemenskapsintresse, inbegripet sammanhållningsmålen. I denna riktning går också olika åtgärder som kommissionen har vidtagit, t.ex. en viss utvidgning av tillämpningsområdet för FoU-stödet, riktlinjerna för licensieringsavtal om tekniköverföring, för omstruktureringsstöd till företag i svårigheter, för utbildningsstöd och för miljöskydd, samt de sektorsövergripande rambestämmelserna för stora investeringsprojekt.
7.3.2 I sin Altmark-dom från juli 2003 slog domstolen fast att statligt stöd i form av ekonomisk ersättning som beviljas vissa företag som fått i uppdrag att sköta tjänster av allmänt ekonomiskt intresse skall undantas, på vissa villkor. Det återstår dock vissa problem, framför allt när det gäller avvägningen mellan statsstöd och tjänster i allmänhetens intresse. De villkor som domstolen fastställt ställer krav på en förbättring av rättssäkerheten, framför allt när det gäller kostnadsberäkningen, ett fastställande av hur tjänsterna skall finansieras [4] och på en bättre beskrivning av kraven på de offentliga tjänster för vilka ersättning kan ges. I grönboken om tjänster av allmänt intresse från maj 2003 erkänns för övrigt behovet av att bedöma om de principer som reglerar tjänsterna av allmänt intresse så småningom behöver konsolideras i en övergripande gemenskapsram, liksom behovet av att fastställa en optimal reglering av sådana tjänster samt åtgärder för att öka rättssäkerheten för alla aktörer.
7.3.3 Kraven på de allmänna tjänsterna kommer, om de inte definieras och finansieras på ett korrekt sätt, att leda till att de företag som lyder under dessa krav drabbas av ökande förluster om konkurrenter dyker upp på de mest lönsamma verksamhetsområdena.
7.3.4 EESK framhåller följaktligen, och i linje med kommitténs yttrande [1] om kommissionens grönbok, behovet av en tydlig lagstiftning om tjänster i allmänhetens intresse i syfte att säkerställa effektiv och rättvis tillgång till tjänster av hög kvalitet som motsvarar användarnas krav. Dessutom rekommenderar kommittén att man, i synnerhet i samband med de sociala tjänsternas funktion och omorganiseringen av dem, främjar en så bred dialog som möjligt med arbetsmarknadsparterna och de icke-statliga organisationerna.
7.4 Fria yrken
7.4.1 Kommissionens grundliga analysarbete om regleringsläget för de fria yrkena i medlemsstaterna har varit till stor nytta eftersom det har gjort det möjligt att med stor effektivitet motivera behovet av att, om än med viss försiktighet, se över de restriktiva bestämmelserna på detta område och att göra de stora befintliga kulturella och kunskapsmässiga resurserna inom sektorn mer produktiva och konkurrenskraftiga. Detta innebär naturligtvis en stor fördel såväl för yrkesmässigt verksamma som för företag och konsumenter.
7.4.2 Det anses nu allmänt att även utbudet av professionella tjänster bör respektera konkurrensbestämmelserna, vilket också är den princip som flera gånger bekräftats av EG-domstolen. Det är visserligen helt korrekt att det ekonomiska kriteriet inte kan utgöra den enda parameter enligt vilken man bedömer det fria yrkenas tjänster, eftersom det inte rör sig om en enkel och repetitiv teknisk tillämpning, utan tjänster som kräver vissa kunskaper i förhållande till problemet, men det är också sant att tillhandahållandet av dessa tjänster utgör en ekonomisk verksamhet som kan producera större välfärd och ge ett viktigt bidrag till Lissabondagordningen om de utvecklas med respekt för konkurrensbestämmelserna.
7.4.2.1 Innehållet i kommissionsrapporten om "konkurrens inom sektorn för professionella tjänster" [6] är betydelsefullt i detta avseende. I rapporten understryker kommissionen å ena sidan den viktiga roll som de fria yrkena kan spela för att förbättra Europas ekonomiska konkurrenskraft, eftersom deras tjänster är av central betydelse för företag och familjer. Å andra sidan framläggs argument, grundade på empirisk forskning, om de negativa effekter som alltför många eller föråldrade restriktiva bestämmelser kan medföra för konsumenterna, exempelvis i fråga om prisreglering, reklam, tillgänglighet och exklusiva rättigheter samt företagsstruktur.
7.4.3 Det är således nödvändigt att genomföra och påskynda reformprocessen. EESK uppmanar i detta syfte kommissionen att respektera de tidigare gjorda åtagandet om att under 2005 offentliggöra en ny rapport om framstegen när det gäller att avskaffa restriktiva och omotiverade bestämmelser. Kommittén påminner för övrigt om att kommissionen i detta sammanhang också har åtagit sig att närmare granska de befintliga kopplingarna mellan regleringsnivån, de ekonomiska resultaten (pris och kvalitet) och konsumenternas tillfredsställelse.
7.4.4 Samtidigt vill kommittén framhäva betydelsen av EG-domstolens dom av den 9 oktober 2003 i målet Consorzio Industrie Fiammiferi, som gör det möjligt för de nationella myndigheterna att upphäva tillämpningen av en nationell lag som tvingar företag att agera i strid mot artikel 81 i EG-fördraget.
7.4.5 Slutligen finns det skäl att främja ett större och mer medvetet deltagande från de berörda aktörerna i reformprocessen.
7.5 Informationsmångfald och konkurrensregler
7.5.1 I sin XXXIII:e rapport om konkurrenspolitiken framhåller kommissionen att det är ett grundläggande mål i allmänhetens intresse för Europeiska unionen att upprätthålla och utveckla mångfalden i media och friheten att tillhandahålla och få information som avgörande värden för den demokratiska processen, men att kontrollen av koncentrationer i mediebranschen i huvudsak skall utövas av medlemsstaterna. Enligt kommissionen skall konkurrensreglerna tillämpas inom mediesektorn endast för att lösa problem till följd av att en dominerande ställning skapas eller förstärks på en viss marknad och för att kontrollera att konkurrenter inte utestängs från denna marknad. EESK menar att denna distinktion mellan EU:s och medlemsstaternas uppgifter dels är mycket vag, dels inte täcker följande viktiga problem:
- Det finns skäl att påminna om att det i de olika medlemsstaterna finns olika regleringar och tillvägagångssätt som kräver en harmonisering. Kommissionen inledde åtgärder i denna riktning 1989, och arbetade vidare 1997 med direktivet "Television utan gränser", som innehöll både målsättningar om ekonomisk effektivitet och respekt för den kulturella mångfalden, skydd av minoriteter, rätten till genmäle osv.
- Dessutom bör man inom medieområdet skilja mellan allmänna antitrustbestämmelser och specifik lagstiftning för skydd av mångfalden i informationsförmedlingen. Att konkurrensreglerna tillämpas är en grundläggande förutsättning, men det får inte leda till minskad mångfald. Till skillnad från ett konkurrenssystem där varje företags marknadskraft står i relation till initiativ och verksamhet inom konkurrerande företag, kräver främjandet och skyddet av mångfalden ett uttryckligt erkännande av medborgarnas rätt att effektivt utnyttja fria informationskällor och alternativ och potentiellt avvikande information, en rätt som skall skyddas på alla nivåer.
- Slutligen gör den successiva konvergensen i fråga om telekommunikationer, IT, radio och television samt förlagsverksamhet det svårt att fastställa vilka strukturella förändringar som äger rum på de olika marknaderna. Om man inte förstår denna process riskerar man samtidigt minskad effektivitet i konkurrensbestämmelserna och en försvagning av mångfaldsprincipen.
7.5.2 Den nya konstitutionen utvidgar avsevärt kommissionens mandat. Europeiska ekonomiska och sociala kommittén är övertygad om att kommissionen kommer att kunna verka med större kraft inom denna nya ram för att försvara och utveckla frihet och mångfald i tillhandahållandet av information.
Bryssel den 9 februari 2005
Europeiska ekonomiska och sociala kommitténs ordförande
Anne-Marie Sigmund
[1] EUT C 80, 30.3.2004.
[2] EUT C 117, 30.4.2004.
[3] Rådets förordning 139/2004 av den 20 januari 2004.
[4] EUT C 157, 28.6.2005.
[5] EUT C 302, 7.12.2004.
[6] KOM(2004) 83 slutlig, 9.2.2004.
--------------------------------------------------
P6_TA(2005)0061
Tillträde till naturgasöverföringsnät ***II
Europaparlamentets lagstiftningsresolution om rådets gemensamma ståndpunkt inför antagandet av Europaparlamentets och rådets förordning om villkor för tillträde till naturgasöverföringsnät (11652/2/2004 - C6-0188/2004 - 2003/0302(COD))
(Medbeslutandeförfarandet: andra behandlingen)
Europaparlamentet utfärdar denna resolution
- med beaktande av rådets gemensamma ståndpunkt (11652/2/2004 - C6-0188/2004),
- med beaktande av parlamentets ståndpunkt vid första behandlingen av ärendet [1], en behandling som avsåg kommissionens förslag till Europaparlamentet och rådet (KOM(2003)0741) [2],
- med beaktande av artikel 251.2 i EG-fördraget,
- med beaktande av artikel 62 i arbetsordningen,
- med beaktande av andrabehandlingsrekommendationen från utskottet för industrifrågor, forskning och energi (A6-0012/2005).
1. Europaparlamentet godkänner den gemensamma ståndpunkten såsom ändrad av parlamentet.
2. Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
[1] Antagna texter sammanträdet den 20.4.2004, P5_TA(2004)0301.
[2] Ännu ej offentliggjort i EUT.
--------------------------------------------------
P6_TA(2005)0128
Bestånden av tunga *
Europaparlamentets lagstiftningsresolution om förslaget till rådets förordning om återhämtningsåtgärder för bestånden av tunga i västra delen av Engelska kanalen och i Biscayabukten (KOM (2003)0819 - C5-0047/2004 - 2003/0327(CNS))
(Samrådsförfarandet)
Europaparlamentet utfärdar denna resolution
- med beaktande av kommissionens förslag till rådet (KOM(2003)0819) [1],
- med beaktande av a/rtikel 37 i EG-fördraget, i enlighet med vilken rådet har hört parlamentet (C5-0047/2004),
- med beaktande av artikel 51 i arbetsordningen,
- med beaktande av betänkandet från fiskeriutskottet (A6-0050/2005).
1. Europaparlamentet godkänner kommissionens förslag såsom ändrat av parlamentet.
2. Europaparlamentet uppmanar kommissionen att ändra sitt förslag i överensstämmelse härmed i enlighet med artikel 250.2 i EG-fördraget.
3. Rådet uppmanas att underrätta Europaparlamentet om rådet har för avsikt att avvika från den text som parlamentet har godkänt.
4. Rådet uppmanas att på nytt höra Europaparlamentet om rådet har för avsikt att väsentligt ändra kommissionens förslag.
5. Europaparlamentet uppdrar åt talmannen att delge rådet och kommissionen parlamentets ståndpunkt.
KOMMISSIONENS FÖRSLAG | PARLAMENTETS ÄNDRINGAR |
Ändring 1
Titel
Förslag till rådets förordning om återhämtningsåtgärder för bestånden av tunga i västra delen av Engelska kanalen och i Biscayabukten | Förslag till rådets förordning om en förvaltningsplan för bestånden av tunga i västra delen av Engelska kanalen och i Biscayabukten (Ändringen innebär att ordet "återhämtning" byts ut mot ordet "förvaltning" i hela texten, förutom i artikel 3.3.) |
Ändring 2
Skäl 1
(1) Av nyligen framlagda vetenskapliga rekommendationer från Internationella havsforskningsrådet (ICES) framgår det att bestånden av tunga i ICES-område VIIe, VIIIa och VIIIb har utsatts för en fiskedödlighet som har minskat mängden lekmogen fisk i havet till en nivå där bestånden inte längre fylls på genom fortplantning, och att dessa bestånd därför hotas av kollaps. | utgår |
Ändring 3
Skäl 2
(2) Åtgärder bör vidtas för att fastställa fleråriga planer för dessa bestånds återhämtning enligt artikel 5 i rådets förordning (EG) nr 2371/2002 av den 20 december 2002 om bevarande och hållbart utnyttjande av fiskeresurserna inom ramen för den gemensamma fiskeripolitiken. | (2) Åtgärder för förvaltning av dessa bestånd bör vidtas i enlighet med artikel 6 i rådets förordning (EG) nr 2371/2002 av den 20 december 2002 om bevarande och hållbart utnyttjande av fiskeresurserna inom ramen för den gemensamma fiskeripolitiken. |
Ändring 4
Skäl 3
(3) Målet för dessa planer skall vara att se till att dessa bestånd åter befinner sig inom säkra biologiska gränser inom fem till tio år. | (3) Målet för dessa planer skall vara att se till att dessa bestånd förblir inom säkra biologiska gränser. |
Ändring 5
Skäl 3a (nytt)
| (3a) Den nya gemensamma fiskeripolitiken har som mål att möjliggöra ett hållbart utnyttjande av de levande akvatiska resurserna genom ett balanserat hänsynstagande till miljömässiga, sociala och ekonomiska faktorer. |
Ändring 6
Skäl 3b (nytt)
| (3b) Kommissionen och medlemsstaterna skall se till att de regionala rådgivande kommittéerna och andra berörda parter medverkar fullt ut i genomförandet av dessa förvaltningsplaner. |
Ändring 7
Skäl 5
(5) De berörda beståndens storlek i absoluta tal, så som de beräknas av STECF och ICES, är alltför osäkra för att användas som mål för återhämtningen, och därför bör målen uttryckas i termer av fiskedödlighet. | utgår |
Ändring 8
Skäl 6
(6) För att detta mål skall kunna uppnås måste fiskedödligheten kontrolleras på ett sätt som gör det högst sannolikt att den minskar år efter år. | utgår |
Ändring 9
Skäl 8
(8) När återhämtningen har uppnåtts bör rådet på kommissionens förslag fatta beslut om uppföljningsåtgärder i enlighet med artikel 6 i förordning (EG) nr 2371/2002. | utgår |
Ändring 10
Artikel 2
Återhämtningsplanens mål är att bestånden av tunga skall öka så att de åter befinner sig inom säkra biologiska gränser. | Förvaltningsplanens mål är att bestånden av tunga skall underhållas så att de åter befinner sig inom säkra biologiska gränser. |
Ändring 12
Artikel 3, punkt 2
2. Om kommissionen på grundval av den årliga utvärderingen finner att något av de berörda bestånden av tunga har uppnått de mål som fastställs i artikel 2 skall rådet med kvalificerad majoritet och på kommissionens förslag fatta beslut om att för det beståndet byta ut den återhämtningsplan som föreskrivs i den här förordningen mot en förvaltningsplan enligt artikel 6 i förordning 2371/2002. | utgår |
Ändring 13
Artikel 3, punkt 3
3. Om kommissionen på grundval av den årliga utvärderingen finner att något av de berörda bestånden av tunga inte visar tillräckliga tecken på återhämtning skall rådet med kvalificerad majoritet och på kommissionens förslag fatta beslut om ytterligare och/eller alternativa åtgärder för att säkerställa de berörda beståndens återhämtning. | 3. Om kommissionen på grundval av den årliga utvärderingen finner att något av de berörda bestånden av tunga hotas av kollaps skall rådet med kvalificerad majoritet och på kommissionens förslag fatta beslut om ytterligare och/eller alternativa åtgärder för att säkerställa de berörda beståndens återhämtning. |
Ändring 14
Artikel 5, punkt 1
1. Om STECF i ljuset av den senaste rapporten från ICES beräknar att fiskedödligheten för ett av de berörda bestånden av tunga ligger över 0,14 per år skall TAC för det beståndet inte överskrida en fångstnivå som enligt en vetenskaplig utvärdering som görs av STECF i ljuset av den senaste rapporten från ICES kommer att resultera i en minskning med a)20 % i fiskedödligheten under det år den tillämpas, jämfört med den fiskedödlighet som beräknats för det föregående året med avseende på beståndet av tunga i område VIIe,b)35 % i fiskedödligheten under det år den tillämpas, jämfört med den fiskedödlighet som beräknats för det föregående året med avseende på beståndet av tunga i område VIIIa och VIIIb. | 1. TAC skall inte överskrida en fångstnivå som, enligt en vetenskaplig utvärdering som görs av STECF i ljuset av den senaste rapporten från ICES, kommer att resultera i en ökning med 15% av mängden lekmogen fisk i havet vid utgången av året för dess tillämpning, i förhållande till de mängder som bedöms ha funnits i havet i början av det aktuella året. |
Ändring 15
Artikel 5, punkt 2
2. Om STECF i ljuset av den senaste rapporten från ICES beräknar att fiskedödligheten för ett av de berörda bestånden av tunga är lika med eller mindre än 0,14 per år skall TAC för det beståndet fastställas på en fångstnivå som enligt en vetenskaplig utvärdering som görs av STECF i ljuset av den senaste rapporten från ICES kommer att resultera i en fiskedödlighet på a)0,11 per år under det år den tillämpas när det gäller beståndet av tunga i område VIIe,b)0,09 per år under det år den tillämpas när det gäller beståndet av tunga i område VIIIa och VIIIb. | 2. Rådet skall inte anta någon TAC för vilken STECF i ljuset av den senaste rapporten från ICES beräknar att den under året för dess tillämpning kommer att leda till en fiskedödlighet som överskrider följande värden: Tunga i Biscayabukten: 0,36 Tunga i västra delen av Engelska kanalen: nivån skall fastställas på grundval av ett senare yttrande från ICES efter införlivandet av uppgiftsserier från vissa länder som hittills inte beaktats. |
Ändring 16
Artikel 6
1. Under det första tillämpningsåret för den här förordningen skall följande bestämmelser gälla: a)Om tillämpningen av artikel 5 leder till en TAC som överskrider det föregående årets TAC med mer än 25 %, skall rådet anta en TAC som inte får vara mer än 25% högre än det årets TAC.b)Om tillämpningen av artikel 5 leder till en TAC som understiger det föregående årets TAC med mer än 25% skall rådet anta en TAC som inte får vara mer än 25% lägre än det årets TAC. | |
2. Från och med det andra tillämpningsåret för den här förordningen skall följande bestämmelser gälla: a)Om tillämpningen av artikel 5 leder till en TAC som överskrider det föregående årets TAC med mer än 15 %, skall rådet anta en TAC som inte får vara mer än 15% högre än det årets TAC.b)Om tillämpningen av artikel 5 leder till en TAC som understiger det föregående årets TAC med mer än 15% skall rådet anta en TAC som inte får vara mer än 15% lägre än det årets TAC. | 2. Från och med det första tillämpningsåret för den här förordningen skall följande bestämmelser gälla: a)Om tillämpningen av artikel 5 leder till en TAC som överskrider det föregående årets TAC med mer än 15 %, skall rådet anta en TAC som inte får vara mer än 15% högre än det årets TAC.b)Om tillämpningen av artikel 5 leder till en TAC som understiger det föregående årets TAC med mer än 15% skall rådet anta en TAC som inte får vara mer än 15% lägre än det årets TAC. |
Ändring 17
Kapitel III
| Detta kapitel utgår. |
Ändring 18
Artikel 16
Genom undantag från artikel 5.2 i kommissionens förordning (EEG) nr 2807/83 av den 22 september 1983 om närmare bestämmelser för registrering av uppgifter om medlemsstaternas fångster av fisk skall den tillåtna toleransmarginalen vid uppskattning av de kvantiteter i kilogram fångst som förvaras ombord vara 5 % av uppgiften i loggboken. | Genom undantag från artikel 5.2 i kommissionens förordning (EEG) nr 2807/83 av den 22 september 1983 om närmare bestämmelser för registrering av uppgifter om medlemsstaternas fångster av fisk skall den tillåtna toleransmarginalen vid uppskattning av de kvantiteter i kilogram färskvikt som förvaras ombord vara 8 % av uppgiften i loggboken. Om ingen omräkningsfaktor fastställts i gemenskapslagstiftningen skall den omräkningsfaktor gälla som har antagits av den medlemsstat vars flagg fartyget för. |
Ändring 19
Artikel 17
De behöriga myndigheterna i en medlemsstat skall se till att alla kvantiteter tunga över 50 kg som fångats i något av de områden som anges i artikel 1 före försäljning vägs med en våg av den typ som används vid fiskauktioner. | De behöriga myndigheterna i en medlemsstat skall se till att alla kvantiteter tunga över 100 kg som fångats i något av de områden som anges i artikel 1 före försäljning vägs med en våg av den typ som används vid fiskauktioner. |
Ändring 20
Artikel 19, punkt 1
1. De behöriga myndigheterna i en medlemsstat får begära att en kvantitet tunga över 50 kg, som har fångats inom något av de geografiska områden som anges i artikel 1 och som först landats i den medlemsstaten, vägs innan den transporteras vidare från den hamn där den först landats. | 1. De behöriga myndigheterna i en medlemsstat får begära att en kvantitet tunga över 100 kg, som har fångats inom något av de geografiska områden som anges i artikel 1 och som först landats i den medlemsstaten, vägs innan den transporteras vidare från den hamn där den först landats. |
Ändring 21
Artikel 19, punkt 2
2. Genom undantag från artikel 13 i förordning (EEG) nr 2847/93 skall kvantiteter över 50 kg av tunga som transporteras någon annanstans än landnings- eller importplats åtföljas av en kopia av en av de deklarationer som anges i artikel 8.1 i förordning (EEG) nr 2847/93 avseende den transporterade kvantiteten tunga. Undantag enligt artikel 13.4 b i rådets förordning (EEG) nr 2847/93 skall inte tillämpas. | 2. Genom undantag från artikel 13 i förordning (EEG) nr 2847/93 skall kvantiteter över 100 kg av tunga som transporteras någon annanstans än landnings- eller importplats åtföljas av en kopia av en av de deklarationer som anges i artikel 8.1 i förordning (EEG) nr 2847/93 avseende den transporterade kvantiteten tunga. Undantag enligt artikel 13.4 b i rådets förordning (EEG) nr 2847/93 skall inte tillämpas. |
Ändring 22
Regionkommitténs yttrande om "En period för eftertanke: strukturen, ämnena och ramen för en utvärdering av debatten om Europeiska unionen"
(2006/C 81/09)
REGIONKOMMITTÉN HAR AVGETT DETTA YTTRANDE
Europaparlamentets beslut av den 6 september 2005 att i enlighet med artikel 265 fjärde stycket i EG-fördraget rådfråga Regionkommittén i ärendet,
Regionkommitténs ordförandes beslut att i enlighet med artikel 40.2 i arbetsordningen utse Franz Schausberger, delstaten Salzburgs företrädare i Regionkommittén (AT–PPE), och Graham Tope, Greater London Authority (UK–ALDE), till huvudföredragande för yttrandet i detta ärende,
Fördraget om upprättande av en konstitution för Europa som undertecknades av stats- och regeringscheferna i Rom den 29 oktober 2004 (CIG 87/04 rev. 1, CIG 87/04 add. 1 rev. 1 och add. 2 rev. 1),
Regionkommitténs yttrande av den 17 november 2004 om Fördraget om upprättande av en konstitution för Europa (CdR 354/2003 fin [1]),
ReK:s rapport av den 6 november 2001 om "Närhetsfrågorna" (CdR 436/2000 fin).
Vid sin 61:a plenarsession den 12– 13 oktober 2005 (sammanträdet den 13 oktober) antog Regionkommittén följande yttrande:
Regionkommitténs synpunkter och rekommendationer
a) Bakgrund
1. För att säkra fred, frihet och välstånd behövs det enligt Regionkommittén ett politiskt starkt och demokratiskt EU, ett kraftfullt europeiskt ledarskap och ett nära samarbete mellan EU-institutionerna i syfte att återlansera det europeiska projektet.
2. Kommittén hyser farhågor för att en alltför lång period för eftertanke kan skada bilden av EU, och uppmanar alla EU-institutioner att arbeta för att återuppta och återlansera den djupare innebörden i det ideal och den plan som ligger bakom det europeiska integrationsprojektet.
3. ReK anser emellertid att det är lämpligt att se reflexionsperioden som ett tillfälle att analysera medborgarnas ståndpunkter beträffande Europeiska unionen, och som en möjlighet att konsolidera EU:s grundläggande mål, värden och principer, t.ex. solidaritet, effektivitet, insyn och samarbete, på grundval av medborgarnas stöd.
4. Kommittén vill i detta sammanhang påminna om betydelsen av de grundläggande rättigheterna inom unionen i enlighet med den stadga som införlivats i det konstitutionella fördraget.
5. ReK anser att Europeiska unionen måste ta resultaten i den franska och den nederländska folkomröstningen på allvar och visa att den gör det. Att fortsätta processen för ratificering av det konstitutionella fördraget utan att ändra den ursprungliga tidsplanen och utan allvarliga diskussioner på europeisk nivå skulle enligt kommitténs åsikt vara detsamma som att ge Europas medborgare en negativ signal och att inbjuda till ytterligare avslag i medlemsstaterna.
6. Kommittén konstaterar dock att skälen till dessa avslag är många och varierade och i vissa fall kanske inte har med själva fördraget att göra. Kommittén anser därför att man i första hand bör koncentrera sig på diskussionens kontext och eftersträva enighet beträffande budgetplanen. Vi vill dock erinra om att mer än hälften av medlemsstaterna redan har ratificerat fördraget på det sätt de själva valt, och besluten i dessa medlemsstater måste väga lika tungt som de negativa folkomröstningsresultaten.
7. Kommittén bekräftar sitt engagemang för det konstitutionella fördraget och dess landvinningar, som innebär en garanti för bättre styresformer i EU tack vare de avsevärda förbättringarna som föreslås, jämfört med de gällande fördragen, i fråga om funktionssätt, enkelhet och insyn i EU.
8. Vi anser att institutionerna i den mer omfattande debatten om Europeiska unionens framtid bör fokusera på de aktuella och potentiella fördelar som medlemskap och medborgarskap i praktiken ger medborgarna.
9. I syfte att återskapa de europeiska medborgarnas förtroende för EU-projektet uppmanar vi EU-institutionerna att
- fatta beslut som är aktuella på de områden där EU-medborgarna tillförs ett verkligt mervärde,
- utforma sin verksamhet på ett mycket mer decentraliserat sätt, med respekt och incitament för subsidiaritetsprincipen,
- aktivt visa att en politisk union inte kommer att undergräva Europas kulturella och språkliga mångfald,
- visa att EU kommer att ge EU-medborgarna möjlighet att utveckla sina professionella och personliga erfarenheter på EU-nivå,
- upprätta en ömsesidig dialog med Europas medborgare,
- utveckla en kultur av ökad öppenhet, framför allt genom att göra rådets arbete mer tillgängligt, så att medborgarna lättare kan förstå EU:s beslutsprocess.
10. Kommittén anser att man bör fullfölja arbetet med att främja tillämpningen av subsidiaritetsprincipen på samtliga områden och utnyttja de fördelar som den ökade närheten till de lokala och regionala myndigheterna innebär för medborgarna.
11. Kommittén uppmanar medlemsstaterna att fördjupa den politiska integrationen i EU, något som utgör en grundläggande förutsättning för att skapa en utvidgad union, samt att ange syfte, potentiella geografiska gränser och långsiktiga mål för EU:s integrationsprocess. EU-medlemskap skall innebära respekt för det lokala och regionala självstyret inom varje stats konstitutionella ramar.
12. Vi uppmanar politiker på såväl medlemsstatsnivå som regional och lokal nivå att ta ansvar för sina handlingar inom de egna ansvarsområdena och att avhålla sig från den utbredda vanan att använda "Bryssel" som syndabock. Vi understryker att Europeiska unionen kan lyckas endast om politikerna på europeisk, nationell, regional och lokal nivå på ett ansvarsfullt sätt delar på åliggandena och erkänner att institutionell respekt är av avgörande betydelse för framgång och en förutsättning för goda styresformer.
b) Debattens struktur
13. Regionkommittén anser att EU-institutionerna måste börja diskutera med de människor och samhällen som de företräder, och att de bör ha samma öppna inställning som rådde i konventet, där fördraget utarbetades av företrädare för nationella parlament, politiska partier, lokala och regionala myndigheter, det civila samhället och arbetsmarknadens parter. I samband med denna diskussion måste medborgarna få klart för sig det politiska, ekonomiska och sociala mervärde som en europeisk union kan ge.
14. Kommittén anser att ReK i sin egenskap av institutionell företrädare för de lokala och regionala myndigheterna i Europeiska unionen måste spela en aktiv roll i de politiska och institutionella initiativen under den reflexionsperiod som stats- och regeringscheferna har inlett. Kommittén föreslår därför en färdplan [2] för att inleda en verklig decentraliserad diskussion i egentlig mening.
15. ReK uppmanar de lokala och regionala myndigheterna att skapa engagemang och informera sina lokalsamhällen om de frågor som är av betydelse för dessa i debatten om Europeiska unionens framtid. De bör på ett bättre sätt förklara processerna i den europeiska integrationen och de praktiska resultaten av denna genom en decentraliserad informationspolicy med regional och lokal bas. Kommittén anser att man inte kan nå ut till den breda allmänheten om debatten förs endast på europeisk nivå. Därför krävs strukturerade debatter med gränsöverskridande inslag på nationell, regional och lokal nivå, med deltagande av kommitténs ledamöter och med stöd av EU-institutionerna.
16. Kommittén vill för övrigt understryka att ReK präglas av arbetssättet nedifrån och upp, och åtar sig att genom sina ledamöter vända sig till och ta upp idéer från organ på regional och lokal nivå när det gäller gemenskapens politik och institutioner samt att överföra budskapet till EU-institutionerna, både vad avser politisk analys och innovativa förslag.
17. ReK rekommenderar att dialogen med medborgarna inte begränsas till enstaka kampanjer eller fokuseras på detaljer i institutionernas verksamhet. Därför uppmanas EU att fokusera på informationsförmedling som har direkt praktisk nytta för medborgarna och hjälper dem att utnyttja de möjligheter som EU erbjuder dem.
18. Kommittén uppmanar EU-institutionerna, medlemsstaterna och de regionala och lokala myndigheterna att skapa nya och kreativa metoder för interaktion med medborgarna på gräsrotsnivå och att i diskussionerna använda moderna elektroniska medier (t.ex. "Europa lyssnar" i Österrike och "Nationellt forum om Europa" i Irland) samt att se till att budskapet förmedlas på medborgarnas modersmål och inte bara på vissa utvalda EU-språk. Det vilar dessutom ett ansvar på institutionerna och medlemsstaterna att bemöta felaktiga fakta om EU som medborgarna kan konfronteras med, framför allt i media.
19. Kommittén konstaterar att lokala och regionala massmedia, och särskilt den lokala pressen, spelar en mycket viktig roll i detta sammanhang, inte minst för att de kan kommunicera direkt med medborgarna med enkla ord på medborgarnas eget språk.
c) Ämnen för reflexion
Allmänna ramar
20. Regionkommittén anser att bestämmelserna i det konstitutionella fördraget om EU:s territoriella dimension och de lokala och regionala myndigheternas medverkan, både institutionellt via ReK och mer generellt, utgör en viktig och positiv utveckling.
21. Kommittén uppmanar EU-institutionerna att hjälpa till att utveckla en verklig "subsidiaritetskultur" i EU, medlemsstaterna och inom de lokala och regionala myndigheterna och att omedelbart börja tillämpa den subsidiaritetsprincip och den proportionalitetsprincip som stadgas i det konstitutionella fördraget. Därigenom kan man på ett enkelt och effektivt sätt kan visa medborgarna att EU endast agerar på de områden där det finns ett tydligt mervärde samt att detta sker i enlighet med principen om bättre lagstiftning.
22. Kommittén skulle vilja att "närhetsbegreppet" tillämpas i EU:s strategier och lagstiftning, eftersom detta tydligt skulle visa en vilja att införa öppnare förfaranden som en omedelbar reaktion på medborgarnas farhågor. I detta sammanhang skulle införandet av ett nytt rättsligt instrument som underlättar mellanregionalt och gränsöverskridande samarbete, inklusive samarbete i ekonomiska och sociala frågor, bland annat kunna betraktas som ett tydligt tecken på ett Europa närmare medborgarna.
23. Dessa komponenter borde ingå i det konstitutionella fördraget, men kommittén vill understryka att många av de åtgärder och skyldigheter som sammanhänger med dessa bestämmelser omedelbart skulle kunna integreras i gemenskapens verksamhet, t.ex. att utvidga konsekvensbedömningarna till att omfatta de ekonomiska och administrativa konsekvenserna av ny EU-lagstiftning för de lokala och regionala myndigheterna.
24. ReK har särskilt välkomnat följande punkter i fördraget som exempel på goda styresformer och skulle vilja försäkra sig om att man under reflexionsperioden verkligen ser till att de kan bibehållas och genomföras:
- Erkännande av de lokala och regionala myndigheternas roll i EU:s styresformer.
- Förbättrat samråd innan lagstiftningsförslag offentliggörs.
- Beaktande av de ekonomiska och administrativa bördor som läggs på de lokala och regionala myndigheterna.
- Breddad definition av subsidiaritetsprincipen: de lokala och regionala myndigheterna skall omfattas.
- Erkännande av att den kulturella och språkliga mångfalden är en källa till välstånd som måste bevaras, samtidigt som de grundläggande principerna om samarbete och integration måste respekteras.
- Förstärkning av Regionkommitténs roll; framför allt skall ReK ges rätt att väcka talan inför EG-domstolen när det gäller kommitténs egna befogenheter och vid brott mot subsidiaritetsprincipen.
- Hänvisning till representativa sammanslutningar (t.ex. lokala och regionala myndigheter).
Aktuella diskussionsfrågor
25. Regionkommittén anser att det är oerhört viktigt att EU har tillräckliga resurser för att genomföra de uppgifter som unionen åläggs. Kommittén upprepar sitt stöd till Europeiska kommissionens förslag till budgetplan för åren 2007–2013.
26. Kommittén anser att det nu är läge att börja diskutera grundvalarna för finansieringen av EU-budgeten på lång sikt och att stärka Europaparlamentets demokratiska kontroll över budgeten.
27. ReK påminner medlemsstaterna om att sammanhållningspolitiken är ett område där EU sedan lång tid tillbaka har uppvisat ett verkligt mervärde, samt att sammanhållningspolitikens synlighet gör det möjligt för medborgarna att i sin vardag uppskatta EU:s konkreta och positiva insatser och att den utgör grunden för europeisk solidaritet och därmed skiljer den europeiska sociala modellen från andra exempel på transnationell integration.
28. ReK upprepar sitt stöd till partnerskapet för tillväxt och sysselsättning (Lissabonstrategin) som en god avvägning mellan ekonomiska målsättningar, hållbar utveckling och den europeiska samhällsmodellens modernisering och framåtskridande.
29. Om EU:s konkurrenskraft skall kunna stärkas måste man enligt ReK:s uppfattning även hjälpa EU-medborgarna att utveckla sina talanger och sin kreativitet över de nationella gränserna. Kommittén är övertygad om att värdet av ett EU med kulturell mångfald kommer att bli mycket mer påtagligt för européerna när de börjar uppleva att deras liv ingår i ett europeiskt sammanhang. För att konkurrenskraften skall stärkas och medborgarna bli delaktiga i Europaprojektet, är det därför nödvändigt att EU även fortsättningsvis underlättar den fria rörligheten för personer och främjar större rörlighet inom EU.
30. ReK bekräftar sitt stöd till EU:s strategi för hållbar utveckling och betonar särskilt att åtgärder och EU-stöd på miljöskyddsområdet kan fungera som motor för ytterligare åtgärder på nationell, regional och lokal nivå.
31. Kommittén erinrar om det europeiska medborgarskapets unika beskaffenhet. Utan att ersätta det nationella medborgarskapet utgör det ett inslag i en europeisk identitet.
32. Kommittén efterlyser mycket större investeringar och samarbete när det gäller utbildning (inklusive möjligheter till livslångt lärande för alla medborgare), forskning och innovation på EU-nivå, eftersom detta är bästa sättet att skapa fler och bättre jobb för Europas medborgare och stärka den europeiska konkurrenskraften inom världsekonomin.
33. ReK är övertygad om att de nationella, regionala och lokala myndigheterna bör involveras i utbildningssatsningarna om man på ett bättre sätt vill förklara vad Europa och EU-politiken innebär. Detta kan ske t.ex. genom att införa specialkurser i skolorna och en europeisk dimension i läroplaner, postgymnasial utbildning och fortbildning för lärare.
34. Regionkommittén är dessutom övertygad om att det är nödvändigt att sprida en EU-positiv kultur bland offentliga tjänstemän på regional och lokal nivå som i sitt dagliga arbete konfronteras med lagar och bestämmelser.
d) Utvärdering
35. Regionkommittén uppmanar EU-institutionerna och medlemsstaterna att lyssna på medborgarna när man utvärderar diskussionsresultaten under reflexionsperioden.
36. Kommittén är medveten om att man under reflexionsperioden kan komma att diskutera olika scenarier, men vänder sig emot att man överger det konstitutionella fördraget till förmån för Nicefördraget. Vi efterlyser ett samförstånd om en ratificering år 2009.
37. Regionkommittén vill aktivt delta i nylanseringen av den konstitutionella processen och stöder Europaparlamentets strävan att uppnå ett framgångsrikt resultat.
Bryssel den 13 oktober 2005
Regionkommitténs
ordförande
Peter Straub
[1] EUT C 71, 22.3.2005, s. 1.
[2] Se bilaga.
--------------------------------------------------
[pic] | EUROPEISKA GEMENSKAPERNAS KOMMISSION |
Bryssel den 23.11.2005
KOM(2005) 585 slutlig
MEDDELANDE FRÅN KOMMISSIONEN
Tredje lagstiftningspaketet om sjösäkerheten i Europeiska unionen
{SEK(2005) 1496}
MEDDELANDE FRÅN KOMMISSIONEN
Tredje lagstiftningspaketet om sjösäkerheten i Europeiska unionen (Text av betydelse för EES)
Prestigeolyckan i november 2002 utlöste starka känslor som utmynnade i en våg av solidaritet genom hela Europa. Unionens institutioner och högsta organ uttryckte sin fasta avsikt att fortsätta och intensifiera det arbete för att höja sjösäkerheten som inleddes efter Erikaolyckan i december 1999.
Under mötet i Köpenhamn den 12 och 13 december 2002, alltså strax efter Prestigeolyckan, erkände Europeiska rådet ”de beslutsamma insatserna inom Europeiska gemenskapen och Internationella sjöfartsorganisationen (IMO) sedan olyckan med Erika för att öka sjösäkerheten och förhindra föroreningar”, och erinrade om unionens fasta avsikt ”att vidta alla åtgärder som är nödvändiga för att undvika att liknande katastrofer upprepas”.
Även Europaparlamentet visade beslutsamhet, och utfärdade den 27 april 2004 en resolution om ökad sjösäkerhet, som byggde på det arbete som utförts av det tillfälliga utskottet för ökad sjösäkerhet (MARE)[1]. Parlamentet bekräftade i resolutionen behovet av att fortsätta sjösäkerhetsarbetet.
Europaparlamentet begär i resolutionen ett antal konkreta åtgärder avsedda att höja sjösäkerheten på internationell nivå och på unionsnivå:
- Inrättandet av ett europeiskt område för sjösäkerhet, grundat på förbud mot fartyg som inte uppfyller normerna, och en ansvarsordning som omfattar hela sjötransportkedjan samt offentliga myndigheter med ansvar för sjösäkerhetsfrågor.
- Utformningen av en beredskapsplan för effektivare insatser vid olyckor som kan begränsa konsekvenserna, inbegripet ett bättre utnyttjande av skyddshamnar.
- En bättre ersättning vid olyckor, bl.a. genom utökad försäkringsplikt och skärpta skadeståndsbestämmelser.
- Stärkt samarbete vid olycksutredningar, och större krav på utredningarnas oberoende.
- Skärpt fartygskontroll, främst genom en strikt tillämpning av hamnstatskontrollen och en bättre kontroll av klassificeringssällskapen.
Erika- och Prestigeolyckorna har alltså lett till en märkbar skärpning av sjösäkerheten på europeisk nivå. Vissa risker har minskats drastiskt, t.ex. riskerna förknippade med transport av tung eldningsolja i enkelskroviga oljetankfartyg.
Arbetet måste fortsätta och intensifieras. Men skärpningarna måste göras på ett sätt som beaktar sjöfartens betydelse för den europeiska konkurrenskraften.
Mot denna bakgrund lägger kommissionen härmed fram sitt tredje lagstiftningspaket för sjösäkerheten i Europeiska unionen. Paketet följer upp Erika I- och Erika II-paketen[2], men innehåller också åtgärder som stärker konkurrenskraften för fartyg under europeisk flagg. Det ligger också i linje med kommissionens strategiska mål för 2005–2009. I EU 2010: Ett partnerskap för Europas förnyelse – Välstånd, solidaritet och säkerhet [3] skissar kommissionen upp sin vision, och betonar att medborgarnas livskvalitet förutsätter en aktiv politik för att minska de risker som medborgarna ställs inför, t.ex. sjöfartsolyckor. Föreliggande förslag har just detta som mål.
I ett vidare perspektiv bidrar paketet till att öka säkerhetsaspekten i den integrerade europeiska sjöfartspolitik som håller på att växa fram. Dess huvuddrag kommer att beskrivas i en kommande grönbok om unionens sjöfartspolitik som skall vara klar under första halvåret 2006, och innehålla ”en europeisk vision om oceaner och hav”. Syftet är att skapa en rättvis balans mellan ekonomiska, arbetsrättsliga och miljö-, skydds- och säkerhetsrelaterade aspekter på utvecklingen av verksamhet som rör haven. Målet är att förena resursbevarande, konkurrenskraft, långsiktig ekonomisk utveckling och högre sysselsättning.
I. EUROPEISKA UNIONEN STÅR FÖR EN KONKURRENSKRAFTIG, SÄKER OCH BRA SJÖFART
Europeiska unionens ekonomiska utveckling är på grund av geografi, historia och handelns tilltagande globalisering helt beroende av sjöfarten. Detta framgår tydligt av följande siffror:
- Nästan 90 % av unionens externa handel och över 40 % den interna handeln beräknat i varuvolym går via sjöfart.
- Varje år kommer ungefär 1 miljard ton olja in i unionen via dess hamnar, eller korsar unionens vatten.
- Rederier som tillhör medborgare i Europeiska unionen kontrollerar nästan 40 % av världsflottan. EU är världens ledande handelsblock, och nästan all extern handel går via fartyg som kontrolleras från unionen.
- Hela sjöfartssektorn, inbegripet varv, hamnar, fisket och kompletterande verksamhet såsom försäkringsbolag och banker, sysselsätter 3 miljoner människor i Europeiska unionen.
Unionen behöver alltså en konkurrenskraftig flotta och en sjöfartssektor som kan säkra sin lönsamhet och sin plats på den internationella marknaden. Unionen har under flera år fört en aktiv politik för att stödja sin flottas konkurrenskraft. Detta har skett på olika sätt:
- Genom lagstiftning: Det statliga stödet till sjöfartssektorn regleras i riktlinjer (reviderade 2004). Riktlinjerna syftar till att försöka få redarna att återigen flagga sina fartyg i unionen, vilket är en förutsättning för högre kvalitet och säkerhet.
- Genom avtal: Bilaterala och internationella avtal erbjuder unionens aktörer fri tillgång utan diskriminering till den internationella transportmarknaden.
- Genom stöd: Unionens ekonomiska stöd utgår främst inom ramen för stödet till de transeuropeiska nätverken i form av stöd till hamnanläggningar och tillfarter, genom stöd till innovativa tjänster via Marco Polo-programmet och genom stödet till havsforskning.
Kvaliteten på aktörernas tjänster har stor betydelse för sektorns konkurrenskraft. Eftersom kommissionens åtgärder i viss mån motiveras av de senaste årens tragiska olyckor med oljetankfartyg måste åtgärderna också syfta till att höja sjöfartssektorns kvalitet. De måste ge de bästa aktörerna tillfälle att konsolidera sin internationella konkurrenskraft.
Med detta paket vill kommissionen främja insynen i sjöfartssektorn, och därmed framväxten av en rättvisare marknad på internationell nivå och unionsnivå, vilket kommer att gynna de europeiska aktörerna. Kommissionen har för avsikt att se till att befintlig lagstiftning följs noga, och kommer även i fortsättningen att främja korsbefruktningen mellan det internationella regelverket och unionslagstiftningen. Med detta vill kommissionen bidra till en rättvis konkurrens på världsmarknaden, vilket är en förutsättning för att de europeiska flaggstaterna skall kunna bibehålla sin kvalitetsnivå. Kommissionen tänker sig följande åtgärder:
- Unionen skall skärpa kontrollen av att dess sjöfartslagstiftning genomförs och följs. Kommissionen kommer att använda sig av de påtryckningsmedel fördraget erbjuder, och har redan inlett överträdelseförfaranden inför EG-domstolen mot stater som inte har fullgjort sina skyldigheter (några förfaranden har redan resulterat i fällande domar).
- Unionen skall delta i det internationella arbetet i större utsträckning.
Kommissionen tänker bl.a. arbeta för och främja en enhetlig och strikt tolkning av IMO:s internationella föreskrifter. Motsvarande åtgärder kommer att vidtas i fråga om ILO:s (Internationella arbetsorganisationen) föreskrifter inom ramen för den pågående omarbetningen av organisationens konventioner. Härvid har det utmärkta samarbetet med arbetsmarknadens parter möjliggjort stora framsteg i arbetet med den nya konvention som kommissionen vill införliva i unionslagstiftningen.
Kommissionen vill även bidra till uppnåendet av Lissabonstrategins mål genom att förbättra och förenkla befintliga texter, t.ex. direktiven om hamnstatskontroll och klassificeringssällskap, som båda har ändrats flera gånger. Målet har i första hand varit att förbättra regelverkets tydlighet och överskådlighet. Detta kommer först och främst medborgarna och de berörda aktörerna till godo.
Genomförandet av paketet kommer i viss mån att involvera Europeiska sjösäkerhetsbyrån, inrättad genom Europaparlamentets och rådets förordning (EG) nr 1406/2002[4]. Vissa av paketets åtgärder nämns redan i förordningen, andra föranleder ändringar. Kommissionen kommer att lägga fram ett förslag om ändring av förordningen under de kommande månaderna.
Sammanfattningsvis: Konsolideringen av gällande lagstiftning, effektiviseringen av sjöfartsmyndigheterna och inriktningen på högriskfartyg med lindrigare kontroller för lågriskfartyg bidrar på ett betydelsefullt sätt till näringslivets konkurrenskraft. Säkerheten går hand i hand med konkurrenskraften.
II. ÅTGÄRDERNA BEHÖVS REDAN FÖR TILLÄMPNINGEN AV BEFINTLIG LAGSTIFTNING
Medlemsstaterna ansvarar för genomförandet av unionens direktiv och förordningar.
I sin resolution av den 27 april 2004 betonade Europaparlamentet ”att i och med lagstiftningen efter katastroferna med Erika och Prestige har viktiga bestämmelser antagits för att göra fartygstrafiken i EU:s farvatten säkrare. Medlemsstaternas snabba och kompletta genomförande och strikta tillämpning av EU-bestämmelserna måste prioriteras.”
Kommissionen är fast besluten att se till att medlemsstaterna tillämpar unionens sjösäkerhetslagstiftning korrekt. Tillsammans med Europeiska sjösäkerhetsbyrån genomför kommissionen ett särskilt program för kontroll av överensstämmelse och tillämpning på sjösäkerhetsområdet under perioden 2005–2007, vilket redan har lett till en ökning av antalet överträdelseförfaranden mot medlemsstater. Per den 30 september 2005 pågick 68 förfaranden rörande sjösäkerhet, inbegripet förfaranden om underlåtenhet att underrätta kommissionen om genomförandeåtgärder samt klagomål.
Genomförandet av Erika I- och II-direktiven har blivit mycket bättre: för närvarande utreder EG-domstolen tre ärenden. För senare lagstiftning är situationen dystrare; 31 förfaranden pågår. Kommissionen är också bekymrad över vissa staters undermåliga genomförandelagstiftning. Detta gäller särskilt texter för genomförandet av direktiven om hamnstatskontroll respektive mottagningsanordningar i hamn för fartygsgenererat avfall och lastrester; 12 förfaranden pågår om detta. För dessa båda direktiv pågår allt som allt 19 förfaranden om bristande tillämpning av nationell lagstiftning.
III. SÄKERHETEN MÅSTE HÖJAS, OCH FÖRORENING FRÅN FARTYG FÖREBYGGAS
Efter Erika- och Prestige-olyckorna agerade Europeiska unionen i vad som kan beskrivas som ett akut läge för att få på plats defensiva åtgärder som kunde skydda Europa från framtida olyckor och utsläpp. Unionen har ibland beskyllts för att vara alltför försiktig jämfört med USA, som genom lagstiftningen OPA 90 (Oil Pollution Act) agerade ensidigt efter Exxon Valdez-olyckan[5]. En sådan anklagelse bortser från det faktum att omständigheterna skiljer sig åt mellan Europa och USA. Det största problemet i Europa gäller fartyg under tredjelands flagg som transiterar unionens vatten, men utanför medlemsstaternas jurisdiktion: ungefär 200 miljoner ton råolja och oljeprodukter[6] transiterar varje år genom våra vatten utan att anlöpa någon hamn, och därmed utan att någon medlemsstat får tillfälle att utöva rätten att genomföra en hamnstatskontroll för fartygen i fråga.
Osäkerheten till sjöss är inte lätt att komma till rätta med, eftersom sjöfarten till sin natur är en riskfylld verksamhet. Det krävs kraftfullare åtgärder om grundförutsättningarna skall kunna ändras och man på ett bestående sätt skall kunna återskapa en rättvis konkurrens för de aktörer som följer de internationella reglerna.
Det finns flera skäl att skärpa alla regler – internationella såväl som unionsrättsliga – som påverkar säkerheten:
- Alla tillgängliga fakta visar att undermåliga fartyg under bekvämlighetsflagg fortfarande har en lönsam marknad. Enligt siffror från OECD bryter 10 till 15 % (dvs. 5 000-7 000 fartyg) av världsflottan mot de internationella säkerhetsnormerna.
- Statistik från Paris MOU[7] visar att allt fler brister upptäcks vid fartygsinspektioner[8], särskilt i fråga om besättningens arbets- och boendeförhållanden ombord och fartygets drift[9]. Siffrorna understryker att viljan att skydda miljön inte får överskugga det höga pris sjöfolket betalar för den bristande säkerheten.
- Varuutbytet med länder utanför unionen via sjöfart har ökat under de senaste fem åren, både i fråga om volym och värde. Fartygstrafiken har ökat i Europa, även om andelen fartyg i transit sjönk i och med utvidgningen. Flera nya sjövägar har kommit till. De nya, stora oljeterminalerna i Ryssland har lett till en spektakulär och hastig ökning av trafiken i Finska viken. År 2000 passerade ca 40 miljoner ton råolja och oljeprodukter genom Finska viken; detta beräknas ha ökat till 100–120 miljoner ton år 2010. - En annan källa till oro är hur man skall kunna skydda Medelhavet från utsläpp från fartygstrafiken från Svarta havet. Under 2002 passerade 122 miljoner ton olja genom Bosporen ombord på 7 400 oljetankfartyg. Även den ökade oljeproduktionen i trakterna kring Kaspiska havet bidrar till den ökade utsläppsrisken. Om alla planerade utvidgnings- och pipelineprojekt förverkligas kommer den genomsnittliga kapaciteten för oljexport från Kaspiska havet till terminalerna vid Svarta havet att nå 2,4 miljoner fat per dag år 2015. Denna utveckling oroar både länderna i norra Europa och Medelhavsländerna, och det är därmed viktigt att diskutera och betona sjösäkerheten inom ramen för dialogen med unionens grannar. Detta bör särskilt ske inom ramen för inrättandet av det gemensamma ekonomiska området för unionen och Ryssland, och den ram för förbindelserna mellan unionen och dess grannar som inrättas genom den europeiska grannskapspolitiken[10]. Handlingsplaner har redan upprättats tillsammans med partnerskapsländerna i Svarta havs- och Medelhavsregionerna, med flera åtgärder avsedda att stärka sjösäkerhetssamarbetet och förbättra genomförandet av hamnstatskontrollen.
- Kommissionens granskningar av klassificeringssällskap erkända på unionsnivå har visat att rutinerna och bestämmelserna måste skärpas om alla fartygs säkerhet skall kunna kontrolleras kontinuerligt.
- Branschens aktörer åläggs endast ett begränsat skadeståndsansvar genom de internationella konventionerna. Så lindriga bestämmelser är sällsynta inom andra branscher, och kan vara en bidragande orsak till att det är så svårt att avgöra vem i aktörskedjan som är ansvarig. De höjningar av ansvarsgränserna som hittills har gjorts har inte varit tillräckliga, även om höjningen – på kommissionens initiativ – av ansvarsgränserna i FIPOL-konventionen[11] från ca 240 miljoner euro till 900 miljoner euro var ett viktigt steg.
IV. DET BEHÖVS ETT BRA SAMARBETE MELLAN UNIONEN OCH INTERNATIONELLA ORGAN
Kommissionen inser till fullo vikten av åtgärder på internationell nivå när det gäller sjösäkerhet. En internationell åtgärd är i allmänhet att föredra framför en regional om den motsvarar unionens behov. Ett närmare samarbete mellan unionens institutioner och organ, medlemsstaterna och internationella organ (IMO) är alltså önskvärt. Tyvärr saknar unionen – trots utvidgningen – ett internationellt inflytande som motsvarar storleken på dess flotta och dess ekonomiska investeringar i sjöfarten. Anledningen är att unionen inte är medlem av och därmed inte kan agera i eget namn inom ramen för IMO. Kommissionen delar därför helhjärtat Europaparlamentets åsikt (uttryckt i MARE-resolutionen) att rådet bör ansluta unionen till IMO (vilket kommissionens föreslog redan 2002).
Slutsats
Detta tredje sjösäkerhetspaket vilar på en helhet av sinsemellan beroende delar. Det omsätter i praktiken de krav som uttryckts av Europaparlamentet, Europeiska rådet och de europeiska ministrarna samlade i rådet (transport) eller vid den mellanstatliga konferensen om hamnstatskontroll som hölls i Vancouver i november 2004.
Kraven är inte bara en reaktion på en viss olycka, utan syftar till en djupare reform av sjöfartens rutiner och visar, med Europaparlamentets ord ur resolutionen av den 27 april 2004, på behovet av en ”övergripande och konsekvent europeisk sjöfartspolitik som syftar till att skapa ett europeiskt område för sjösäkerhet.” I likhet med föregående paket bidrar det till förverkligandet av de mål som uppställs i den tematiska strategin för skydd av havsmiljöer, i enlighet med Sjätte miljöhandlingsprogrammet.
Åtgärderna i detta tredje paket bidrar till detta, och ingår i en övergripande politik avsedd att lyfta fram en effektiv och bra sjöfart som respekterar människor och miljö. Europeiska unionens samlade insatser, av nationella myndigheter och näringsliv, för att främja en hållbar och lönsam sjöfart kommer att gynna de aktörer som följer säkerhetsnormerna. Paketet skapar rättvisa konkurrensförhållanden som unionens sjöfartsbransch – som bidrar till Europas tillväxt och framgång – kan dra full nytta av.
Europeiska unionen arbetar med en ambitiös politik för att skapa höghastighetsleder till sjöss[12]. Nu behövs tydliga och förutsebara bestämmelser som kan ligga till grund för de investeringar som behövs för detta.
[1] http://www.europarl.eu.int/comparl/tempcom/mare/default_en.htm
[2] KOM(2000) 142 och KOM(2000) 802. Både Erika I och II siktar i första hand på att skärpa befintlig lagstiftning (främst om hamnstatskontroll) men innehåller också helt nya åtgärder, t.ex. om en snabbare utfasning av fartyg med enkelskrov, trafikövervakning, skadestånd vid utsläpp och inrättandet av en europeisk sjösäkerhetsbyrå (med uppgift att bistå kommissionen och medlemsstaterna vid genomförandet av gemenskapslagstiftningen).
[3] KOM(2005) 12, 26.1.2005.
[4] EGT L 208, 5.8.2002, s. 1.
[5] Grundstötningen av det amerikanska oljetankfartyget Exxon-Valdez den 24 mars 1989 ledde till att 40 000 ton råolja släpptes ut utanför Alaskas kust.
[6] Dvs. en fjärdedel av den europeiska importen via sjöfart (som uppgår till 800 miljoner ton och motsvarar 90 % av den totala importen).
[7] http://www.parismou.org
[8] Nästan 72 000 år 2003 mot färre än 58 000 år 1998.
[9] Mellan 2001 och 2003 ökade anmärkningarna om besättningens utbildning och certifiering med 152 %, och anmärkningarna om säkerhetsrutinerna (ISM) med 186 %.
[10] KOM(2004) 373, 12.5.2004.
[11] 1992 års internationella konvention om upprättande av en internationell fond för ersättning av skada orsakad av föroreningar genom olja (http://en.iopcfund.org/).
[12] I kommissionens vitbok om Den gemensamma transportpolitiken fram till 2010: Vägval inför framtiden - KOM(2001) 370 - föreslås att unionen skall försöka skapa höghastighetsleder till sjöss mellan europeiska hamnar, för att ge ett konkurrenskraftigt alternativ till landtransporterna.
P6_TA(2005)0194
Ramavtal om förbindelserna mellan Europaparlamentet och kommissionen
Europaparlamentets beslut om översynen av ramavtalet mellan Europaparlamentet och kommissionen (2005/2076(ACI))
Europaparlamentet fattar detta beslut
- med beaktande av artikel 10 i Fördraget om upprättandet av Europeiska gemenskapen och förklaring 3 som är fogad till slutakten från den regeringskonferens som fastställde Nicefördraget,
- med beaktande av artikel III-397 i Fördraget om upprättande av en konstitution för Europa,
- med beaktande av ramavtalet om förbindelserna mellan Europaparlamentet och kommissionen av den 5 juli 2000 [1],
- med beaktande av sin resolution av den 18 november 2004 om val av den nya kommissionen [2],
- med beaktande av talmanskonferensens beslut av den 14 april 2005,
- med beaktande av förslaget till ramavtal om förbindelserna mellan Europaparlamentet och kommissionen (nedan kallat avtalet),
- med beaktande av artikel 24.3 och artikel 120 i arbetsordningen samt punkt XVIII.4 i bilaga VI till arbetsordningen,
- med beaktande av betänkandet från utskottet för konstitutionella frågor (A6-0147/2005), och av följande skäl:
A. Fördjupningen av demokratin i Europeiska unionen, som undertecknandet av Fördraget om upprättande av en konstitution för Europa är ett bevis på, innebär att förbindelserna mellan Europaparlamentet och kommissionen bör stärkas och att den parlamentariska kontrollen över den verkställande myndigheten bör förbättras.
B. Processen för att tillsätta den nuvarande kommissionen förstärkte den demokratiska legitimiteten i EU:s institutionella system och underströk den politiska dimensionen i förbindelserna mellan de båda institutionerna.
C. Det nya avtal som förelagts parlamentet återspeglar denna utveckling.
D. Nedanstående förtydliganden behöver göras i detta avtal.
E. Mot bakgrund av förloppet hos de förhandlingar som ledde till en politisk överenskommelse är det viktigt att förhandlingarna i fortsättningen anförtros åt personer med ett politiskt mandat.
F. Interinstitutionella avtal och ramavtal har långtgående konsekvenser, och för att öka tillgängligheten och säkra öppenheten är det därför nödvändigt att sammanställa alla befintliga avtal och offentliggöra dessa som bilagor till parlamentets arbetsordning.
1. Förutom den ökade konsekvensen och förenklingen av strukturen välkomnar Europaparlamentet också följande positiva punkter i förslaget till nytt avtal.
a) De nya bestämmelserna om eventuella intressekonflikter (punkt 2).
b) Förfaranden i händelse av att en ledamot av kommissionen byts ut under kommissionens mandattid (punkt 4).
c) Utfästelsen om att alla relevanta uppgifter kommer att lämnas av de nominerade kommissionsledamöterna vid förfarandet för godkännande av kommissionen (punkt 7).
d) Inrättandet av en löpande dialog på högsta nivå mellan kommissionens ordförande och talmanskonferensen (punkt 10).
e) Gemensamt fastställande av särskilt viktiga förslag och initiativ utifrån kommissionens lagstiftnings- och arbetsprogram, den fleråriga interinstitutionella programplaneringen och garantin om att parlamentet informeras på samma sätt som rådet om all kommissionens verksamhet (punkterna 8 och 12).
f) Bättre information från kommissionen om uppföljningen och beaktandet av parlamentets ståndpunkter (punkterna 14 och 31).
g) Offentliggörande av relevant information om kommissionens expertgrupper (punkt 16), med förbehåll för att punkt 2 i detta beslut beaktas.
h) Bekräftelsen av bestämmelserna om parlamentets deltagande i internationella konferenser och nya särskilda hänvisningar till givarkonferenser och valobservation (punkterna 19-25), med förbehåll för den begäran som anges i punkt 4 i detta beslut.
i) Införandet i avtalet (artikel 35) av de åtaganden som kommissionen gjort beträffande genomförandeåtgärderna avseende värdepappers-, bank- och försäkringssektorn ("Lamfalussy-förfarandet") och av överenskommelsen mellan Europaparlamentet och kommissionen om tillämpningsföreskrifter till beslutet om kommittésystemet [3], med förbehåll för kommentarerna i punkt 3 i detta beslut.
j) De åtaganden som gjorts om kommissionens deltagande i parlamentets arbete (punkterna 37-39).
k) Införandet av en bestämmelse om översyn av avtalet (punkt 43) efter det att Fördraget om upprättande av en konstitution för Europa trätt i kraft.
2. Europaparlamentet betonar att det anser att det är viktigt med full insyn när det gäller kommissionens expertgruppers sammansättning och verksamhet (punkt 16 i avtalet) och begär att kommissionen skall tilllämpa avtalet i denna anda.
3. Europaparlamentet uppmanar kommissionen att mot bakgrund av dess förslag av den 11 december 2002 beakta de politiska riktlinjer som parlamentet beslutar om när det utövar sina befogenheter att behandla dokument i kommittéförfarandet.
4. När det handlar om parlamentsledamöters deltagande i delegationer till internationella konferenser och andra internationella förhandlingar anser Europaparlamentet att det är viktigt att parlamentets ledamöter skall få närvara vid EU-interna samordningsmöten, varvid parlamentet förpliktar sig att följa de sekretessregler som gäller för dessa möten. Parlamentet uppmanar därför kommissionen att gentemot rådet stödja sådana önskningar från parlamentets sida.
5. Europaparlamentet insisterar på att kommissionen avsätter en period på minst två månader vid framläggandet av de integrerade riktlinjerna för ekonomi och sysselsättning så att ett ändamålsenligt samråd med Europaparlamentet kan äga rum.
6. Europaparlamentet godkänner det bifogade avtalet.
7. Europaparlamentet beslutar att foga detta avtal som bilaga till arbetsordningen och att det skall ersätta bilagorna XIII och XIV till denna.
8. Europaparlamentet uppdrar åt talmannen att översända detta beslut med bilaga till kommissionen och rådet samt till medlemsstaternas parlament.
[1] EGT C 121, 24.4.2001, s. 122.
[2] Antagna texter, P6_TA(2004)0063.
[3] Rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter (EGT L 184, 17.7.1999, s. 23).
--------------------------------------------------
P6_TA(2005)0057
Togo
Europaparlamentets resolution om Togo
Europaparlamentet utfärdar denna resolution
- med beaktande av ordförandeskapets förklaring på EU:s vägnar av den 9 februari 2005 om den politiska situationen i Togo efter president Eyadémas död,
- med beaktande av det uttalande som ordförandena för den parlamentariska församlingen AVS-EU gjorde den 8 februari 2005 med anledning de händelser som följde president Eyadémas död den 5 februari 2005,
- med beaktande av de uttalanden som ECOWAS, Afrikanska unionen och många afrikanska ledare gjort om situationen i Togo,
- med beaktande av förklaringen av "Organisation Internationale de la Francophonie",
- med beaktande av den afrikanska stadgan om människors och folks rättigheter,
- med beaktande av artikel 65 i Togos grundlag som föreskriver att om republikens president avlider skall presidentämbetets funktioner tillfälligtvis utövas av nationalförsamlingens talman,
- med beaktande av artikel 76 i samma grundlag som föreskriver att personer som utövar regeringsfunktioner inte på några villkor får inneha parlamentariskt mandat,
- med beaktande av artikel 144 i samma grundlag som föreskriver att under interimperioder får inga översynsförfaranden inledas eller fullföljas,
- med beaktande av artikel 115.5 i arbetsordningen, och av följande skäl:
A. Efter president Gnassingbe Eyadémas plötsliga död den 5 februari 2005, efter 38 år vid makten, installerade Togos väpnade styrkor dennes 39-årige son Faure Gnassingbé som president.
B. Enligt landets grundlag skulle talmannen i Togos nationalförsamling, Fambare Ouattara Natchaba, ha utnämnts till interimpresident med uppgift att anordna presidentval inom 60 dagar.
C. Togos nationalförsamling som domineras av Eyadémas parti Rassemblement du Peuple Togolais (RPT) sammankallades hastigt den 6 februari 2005 för att i efterhand legitimera Gnassingbés gripande av makten och ändra landets grundlag för att Gnassingbé skall kunna regera under de återstående tre åren av hans faders mandat.
D. Även om nationalförsamlingen har återupprättat den grundlag som gällde före hans faders död har Faure Gnassingbé ännu inte reagerat på det internationella samfundets uppmaningar att avgå, så att en interimpresident kan på ett effektivt sätt anordna de presidentval som enligt grundlagen skall hållas inom 60 dagar.
E. EU kommer aldrig att erkänna som giltigt ett val anordnat av en olaglig president som tillsatts genom en militärkupp.
F. Vid sitt möte i Niamey (Niger) den 9 februari 2005 förkastade stats- och regeringscheferna för ECOWAS-länderna i starka ordalag den militära intervention som en statskupp varigenom Faure Gnassingbé installerades som president, fördömde nationalförsamlingens lagstridiga hantering av grundlagen och begärde att de togolesiska myndigheterna återupprättar den föregående grundlagen så att presidentval kan hållas inom två månader, med hot om att annars utsättas för sanktioner.
G. Afrikanska unionens ordförande Alpha Oumar Konaré har i ett uttalande slagit fast att Afrikanska unionen inte kan godta att man tilltvingar sig makten med våld.
H. Även "Organisation Internationale de la Francophonie" har i mycket kraftiga ordalag fördömt statskuppen och har beslutat utesluta Togo ur alla sina organ liksom att avbryta allt multilateralt samarbete med landet, med undantag för de program som direkt gynnar civilbefolkningen och som kan bidra till att demokratin återupprättas.
I. EG:s samarbete med Togo avbröts 1993.
1. Europaparlamentet fördömer den statskupp varmed militären möjliggjorde Faure Gnassingbés övertagande av presidentmakten på bekostnad av nationalförsamlingens talman Fambare Ouattara Natchaba.
2. Europaparlamentet kräver att Faure Gnassingbé omedelbart träder tillbaka.
3. Europaparlamentet noterar att grundlagen ändrades den 21 februari 2005, men understryker att en återgång till den konstitutionella ordningen inte säkrats förrän nationalförsamlingens talman Fambare Ouattara Natchaba installerats som interimpresident med uppgift att anordna presidentval i enlighet med landets grundlag.
4. Europaparlamentet välkomnar de sanktioner som ECOWAS införde mot Togo efter tio dagars fruktlösa medlingsförsök, då man bland annat uteslöt Togo ur ECOWAS, återkallade sina ambassadörer och införde ett förbud mot vapenhandel och utfärdande av visum.
5. Europaparlamentet välkomnar de likartade uttalanden och beslut som går i samma riktning av FN, Afrikanska unionen, EU och "Organisation Internationale de la Francophonie".
6. Europaparlamentet uppmanar Togos nationalförsamling och andra myndigheter att omedelbart vidta åtgärder för att lösa den uppkomna situationen och se till att fria och rättvisa val hålls inom två månader, i enlighet med landets grundlag, och att internationella observatörer ges fritt tillträde till dessa.
7. Europaparlamentet upprepar sin övertygelse att återgången till en grundlagsenlig ordning förutsätter en dialog mellan Togos politiska krafter och en översyn av vallagen utifrån principen om samförstånd och i syfte att hålla fria och demokratiska val med full insyn i valprocessen.
8. Europaparlamentet fördömer beslutet att förbjuda alla folkliga demonstrationer under två månader, nedläggningen av åtta privata TV- och radiostationer samt militärens obefogade påtryckningar på oberoende medier i form av hot riktade mot journalister med anledning av deras nyhetsbevakning. Parlamentet uppmanar Togos väpnade styrkor att förbli i sina kaserner och att avstå från handlingar som skulle kunna leda till ytterligare oro.
9. Europaparlamentet kräver att rätten att anordna fredliga demonstrationer och delta i politiska kampanjer skall garanteras, och att de ansvariga för mord och andra brott mot de mänskliga rättigheterna riktade mot människor som deltagit i demonstrationer mot den militära statskuppen ställs inför rätta och straffas.
10. Europaparlamentet erinrar om att de självutnämnda togolesiska myndigheterna måste påta sig det fulla ansvaret för alla angrepp mot civilbefolkningens fysiska säkerhet, i synnerhet angrepp riktade mot representanter för oppositionspartier, människorättsaktivister och journalister.
11. Europaparlamentet uppmanar kommissionen att inte återuppta förhandlingar i syfte att gradvis återupprätta samarbetet tills dess att fria president- och parlamentsval hållits med full insyn.
12. Europaparlamentet uppmanar kommissionen att föreslå riktade sanktioner mot de som står bakom statskuppen.
13. Europaparlamentet uppdrar åt talmannen att översända denna resolution till rådet, kommissionen, generalsekreterarna för FN, Afrikanska unionen och ECOWAS, ordförandena för den parlamentariska församlingen AVS-EU samt till Togos president, regering och nationalförsamling.
--------------------------------------------------
P6_TA(2005)0076
Situationen i Libanon
Europaparlamentets resolution om situationen i Libanon
Europaparlamentet utfärdar denna resolution
- med beaktande av sin resolution av den 16 januari 2003 om ingåendet av ett associeringsavtal med Republiken Libanon [1],
- med beaktande av sina tidigare resolutioner om Europa-Medelhavspartnerskapet, särskilt resolutionen av den 23 februari 2005 [2],
- med beaktande av FN:s säkerhetsråds resolution 1559 om Libanon av den 2 september 2004,
- med beaktande av förklaringen om Libanonn av den 15 februari 2005 från ordföranden i FN:s säkerhetsråd,
- med beaktande av rådets slutsatser om fredsprocessen i Mellanöstern av den 21 februari 2005,
- med beaktande av sin resolution av den 20 november 2003 om ett utvidgat europeiskt grannskap: En ny ram för förbindelserna med våra grannländer i öster och söder [3],
- med beaktande av sin resolution av den 12 februari 2004 om stärkande av EU:s åtgärder för mänskliga rättigheter och demokratisering i samarbete med Medelhavspartnerna [4],
- med beaktande av artikel 103.4 i arbetsordningen, och av följande skäl:
A. Europaparlamentet är djupt chockat över attentatet i Beirut den 14 februari 2005 då Libanons förre premiärminister Rafiq Hariri och andra oskyldiga civila dödades.
B. Rafiq Hariri var en de mest inflytelserika politikerna och en av mest hängivna i Libanons försoningsprocess. Han var också en stark förespråkare av att utländska trupper skulle dra sig tillbaka från hans land.
C. Libanon är ett land med starka historiska, kulturella och ekonomiska band till Europa. Landet är en viktig partner för EU i Mellanöstern och en deltagare i den Europeiska grannskapspolitiken. Denna tragedi utgör ett brott mot de demokratiska principer som både Libanon och Europeiska unionen värnar om.
D. Europaparlamentet gläds åt omfattningen av de senaste dagarnas fredliga och demokratiska folkliga demonstrationer, som har visat att det finns stor nationell enighet mellan människor från de olika politiska och religiösa grupperna i landet.
E. Europaparlamentet välkomnar FN:s generalsekreterare Kofi Annans beslut att tillsätta en undersökningsgrupp som skall ha i uppdrag att utreda "omständigheterna kring, orsakerna till och effekterna av" Libanons tidigare premiärminister Rafiq Hariris död.
F. Den 28 februari 2005 avgick Libanons premiärminister Omar Karami sedan oppositionen inlett en debatt i parlamentet om ett förslag till betänkande om misstroendevotum mot regeringen och som en följd av den folkstorm som kom till uttryck genom de stora folkmassor som oppositionen samlat till demonstrationer för att kräva att de syrianska trupperna skulle dras tillbaka.
G. Enligt planerna skall ett parlamentsval i Libanon hållas i maj 2005, och Libanons folk vill och bör själva avgöra sin politiska framtid.
H. Syriens och Libanons presidenter har beslutat att de syrianska trupperna skall dras tillbaka till östra Bekaadalen. Detta trots att det internationella samfundet krävde en snabb och fullständig reträtt från Libanon.
I. Samtalen mellan Israels regering och den palestinska nationella myndigheten har tagits upp igen, vilket gör det ännu mer angeläget att involvera Syrien och Libanon i processen för att nå en övergripande och varaktig lösning på Mellanösternkonflikten.
J. Syrien skall inom kort underteckna ett associeringsavtal med EU. Därmed åtar sig landet att delta i en politisk dialog som bygger på stöd för demokrati, mänskliga rättigheter, rättsstatsprincipen och respekt för folkrätten.
K. Det är viktigt att hindra att Libanon faller tillbaka i en ny orolig period. Landets sköra demokratiska institutioner måste stödjas och stärkas, och återuppbyggnadsprocessen måste gå vidare.
L. Ett fullständigt demokratiskt och suveränt Libanon kan spela en viktig roll i utvecklingen av Europa-Medelhavspartnerskapet och inom ramen för den europeiska grannskapspolitiken.
1. Europaparlamentet fördömer otvetydigt bombattentatet i Beirut den 14 februari 2005 som orsakade Libanons premiärminister Rafiq Hariris och andra oskyldiga civilpersoners död. Parlamentet ser med förfäran och indignation på denna barbariska handling och uttrycker sitt djupaste deltagande till Hariris anhöriga och till de övriga offrens familjer.
2. Europaparlamentet önskar i enlighet med förklaringen av ordföranden i FN:s säkerhetsråd av den 15 februari 2005 att med all tilgänglig kraft utreda orsakerna till, omständigheterna kring och följderna av detta attentat. Parlamentet uppmanar de libanesiska myndigheterna att fortsätta samarbeta med FN:s utredningsgrupp.
3. Europaparlamentet hoppas att detta brott inte kommer att underminera valprocessen i Libanon och betonar vikten av att fria, demokratiska och öppna parlamentsval hålls i landet. Europaparlamentet upprepar sitt krav att unionen skall sända en delegation med observatörer för att övervaka parlamentsvalet i Libanon, och uppmanar kommissionen att vidta alla åtgärder som behövs i denna fråga.
4. Europaparlamentet uppmanar kommissionen att omedelbart inleda ett samarbete genom att stödja det civila samhället och de oberoende icke-statliga organisationerna via Meda-programmet och det europeiska initiativet för demokrati och mänskliga rättigheter.
5. Europaparlamentet uppmanar kommissionen att färdigställa handlingsplanen för Libanon, vilken bör omfatta alla frågor om politisk stabilitet i landet, förstärkning av landets demokratiska institutioner och påskyndande av återuppbyggnadsprocessen.
6. Europaparlamentet välkomnar varmt den positiva utvecklingen i Mellanöstern de senaste veckorna, även den upplivade förhandlingsprocessen mellan Israel och Palestina, och uppmanar Syrien att inte tolerera någon form av terrorism, vilket även omfattar stöd till Hizbollah och till andra väpnade grupper.
7. Det finns klara bevis för Hizbollahs terroristaktiviteter. Enligt Europaparlamentet är det därför nödvändigt att rådet vidtar alla åtgärder som behövs för att stoppa gruppens terrordåd.
8. Europaparlamentet anser att det i detta sammanhang är viktigt att Syrien och Israel återupptar en direkt dialog för att skapa fred och säkerhet och trygga ländernas suveränitet och integritet i överensstämmelse med FN:s säkerhetsråds resolutioner.
9. Europaparlamentet uppmanar Syrien att samarbeta fullt ut med Europeiska unionen inom ramen för grannskapspolitiken för att trygga fred och stabilitet i regionen, och påminner om hur betydelsefullt det är att resolution 1559 genomförs, i vilken det internationella samfundets stöd för Libanons territoriella integritet, suveränitet och oberoende bekräftas. Parlamentet uppmanar även Syrien att avhålla sig från all form av inblandning i Libanons inre angelägenheter. Parlamentet noterar beslutet om att de syrianska trupperna skall dras tillbaka före slutet av mars, men begär en total reträtt från Libanon av de syrianska trupperna och Syriens underrättelsetjänst i enlighet med FN:s säkerhetsråds resolutioner. Parlamentet anser att associeringsavtalet och fortsatt utveckling a
P6_TA(2005)0116
Ekonomiska följder av Rumäniens och Bulgariens anslutning
Europaparlamentets resolution om de ekonomiska följderna av Bulgariens och Rumäniens anslutning(2005/2031(INI))
Europaparlamentet utfärdar denna resolution
- med beaktande av artikel 272 i EG-fördraget,
- med beaktande av det interinstitutionella avtalet av den 6 maj 1999 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och förbättring av budgetförfarandet [1], särskilt punkterna 27 och 30,
- med beaktande av resultatet av förhandlingarna med rådets ordförandeskap och trepartsmötena den 5 och 13 april 2005,
- med beaktande av artikel 45 i arbetsordningen,
- med beaktande av budgetutskottets betänkande (A6-0090/2005), och av följande skäl:
A. EG-fördraget, särskilt artikel 272, och det interinstitutionella avtalet av den 6 maj 1999, särskilt punkterna 27 och 30, innehåller bestämmelser som fastslår budgetmyndighetens befogenheter och förfaranden när det gäller klassificering av utgifter och ansvarig myndighet.
1. Europaparlamentet godkänner det gemensamma uttalande som bifogas denna resolution.
2. Europaparlamentet uppdrar åt talmannen att översända denna resolution tillsammans med det gemensamma uttalandet till rådet och kommissionen.
[1] EGT C 172, 18.6.1999, s. 1. Avtalet ändrat genom beslut 2003/429/EG (EUT L 147, 14.6.2003, s. 25).
--------------------------------------------------
[pic] | EUROPEISKA GEMENSKAPERNAS KOMMISSION |
Bryssel den 08.04.2005
KOM(2005)131 slutlig
2005/0031(CNS)
Förslag till
RÅDETS BESLUT
om undertecknandet av ett protokoll till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge
Förslag till
RÅDETS BESLUT
om ingåendet av ett protokoll till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge
(framlagda av Komissionen)
MOTIVERING
politisk och rättslig ram
Den 19 januari 2001 ingick Europeiska gemenskapen ett avtal med Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge. I artikel 12 i detta avtal anges att Danmark kan begära att få ansluta sig till detta avtal och att gemenskapen, Norge och Island, med Danmarks medgivande, fastställer villkoren för detta i ett protokoll till avtalet.
I enlighet med artiklarna 1 och 2 i protokollet om Danmarks ställning som är fogat till Fördraget om Europeiska unionen och Fördraget om upprättandet av Europeiska gemenskapen deltog Danmark inte i rådets antagande av förordning (EG) nr 343/2003 om kriterier och mekanismer för att avgöra vilken medlemsstat som har ansvaret för att pröva en asylansökan som en medborgare i tredje land har gett in i någon medlemsstat (Dublin II-förordningen) och förordning (EG) nr 2725/2000 om inrättande av Eurodac för jämförelse av fingeravtryck för en effektiv tillämpning av Dublinkonventionen (Eurodac-förordningen). Danmark är part i konventionen rörande bestämmandet av den ansvariga staten för prövningen av en ansökan om asyl som framställts i en av medlemsstaterna i de Europeiska gemenskaperna (Dublinkonventionen), som undertecknades i Dublin den 15 juni 1990.
Den 16 februari 2001 begärde Danmark att få delta i avtalet mellan Europeiska gemenskapen, Danmark och Norge.
Genom sitt beslut av den 6 maj 2003 bemyndigade rådet kommissionen att inleda förhandlingar om ett protokoll till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge i enlighet med artikel 12 i avtalet.
Förhandlingarna om ingående av ett protokoll till avtalet med Norge och Island slutfördes i och med att texten paraferades den 12 januari 2005.
Bifogade förslag utgör de rättsliga instrumenten för undertecknandet respektive ingåendet av protokollet. Vad gäller gemenskapen är den rättsliga grunden för beslutet om undertecknande artikel 63.1 a jämförd med artikel 300.2 första stycket första meningen och för beslutet om ingående artikel 63.1 a jämförd med artikel 300.2 första stycket första meningen och artikel 300.3 första stycket. Detta innebär att rådet skall besluta med kvalificerad majoritet efter att ha hört Europaparlamentet om ingåendet av protokollet.
II. resultaten av förhandlingarna
Kommissionen anser att de mål som rådet fastställde i sina förhandlingsdirektiv är uppnådda och att förslaget till protokoll är godtagbart för gemenskapen. Avtalet består av sammanlagt sex artiklar. Det innehåller också en bilaga som är en integrerad del av avtalet.
Det slutliga innehållet i protokollet kan sammanfattas enligt följande:
- Genom protokollet skall bestämmelserna i de så kallade Dublin II- och Eurodacförordningarna och dessas tillämpningsförordningar tillämpas i förbindelserna mellan Konungariket Danmark, å ena sidan, och Republiken Island och Konungariket Norge, å andra sidan. Genom protokollet skall även kommande ändringar eller nya tillämpningsföreskrifter vara tillämpliga i dessa länder.
- Island och Norge ges rätt att lägga fram inlagor eller andra skriftliga synpunkter till EG-domstolen om en dansk domstol begär förhandsavgörande från denna om tolkningen av en bestämmelse i avtalet mellan Europeiska gemenskapen och Danmark.
- En förlikningsmekanism föreskrivs för det fall då oenighet föreligger mellan Danmark, å ena sidan, och Island eller Norge, å andra sidan, om tolkningen eller tillämpningen av protokollet.
- Protokollet innehåller bestämmelser om upphörande.
III. SLUTSATSER
Mot bakgrund av ovan nämnda resultat förslår kommissionen att rådet
- beslutar att protokollet skall undertecknas på gemenskapens vägnar och bemyndigar rådets ordförande att utse den eller de personer som skall ha behörighet att underteckna avtalet på gemenskapens vägnar, och
- efter att ha hört Europaparlamentet, godkänner protokollet till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge.
Förslag till
RÅDETS BESLUT
om undertecknandet av ett protokoll till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge
(Text av betydelse för EES)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 63.1 a, jämförd med artikel 300.2 första stycket första meningen i detta,
med beaktande av kommissionens förslag[1], och
av följande skäl:
(1) Genom sitt beslut av den 6 maj 2003 bemyndigade rådet kommissionen att inleda förhandlingar om ett protokoll till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge.
(2) Förhandlingarna om undertecknandet av avtalet ägde rum under perioden juni 2004–januari 2005.
(3) Avtalet, som paraferades i Bryssel den 12 januari 2005, bör undertecknas med förbehåll för att det ingås.
(4) I enlighet med artikel 3 i protokollet om Förenade kungarikets och Irlands ställning som är fogat till Fördraget om Europeiska unionen och Fördraget om upprättandet av Europeiska gemenskapen, deltar Förenade kungariket och Irland i antagandet och tillämpningen av detta beslut.
(5) I enlighet med artiklarna 1 och 2 i protokollet om Danmarks ställning, fogat till Fördraget om Europeiska unionen och Fördraget om upprättandet av Europeiska gemenskapen, deltar Danmark inte i antagandet av detta beslut som därför inte är bindande för eller tillämpligt i Danmark.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Enda artikel
Med förbehåll för att protokollet ingås bemyndigas rådets ordförande att utse den eller de personer som skall ges befogenhet att på Europeiska gemenskapens vägnar underteckna protokollet till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge.
[pic] | EUROPEISKA GEMENSKAPERNAS KOMMISSION |
Bryssel den 08.04.2005
KOM(2005)131 slutlig
2005/0031(CNS)
Förslag till
RÅDETS BESLUT
om undertecknandet av ett protokoll till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge
Förslag till
RÅDETS BESLUT
om ingåendet av ett protokoll till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge
(framlagda av Komissionen)
MOTIVERING
politisk och rättslig ram
Den 19 januari 2001 ingick Europeiska gemenskapen ett avtal med Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge. I artikel 12 i detta avtal anges att Danmark kan begära att få ansluta sig till detta avtal och att gemenskapen, Norge och Island, med Danmarks medgivande, fastställer villkoren för detta i ett protokoll till avtalet.
I enlighet med artiklarna 1 och 2 i protokollet om Danmarks ställning som är fogat till Fördraget om Europeiska unionen och Fördraget om upprättandet av Europeiska gemenskapen deltog Danmark inte i rådets antagande av förordning (EG) nr 343/2003 om kriterier och mekanismer för att avgöra vilken medlemsstat som har ansvaret för att pröva en asylansökan som en medborgare i tredje land har gett in i någon medlemsstat (Dublin II-förordningen) och förordning (EG) nr 2725/2000 om inrättande av Eurodac för jämförelse av fingeravtryck för en effektiv tillämpning av Dublinkonventionen (Eurodac-förordningen). Danmark är part i konventionen rörande bestämmandet av den ansvariga staten för prövningen av en ansökan om asyl som framställts i en av medlemsstaterna i de Europeiska gemenskaperna (Dublinkonventionen), som undertecknades i Dublin den 15 juni 1990.
Den 16 februari 2001 begärde Danmark att få delta i avtalet mellan Europeiska gemenskapen, Danmark och Norge.
Genom sitt beslut av den 6 maj 2003 bemyndigade rådet kommissionen att inleda förhandlingar om ett protokoll till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge i enlighet med artikel 12 i avtalet.
Förhandlingarna om ingående av ett protokoll till avtalet med Norge och Island slutfördes i och med att texten paraferades den 12 januari 2005.
Bifogade förslag utgör de rättsliga instrumenten för undertecknandet respektive ingåendet av protokollet. Vad gäller gemenskapen är den rättsliga grunden för beslutet om undertecknande artikel 63.1 a jämförd med artikel 300.2 första stycket första meningen och för beslutet om ingående artikel 63.1 a jämförd med artikel 300.2 första stycket första meningen och artikel 300.3 första stycket. Detta innebär att rådet skall besluta med kvalificerad majoritet efter att ha hört Europaparlamentet om ingåendet av protokollet.
II. resultaten av förhandlingarna
Kommissionen anser att de mål som rådet fastställde i sina förhandlingsdirektiv är uppnådda och att förslaget till protokoll är godtagbart för gemenskapen. Avtalet består av sammanlagt sex artiklar. Det innehåller också en bilaga som är en integrerad del av avtalet.
Det slutliga innehållet i protokollet kan sammanfattas enligt följande:
- Genom protokollet skall bestämmelserna i de så kallade Dublin II- och Eurodacförordningarna och dessas tillämpningsförordningar tillämpas i förbindelserna mellan Konungariket Danmark, å ena sidan, och Republiken Island och Konungariket Norge, å andra sidan. Genom protokollet skall även kommande ändringar eller nya tillämpningsföreskrifter vara tillämpliga i dessa länder.
- Island och Norge ges rätt att lägga fram inlagor eller andra skriftliga synpunkter till EG-domstolen om en dansk domstol begär förhandsavgörande från denna om tolkningen av en bestämmelse i avtalet mellan Europeiska gemenskapen och Danmark.
- En förlikningsmekanism föreskrivs för det fall då oenighet föreligger mellan Danmark, å ena sidan, och Island eller Norge, å andra sidan, om tolkningen eller tillämpningen av protokollet.
- Protokollet innehåller bestämmelser om upphörande.
III. SLUTSATSER
Mot bakgrund av ovan nämnda resultat förslår kommissionen att rådet
- beslutar att protokollet skall undertecknas på gemenskapens vägnar och bemyndigar rådets ordförande att utse den eller de personer som skall ha behörighet att underteckna avtalet på gemenskapens vägnar, och
- efter att ha hört Europaparlamentet, godkänner protokollet till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge.
Förslag till
RÅDETS BESLUT
om undertecknandet av ett protokoll till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge
(Text av betydelse för EES)
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 63.1 a, jämförd med artikel 300.2 första stycket första meningen i detta,
med beaktande av kommissionens förslag[1], och
av följande skäl:
(1) Genom sitt beslut av den 6 maj 2003 bemyndigade rådet kommissionen att inleda förhandlingar om ett protokoll till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge.
(2) Förhandlingarna om undertecknandet av avtalet ägde rum under perioden juni 2004–januari 2005.
(3) Avtalet, som paraferades i Bryssel den 12 januari 2005, bör undertecknas med förbehåll för att det ingås.
(4) I enlighet med artikel 3 i protokollet om Förenade kungarikets och Irlands ställning som är fogat till Fördraget om Europeiska unionen och Fördraget om upprättandet av Europeiska gemenskapen, deltar Förenade kungariket och Irland i antagandet och tillämpningen av detta beslut.
(5) I enlighet med artiklarna 1 och 2 i protokollet om Danmarks ställning, fogat till Fördraget om Europeiska unionen och Fördraget om upprättandet av Europeiska gemenskapen, deltar Danmark inte i antagandet av detta beslut som därför inte är bindande för eller tillämpligt i Danmark.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Enda artikel
Med förbehåll för att protokollet ingås bemyndigas rådets ordförande att utse den eller de personer som skall ges befogenhet att på Europeiska gemenskapens vägnar underteckna protokollet till avtalet mellan Europeiska gemenskapen och Republiken Island och Konungariket Norge om kriterier och mekanismer för att fastställa vilken stat som skall ansvara för handläggningen av en asylansökan som görs i en medlemsstat eller i Island eller Norge.
[pic] | EUROPEISKA GEMENSKAPERNAS KOMMISSION |
Bryssel den 13.05.2005
KOM(2005) 190 slutlig
2005/0072 (COD)
2005/0073 (COD)
2005/0074 (COD)
2005/0075 (COD)
2005/0076 (COD)
2005/0077 (CNS)
2005/0078 (CNS)
2005/0079 (CNS)
2005/0080 (CNS)
2005/0081 (COD)
2005/0082 (COD)
2005/0083 (COD)
2005/0084 (CNS)
2005/0085 (COD)
2005/0086 (COD)
2005/0087 (COD)
2005/0088 (COD)
2005/0089 (CNS)
Förslag till
EUROPAPARLAMENTETS OCH RÅDETS FÖRORDNING
om ändring av förordning (EEG) nr 1210/90 om inrättande av Europeiska miljöbyrån och Europeiska nätverket för miljöinformation och miljöövervakning, vad beträffar mandatperioden för den verkställande direktören
Förslag till
EUROPAPARLAMENTETS OCH RÅDETS FÖRORDNING
om ändring av förordning (EEG) nr 337/75 om uppbyggnaden av ett europeiskt centrum för utveckling av yrkesutbildning, vad beträffar mandatperioden för direktören
Förslag till
EUROPAPARLAMENTETS OCH RÅDETS FÖRORDNING
om ändring av förordning (EEG) nr 1365/75 om bildande av en europeisk fond för förbättring av levnads- och arbetsvillkor, vad beträffar mandatperioden för den verkställande direktören och den vice verkställande direktören
Förslag till
EUROPAPARLAMENTETS OCH RÅDETS FÖRORDNING
om ändring av förordning (EEG) nr 1360/90 om inrättandet av en europeisk yrkesutbildningsstiftelse vad direktörens ämbetsperiod avser
Förslag till
EUROPAPARLAMENTETS OCH RÅDETS FÖRORDNING
om ändring av förordning (EEG) nr 302/93 om upprättande av ett europeiskt centrum för kontroll av narkotika och narkotikamissbruk, vad beträffar mandatperioden för direktören
MOTIVERING
1. FÖRSLAGETS SYFTEN
I Europeiska unionen finns det för närvarande 20 decentraliserade organ som kan inordnas under beteckningen gemenskapsorgan (eller byråer). Dessa har vissa gemensamma kännetecken, t.ex. att varje organ har inrättats genom att det har antagits en förordning som rättslig grund för organet i fråga och att de har ställning som juridisk person, autonomi i administrativt och finansiellt hänseende och ett tydligt avgränsat behörighets- och verksamhetsområde.
Ledaren för ett gemenskapsorgan har i regel titeln direktör. I vissa organ finns det även en eller flera vice direktörer. Varaktigheten för dessa personers mandat är i allmänhet 4-5 år. Enligt de flesta grundförordningarna kan en direktörs (eller i förekommande fall vice direktörs) mandat emellertid förlängas med en eller flera perioder. Villkoren för utseende av direktören och varaktigheten för dennes mandat anges i grundförordningen för varje gemenskapsorgan.
De organ som är behöriga för utseendet valde fram till de senaste åren att förlänga mandatet för en tjänstgörande direktör helt enkelt genom att fatta ett beslut. Kommissionen kom efter att ha företagit en ingående prövning av bestämmelserna i grundförordningarna fram till att det tillvägagångssättet innebar ett juridiskt problem.
I de franskspråkiga versionerna av grundförordningarna för gemenskapsorganen används (utom i de franskspråkiga versionerna av förordning (EEG) nr 1360/90 om inrättandet av en europeisk yrkesutbildningsstiftelse och förordning (EG) nr 851/2004 om inrättande av ett europeiskt centrum för förebyggande och kontroll av sjukdomar) begreppen renouvelable och renouvellement när texterna handlar om möjligheterna att förlänga mandatet för en direktör eller motsvarande (i de svenskspråkiga versionerna talas det i regel om att ett mandat kan förnyas eller förlängas). I artikel 214.1 (som handlar om hur ledamöterna av kommissionen utses) och artiklarna 223 och 224 (som handlar om hur bl.a. domarna i EG-domstolen utses) i Fördraget om upprättandet av Europeiska gemenskapen finns analoga bestämmelser. I båda fallen har det fastställts att möjligheten till renouvellement (förnyelse) av ett mandat inte innebär att ett förenklat utseendeförfarande tillämpas och att mandatet kan förlängas utan att det i fördraget angivna utseendeförfarandet behöver iakttas.
Under dessa omständigheter kan möjligheten till förnyelse av mandatet inte tolkas på annat sätt än att innehavaren av tjänsten när mandatet löper ut åter måste anmäla sig som kandidat.
Om detta tillämpas på gemenskapsorganen, leder det till slutsatsen att möjligheten att förnya mandatet för direktören inte innebär en befrielse från tillämpning av det i grundförordningen angivna utseendeförfarandet.
En direktör eller vice direktör är för övrigt inte bara innehavare av ett mandat, utan även medlem av personalen i gemenskapsorganet och anställd på kontrakt som tillfälligt anställd. Tjänsten som direktör eller vice direktör omfattas därmed av de s.k. anställningsvillkoren för övriga anställda i Europeiska gemenskaperna.
Utseendeförfarandet måste därför omfatta bl.a. offentliggörande av tjänsten i samtliga medlemsstater och ett urvalsförfarande som är förenligt med reglerna i grundförordningen och i anställningsvillkoren för övriga anställda i Europeiska gemenskaperna.
Dessa förfaranden är i allmänhet långdragna och relativt kostsamma. Om de måste tillämpas och en tjänstgörande direktör beslutar sig för att åter anmäla sig som kandidat, kan följden också bli att gemenskapsorganets verksamhet avtar eller störs under den tid förfarandena pågår.
Med beaktande av gemenskapsorganens specifika behov och av tillvägagångssättet under de senaste åren förefaller det inte vara lämpligt att tvinga gemenskapsorganen att genomföra ett urvalsförfarande varje gång det första mandatet för en direktör (eller en annan berörd befattningshavare) löper ut. De organ som är behöriga för utseendet borde ha möjlighet att välja mellan en förlängning av det första mandatet och ett nytt urvalsförfarande.
Det bör även beaktas att direktören inte bara är ansvarig för förvaltningen utan även har en viktig roll att spela i arbetet i gemenskapsorganet och när det gäller att uppnå organets mål. Den utseende myndigheten måste när den fattar sitt beslut ta hänsyn såväl till behovet av att sörja för kontinuitet i den administrativa ledningen av gemenskapsorganet som till betydelsen av att organet utvecklas i riktning mot nya idéer och strategier.
Därför bör ett beslut om att förlänga mandatet för en tjänstgörande direktör fattas på grundval av en utvärdering (som utförts av den myndighet som vid ett urvalsförfarande föreslår den utseende myndigheten kandidater) av de resultat som direktören har uppnått och av gemenskapsorganets behov och bör en förlängning medges endast en gång och för en tid som inte överstiger den som anges för det första mandatet.
Kommissionen föreslår att grundförordningarna för 18 gemenskapsorgan ändras och lägger därför fram sammanlagt 18 förslag till förordningar om ändring av de artiklar i grundförordningarna som handlar om hur ledarna för organen utses.
Grundförordningarna för två gemenskapsorgan behöver inte ändras: rådets förordning (EG) nr 2667/2000 av den 5 december 2000 om Europeiska byrån för återuppbyggnad[1] och Europaparlamentets och rådets förordning (EG) nr 460/2004 av den 10 mars 2004 om inrättandet av den europeiska byrån för nät- och informationssäkerhet[2]. I de förordningarna finns det nämligen inga bestämmelser om en eventuell förnyelse av mandatet för direktören, eftersom de berörda gemenskapsorganen har inrättats för att verka enbart under en begränsad tid.
Det läggs inte heller fram några förslag till ändring av de rättsakter genom vilka de organ som omfattas av andra och tredje pelaren inrättades.
Vad beträffar de båda (ännu icke inrättade) gemenskapsorgan som har varit föremål för förordningsförslag som är under prövning eller håller på att antas (Europeiska kemikaliemyndigheten[3] och Gemenskapens kontrollorgan för fiske[4]) kommer kommissionen vid behov att lägga fram ändringsförslag i syfte att sörja för harmonisering av texterna för samtliga gemenskapsorgan.
2. RÄTTSLIG GRUND OCH ANTAGANDEFÖRFARANDE
Varje förordning om inrättande av ett gemenskapsorgan grundar sig i princip på en fördragsartikel som handlar om ett ämnesområde som har att göra med det berörda organets behörighets- och verksamhetsområde och av vilken det framgår vilket förfarande som är tillämpligt för antagandet av åtgärder på ämnesområdet i fråga.
Av denna anledning förefaller det nödvändigt att anta en ändringsförordning för var och en av de grundförordningar om inrättande av ett gemenskapsorgan som skall ändras.
Vad beträffar förfarandet för antagandet av de enskilda ändringsförordningarna bör det förfarande som gällde vid tidpunkten för antagandet av grundförordningen iakttas men bör även sådana förändringar – ändringar av Europaparlamentets befogenheter enligt fördraget eller ändringar av den rättsliga grunden för antagande av åtgärder inom det berörda ämnesområdet – som inträffat efter antagandet av grundförordningen beaktas.
Detta gäller för ändringen av grundförordningen för Europeiska miljöbyrån men även för ändringen av fem grundförordningar för vilka den rättsliga grunden för antagande av åtgärder inte längre är artikel 308 (f.d. artikel 235) i fördraget utan fördragsartiklar som har ett närmare samband med de berörda organens behörighets- och verksamhetsområden.
Det rör sig här å ena sidan om ändringen av grundförordningen för Europeiska centrumet för kontroll av narkotika och narkotikamissbruk, vilken förordning för närvarande är föremål för kodifiering (rådets uppfattning i samband med detta arbete är att artikel 152 i fördraget nu bör användas som rättslig grund och kommissionen har godtagit detta), och å andra sidan om ändringen av förordningen för Europeiskt centrum för utveckling av yrkesutbildning (artikel 150 används som rättslig grund för ändringsförordningen), för Europeiska fonden för förbättring av levnads- och arbetsvillkor (artikel 137.1 a och b), för Europeiska yrkesutbildningsstiftelsen (artikel 150) och för Europeiska arbetsmiljöbyrån (artikel 137.1 a).
3. FÖRORDNINGSFÖRSLAGENS UTFORMNING
3.1. De tre skälen i ingressen har samma utformning i alla förordningsförslag:
Det är nödvändigt att harmonisera reglerna rörande villkoren och förfarandena för förlängning av mandatperioden för, alltefter omständigheterna, direktören, vice direktören eller ordföranden i vissa gemenskapsorgan.
Det bör föreskrivas att mandatperioden skall kunna förlängas en gång efter det att en lämplig utvärdering har gjorts.
… förordning (…) nr …/… … [titeln på den förordning genom vilken gemenskapsorganet inrättas] bör därför ändras.
3.2. För de förordningar som ändras föreslås som regel följande standardformulering:
Xxx [beteckningen på gemenskapsorganet, t.ex. Byrån] skall ledas av en yyy [beteckningen på den som leder gemenskapsorganet, t.ex. direktör] som på förslag av kommissionen** utnämns av styrelsen* för en period av fem år, vilken period på förslag av kommissionen** och efter det att en utvärdering har gjorts kan förlängas en gång, med högst fem år.
Inom ramen för utvärderingen skall kommissionen** särskilt bedöma
- de resultat som har uppnåtts under den första mandatperioden och det sätt på vilket resultaten har uppnåtts, och
- xxxs uppgifter och behov under de närmaste åren.
* Ledaren för följande gemenskapsorgan utnämns av rådet: Gemenskapens växtsortsmyndighet (CPVO) och Kontoret för harmonisering inom den inre marknaden (varumärken och mönster) (KHIM). Ledaren för följande gemenskapsorgan utnämns av kommissionen: Europeiskt centrum för utveckling av yrkesutbildning (Cedefop) och Europeiska fonden för förbättring av levnads- och arbetsvillkor (Eurofound).
** Styrelsen, vad KHIM, Cedefop och Eurofound beträffar.
3.3. De föreslagna ändringarna rör följande gemenskapsorgan och förordningar:
- Europeiskt centrum för utveckling av yrkesutbildning (Cedefop): rådets förordning (EEG) nr 337/75 av den 10 februari 1975 om uppbyggnaden av ett europeiskt centrum för utveckling av yrkesutbildning (artikel 6.2).
- Europeiska fonden för förbättring av levnads- och arbetsvillkor (Eurofound): rådets förordning (EEG) nr 1365/75 av den 26 maj 1975 om bildande av en europeisk fond för förbättring av levnads- och arbetsvillkor (artikel 8.3).
- Europeiska miljöbyrån (EEA): rådets förordning (EEG) nr 1210/90 av den 7 maj 1990 om inrättande av Europeiska miljöbyrån och Europeiska nätverket för miljöinformation och miljöövervakning (artikel 9.1).
- Europeiska yrkesutbildningsstiftelsen (ETF): rådets förordning (EEG) nr 1360/90 av den 7 maj 1990 om inrättandet av en europeisk yrkesutbildningsstiftelse (artikel 7.1), ändrat genom rådets förordning (EG) nr 1572/98 av den 17 juli 1998.
- Europeiska centrumet för kontroll av narkotika och narkotikamissbruk (ECNN): rådets förordning (EEG) nr 302/93 av den 8 februari 1993 om upprättande av ett europeiskt centrum för kontroll av narkotika och narkotikamissbruk (artikel 9.1).
- Kontoret för harmonisering inom den inre marknaden (varumärken och mönster) (KHIM): rådets förordning (EG) nr 40/94 av den 20 december 1993 om gemenskapsvarumärken (artikel 120.2).
- Europeiska arbetsmiljöbyrån (OSHA): rådets förordning (EG) nr 2062/94 av den 18 juli 1994 om upprättande av en europeisk arbetsmiljöbyrå (artikel 11.1).
- Gemenskapens växtsortsmyndighet (CPVO): rådets förordning (EG) nr 2100/94 av den 27 juli 1994 om gemenskapens växtförädlarrätt (artikel 43.2).
- Översättningscentrum för Europeiska unionens organ (CdT): rådets förordning (EG) nr 2965/94 av den 28 november 1994 om upprättande av ett översättningscentrum för Europeiska unionens organ (artikel 9.1).
- Europeiskt centrum för övervakning av rasism och främlingsfientlighet (EUMC): rådets förordning (EG) nr 1035/97 av den 2 juni 1997 om inrättande av ett europeiskt centrum för övervakning av rasism och främlingsfientlighet (artikel 10.1).
- Europeiska myndigheten för livsmedelssäkerhet (EFSA): Europaparlamentets och rådets förordning (EG) nr 178/2002 av den 28 januari 2002 om allmänna principer och krav för livsmedelslagstiftning, om inrättande av Europeiska myndigheten för livsmedelssäkerhet och om förfaranden i frågor som gäller livsmedelssäkerhet (artikel 26.1).
- Europeiska sjösäkerhetsbyrån (EMSA): Europaparlamentets och rådets förordning (EG) nr 1406/2002 av den 27 juni 2002 om inrättande av en europeisk sjösäkerhetsbyrå (artikel 16.2).
- Europeiska byrån för luftfartssäkerhet (EASA): Europaparlamentets och rådets förordning (EG) nr 1592/2002 av den 15 juli 2002 om fastställande av gemensamma bestämmelser på det civila luftfartsområdet och inrättande av en europeisk byrå för luftfartssäkerhet (artikel 30.4).
- Europeiskt centrum för förebyggande och kontroll av sjukdomar (ECDPC): Europaparlamentets och rådets förordning (EG) nr 851/2004 av den 21 april 2004 om inrättande av ett europeiskt centrum för förebyggande och kontroll av sjukdomar (artikel 17.1).
- Europeiska läkemedelsmyndigheten (EMEA): Europaparlamentets och rådets förordning (EG) nr 726/2004 av den 31 mars 2004 om inrättande av gemenskapsförfaranden för godkännande av och tillsyn över humanläkemedel och veterinärmedicinska läkemedel samt om inrättande av en europeisk läkemedelsmyndighet (artikel 64.1).
- Europeiska järnvägsbyrån (ERA): Europaparlamentets och rådets förordning (EG) nr 881/2004 av den 29 april 2004 om inrättande av en europeisk järnvägsbyrå (artikel 31.3).
- Europeiska tillsynsmyndigheten för GNSS: rådets förordning (EG) nr 1321/2004 av den 12 juli 2004 om inrättandet av strukturer för förvaltningen av de europeiska programmen för satellitbaserad radionavigering (artikel 7.2 tredje stycket).
- Europeiska byrån för förvaltningen av det operativa samarbetet vid de yttre gränserna: rådets förordning (EG) nr 2007/2004 av den 26 oktober 2004 om inrättande av en europeisk byrå för förvaltningen av det operativa samarbetet vid Europeiska unionens medlemsstaters yttre gränser (artikel 26.5).
2005/0072 (COD)
Förslag till
EUROPAPARLAMENTETS OCH RÅDETS FÖRORDNING
om ändring av förordning (EEG) nr 1210/90 om inrättande av Europeiska miljöbyrån och Europeiska nätverket för miljöinformation och miljöövervakning, vad beträffar mandatperioden för den verkställande direktören
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av Fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 175 i detta,
med beaktande av kommissionens förslag[5],
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande[6],
med beaktande av Regionkommitténs yttrande[7],
i enlighet med förfarandet i artikel 251 i EG-fördraget[8], och
av följande skäl:
(1) Det är nödvändigt att harmonisera reglerna rörande villkoren och förfarandena för förlängning av mandatperioden för, alltefter omständigheterna, direktören, vice direktören eller ordföranden i vissa gemenskapsorgan.
(2) Det bör föreskrivas att mandatperioden skall kunna förlängas en gång efter det att en lämplig utvärdering har gjorts.
(3) Rådets förordning (EEG) nr 1210/90 av den 7 maj 1990 om inrättande av Europeiska miljöbyrån och Europeiska nätverket för miljöinformation och miljöövervakning[9] bör därför ändras.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Artikel 9.1 första meningen i förordning (EEG) nr 1210/90 skall ersättas med följande:
”1. Byrån skall ledas av en verkställande direktör som på förslag av kommissionen utnämns av styrelsen för en period av fem år, vilken period på förslag av kommissionen och efter det att en utvärdering har gjorts kan förlängas en gång, med högst fem år.
Inom ramen för utvärderingen skall kommissionen särskilt bedöma
- de resultat som har uppnåtts under den första mandatperioden och det sätt på vilket resultaten har uppnåtts, och
- byråns uppgifter och behov under de närmaste åren.”
Artikel 2
Denna förordning träder i kraft den […] dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning .
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
[pic] | EUROPEISKA GEMENSKAPERNAS KOMMISSION |
Bryssel den 11.3.2005
SEK(2005) 332 slutlig
Utkast till
GEMENSAMMA EES-KOMMITTÉNS BESLUT
om ändring av protokoll 31till EES-avtalet om samarbete inom särskilda områden vid sidan om de fyra friheterna
- Utkast till gemenskapens gemensamma ståndpunkt - (framlagt av kommissionen)
MOTIVERING
1. Protokoll 31 till EES-avtalet innehåller särskilda bestämmelser om samarbetet mellan gemenskapen och Eftastaterna i EES vid sidan om de fyra friheterna.
2. Syftet med bifogade utkast till beslut av Gemensamma EES-kommittén är att ändra i syfte att utvidga protokoll 31 samarbetet inom miljöområdet. Genom beslutet tillhandahålls en ram för samarbetet och anges formerna för hur Eftastaterna i EES kan delta i gemenskapens program och åtgärder på detta område genom införlivande av:
- 32002 D 1600 : Europaparlamentets och rådets beslut nr 1600/2002/EG av den 22 juli 2002 om fastställande av gemenskapens sjätte miljöhandlingsprogram.
3. Enligt artikel 1.3 b i rådets förordning (EG) nr 2894/94 rörande formerna för genomförandet av EES-avtalet skall rådet när det gäller denna typ av beslut fastställa gemenskapens ståndpunkt på förslag av kommissionen.
4. Utkastet till Gemensamma EES-kommitténs beslut överlämnas till rådet för godkännande. Kommissionen har för avsikt att lägga fram gemenskapens ståndpunkt i Gemensamma EES-kommittén så snart som möjligt.
Utkast till
GEMENSAMMA EES-KOMMITTÉNS BESLUT
om ändring av protokoll 31till EES-avtalet om samarbete inom särskilda områden vid sidan om de fyra friheterna
GEMENSAMMA EES-KOMMITTÉN HAR BESLUTAT FÖLJANDE
med beaktande av avtalet om Europeiska ekonomiska samarbetsområdet, ändrat genom protokollet med justeringar av avtalet om Europeiska ekonomiska samarbetsområdet, nedan kallat ”avtalet”, särskilt artiklarna 86 och 98 i detta, och
av följande skäl:
(1) Protokoll 31 till avtalet ändrades genom Gemensamma EES-kommitténs beslut nr ... av den .....[1].
(2) Samarbetet mellan parterna i avtalet bör utvidgas till att omfatta Europaparlamentets och rådets beslut nr 1600/2002/EG av den 22 juli 2002 om fastställande av gemenskapens sjätte miljöhandlingsprogram[2].
(3) Protokoll 31 till avtalet bör därför ändras så att detta utvidgade samarbete kan äga rum med verkan från och med den 1 januari 2005.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Följande skall läggas till i artikel 3.7 i protokoll 31 till avtalet:
”d) Gemenskapsrättsakter som skall gälla från och med den 1 januari 2005:
- 32002 D 1600 : Europaparlamentets och rådets beslut nr 1600/2002/EG av den 22 juli 2002 om fastställande av gemenskapens sjätte miljöhandlingsprogram (EUT L 242, 10.9.2002, s. 1.)’.
Artikel 2
Detta beslut träder i kraft dagen efter det att den sista anmälan enligt artikel 103.1 i avtalet har gjorts till Gemensamma EES-kommittén*.
Det skall tillämpas från och med den 1 januari 2005.
Artikel 3
Detta beslut skall offentliggöras i EES-delen av och EES-supplementet till Europeiska unionens officiella tidning .
Statistik över tekniska bestämmelser som anmälts under 2004 inom ramen för anmälningsförfarandet 98/34
Uppgifter från kommissionen i enlighet med artikel 11 i Europaparlamentets och rådets direktiv 98/34/EG om ett informationsförfarande beträffande tekniska standarder och föreskrifter och beträffande föreskrifter för informationssamhällets tjänster [1]
(2005/C 158/05)
(Text av betydelse för EES)
I. TABELL ÖVER DE OLIKA SLAGEN AV REAKTIONER RIKTADE MOT EG:S MEDLEMSSTATER AVSEENDE FÖRSLAG SOM ANMÄLTS AV VAR OCH EN AV DESSA
Medlemsstater | Anmäningar | Anmärkningar | Detaljerade yttranden | Förslag till gemenskapsrättsakter |
Medlemsstaterna | Kommissionen | EFTA | Medlemsstaterna | Kommissionen | 9.3 | 9.4 |
Belgien | 18 | 4 | 4 | | 3 | 4 | 0 | 0 |
Danmark | 40 | 8 | 19 | | 1 | 2 | 0 | 0 |
Tyskland | 99 | 40 | 46 | | 19 | 13 | 0 | 0 |
Spanien | 24 | 4 | 13 | | 3 | 2 | 0 | 0 |
Finland | 21 | 10 | 11 | | 2 | 3 | 0 | 0 |
Frankrike | 37 | 6 | 12 | | 2 | 2 | 0 | 0 |
Grekland | 34 | 7 | 33 | | 0 | 5 | 0 | 0 |
Irland | 6 | 1 | 2 | | 1 | 0 | 0 | 0 |
Italien | 28 | 20 | 10 | 1 | 10 | 5 | 0 | 0 |
Luxemburg | 4 | 1 | 2 | | 0 | 1 | 0 | 0 |
Nederländerna | 54 | 12 | 17 | | 7 | 3 | 0 | 0 |
Österrike | 50 | 8 | 10 | | 3 | 4 | 0 | 0 |
Portugal | 3 | 2 | 2 | | 0 | 1 | 0 | 0 |
Sverige | 23 | 6 | 8 | | 2 | 2 | 0 | 0 |
Förenade kungariket | 52 | 16 | 16 | | 1 | 6 | 1 | 0 |
Lettland | 13 | 11 | 5 | | 2 | 4 | 0 | 0 |
Malta | 2 | 1 | 1 | | 0 | 1 | 0 | 0 |
Cypern | 1 | 0 | 0 | | 0 | 1 | 0 | 0 |
Republiken Tjeckien | 14 | 7 | 6 | | 2 | 3 | 0 | 0 |
Ungern | 4 | 2 | 0 | | 0 | 0 | 0 | 0 |
Litauen | 4 | 4 | 4 | | 0 | 0 | 0 | 0 |
Estland | 0 | 0 | 0 | | 0 | 0 | 0 | 0 |
Slovenien | 12 | 2 | 1 | | 1 | 2 | 0 | 0 |
Polen | 8 | 5 | 3 | | 0 | 1 | 0 | 0 |
Slovakien | 6 | 1 | 4 | | 1 | 1 | 0 | 0 |
Totalt | 557 | 178 | 229 | 1 | 60 | 66 | 1 | 0 |
II. TABELL ÖVER FÖRDELNINGEN PER SEKTOR AV FÖRSLAG ANMÄLDA AV EG:S MEDLEMSSTATER
Sektor | BE | DK | DE | ES | FI | FR | GR | IE | IT | LU | NL | AT | PT | SE | UK | LT | MT | CY | CZ | HU | LV | EE | SI | PL | SK | EG totalt |
Byggnad och anläggning | 2 | 6 | 23 | 3 | 10 | 4 | | 1 | 2 | | 2 | 26 | | | 6 | | | | 1 | | | | 10 | | 1 | 97 |
Livsmedels och jordbruksprodukter | 6 | 5 | 6 | 6 | 1 | 10 | 1 | 2 | 13 | 1 | 11 | 7 | 1 | 4 | 17 | 4 | | | 4 | 2 | 3 | | 1 | 2 | 2 | 110 |
Kemiska produkter | 1 | 4 | 4 | 1 | | 1 | 1 | | 1 | | 3 | | | 2 | 2 | | | | | | 1 | | | | | 21 |
Läkemedelsprodukter | | | 4 | | 1 | 2 | | | | | | 1 | | 1 | 3 | | | | | | 1 | | | | | 13 |
Hem- och fritidsutrustning | 2 | | | 3 | | | | | | | | | 1 | 1 | | | | | 1 | | | | | 1 | | 9 |
Mekanik | 1 | 3 | | 3 | | 4 | | | 3 | | 4 | 1 | | 1 | 3 | | | | 1 | | 4 | | | | | 28 |
Energi, mineraler, trä | 1 | 2 | | 2 | 1 | | 1 | | 1 | | 5 | 2 | | 2 | | | | | | | 2 | | | 1 | | 20 |
Miljö, paketering | 1 | 2 | 6 | | 1 | 1 | | | 2 | | 8 | 3 | | 3 | 2 | | | | 5 | | 1 | | | 3 | | 38 |
Hälsovård, medicinsk utrustning | 1 | | | | | 3 | | | | | | | | 2 | | | | | | | | | | | | 6 |
Transport | 1 | 14 | 7 | 2 | 4 | 2 | | 3 | 1 | | 7 | 2 | | 5 | 16 | | 1 | | 1 | | | | | | | 66 |
Telekommunikationer | | 2 | 45 | 1 | 1 | 7 | 30 | | | | 6 | 3 | | 2 | 3 | | | | | | | | 1 | | 1 | 102 |
Övriga produkter | 2 | 2 | 2 | 1 | | 2 | 1 | | 1 | 1 | 4 | 2 | | | | | 1 | 1 | | 2 | 1 | | | 1 | 2 | 26 |
Informationssamhällets tjänster | | | 2 | 2 | 2 | 1 | | | 4 | 1 | 4 | 3 | 1 | | | | | | 1 | | | | | | | 21 |
Totalt per medlemsstat | 18 | 40 | 99 | 24 | 21 | 37 | 34 | 6 | 28 | 3 | 54 | 50 | 3 | 23 | 52 | 4 | 2 | 1 | 14 | 4 | 13 | | 12 | 8 | 6 | 557 |
III. TABELL ÖVER ANMÄRKNINGAR AVSEENDE FÖRSLAG ANMÄLDA AV ISLAND, LIECHTENSTEIN, NORGE [7] OCH SCHWEIZ [8]
Land | Anmälningar | EG-anmärkningar |
Island | 11 | 4 |
Liechtenstein | 3 | 2 |
Norge | 23 | 13 |
Schweiz | 15 | 9 |
Totalt | 52 | 28 |
IV. TABELL ÖVER FÖRDELNINGEN PER SEKTOR AV FÖRSLAG ANMÄLDA AV ISLAND, LIECHTENSTEIN, NORGE OCH SCHWEIZ
Sektor | Island | Liechtenstein | Norge | Schweiz | Totalt per sektor |
Byggnad och anläggning | | 1 | | | 1 |
Livsmedels- och jordbruksprodukter | 4 | 1 | 4 | 5 | 14 |
Kemiska produkter | | | 2 | 4 | 6 |
Läkemedelsprodukter | | | 1 | | 1 |
Hem- och fritidsutrustning | 2 | | | | 2 |
Mekanik | 1 | | 1 | 1 | 3 |
Miljö, paketering | 1 | | 1 | 1 | 3 |
Energi, mineraler, trä | | | 1 | | 1 |
Transport | 2 | | 9 | 2 | 13 |
Telekommunikationer | | | 2 | 2 | 4 |
Övriga produkter | 1 | | 1 | | 2 |
Informationssamhällets tjänster | | 1 | 1 | | |
Totalt per land | 11 | 3 | 23 | 15 | 52 |
V. TABELL ÖVER FÖRDELNINGEN PER SEKTOR FÖR ANMÄLDA FÖRSLAG FRÅN TURKIET OCH SYNPUNKTER PÅ DESSA FÖRSLAG
Turkiet | Sektorer | Synpunkter EG |
| Livsmedels- och jordbruksprodukter | 1 |
| Telekommunikation | 1 |
| Diverse produkter, textil | 1 |
Summa 3 | | 3 |
VI. TABELL ÖVER FÖRDELNINGEN PER SEKTOR FÖR ANMÄLDA FÖRSLAG FRÅN NYA MEDLEMSSTATER FÖRE UTVIDGNINGEN DEN 1 MAJ 2004 OCH SYNPUNKTER PÅ DESSA FÖRSLAG
Land | Sektorer | Synpunkter EG |
Malta | Energi, elektricitet | 1 |
Summa 1 | | 1 |
VII. STATISTIK ÖVER PÅGÅENDE ÖVERTRÄDELSEFÖRFARANDEN 2004 PÅ GRUNDVAL AV ARTIKEL 226 I EG-FÖRDRAGET SOM GÄLLER NATIONELLA TEKNISKA BESTÄMMELSER, SOM ANTAGITS I STRID MED BESTÄMMELSERNA I DIREKTIV 98/34/EG.
(Tabell över antalet överträdelseförfaranden per medlemsstat) |
Land | Antal |
Belgien | 2 |
Tyskland | 1 |
Spanien | 1 |
Frankrike | 1 |
Irland | 1 |
Italien | 4 |
Luxemburg | 1 |
Nederländerna | 1 |
Portugal | 2 |
EG totalt | 14 |
[1] Direktiv 98/34/EG av den 22 juni 1998 (EGT L 204, 21.7.1998) kodifierar direktiv 83/189/EEG med de förändringar som tillförts främst genom direktiv 88/182/EEG och 94/10/EG. För att kunna utvidga direktivets tillämpningsområde till att omfatta även informationssamhällets tjänster har det har ändrats genom direktiv 98/48/EG av den 20 juli 1998 (EGT L 217, 5.8.1998). Utvidgningen trädde i kraft den 5 augusti 1999.
[7] EES-avtalet (se not 4) föreskriver att det är nödvändigt att de EFTA-länder som anslutit sig till detta avtal anmäler förslag till tekniska bestämmelser till kommissionen.
[8] På grundval av det informella avtalet om informationsutbyte inom området för tekniska föreskrifter (se not 4) överlämnar Schweiz sina förslag till tekniska föreskrifter till kommissionen.
--------------------------------------------------
Offentliggörande av en ansökan om registrering i enlighet med artikel 6.2 i rådets förordning (EEG) nr 2081/92 om skydd för geografiska beteckningar och ursprungsbeteckningar
(2005/C 172/06)
Genom detta offentliggörande tillgodoses den rätt till invändningar som fastställs genom artiklarna 7 och 12d i ovan nämnda förordning. Alla invändningar mot ansökan skall göras genom den behöriga myndigheten i medlemsstaten, i ett WTO-land eller i ett tredjeland som godkänts i enlighet med artikel 12.3 inom sex månader efter detta offentliggörande, som sker av de motiv som anges nedan, särskilt punkt 4.6, genom vilka ansökan bedöms kunna godtas enligt förordning (EEG) nr 2081/92.
SAMMANFATTNING
RÅDETS FÖRORDNING (EEG) nr 2081/92
"ACEITE DE LA RIOJA"
EG-NUMMER: ES/00327/ 21.08.2003
SUB ( X ) SGB ( )
Denna sammanfattning har tagits fram i informationssyfte. För fullständig information, särskilt för nya producenter av de produkter som omfattas av den skyddade ursprungsbeteckningen eller den skyddade geografiska beteckningen i fråga, är det bäst att använda den fullständiga versionen av produktspecifikationen. Denna kan erhållas antingen hos nationella myndigheter eller hos Europeiska kommissionen [1].
1 Behörig myndighet i medlemsstaten:
Namn: | Subdirección General de Sistemas de Calidad Diferenciada – Dirección General de Alimentación Secretaría General de Agricultura y Alimentación del Ministerio de Agricultura, Pesca y Alimentación de España |
Adress: | Infanta Isabel, 1, E28071 Madrid |
Telefon: | +34-941 - 347 53 94 |
Fax: | +34-941 - 347 54 10 |
2. Grupp:
2.1.Namn: | "Asolrioja" Asociación de Trujales y Olivicultores de La Rioja |
2.2.Adress: | C/ Gran Vía, no 14, 8oA. Logroño La Rioja |
Tfn | 655 93 89 80 |
2.3.Sammansättning: | Producent/bearbetningsföretag (X) annan ( ) |
3. Produkttyp:
Extra jungfruolja: Klass 1.5: Oljor och fetter (smör, margarin, oljor etc.)
4. Produktspecifikation:
(Sammanfattning av kraven i artikel 4.2)
Namn: "Aceite de La Rioja"
Beskrivning:
Produkten utvinns ur olivträdets frukt (oliver) med helt mekaniska metoder eller processer, inklusive pressning, under förhållanden (särskilt temperatur) som inte medför förändringar i oljan. Oljan har en oklanderlig smak och oljans halt av fria fettsyror uttryckt i oljesyra överstiger inte 0,8 gram per 100 gram olja. I tillverkningen får inga lösningsmedel eller återförestring användas och oljan får inte på något sätt blandas med andra typer av oljor eller olivolja som utvunnits på annat sätt.
De skyddade oljorna är av typen extra jungfruolja och har ett klart utseende, utan tecken på slöja, grumlighet eller orenheter som stör klarheten. Oljan är grön med vissa nyanser som kan variera från intensivt ljusgrönt till intensivt mörkgrönt. Oljan har inga defekter och den har tillfredsställande positiva egenskaper. Den är fruktig i början av säsongen och har en mild mandelliknande smak utan bitterhet. Den är mjuk och lätt pepprig.
Efter mognaden har Aceite de La Rioja följande fysikalisk-kemiska egenskaper: syrahalt högst 0,8, UV-absorption (K 270), högst 0,20, UV-absorption (K 232) högst 2,50, peroxidvärde högst 15 mEq O2, fukthalt och flyktiga material efter torkning i ugn vid 105° C högst 0,1 %, föroreningar som är olösliga i petroleter högst 0,1 %, organoleptisk utvärdering, medianvärde för defekter (Md), Md = 0 och organoleptisk utvärdering, medianvärde för fruktighet (Mf), Mf %lt% 0.
Geografiskt område: Produktionsområdet sammanfaller med området för förvaring, utvinning och buteljering, och omfattar de 503388 hektar som utgör regionen Rioja.
Bevis på ursprung:
Gårdarna och/eller odlingarna, oljekvarnarna och buteljeringsanläggningarna inom det avgränsade område där råvaran kommer från och dit den förs för bearbetning, måste vara registrerade hos organisationen Asolrioja.
Dessa gårdar och odlingar, oljekvarnar och buteljeringsanläggningar måste ha ett internt kontrollsystem. Dessutom skall de genomgå extern kontroll som görs av ICAR (Instituto de Calidad Agroalimentaria de la Rioja) och/eller ett utomstående kontrollorgan som utses av organisationen Asolrioja. Detta skall vara godkänt av den behöriga myndigheten (Consejería de Agricultura, Ganadería y Desarrollo Rural del Gobierno de La Rioja) i fråga om uppfyllandet av normen UNE EN 45.004. På detta sätt intygas på ett opartiskt sätt att den skyddade extra jungfruoljan uppfyller kraven enligt förordningen och produktspecifikationen.
Varje gård och odling, olivkvarn och buteljeringsanläggning måste begära av organisationen att bli registrerad i kontrollsystemet. ICAR och/eller det auktoriserade utomstående kontrollorganet utvärderar produktionsenheten genom ett granskningsförfarande. Efter godkännande förs produktionsenheten in i organisationens register. Organisationen har ansvaret för underhållet av registret. Därefter fastställer ICAR och/eller det utomstående kontrollorganet ett granskningssystem och en rapport lämnas för utvärdering till ICAR. Om rapporten godkänns utfärdas en produktcertifiering om att endast extra jungfruolja som godkänts i alla steg av produktionsprocessen får saluföras med garanti om ursprung. Det skall också finnas ett samordningsråd som skall se till att organisationen, ICAR och/eller det auktoriserade utomstående kontrollorganet fungerar opartiskt.
Produktens spårbarhet garanteras genom märkning i varje produktions- och saluföringssteg.
Framställningsmetod:
Friska oliver, lämplig tidpunkt för skörd och de allt modernare bearbetningsteknikerna innebär att oliverna inom produktionsområdet är av god kvalitet, vilket är grunden för god kvalitet på den olja som utvinns ur dem. Olivträdets produktionsbelastning och grad av skugga anpassas till odlingarnas vegetativa stadium. Skörden genomförs alltid varsamt och endast friska oliver som har skördats direkt från trädet och har en lämplig mognadsgrad används för tillverkning av de skyddade olivoljorna.
Alla olivkvarnar och buteljeringsanläggningar har system för att se till att oliverna som är avsedda för tillverkning av extra jungfruoljan "Aceite de La Rioja" eller av denna olja och övriga hanteras separat för att undvika eventuella blandningar. Det finns även anpassade utrymmen för förvaring av oliverna eller den skyddade oljan före bearbetningen. Oliverna krossas högst 48 timmar efter skörden för att undvika att förändringar inträder som ger upphov till förhöjd syrahalt i oliverna. Under oljeutvinningen får temperaturen inte överstiga 30° C vid pressningen och 45° C vid centrifugeringen.
Blandningen får ta högst 60 minuter, temperaturen får stiga till högst 30° C och endast en cykel får genomföras.
Den extra jungfruoljan "Aceite de La Rioja" är aldrig raffinerad.
Oljan lagras i förhållanden som garanterar bästa hållbarhet, helst i behållare av rostfritt stål eller i oljepressar och/eller metallbehållare som invändigt är beklädda med keramiskt material, epoxihartser eller något annat inre material som lämpar sig för livsmedel. Behållarna är hermetiskt tillslutna och hålls vid en mild och konstant temperatur som inte får överskrida 22° C.
Oljan buteljeras endast när den uppfyller de fysikalisk-kemiska kraven enligt punkt 4.2 och har fått organoleptiskt godkännande av en provsmakningskommitté.
För att trygga kvaliteten och garantera produktens spårbarhet och kontrollen av den sker all produktion, mottagning, bearbetning och buteljering inom det avgränsade geografiska området.
Samband med området:
Historiskt samband: Olivoljan, idag ett uppskattat inslag i Medelhavskosten, har länge använts som födoämne i Rioja. Den har även använts för kosmetiska ändamål och massage. De fromma använde oljan i helgedomarnas lampor och för helande massage som gjordes i helgonens namn. Jordbrukarna i Rioja har i åratal använt krossade och smaksatta oliver som aperitif och mellanmål, konserverade i enbärslag med salt, timjan, vitlök och apelsinskal.
Romarna var dock de första i Rioja som utvann olja ur oliver genom pressning. Bevis på detta är den romerska motvikt som hittades i Murillo de Río Leza och en oljebehållare som hittades i ett oljepressningshus (torcularium) i Alfaro där man kan se två stora oljefläckar.
Det finns skriftliga hänvisningar ända från 1700-talet om olivodlingar i provinsen, de enda odlingar som reglerades av dekret, och om de oljepressar som användes. Enligt dessa källor fanns det i La Rioja 42 pressar som 1861 hade minskat till 39 för att 1945 ha ökat till 64 och 1953 till 81. Dessutom fanns en anläggning för utvinning av olja ur pressrester, fyra fabriker för industritvål och sex fabriker för vanlig tvål som tillverkades av olivolja. Under samma århundrade hade även Berceo stor betydelse, det vill säga den olja från La Rioja som exporterades till Väst- och Ostindien.
I verket Madoz, Diccionario Geográfico Estadístico Histórico de España y sus Posesiones de Ultramar konstateras att exporten av olivolja under åren 1846–1850 i Alfaro var viktig.
Samband med området: Olivodlingarna i La Rioja ligger huvudsakligen på brun mark med ett humusfattigt toppskikt och med en hög halt av kalksten, lera, gyttja och sand. Marken saknar ogenomträngliga skikt, vilket ger rätt sorts dränering och därmed begränsad tillväxt, särskilt under vilofasen. På så sätt uppnås rätt hormonbalans som inverkar på olivoljornas kvalitet genom att oliverna får en högre halt av olja, polyfenoler, antocyaner och aromer och ett lägre pH samt en lägre halt av äppelsyra, kalium och mindre grässmak. Om marken vore bördigare skulle träden växa för mycket och, vilket är särskilt negativt, fortsätta växa medan oliverna mognar, vilket skulle leda till att oliverna inte blir gröna i tid och inte hinner mogna tillräckligt. Problemen med skugga skulle dessutom vara större på grund av tätare bladverk, lummigare vegetation och fler kryptogamiska sjukdomar, vilket skulle leda till sämre kvalitet.
I det avgränsade geografiska området råder ett milt Medelhavsklimat med vissa inslag av kontinentalklimat med milda vintrar och långa varma somrar med lite nederbörd som ändå är tillräcklig för att odlingarna skall kunna utvecklas. Sommaren innebär mycket ljus och små temperaturvariationer mellan dag och natt, och i dessa idealiska förhållanden utvecklas oliverna på rätt sätt, med en ökning av oljehalten och aromen och en minskning av den totala syrahalten.
De låga temperaturerna under vinterdygnens kalla timmar behövs å andra sidan för att olivträdet skall kunna blomma och bära frukt. Under vintern vilar trädet utan blad och utan frukt, och det tål temperaturer på ned till -10° C. Efter vintervilan behöver olivträdet ljus och temperaturer på mellan 10 och 25° C för att utvecklas rätt. Det avgränsade områdets Medelhavsklimat tryggar tillräckligt med ljus och värme. Hettan blir dock inte så stark att fotosyntesen stoppas och bladen börjar vissna på grund av att vattenförsörjningen från rötterna inte räcker till för att kompensera avdunstningen från bladen.
Även den temperaturskillnad som normalt endast förekommer under olivernas mognadsperiod har en positiv inverkan på antocyanbildningen.
En annan mycket viktig faktor för en god skörd och därmed en god olivolja är olivodlarna, som genom sitt omsorgsfulla arbete och anpassade metoder tar vara på det som regionens natur har att erbjuda. Områdets olivodlare har ingående kunskaper om olivträd och använder traditionella odlingstekniker inriktade på balanserade olivlundar med tydlig inriktning på tillverkning av olivolja av hög kvalitet.
Namn: | Instituto de Calidad Agroalimentaria de La Rioja (ICAR) |
Adress: | Avda. de La Paz, 8–10, 26071, Logroño (La Rioja) |
Tfn | 941 29 16 00 |
Fax | 941 29 16 02 |
Märkning: Märkningen skall innehålla frasen "Denominación de origen Protegida Aceite de La Rioja".
- Lag 3/1982, av den 9 juni 1982, Estatuto de Autonomía de La Rioja (ändrad genom lagarna 3/1994 av den 24 mars 1994 och 2/1999 av den 7 januari 1999)
- Lag 3/1995 av den 8 mars 1995, Régimen Jurídico del Gobierno y la Administración Pública de la Comunidad Autónoma de La Rioja
- Lag 30/1992 av den 26 november, Régimen Jurídico de las Administraciones Públicas y del Procedimiento Administrativo Común
- Dekret av den 25 januari 1994 om fastställande av överensstämmelse mellan den spanska lagstiftningen och förordning (EEG) nr 2081/92 om skydd för geografiska och ursprungsbeteckningar för jordbruksprodukter och livsmedel
- Kungligt dekret nr 1643/1999 av den 22 oktober 1999 om handläggningsförfarandet för ansökningar om införande av gemenskapens register över skyddade ursprungsbeteckningar och skyddade geografiska beteckningar
[1] Europeiska kommissionen - Generaldirektoratet för Jordbruk - Kvalitetspolitik för jordbruksprodukter - B-1049 Bryssel.
--------------------------------------------------
Meddelande om att vissa antidumpningsåtgärder upphör att gälla
(2005/C 235/02)
Sedan kommissionen offentliggjort ett tillkännagivande om att åtgärdernas giltighetstid snart kommer att löpa ut [1] och inte mottagit någon begäran om översyn till följd av detta, tillkännager kommissionen härmed att de nedanstående antidumpningsåtgärderna snart kommer att upphöra att gälla. Detta meddelande offentliggörs i enlighet med artikel 11.2 i rådets förordning (EG) nr 384/96 [2] av den 22 december 1995 om skydd mot dumpad import från länder som inte är medlemmar i Europeiska gemenskapen.
Produkt | Ursprungs- eller exportland/länder | Åtgärd | Hänvisning | Utgångsdatum |
Flusspat | Folkrepubliken Kina | Antidumpningstull | Rådets förordning (EG) nr 2011/2000 (EGT L 241, 26.9.2000, s. 5) | 27.9.2005 |
[1] EGT C 309, 15.12.2004, s. 2.
[2] EGT L 56, 6.3.1996, s. 1. Förordning senast ändrad genom rådets förordning (EG) nr. 461/2004 (EGT L 77, 13.3.2004, s. 12)
--------------------------------------------------
Förlängning och ändring av bestämmelserna om allmän trafikplikt för regelbunden lufttrafik inom Grekland i enlighet med rådets förordning (EEG) nr 2408/92
(2005/C 266/02)
(Text av betydelse för EES)
1. I enlighet med artikel 4.1 a i rådets förordning (EEG) nr 2408/92 av den 23 juli 1992 om EG-lufttrafikföretags tillträde till flyglinjer inom gemenskapen har Grekland beslutat att från och med den 1 april 2006 förlänga och ändra de bestämmelser om allmän trafikplikt för regelbunden lufttrafik inom Grekland, som offentliggjordes i Europeiska gemenskapernas officiella tidning C 164 av den 10 juli 2002.
2. Ändringarna av den allmänna trafikplikten omfattar följande:
Minsta antal flygningar och minsta antal platser tillgängliga per vecka för följande sträckor:
- Athen–Κarpathos
- Athen–Sitia
- Thessaloniki–Korfu
Athen–Karpathos
Tre flygningar tur och retur per vecka, med sammanlagt 150 platser per vecka i båda riktningar under vinterhalvåret.
Sju flygningar tur och retur per vecka, med sammanlagt 350 platser per vecka i båda riktningar under sommarhalvåret.
Athen–Sitia
Tre flygningar tur och retur per vecka, med sammanlagt 90 platser per vecka i båda riktningar under vinterhalvåret.
Fyra flygningar tur och retur per vecka, med sammanlagt 120 platser per vecka i båda riktningar under sommarhalvåret.
Thessaloniki–Korfu
Tre flygningar tur och retur per vecka, med sammanlagt 180 platser per vecka i båda riktningar under vinterhalvåret.
Fyra flygningar tur och retur per vecka, med sammanlagt 240 platser per vecka i båda riktningar under sommarhalvåret.
--------------------------------------------------
Medlemsstaternas uppgifter om statligt stöd som beviljats med stöd av kommissionens förordning (EG) nr 70/2001 av den 12 januari 2001 om tillämpningen av artiklarna 87 och 88 i EG-fördraget på statligt stöd till små och medelstora företag
(2005/C 268/06)
(Text av betydelse för EES)
Stöd nummer: XS 125/03
Medlemsstat: Tyskland
Region: Sachsen-Anhalt
Stödordningens namn: Särskilt program för uppbyggnad av informationssamhället i Sachsen-Anhalt
- Landeshaushaltsordnung (LHO) vom 30.4.1991 (GVBl. LSA S. 45), insbesondere die Verwaltungsvorschriften zu § 44 LHO des Landes Sachsen-Anhalt;
- Verordnung (EG) Nr. 70/2001 der Kommission vom 12.1.2001 über die Anwendung der Artikel 87 und 88 EG-Vertrag auf staatliche Beihilfen an kleine und mittlere Unternehmen (ABl. L 10 vom 13.1.2002, S. 33) Stödordningens beräknade utgifter per år: C:a 2,5 miljoner EUR
— Investeringsbidrag
Stödnivån är begränsad till högst 50 % brutto (35 % brutto regionalstöd och 15 % brutto i tillägg för små och medelstora företag).
— Rådgivningsstöd
För utgifter för rådgivning från externa rådgivare till befintliga eller nya små och medelstora företag, samt till utgifter för genomförbarhetsstudier. Stödet begränsas till 50 % brutto av de stödberättigande utgifterna
Datum för genomförande: Från och med den 1 januari 2003
Stödordningens varaktighet: Till och med den 31 december 2004
- Ge stöd till små och mellanstora företag vid utveckling, tillämpning och användning av digital informations-, kommunikations- och medieteknologi.
- Förbättra konkurrensvillkoren för små och medelstora företag.
- Ge stöd till utveckling av regionala företagsnätverk inom teknologiorienterade branscher.
- Göra regionen attraktivare för företag.
- Ge impulser till ökad jämställdhet mellan kvinnor, män och missgynnade personer vid utbildning och på arbetsmarknaden
- Verksamheter i samband med produktion, bearbetning eller marknadsföring av de produkter som förtecknas i bilaga I till fördraget.
- Stöd till exportrelaterad verksamhet.
- Stöd som förutsätter att inhemska produkter används på bekostnad av importerade produkter.
- Stöd till stål-, syntetfiber-, motorfordons- och varvsindustrin.
Eftersom särskilda bestämmelser gäller för jordbruk, fiske och vattenbruk och det finns risk för att även små stödbelopp uppfyller kriterierna i artikel 87.1 i EG-fördraget, är dessa sektorer undantagna från stödet.
På grund av avtalen om lämpliga åtgärder på området för regionalt investeringsstöd är stål-, konstfiber-, motorfordons- och varvssektorerna också undantagna
Den beviljande myndighetens namn och adress Landesförderinstitut Sachsen-Anhalt
Gruppe Sonderprogramm
Domplatz 12
DE-39104 Magdeburg
Övriga upplysningar Ministerium für Wirtschaft und Arbeit
Referat 35
Hasselbachstraße 4
DE-39104 Magdeburg
--------------------------------------------------
Statligt stöd – Nederländerna
Statligt stöd nr C 35/2005 (f.d. N 59/2005)
Bredbandsutbyggnad i Appingedam
Uppmaning att inkomma med synpunkter enligt artikel 88.2 i EG-fördraget
(2005/C 321/07)
(Text av betydelse för EES)
Genom den skrivelse, daterad den 20.10.2005, som återges på det giltiga språket på de sidor som följer på denna sammanfattning, underrättade kommissionen Nederländerna om sitt beslut att inleda det förfarande som anges i artikel 88.2 i EG-fördraget avseende ovannämnda stödåtgärd.
Berörda parter kan inkomma med sina synpunkter på finansieringen av projektet för bredbandsutbyggnad i Appingedam inom en månad från dagen för offentliggörandet av denna sammanfattning och den därpå följande skrivelsen. Synpunkterna skall sändas till följande adress:
Europeiska kommissionen
Generaldirektoratet för konkurrens
Registreringsenheten för statligt stöd
Kontor SPA 3 06/05
B-1049 Bryssel
Fax: (32-2) 296 12 42
Synpunkterna kommer att meddelas Nederländerna. Den tredje part som inkommer med synpunkter kan skriftligen begära konfidentiell behandling av sin identitet, med angivande av skälen för begäran.
SAMMANFATTNING
Förfarande
I november 2004 lämnade kabeloperatören Essent in ett klagomål till kommissionen om den offentliga finansieringen av ett fiberaccessnät i Appingedam, Nederländerna. Essent hade redan i september 2004 väckt talan i en nederländsk domstol. Domstolen förpliktade kommunen att anmäla planerna att bevilja stöd till kommissionen och att avbryta den fortsatta utbyggnaden av nätet [1]. I februari 2005 anmälde de nederländska myndigheterna åtgärden till kommissionen, men hävdade samtidigt att det inte var fråga om stöd. Kommissionen begärde ytterligare upplysningar från de nederländska myndigheterna i mars 2005. Myndigheterna svarade i augusti 2005 efter en förlängning av tidsfristen.
Beskrivning av åtgärden
Appingedams kommun anser att det krävs offentliga insatser för att förbättra det otillräckliga utbudet av avancerade bredbandstjänster till företag och allmänhet genom att stödja utbyggnad av ett fiberaccessnät (Fibre to the Home, FTTH). Kommunen beslutade att delta i finansieringen av projektet, eftersom marknadsaktörerna inte visat något intresse för att delta i projektet på marknadsvillkor.
Det planerade fibernätet är uppdelat i en passiv och en aktiv del. Den passiva delen kommer att ägas och finansieras av en offentlig stiftelse som kommunen kommer att bilda och kontrollera. Den aktiva delen kommer att ägas och finansieras av en enhet som bildas av privata investerare (Damsternet). Damsternet självt kommer endast att tillhandahålla grossisttjänster till tjänsteleverantörer som tillhandahåller bredbandstjänster till slutkunder (hushåll och företag).
Bedömning av åtgärden
Det är fråga om statliga medel eftersom den passiva delen av nätet finansieras av Appingedams kommun. Stiftelsen, Damsternet och de tjänsteleverantörer som levererar till slutkunder får en ekonomisk fördel, eftersom de kommer att tillhandahålla och ha tillgång till infrastruktur på villkor som är mer förmånliga än marknadsvillkoren. Den statliga åtgärden snedvrider konkurrensen, eftersom den ändrar de gällande marknadsvilkoren genom att möjliggöra inträde på grossistmarknaden för snabba bredbandstjänster (Damsternet) och genom att ge tjänsteleverantörer möjlighet att gå in på marknaderna i efterföljande led, dvs. tillhandahållande av bredbands- och teletjänster till slutkunder. Denna statliga åtgärd påverkar handeln mellan medlemsstater, eftersom den kan påverka leverantörer av elektroniska kommunikationstjänster i andra medlemsstater.
En bedömning av åtgärdens förenlighet med den gemensamma marknaden kan endast göras på grundval av artikel 87.3 c i EG-fördraget. Enligt den artikeln skall åtgärden vara nödvändig och proportionerlig för att främja genomförandet av ett mål av gemensamt intresse, dvs. att avhjälpa ett marknadsmisslyckande eller att uppnå ett godkänt mål som syftar till sammanhållning eller omfördelning.
Nödvändighet och proportionalitet
Bredbandsanslutning är en typ av tjänst som kan påverka produktiviteten och tillväxten. I andra fall har kommissionen funnit att stöd till infrastruktur kan vara ett lämpligt och proportionerligt instrument för att angripa marknadsmisslyckanden och rättviseproblem. Även det nu aktuella projektet har vissa av de egenskaper som har bedömts positivt i tidigare kommissionsbeslut om offentlig finansiering av bredbandsprojekt (öppen anbudsinfordran, allmän access osv.). Eftersom FTTH-nätens tekniska egenskaper gör det möjligt att tillhandahålla mer avancerade tjänster än genom traditionella koppar- eller kabelnät [2], skulle man kunna hävda att statligt stöd är ett lämpligt sätt att påskynda innovationstakten, även om det innebär att den privata sektorns redan gjorda investeringar riskeras och att den privata sektorn avskräcks från att investera i framtiden.
Kommissionen har hittills bara godkänt ärenden där marknaden inte tillhandahöll ett konkurrenskraftigt utbud av bredbandstjänster. I detta ärende är det fråga om en åtgärd som görs i ett område där bredbandstjänster till slutkund (KPN och Essent) och i viss mån även infrastruktur för att tillhandahålla grossistjänster (KPN) redan finns tillgängliga till priser som är jämförbara med priserna i andra regioner. Det finns en stor överlappning med befintliga nät när det gäller nättäckning och tjänstevillkor och det finns därför en stor risk för att en statlig åtgärd skulle tränga ut marknadsaktörernas nuvarande och framtida investeringar.
Kommissionen har beslutat att inleda förfarandet enligt artikel 88.2 i EG-fördraget om den omstridda åtgärden, eftersom kommissionen inte är övertygad om att åtgärden är förenlig med den gemensamma marknaden i enlighet med artikel 87.3 c i EG-fördraget.
Enligt artikel 14 i rådets förordning (EG) nr 659/1999 kan allt olagligt stöd komma att återkrävas från mottagaren.
SJÄLVA SKRIVELSEN
%quot%Met dit schrijven stelt de Commissie Nederland ervan in kennis dat zij, na onderzoek van de door uw autoriteiten verstrekte inlichtingen betreffende bovengenoemde steunmaatregel, heeft besloten de procedure van artikel 88, lid 2, van het EG-Verdrag in te leiden.
I. Procedure
1. Bij schrijven van 2 november 2004 (dat op 18 november 2004 geregistreerd werd onder nummer CP 212/2004) diende kabelexploitant Essent Kabelcom (hierna: Essent), een informele klacht in bij de Commissie. De klacht betreft overheidsfinanciering voor een glasvezelaansluitnetwerk (Fibre-to-the-Home, FTTH) in Appingedam, een stad in Noord-Nederland. Essent heeft intussen bevestigd dat de klacht als een formele klacht dient te worden beschouwd.
2. Essent, die de op een na grootste kabelexploitant van Nederland is en die ook een kabelnetwerk in Appingedam exploiteert, had de zaak in september 2004 al aanhangig gemaakt bij een Nederlandse rechtbank. De rechtbank heeft de gemeente op grond van artikel 88, lid 3, EG-Verdrag opgedragen het steunvoornemen aan te melden bij de Commissie en de verdere aanleg van het netwerk te staken.
3. Bij een schrijven dat op 3 februari 2005 werd geregistreerd, meldden de Nederlandse autoriteiten de maatregel bij de Commissie aan om redenen van rechtszekerheid, waarbij ze aanvoerden dat de maatregel geen steun behelsde. Op 31 maart 2005 verzocht de Commissie de Nederlandse autoriteiten om verdere informatie. Na een verlenging van de termijn antwoordden zij hierop bij brief van 4 augustus 2005, die op 16 augustus 2005 werd geregistreerd. De informatie in deze brief verschilt aanzienlijk van de informatie die bij de oorspronkelijke aanmelding werd verstrekt.
II. Uitvoerige beschrijving van de maatregel
Achtergrond
4. De gemeente Appingedam vindt dat de tussenkomst van de overheid nodig is om te voorzien in de algemene beschikbaarheid van geavanceerde breedbanddiensten voor ondernemingen en particulieren door uitrol van een glasvezelaansluitnetwerk (Fibre-to-the-Home, FTTH) in Appingedam te steunen. Volgens de gemeente bieden Essent en telecommunicatie-exploitant KPN in Appingedam weliswaar internettoegang maar geen geavanceerde breedbanddiensten. De gemeente heeft besloten financieel deel te nemen in het project nadat gebleken was dat de marktpartijen geen belangstelling hadden om hierin op marktvoorwaarden deel te nemen.
De componenten van het netwerk
5. De passieve laag van het glasvezelnetwerk (graafrechten, buizen, glasvezels, enz.) zal het eigendom worden van een openbare stichting (%quot%Stichting Glasvezelnet Appingedam%quot%, hierna: de stichting), op te richten door en onder toezicht van de gemeente. De investering in de passieve laag wordt op 4,9 miljoen EUR geschat. Aanvankelijk was niet voorzien dat de aanleg van de passieve laag openbaar zou worden aanbesteed. Er is evenwel besloten, zoals in de brief van 4 augustus 2005 wordt verklaard, om dit wel te doen.
6. De kosten van de actieve laag (telecommunicatieapparatuur, netwerkbeheer, enz.) worden op 1 tot 1,3 miljoen EUR geschat. De actieve componenten hebben een geschatte economische levensduur van 5 tot 8 jaar. De exploitant van de actieve laag zal alleen wholesale-diensten aanbieden aan service providers die breedbanddiensten aan de eindgebruikers (huishoudens en bedrijven) zullen verstrekken.
7. De autoriteiten verklaarden aanvankelijk dat de actieve laag eigendom zou worden van en gefinancierd zou worden door een entiteit (%quot%Stichting Damsternet%quot%, hierna: Damsternet) die door bepaalde particuliere investeerders zou worden opgericht. Niet alle particuliere partijen waren bekend. Volgens de autoriteiten hebben NKF (een kabelfabrikant), Nacap (de pijpleidingdivisie van een internationaal actieve bouwonderneming, genaamd Koop Holding) en Ericsson Telecommunications belangstelling getoond. In de brief van 4 augustus 2005 hebben de autoriteiten evenwel verklaard dat de gemeente het gebruiksrecht van het actieve netwerk uiteindelijk openbaar zou aanbesteden. In dit stadium is het bovendien niet duidelijk op basis van welke financiële voorwaarden het gebruiksrecht zou worden gegund. In de concept-gebruiksovereenkomst wordt bepaald dat de houder van het gebruiksrecht jaarlijks een gebruiksvergoeding aan de stichting zal betalen. De stichting zal echter %quot%maximaal een bedrag opeisen dat overeenkomt met 80 % van de in dat jaar gegenereerde cashflow%quot%. Indien deze cashflow negatief is, zal de stichting geen vergoeding opeisen. In een dergelijk geval zullen zij slechts een minimale betaling verlangen, zoals aangegeven in een bijlage bij de gebruiksovereenkomst. In de bijlage wordt evenwel nog niet bepaald welke betaling voorzien is.
III. Het standpunt van de Nederlandse autoriteiten
8. De Nederlandse autoriteiten stellen dat er geen sprake is van een steunmaatregel en voeren hiervoor verschillende argumenten aan.
9. Allereerst beroepen zij zich op een %quot%marktfalen%quot%, d.w.z. dat de markt niet de diensten verschaft die door de autoriteiten essentieel worden geacht voor de bevolking. Marktinvesteerders zijn niet bereid om in het project te investeren omdat het geen marktconform financieel rendement zou opleveren. Doordat de markt niet in het project investeert, ziet Appingedam zich genoodzaakt dit glasvezelnetwerk aan te leggen als een %quot%publieke infrastructuur%quot%. De Nederlandse autoriteiten voeren daarom aan dat de gemeente Appingedam enkel steun verleent voor de aanleg van een %quot%publieke infrastructuur%quot% die voor alle partijen openstaat op vergelijkbare voorwaarden.
10. In de tweede plaats betogen de autoriteiten dat er geen steun gemoeid is met dit project op de vier niveaus die daarbij kunnen worden onderscheiden. Er is geen sprake van een voordeel voor de stichting en zelfs wanneer dat het geval zou zijn, zou dat niet van invloed zijn op het handelsverkeer tussen de lidstaten. Er wordt ook geen steun verleend aan de exploitant van de actieve laag. De Commissie merkt op dat de autoriteiten evenwel geen argumenten aanvoeren om deze beweringen te staven. Voorts zijn de autoriteiten van mening dat er geen steun wordt verleend aan de dienstenaanbieders. De exploitant zou een marktconforme wholesale-prijs moeten aanrekenen aan de providers die retail-diensten aanbieden die zij reeds via bestaande infrastructuur aanboden. Indien de Commissie garanties van de gemeente zou verlangen dat de exploitant marktconforme prijzen aanrekent, zal de gemeente dit vastleggen in de overeenkomst tussen de stichting en de exploitant. Tenslotte betogen de autoriteiten dat, in tegenstelling tot de zaak ATLAS [3], het netwerk in Appingedam hoofdzakelijk zou worden gebruikt om diensten te verlenen aan huishoudens/particulieren die geen economische activiteiten verrichten. Voorzover er sprake is van steun aan ondernemingen in Appingedam, blijft deze onder de toegestane steunintensiteit die is vastgelegd in Verordening (EG) nr. 69/2001 (%quot%de minimis-steun%quot%) en bovendien valt deze onder de kaderregeling voor steun aan kleine en middelgrote ondernemingen (MKB).
11. De Nederlandse autoriteiten betogen dat indien de Commissie tot de conclusie komt dat de maatregel steun vormt, de maatregel verenigbaar is omdat deze zowel noodzakelijk als evenredig is. De maatregel is nodig omdat particuliere investeerders niet willen investeren in Appingedam, een perifeer gebied met een sociaal-economische achterstand. Voor zover er breedbanddiensten beschikbaar zijn, zijn de huidige prijzen ervan hoger dan in andere gebieden van Nederland. Aangezien alle exploitanten open toegang tot het netwerk zullen krijgen op gelijke voorwaarden, is de mededinging gewaarborgd en zal geen enkele exploitant een selectief voordeel genieten. De autoriteiten stellen ook dat de maatregel evenredig is. De stichting is niet betrokken bij de exploitatie van de actieve laag. De operator zal een niet-discriminerende, open toegang bieden en niet met dienstenaanbieders concurreren. De aanleg van het netwerk zal plaatsvinden op marktvoorwaarden.
IV. Beoordeling van de maatregel/steun
12. Op grond van het Verdrag en geconsolideerde rechtspraak is er sprake van staatssteun in de zin van artikel 87, lid 1, wanneer door overheidsbemoeienis of door met staatsmiddelen bekostigde maatregelen een voordeel wordt verleend aan de begunstigde, welke de mededinging vervalst of dreigt te vervalsen en het handelsverkeer tussen de lidstaten ongunstig dreigt te beïnvloeden.
Staatsmiddelen
13. De gemeente Appingedam zal ofwel een lening ofwel een garantie voor een lening verstrekken. Bijgevolg zijn de middelen voor de financiering van de passieve laag van dit netwerk afkomstig van de gemeente Appingedam. Deze middelen moeten daarom als staatsmiddelen worden beschouwd.
Economisch voordeel
14. De autoriteiten hebben verschillende argumenten aangevoerd als zou de maatregel geen steun behelzen, ofwel omdat deze geen voordeel meebrengt ofwel omdat deze niet van invloed is op het handelsverkeer tussen de lidstaten. Op deze argumenten zal hierna worden ingegaan.
15. Volgens de Nederlandse autoriteiten valt een dergelijke vorm van overheidsbemoeienis niet onder artikel 87, lid 1, EG-Verdrag, maar dient deze veeleer te worden gezien als een typische overheidstaak, aangezien algemene infrastructuur wordt aangelegd.
16. De Commissie is echter niet overtuigd dat dit project kan worden beschouwd als het verschaffen van een algemene infrastructuur. Overeenkomstig de bevindingen van de Commissie in de zaak ATLAS [4] bieden het passieve netwerk en de actieve componenten geen dienst aan eindgebruikers, maar voorzieningen voor bedrijven die breedbanddiensten aanbieden. Zoals uit de aanwezigheid van KPN en Essent in Appingedam blijkt, is het verschaffen van dit soort infrastructuur geen typische overheidstaak, maar een activiteit die gewoonlijk wordt verricht door marktpartijen die de uiteindelijke dienst aan huishoudens en bedrijven verstrekken. Het project overlapt daarmee tot op zekere hoogte marktinitiatieven of voorziet in de verstrekking van diensten die al beschikbaar zijn, hoewel de door de stichting aan te leggen infrastructuur graafwerkzaamheden en passieve elementen behelst. De Commissie is derhalve in dit stadium van mening dat het project in Appingedam onder de staatssteunregels valt en niet als algemene infrastructuur kan worden aangemerkt die tot de gewone verantwoordelijkheden van de staat jegens de bevolking behoort.
Voordeel voor de stichting
17. De stichting die eigenaar is van de passieve infrastructuur, is opgericht door de gemeente en staat onder haar toezicht. De stichting stelt de passieve laag ter beschikking van de exploitant. Dit kan als een economische activiteit worden beschouwd en de stichting kan derhalve worden aangemerkt als een onderneming in de zin van artikel 87, lid 1, EG-Verdrag. De passieve laag wordt door de gemeente gefinancierd zonder enige vergoeding van de stichting. Dit komt neer op een economisch voordeel voor de stichting in de zin van artikel 87, lid 1, EG-Verdrag.
Voordeel voor de exploitant
18. De bewering dat er geen steun wordt verleend aan de exploitant, wordt niet door de autoriteiten gestaafd.
19. De autoriteiten hebben bevestigd dat het gebruiksrecht openbaar zal worden aanbesteed. Indien dat gebeurt, kan de aanbesteding in principe het economische voordeel voor de winnende leverancier tot een minimum worden beperkt in de zin van artikel 87, lid 1, EG-Verdrag. Het valt evenwel te betwijfelen of de passieve laag op dezelfde voorwaarden zal worden aangelegd als bij een particuliere investering. Volgens de autoriteiten kon het project niet door particuliere investeerders worden uitgevoerd en waren banken evenmin bereid om geld te steken in dit project. De gemeente heeft verschillende banken gevraagd om dit project te financieren, maar met uitzondering van de Bank Nederlandse Gemeenten (BNG) hebben zij dit allemaal geweigerd. BNG is bereid de gemeente een lening te verstrekken omdat zij, aldus de gemeente, alleen de kredietwaardigheid van de begunstigde van de lening, in casu de gemeente, maar niet de aanleg van het FTTH-netwerk door de stichting of het project als zodanig heeft beoordeeld.
Voordeel voor internetaanbieders (ISP's) en andere aanbieders van elektronische communicatiediensten
20. Zelfs wanneer de toegang tot het optische netwerk via de exploitant op transparante en gelijke voorwaarden aan alle geïnteresseerde ISP's en andere exploitanten zal worden verleend, zal de tarifering van deze toegang waarschijnlijk ruim onder de onderliggende kosten liggen als gevolg van de overheidsbemoeienis en niet gebaseerd zijn op de markttarieven voor vergelijkbare wholesale-breedbanddiensten. De dienstenaanbieders zal daarom een voordeel worden verleend aangezien zij de kans krijgen om tot de markt voor snelle retail-breedbanddiensten toe te treden en bedrijfsactiviteiten te ontwikkelen tegen voorwaarden die anders niet op de markt kunnen worden verkregen.
Voordeel voor de eindgebruikers
21. Het voorgaande suggereert dat het voordeel dat aan de exploitant, dienstenaanbieders en andere aanbieders van telecommunicatiediensten wordt verleend, zich ook zou kunnen vertalen in een voordeel voor de huishoudens en ondernemingen in Appingedam. Particuliere gebruikers vallen niet onder de staatssteunregels. Echter ondernemingen in het beoogde gebied zouden wellicht kunnen profiteren van een dienstverlening die verder reikt en lager geprijsd is dan wat op louter commerciële basis zou worden aangeboden gezien de huidige aanbiedingen voor huurlijnen en satellietverbindingen. Bovendien zouden zij een voordeel kunnen genieten in vergelijking met bedrijven in andere regio's van Nederland. De autoriteiten hebben bij herhaling aangevoerd dat, indien er sprake is van steun voor ondernemingen in Appingedam, het steunniveau onder de toegestane steunintensiteit ligt, zoals bepaald bij Verordening (EG) nr. 69/2001 (%quot%de minimis-steun%quot%), en dat de maatregel bovendien onder de kaderregeling inzake overheidssteun voor kleine en middelgrote ondernemingen (KMO's) valt. De Commissie erkent dat het voordeel voor elk van de zakelijke eindgebruikers onder de drempel voor de minimis-steun zou kunnen liggen. Er kan in dit stadium echter niet worden uitgesloten dat de steun wel de in deze verordening vastgelegde plafonds overschrijdt.
Concurrentievervalsing
22. Door deze tussenkomst van de overheid worden de bestaande marktvoorwaarden in Appingedam gewijzigd doordat de gesubsidieerde toegang van de exploitant tot de wholesale-markt voor snelle breedbanddiensten alsmede de toegang van dienstenaanbieders tot de downstream-markten van onder andere retail-breedband- en retail-telecommunicatiediensten mogelijk wordt gemaakt. De bestaande exploitanten, Essent en KPN, hebben bij hun beslissingen inzake infrastructuurinvesteringen en -onderhoud, hun berekeningen gebaseerd op de veronderstelling dat andere exploitanten de kosten van nieuwe infrastructuur zouden moeten dragen of een marktprijs zouden moeten betalen voor de toegang tot wholesale-diensten, hetgeen niet langer het geval lijkt te zijn als er overheidssteun wordt verleend. Het feit dat er nieuwe infrastructuur beschikbaar komt tegen voorwaarden die op het eerste gezicht niet marktconform zijn, heeft tot gevolg dat de concurrentie wordt vervalst, ook op de downstream-markten van retail-breedband- en andere retail-elektronische communicatiediensten.
Gevolgen voor het handelsverkeer
23. Voor zover de overheidsmaatregelen gevolgen kunnen hebben voor telecommunicatiebedrijven en dienstenaanbieders in andere lidstaten, zijn deze van invloed op het handelsverkeer. De telecommunicatiemarkt staat steeds meer open voor concurrentie tussen exploitanten en dienstenaanbieders, die zich over het algemeen bezighouden met activiteiten waarvoor handelsverkeer bestaat tussen de lidstaten.
Conclusie
24. In het licht van het voorgaande is de Commissie van mening dat het met staatsmiddelen gefinancierde project een economisch voordeel verleent aan de stichting, de exploitant en de dienstenaanbieders, hetgeen zich tenminste ten dele zou kunnen vertalen in een economisch voordeel voor ondernemingen in Appingedam. Voorts is het project concurrentievervalsend en van invloed op het handelsverkeer tussen de lidstaten.
V. Beoordeling van de steunmaatregel: verenigbaarheid
25. Na de vaststelling dat er sprake is van staatssteun in de zin van artikel 87, lid 1, van het EG-Verdrag, dient te worden nagegaan of de maatregel verenigbaar met de gemeenschappelijke markt kan worden geacht.
26. Wanneer staatsmiddelen enkel worden verleend ter compensatie van de verstrekking van een dienst van algemeen economisch belang (hierna: DAEB), dan hoeft hiermee geen staatssteun te zijn gemoeid. Het Hof van Justitie heeft te kennen gegeven dat de compensatie van kosten die voortvloeien uit openbare dienstverplichtingen, niet onder de werkingssfeer van artikel 87, lid 1, van het Verdrag vallen indien aan een aantal voorwaarden is voldaan. Deze voorwaarden worden beschreven in het Altmark-arrest van 24 juli 2003 [5]. De autoriteiten hebben zich evenwel niet beroepen op de voorwaarden die zijn vastgelegd in het Altmark-arrest en hebben evenmin het bestaan van een DAEB aangevoerd, zelfs niet impliciet. Er zijn geen aanwijzingen dat de overheidsmaatregel moet worden beschouwd als compensatie voor de diensten die door de begunstigde ondernemingen worden verstrekt. Daarom heeft de Commissie in dit stadium de aangemelde maatregel niet bezien tegen deze achtergrond of getoetst aan het bepaalde in artikel 86, lid 2, van het EG-Verdrag.
27. De Commissie merkt op dat met het voorgenomen project wordt beoogd de ruime beschikbaarheid en het ruime gebruik van snelle breedbanddiensten te verzekeren tegen voorwaarden die meer overeenkomen met minder afgelegen gebieden die dichter bevolkt zijn en relatief meer bedrijven tellen. Voorts wordt erkend dat de bestaande kaderregelingen en richtsnoeren niet kunnen worden toegepast voor de beoordeling van steunmaatregelen die dit specifiek tot doel hebben. De Commissie is derhalve van mening dat de toetsing van de verenigbaarheid van de maatregel met de gemeenschappelijke markt rechtstreeks op artikel 87, lid 3, onder c), van het EG-Verdrag dient te worden gebaseerd [6].
28. In artikel 87, lid 3, onder c), EG-Verdrag wordt bepaald dat:
%quot%steunmaatregelen om de ontwikkeling van bepaalde vormen van economische bedrijvigheid of van bepaalde regionale economieën te vergemakkelijken, mits de voorwaarden waaronder het handelsverkeer plaatsvindt daardoor niet zodanig worden veranderd dat het gemeenschappelijke belang wordt geschaad, als verenigbaar met de gemeenschappelijke markt kunnen worden beschouwd%quot%.
29. In het kader van een toetsing aan artikel 87, lid 3, onder c), van het EG-Verdrag houdt dit in dat de overheidsmaatregel noodzakelijk moet zijn en in verhouding dient te staan tot het beoogde doel van algemeen belang, d.w.z. de correctie van een gebrekkige marktwerking.
Noodzakelijkheid
30. De toegang tot een breedbandnetwerk is een voorziening die door zijn aard een positieve invloed kan hebben op de productiviteit en de groei van een groot aantal sectoren en activiteiten [7]. Er zijn aanwijzingen dat een grotere beschikbaarheid van breedbandnetwerken ten goede kan komen aan de regionale economische ontwikkeling en de schepping en het behoud van werkgelegenheid, alsook verbeterde gezondheids- en onderwijsvoorzieningen [8].
31. De autoriteiten stellen dat de maatregel gericht is tegen een gebrekkige marktwerking: Appingedam is een achterstandsgebied waar de netwerkeigenaren Essent en KPN niet hun netwerken willen upgraden noch toegang willen verlenen tot hun core-netwerken of %quot%dark fibre%quot% aan providers die FTTH willen aanbieden. De autoriteiten hebben ook verklaard dat Essent en KPN pas na de aankondiging van de gemeente dat zij haar eigen FTTH-initiatief zou lanceren, hun netwerken hebben geüpgraded teneinde breedbanddiensten aan te bieden.
32. Het is evenwel de vraag of er bij de situatie in Appingedam wel sprake is van een %quot%gebrekkige marktwerking%quot%. In de eerste plaats voorziet de markt, aldus de autoriteiten, niet in de FTTH-infrastructuur omdat het verwachte rendement op de investering onvoldoende was om een investering tegen marktvoorwaarden te rechtvaardigen. Dit kan worden verklaard door een lage vraag naar breedbanddiensten alsook de hoge kapitaaluitgaven voor de aanleg van de infrastructuur.
33. In de tweede plaats is, aldus de Commissie, de toegang tot een breedbandnetwerk al beschikbaar in Appingedam hoewel de diensten die thans worden verstrekt, niet geheel vergelijkbaar zijn met de diensten die met het geplande netwerk zouden kunnen worden aangeboden. KPN en Essent bieden allebei retail-breedbanddiensten aan tot 8Mbit/s en KPN biedt tot op zekere hoogte ook wholesale-toegang tot infrastructuur en diensten. Bijgevolg is er een aanzienlijke overlapping van netwerkdekking en dienstverlening, die tot de beste in de Europese Unie behoren, en daarom valt het te betwijfelen of er sprake is van een %quot%marktfalen%quot%, die met deze maatregel kan worden verholpen.
Evenredigheid
34. Om te bepalen of de maatregel verenigbaar is met de gemeenschappelijke markt, dient ook de evenredigheid van de maatregel te worden onderzocht. De maatregel dient in verhouding te staan tot het beoogde doel en mag de concurrentie niet zo zeer vervalsen dat het gemeenschappelijke belang wordt geschaad.
35. Er dient te worden erkend dat de technische kenmerken van bijvoorbeeld glasvezelaansluitnetwerken verschillen van de bestaande kabel- en telecommunicatienetwerken in Appingedam. Er kan worden aangevoerd dat de nieuwe generatie netwerken niet te vergelijken valt met de bestaande netwerken omdat zij andere en veel geavanceerdere diensten mogelijk maken dan de bestaande netwerken. Volgens degenen die zich hierop beroepen kan overheidssteun voor de volgende generatie van openbaar toegankelijke, lokale aansluitnetwerken een positief effect hebben op de economische ontwikkeling vanwege de positieve externe effecten die deze netwerken zullen hebben op innovatie en groei. Bovendien hebben de bestaande exploitanten van elektronische communicatienetwerken (nog) niet in deze infrastructuur geïnvesteerd vanwege de hoge kapitaaluitgaven en omdat hun bestaande investeringen daardoor niet meer van nut zouden zijn. Wanneer deze redenering wordt doorgetrokken, zou staatssteun voor de nieuwe generatie netwerken een gewenst middel kunnen zijn om het tempo van innovatie en economische ontwikkeling te versnellen, zelfs tegen de prijs dat in het verleden gedane investeringen mogelijk worden ondermijnd en toekomstige investeringen ontmoedigd.
36. In dit stadium valt evenwel moeilijk te bezien welke toepassingen of diensten aan particulieren en bedrijven kunnen worden aangeboden die niet met behulp van breedbanddiensten via de bestaande netwerken kunnen worden verschaft. Dit betekent dat er sprake is van een hoge substitueerbaarheid tussen enerzijds de retail en wholesale-diensten die via het geplande FTTH-netwerk worden verstrekt en anderzijds de diensten die via de bestaande netwerken worden verstrekt, waardoor de maatregel de mededinging in de nabije toekomst ernstig zou kunnen vervalsen. Dit geldt des te meer in het licht van een aantal geplande ontwikkelingen. KPN heeft aangekondigd dat zij de capaciteit van haar dienstverlening zal verhogen en Essent onderzoekt de mogelijkheid om de superbreedbandverbinding ETTH (Ethernet to the home) via haar bestaande netwerken aan te bieden, waardoor de capaciteit van haar netwerk aanzienlijk wordt vergroot. De maatregel die door de autoriteiten wordt voorzien, houdt daarom een ernstig risico in van verdringing van bestaande en toekomstige investeringen door marktpartijen als gevolg van de overheidssteun. Onder de gegeven omstandigheden is het daarom de vraag of de geplande maatregel en het gebruik als zodanig van het steuninstrument als evenredig kunnen worden beschouwd.
Conclusie
37. Op grond van het voorgaande en de informatie die in dit stadium beschikbaar is, betwijfelt de Commissie of de betwiste maatregel verenigbaar is met de gemeenschappelijke markt in overeenstemming met artikel 87, lid 3, onder c), van het EG-Verdrag.
VI. Besluit
38. In het licht van het voorgaande heeft de Commissie besloten de procedure van artikel 88, lid 2, van het EG-Verdrag in te leiden ten aanzien van de betwiste maatregel omdat zij betwijfelt of deze verenigbaar is met de gemeenschappelijke markt in overeenstemming met artikel 87, lid 3, onder c), van het EG-Verdrag.
Gelet op de bovenstaande overwegingen verzoekt de Commissie Nederland in het kader van de procedure van artikel 88, lid 2, van het EG-Verdrag binnen een maand vanaf de datum van ontvangst van dit schrijven zijn opmerkingen te maken en alle dienstige inlichtingen te verstrekken voor de beoordeling van de steunmaatregel. Zij verzoekt uw autoriteiten onverwijld een afschrift van deze brief aan de potentiële begunstigden van de steunmaatregel te doen toekomen.
De Commissie wijst Nederland op de schorsende werking van artikel 88, lid 3, van het EG-Verdrag. Zij verwijst naar artikel 14 van Verordening (EG) nr. 659/1999, volgens hetwelk elke onrechtmatige steun van de begunstigden kan worden teruggevorderd.
Voorts deelt de Commissie Nederland mee, dat zij de belanghebbenden door de bekendmaking van dit schrijven en van een samenvatting ervan in het Publicatieblad van de Europese Unie in kennis zal stellen. Tevens zal zij de belanghebbenden in de lidstaten van de EVA die partij zijn bij de EER-Overeenkomst door de bekendmaking van een mededeling in het EER-supplement van het Publicatieblad in kennis stellen, alsmede de Toezichthoudende Autoriteit van de EVA door haar een afschrift van dit schrijven toe te zenden. Alle bovengenoemde belanghebbenden zal worden verzocht hun opmerkingen te maken binnen een maand vanaf de datum van deze bekendmaking.%quot%
[1] På begäran av Essent förpliktade distriktsdomstolen i Groningen kommunen att anmäla planerna till kommissionen enligt artikel 88.3 i EG-fördraget.
[2] Det finns de som hävdar att den nya generationens nät inte är jämförbara med dagens koppar- eller kabelnät och att statliga åtgärder till förmån för den nya generationens allmänna, offentliga lokala accessnät kan påverka den ekonomiska utvecklingen positivt på grund av nätens positiva effekter på innovation och tillväxt. De företag som i dag driver elektroniska kommunikationsnät har ännu inte börjat investera i dessa infrastrukturer på grund av de höga kapitalkostnaderna och på grund av att det skulle göra deras befintliga nät föråldrade (motstridiga intressen).
[3] Zie beschikking van de Commissie van 9 september 2004 in zaak N 213/03: steunmaatregel N 213/2003 — ATLAS-project in het Verenigd Koninkrijk; regeling breedbandinfrastructuur voor bedrijventerreinen (Corrigendum).
[4] Zie 3.
[5] Arrest van het Hof van Justitie van 24 juli 2003, in zaak C-280/00, Altmark Trans, Jurispr. 2003, blz. I-7747 .
[6] Zie de beschikkingen van de Commissie in de zaken N 213/03, %quot%ATLAS-project%quot%, en bijv. N 126/04 %quot%Breedbanddiensten voor KMO's in Lincolnshire%quot% en N 307/04, %quot%Breedbanddiensten in Schotland — afgelegen en plattelandsgebieden%quot%.
[7] Zie bijvoorbeeld: Lehr, Osorio, Gillet en Sirbu: %quot%Measuring Broadband's Economic Impact%quot%, 2005.
[8] OESO %quot%Broadband Driving Growth: Policy Responses%quot%, oktober 2003; Orazem, Peter, University of Kansas Business School, %quot%The Impact of High-Speed Internet Access on Local Economic Growth%quot%, augustus 2005.
--------------------------------------------------
Meddelande av den 21 januari 2005 från Maltas regering i enlighet med Europaparlamentets och rådets direktiv 94/22/EG av den 30 maj 1994 (om villkoren för beviljande och utnyttjande av tillstånd för prospektering efter samt undersökning och utvinning av kolväten) [1]
(2005/C 62/06)
(Text av betydelse för EES)
I enlighet med artikel 3.3 i ovannämnda direktiv underrättar Republiken Maltas ministerium för resurser och infrastruktur (Ministry for Resources and Infrastructure of the Republic of Malta – l-Ministeru tar-Riÿorsi u l-Infrastruttura tar-Repubblika ta' Malta) härmed att följande offshoreområden, eller block inom dem, är aktuella för beviljande av tillstånd, antingen för enbart prospektering eller för både prospektering och produktion:
(i) Område 1
(ii) Område 3 (utom för nedan angivna block)
(iii) Område 4 (utom för nedan angivna block)
(iv) Område 6
För följande områden eller block finns tillstånd som beviljats före den 1 maj 2004. Nya tillstånd får således inte beviljas innan annat meddelas.
(i) Område 2
(ii) Block 4 och 5 i område 3
(iii) Block 3 i område 4
(iv) Område 5
(v) Område 7
Sökande skall inkomma med uppgifter som skall fyllas i på den blankett som publiceras i Republiken Maltas bestämmelser om oljeproduktion (rättsliga meddelanden nr 320 av den 1 december 2001) (Petroleum [Production] Regulations [Legal Notice 320, 1st December 2001] – Regolamenti dwar iÿ-ÿejt [Produzzjoni], 2001 [Avviÿ Legali 320 ta' l-2001, 1 ta' Diÿembru 2001]).
De områden eller block som är aktuella för beviljande av tillstånd, liksom de områden eller block för vilka tillstånd redan beviljats, begränsas av geografiska koordinater. Ni kan erhålla uppgift om dessa, liksom annan information, genom att kontakta byrån för oljeprospektering vid ministeriet för resurser och infrastruktur (Oil Exploration Department at the Ministry for Resources and Infrastructure – mid-Dipartiment ta' l-Esplorazzjoni gÿaÿ-ÿejt fil-Ministeru tar-Riÿorsi u l-Infrastruttura), adress Blokk B, il-Furjana CMR 02, Malta (tfn (356) 21 23 79 21).
[1] EGT L 164, 30.6.1994, s. 3.
--------------------------------------------------
Administrativa kommissionen för social trygghet för migrerande arbetare
(2005/C 232/03)
Vid beräkningen av de genomsnittliga årskostnaderna tas inte hänsyn till den minskning med 20 % som föreskrivs i artiklarna 94.2 och 95.2 i rådets förordning (EEG) nr 574/72.
De genomsnittliga nettokostnaderna per månad har däremot minskats med 20 %.
GENOMSNITTLIGA KOSTNADER FÖR VÅRDFÖRMÅNER – 2001 [1]
I. Tillämpning av artikel 94 i rådets förordning (EEG) nr 574/72
De belopp som skall återbetalas för vårdförmåner som utgetts under 2001 till familjemedlemmar i enlighet med artikel 19.2 i rådets förordning (EEG) nr 1408/71 kommer att fastställas på grundval av följande genomsnittliga kostnader:
| Årskostnad | Netto per månad |
Irland | EUR 2649,76 | EUR 176,65 |
II. Tillämpning av artikel 95 i rådets förordning (EEG) nr 574/72
De belopp som skall återbetalas för vårdförmåner som utgetts under 2001 i enlighet med artiklarna 28 och 28a i rådets förordning (EEG) nr 1408/71 kommer att fastställas på grundval av följande genomsnittliga kostnader:
| Årskostnad | Netto per månad |
Irland | | |
—per familj | EUR 6149,54 | EUR 409,97 |
—per person | EUR 4978,20 | EUR 331,88 |
GENOMSNITTLIGA KOSTNADER FÖR VÅRDFÖRMÅNER – 2002 [2]
I. Tillämpning av artikel 94 i rådets förordning (EEG) nr 574/72
De belopp som skall återbetalas för vårdförmåner som utgetts under 2002 till familjemedlemmar i enlighet med artikel 19.2 i rådets förordning (EEG) nr 1408/71 kommer att fastställas på grundval av följande genomsnittliga kostnader:
| Årskostnad | Netto per månad |
Förenade kungariket | GBP 1554,78 | GBP 103,65 |
Italien | EUR 1898,61 | EUR 126,57 |
Tyskland | | |
—per person | EUR 1023,93 | EUR 68,26 |
II. Tillämpning av artikel 95 i rådets förordning (EEG) nr 574/72
De belopp som skall återbetalas för vårdförmåner som utgetts under 2002 i enlighet med artiklarna 28 och 28a i rådets förordning (EEG) nr 1408/71 kommer att fastställas på grundval av följande genomsnittliga kostnader (endast per person från 2002):
| Årskostnad | Netto per månad |
Förenade kungariket | GBP 2379,72 | GBP 158,65 |
Italien | EUR 2240,74 | EUR 149,38 |
Tyskland | EUR 4084,27 | EUR 272,28 |
GENOMSNITTLIGA KOSTNADER FÖR VÅRDFÖRMÅNER – 2003 [3]
I. Tillämpning av artikel 94 i rådets förordning (EEG) nr 574/72
De belopp som skall återbetalas för vårdförmåner som utgetts under 2003 till familjemedlemmar i enlighet med artikel 19.2 i rådets förordning (EEG) nr 1408/71 kommer att fastställas på grundval av följande genomsnittliga kostnader:
| Årskostnad | Netto per månad |
Nederländerna
—försäkrade och pensionstagare under 65 år | EUR 1651,65 | EUR 110,11 |
Tyskland
—per person | EUR 1043,67 | EUR 69,58 |
Frankrike
—per familj | EUR 1792,50 | EUR 119,50 |
II. Tillämpning av artikel 95 i rådets förordning (EEG) nr 574/72
De belopp som skall återbetalas för vårdförmåner som utgetts under 2003 i enlighet med artiklarna 28 och 28a i rådets förordning (EEG) nr 1408/71 kommer att fastställas på grundval av följande genomsnittliga kostnader (endast per person från 2002):
| Årskostnad | Netto per månad |
Nederländerna | | |
—pensionstagare 65 år och över och deras familjemedlemmar | EUR 8600,13 | EUR 573,34 |
Tyskland | EUR 4262,70 | EUR 284,18 |
Frankrike | EUR 4349,29 | EUR 289,95 |
GENOMSNITTLIGA KOSTNADER FÖR VÅRDFÖRMÅNER – 2004
I. Tillämpning av artikel 94 i rådets förordning (EEG) nr 574/72
De belopp som skall återbetalas för vårdförmåner som utgetts under 2004 till familjemedlemmar i enlighet med artikel 19.2 i rådets förordning (EEG) nr 1408/71 kommer att fastställas på grundval av följande genomsnittliga kostnader:
| Årskostnad | Netto per månad |
Lettland | LVL 132,42 | LVL 8,83 |
II. Tillämpning av artikel 95 i rådets förordning (EEG) nr 574/72
De belopp som skall återbetalas för vårdförmåner som utgetts under 2004 i enlighet med artiklarna 28 och 28a i rådets förordning (EEG) nr 1408/71 kommer att fastställas på grundval av följande genomsnittliga kostnader (endast per person från 2002):
| Årskostnad | Netto per månad |
Lettland | LVL 141,60 | LVL 9,44 |
[1] Genomsnittliga kostnader 2001:
- Spanien och Österrike (EGT C 3, 8.1.2003).
- Sverige (EUT C 163, 12.7.2003).
- Belgien, Tyskland, Grekland, Frankrike, Luxemburg, Nederländerna och Portugal (EUT C 37, 11.2.2004).
- Norge (EUT C 27, 3.2.2005).
[2] Genomsnittliga kostnader 2002:
- Luxemburg och Österrike (EUT C 37, 11.2.2004).
- Belgien, Frankrike, Portugal, Sverige (EUT C 27, 3.2.2005, s. 4).
[3] Genomsnittliga kostnader 2003:
- Österrike, Spanien och Schweiz (EUT C 27, 3.2.2005, s. 4)
--------------------------------------------------
Meddelande från de franska myndigheterna om tillämpning av Europaparlamentets och rådets direktiv 94/22/EG av den 30 maj 1994 om villkoren för beviljande och utnyttjande av tillstånd för prospektering efter samt undersökning och utvinning av kolväten [1]
(Yttrande över en ansökan om ett exklusivt tillstånd för prospektering efter flytande kolväten eller kolväten i gasform (Claracq-tillstånd)
(2005/C 331/03)
(Text av betydelse för EES)
Den 15 februari 2005 lämnade företaget Celtique Energie Limited (huvudkontorets adress: 36 Sekforde Street, London (England)) in en ansökan om ett treårigt exklusivt tillstånd för prospektering efter flytande kolväten och kolväten i gasform ("Claracq-tillstånd") i ett ungefär 726 kvadratkilometer stort område, i de franska departementen Pyrénées Atlantiques och Landes.
Ansökan avser ett område som avgränsas av linjer mellan de punkter på längd- och breddgrader, vars geografiska koordinater anges nedan och som successivt sammanbinds. Parismeridianen räknas som nollmeridian. (Greenwich-graderna anges i informationssyfte):
Punkt | Y( Latitud) | X( Longitud) |
A | 48,50 gr N | 3,30 gr V |
B | 48,50 gr N | 3,05 gr V |
C | 48,47 gr N | 3,05 gr V |
D | 48,47 gr N | 2,93 gr V |
E | 48,50 gr N | 2,93 gr V |
F | 48,50 gr N | 2,90 gr V |
G | 48,35 gr N | 2,90 gr V |
H | 48,35 gr N | 2,87 gr V |
I | 48,34 gr N | 2,87 gr V |
J | 48,34 gr N | 2,85 gr V |
K | 48,33 gr N | 2,85 gr V |
L | 48,33 gr N | 2,80 gr V |
M | 48,20 gr N | 2,80 gr V |
N | 48,20 gr N | 3,10 gr V |
O | 48,30 gr N | 3,10 gr V |
P | 48,30 gr N | 3,13 gr V |
Q | 48,33 gr N | 3,13 gr V |
R | 48,33 gr N | 3,17 gr V |
S | 48,35 gr N | 3,17 gr V |
T | 48,35 gr N | 3,25 gr V |
U | 48,40 gr N | 3,25 gr V |
V | 48,40 gr N | 3,30 gr V |
Inlämnande av ansökningar
De företag som lämnat in den ursprungliga ansökan samt de som lämnar in en konkurrerande ansökan skall visa att villkoren för beviljande av licensen är uppfyllda. Dessa villkor anges i artiklarna 3–5 i det ändrade dekretet 95-427 av den 19 april 1995 om gruvdriftslicenser.
Intresserade företag kan lämna in en konkurrerande ansökan inom 90 dagar räknat från offentliggörandet av detta tillkännagivande i enlighet med det förfarande som anges i tillkännagivandet om ansökningsförfarande för gruvdriftslicenser för kolväten i Frankrike (offentliggjort i Europeiska gemenskapernas officiella tidning C 374 av den 30 december 1994, sidan 11) och som fastställs genom dekret 95-427 av den 19 april 1995 om brytningsrättigheter ("Journal officiel de la République française" av den 22 april 1995).
Konkurrerande ansökningar skall skickas till den minister som ansvarar för gruvor, på nedan angivna adress. Beslutet om beviljande av licens till det ansökande företaget eller ett konkurrerande företag kommer att fattas inom två år räknat från det att de franska myndigheterna tog emot den första ansökningen, dvs. senast den 15 februari 2007.
Villkor och krav beträffande utövande och avslutande av verksamheten
De sökande hänvisas till artikel 79 och artikel 79.1 i gruvlagstiftningen och till det ändrade dekretet nr 95-696 av den 9 maj 1995 (décret relatif à l'ouverture des travaux miniers et à la police des mines) som offentliggjorts i "Journal officiel de la République française" av den 11 maj 1995.
Ytterligare information kan erhållas från följande adress: Ministère de l'économie, des finances et de l'industrie (direction générale de l'énergie et des matières premières, direction des ressources énergétiques et minérales, bureau de la législation minière), 61, Boulevard Vincent Auriol, Teledoc 133, F-75703 Paris, Cedex 13, (tfn (33-1) 44 97 23 02, fax (33-1) 44 97 05 70).
De lagar och andra bestämmelser som anges ovan finns tillgängliga på följande webbplats: http:// www.legifrance.gouv.fr
[1] EGT L 164 av den 30 juni 1994, s. 3.
--------------------------------------------------
Gemensam ståndpunkt (EG) nr 9/2006
antagen av rådet den 9 mars 2006
inför antagandet av Europaparlamentets och rådets förordning (EG) nr 000/2006 av den … om ändring av rådets förordning (EEG) nr 3922/91 om harmonisering av tekniska krav och administrativa förfaranden inom området civil luftfart
(2006/C 179 E/01)
(Text av betydelse för EES)
EUROPAPARLAMENTET OCH EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 80.2,
med beaktande av kommissionens förslag,
med beaktande av Europeiska ekonomiska och sociala kommitténs yttrande [1],
efter att ha hört Regionkommittén,
i enlighet med förfarandet i artikel 251 i fördraget [2], och
av följande skäl:
(1) I förordning (EEG) nr 3922/91 [3] fastställdes gemensamma säkerhetsnormer förtecknade i bilaga II till den förordningen, särskilt med avseende på konstruktion, tillverkning, drift och underhåll av luftfartyg samt personer och organisationer som sysslar med dessa uppgifter. Dessa harmoniserade säkerhetsnormer gällde samtliga luftfartyg som drivs av gemenskapens operatörer, vare sig luftfartygen är registrerade i en medlemsstat eller i ett tredjeland.
(2) Vad avser områden som inte fanns förtecknade i bilaga II till den förordningen skall det, enligt artikel 4.1 i den förordningen, antas gemensamma tekniska krav och administrativa förfaranden på grundval av artikel 80.2 i fördraget.
(3) I artikel 9 i förordning (EEG) nr 2407/92 av den 23 juli 1992 om utfärdande av tillstånd för lufttrafikföretag [4] föreskrivs att det alltid skall vara ett villkor för utfärdandet av en operativ licens och för dess giltighet att det berörda företaget har ett gällande drifttillstånd att utöva trafikrättigheter som täcker den verksamhet som den operativa licensen omfattar och som uppfyllde krav som skall fastställas i en framtida förordning. Det är nu lämpligt att fastställa sådana krav.
(4) De gemensamma luftfartsmyndigheterna, JAA (Joint Aviation Authorities), har antagit ett antal harmoniserade bestämmelser för kommersiell luftfart med flygplan, Gemensamma luftfartsbestämmelser - kommersiella flygtransporter (flygplan) (JAR-OPS 1) i dess ändrade version. I dessa bestämmelser (ändring 8 av den 1 januari 2005) fastställs en lägsta säkerhetsnivå, och de utgör därför ett bra underlag för gemenskapslagstiftning om drift av flygplan. Ändringar av JAR-OPS 1 måste dock göras, så att den blir förenlig med gemenskapens lagstiftning och politik, med hänsyn till dess betydelse för den ekonomiska och sociala sektorn. Den nya texten kan inte införlivas med gemenskapsrätten enbart genom en enkel hänvisning till JAR-OPS 1 i förordning (EEG) nr 3922/91. Således bör en ny bilaga med de gemensamma bestämmelserna fogas till den förordningen.
(5) Villkoren för lufttransportföretag bör vara tillräckligt flexibla så att de kan hantera oförutsedda brådskande driftsrelaterade omständigheter, driftsrelaterade behov av begränsad varaktighet eller visa att de kan uppnå motsvarande säkerhetsnivå genom andra åtgärder än tillämpning av de gemensamma bestämmelserna i bilagan (nedan kallad "bilaga III"). Medlemsstaterna bör därför ha rätt att bevilja undantag från eller införa varianter av de gemensamma tekniska kraven och administrativa förfarandena. Eftersom sådana undantag och varianter i vissa fall kan urholka de gemensamma säkerhetsnormerna eller förorsaka en snedvridning av marknaden, bör deras tillämpningsområde snävt begränsas och gemenskapen bör på lämpligt sätt kontrollera beviljandet. Kommissionen bör ges befogenhet att besluta om skyddsåtgärder i detta avseende.
(6) Det finns klart angivna fall då medlemsstaterna bör få anta eller behålla nationella bestämmelser om flyg- och tjänstgöringstidsbegränsningar och kraven på vila, under förutsättning att de överensstämmer med allmänt etablerade förfaranden och till dess att gemenskapsbestämmelser har fastställts på grundval av vetenskapliga rön och bästa praxis.
(7) Bestämmelserna om kommittéförfarandet i förordning (EEG) nr 3922/91 bör anpassas, så att hänsyn tas till rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter [5].
(8) Bestämmelserna i förordning (EEG) nr 3922/91 om tillämpningsområdet bör anpassas, så att hänsyn tas till Europaparlamentets och rådets förordning (EG) nr 1592/2002 av den 15 juli 2002 om fastställande av gemensamma bestämmelser på det civila luftfartsområdet och inrättande av en europeisk byrå för luftfartssäkerhet [6] samt till tillämpningsföreskrifterna till denna i kommissionens förordning (EG) nr 1702/2003 av den 24 september 2003 om fastställande av tillämpningsföreskrifter för luftvärdighets- och miljöcertifiering av luftfartyg och tillhörande produkter, delar och utrustningar samt för certifiering av konstruktions- och tillverkningsorganisationer [7] och i kommissionens förordning (EG) nr 2042/2003 av den 20 november 2003 om fortsatt luftvärdighet för luftfartyg och luftfartygsprodukter, delar och utrustning och om godkännande av organisationer och personal som arbetar med dessa arbetsuppgifter [8].
(9) I denna förordning, särskilt i bestämmelserna om flyg- och tjänstgöringstidsbegränsningar och kraven på vila i kapitel Q i bilaga III, beaktas de begränsningar och miniminormer som redan har fastställts i direktiv 2000/79/EG [9]. De begränsningar som fastställs i det direktivet bör alltid iakttas för flygpersonal inom civil luftfart. Inte i något avseende bör bestämmelserna i kapitel Q i bilaga III och andra bestämmelser som godkänns enligt denna förordning vara vidare och därigenom ge den personalen mindre skydd.
(10) Medlemsstaterna bör kunna fortsätta att tillämpa nationella bestämmelser om flyg- och tjänstgöringstidsbegränsningar och krav på vila för besättningsmedlemmar, under förutsättning att de gränser som fastställs i sådana nationella bestämmelser ligger mellan de undre och övre gränser som anges i kapitel Q i bilaga III.
(11) Medlemsstaterna bör kunna fortsätta att tillämpa nationella bestämmelser om flyg- och tjänstgöringstidsbegränsningar och krav på vila för besättningsmedlemmar på områden som för närvarande inte omfattas av kapitel Q i bilaga III, t.ex. maximala dagliga flygtjänstgöringsperioder för enpilotverksamhet och brådskande medicinska transporter samt bestämmelser om minskning av flygtjänstgöringsperioder eller ökning av viloperioder vid flygningar över flera tidszoner.
(12) En vetenskaplig och medicinsk utvärdering av bestämmelserna om flyg- och tjänstgöringstidsbegränsningar och kraven på vila samt, om så behövs, av bestämmelserna om kabinbesättningar bör genomföras inom tre år efter det att denna förordning har trätt i kraft.
(13) Denna förordning bör inte påverka tillämpningen av de bestämmelser om inspektioner som fastställs i 1944 års Chicagokonvention angående internationell civil luftfart och i Europaparlamentets och rådets direktiv 2004/36/EG av den 21 april 2004 om säkerheten i fråga om luftfartyg från tredje land som använder flygplatser i gemenskapen [10].
(14) En överenskommelse om utökat samarbete i fråga om användningen av flygplatsen i Gibraltar träffades i London den 2 december 1987 mellan Konungariket Spanien och Förenade kungariket genom en gemensam förklaring från de båda ländernas utrikesministrar. Denna överenskommelse har ännu inte trätt i kraft.
(15) Förordning (EEG) nr 3922/91 bör därför ändras i enlighet med detta.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Förordning (EEG) nr 3922/91 skall ändras på följande sätt:
1. Det sista skälet skall ersättas med följande skäl:
"De åtgärder som är nödvändiga för att genomföra denna förordning bör antas i enlighet med rådets beslut 1999/468/EG av den 28 juni 1999 om de förfaranden som skall tillämpas vid utövandet av kommissionens genomförandebefogenheter [11]."
2. Artikel 1 skall ändras på följande sätt:
a) Punkt 1 skall ersättas med följande:
"1. Denna förordning skall tillämpas på harmoniseringen av sådana tekniska krav och administrativa förfaranden inom den civila luftfarten som avser drift och underhåll av luftfartyg, och personal och organisationer som sysslar med sådan verksamhet."
b) Följande punkter skall läggas till:
"3. Tillämpningen av denna förordning på flygplatsen i Gibraltar skall inte anses påverka Konungariket Spaniens respektive Förenade kungarikets rättsliga ståndpunkter i tvisten om överhögheten över det territorium där flygplatsen är belägen.
4. Tillämpningen av denna förordning på flygplatsen i Gibraltar skall uppskjutas tills överenskommelsen enligt den gemensamma förklaringen från Konungariket Spaniens och Förenade kungarikets utrikesministrar den 2 december 1987 har trätt i kraft. Konungariket Spaniens och Förenade kungarikets regeringar skall informera rådet om när detta sker."
3. Följande definition skall läggas till i artikel 2:
"i) myndighet: i bilaga III den behöriga myndighet som har beviljat lufttrafikföretagets drifttillstånd (AOC)."
4. Artikel 3 skall ersättas med följande:
"Artikel 3
1. Utan att det påverkar tillämpningen av artikel 11 skall de gemensamma tekniska krav och administrativa förfaranden som är tillämpliga inom gemenskapen vad gäller kommersiella transporter med flygplan vara de som anges i bilaga III.
2. Hänvisningar till kapitel M i bilaga III eller någon av bestämmelserna i det skall avse del-M i kommissionens förordning (EG) nr 2042/2003 av den 20 november 2003 om fortsatt luftvärdighet för luftfartyg och luftfartygsprodukter, delar och utrustning och om godkännande av organisationer och personal som arbetar med dessa arbetsuppgifter [12] eller relevanta bestämmelser i denna."
5. Artikel 4.1 skall ersättas med följande:
"1. Vad avser områden som inte omfattas av bilaga III skall gemensamma tekniska krav och administrativa förfaranden antas på grundval av artikel 80.2 i fördraget. Kommissionen skall i förekommande fall och så snart som möjligt lägga fram lämpliga förslag inom dessa områden."
6. Artikel 6 skall ersättas med följande:
"Artikel 6
Ett luftfartyg som är i drift enligt ett godkännande som beviljats av en medlemsstat i enlighet med de gemensamma tekniska kraven och administrativa förfarandena får tas i drift på samma villkor i övriga medlemsstater, utan ytterligare tekniska krav eller utvärderingar i dessa medlemsstater."
7. Artikel 7 skall ersättas med följande:
"Artikel 7
Medlemsstaterna skall erkänna en certifiering av organ eller personer under dess jurisdiktion och myndighet, vilka sysslar med underhåll av produkter och drift av luftfartyg, när denna utfärdats enligt denna förordning av en annan medlemsstat eller av ett organ som handlar på dess uppdrag."
8. Artikel 8 skall ersättas med följande:
"Artikel 8
1. Bestämmelserna i artiklarna 3–7 får inte hindra en medlemsstat från att omedelbart reagera om det uppstår ett säkerhetsproblem som rör en produkt, person eller organisation som omfattas av denna förordning.
Om säkerhetsproblemet är ett resultat av en otillräcklig säkerhetsnivå som beror på de gemensamma tekniska kraven och administrativa förfarandena, eller på brister i dessa tekniska krav och förfaranden, skall medlemsstaten omedelbart meddela kommissionen och de övriga medlemsstaterna vilka åtgärder som vidtagits och skälen till detta.
Kommissionen skall i enlighet med förfarandet i artikel 12.2 besluta om huruvida en otillräcklig säkerhetsnivå eller en brist i de gemensamma tekniska kraven och administrativa förfarandena gör fortsatt tillämpning av de åtgärder som vidtagits i enlighet med första stycket i denna punkt motiverad. Kommissionen skall i så fall vidta nödvändiga åtgärder för att ändra de berörda gemensamma tekniska kraven och administrativa förfarandena i enlighet med artikel 4 eller artikel 11. Om det visar sig att medlemsstatens åtgärder inte är motiverade, skall den återkalla åtgärderna.
2. En medlemsstat får bevilja undantag från de tekniska krav och administrativa förfaranden som anges i denna förordning vid oförutsedda brådskande driftsrelaterade omständigheter eller driftsrelaterade behov av begränsad varaktighet.
Kommissionen och de övriga medlemsstaterna skall underrättas om de beviljade undantagen, om dessa upprepas eller om de har beviljats för en period som är längre än två månader.
När kommissionen och övriga medlemsstater underrättas om undantag som beviljats av en medlemsstat i enlighet med andra stycket skall kommissionen undersöka huruvida undantagen är förenliga med säkerhetsmålen i denna förordning eller andra bestämmelser i gemenskapsrätten.
Om kommissionen finner att de beviljade undantagen inte är förenliga med säkerhetsmålen i denna förordning eller andra bestämmelser i gemenskapsrätten, skall kommissionen besluta om skyddsåtgärder i enlighet med förfarandet i artikel 12a.
Den berörda medlemsstaten skall i så fall upphäva undantaget.
3. Där det är möjligt att med andra medel uppnå en säkerhetsnivå som motsvarar den nivå som uppnås genom tillämpning av de gemensamma tekniska kraven och administrativa förfarandena i bilaga III, får medlemsstaterna, utan diskriminering på grund av sökandens nationalitet och med beaktande av behovet av att inte snedvrida konkurrensen, bevilja ett godkännande med avvikelse från dessa bestämmelser.
Den berörda medlemsstaten skall i så fall till kommissionen anmäla sin avsikt att bevilja ett sådant godkännande, skälen till detta och villkoren för att säkerställa att en motsvarande säkerhetsnivå uppnås.
Inom tre månader efter det att en medlemsstat lämnat in en anmälan skall kommissionen inleda det förfarande som avses i artikel 12.2 i syfte att besluta huruvida det föreslagna godkännandet av åtgärden kan beviljas.
I så fall skall kommissionen meddela samtliga medlemsstater sitt beslut, och de skall därvid ha rätt att tillämpa åtgärden. Tillämpliga bestämmelser i bilaga III får också ändras för att återspegla en sådan åtgärd.
Bestämmelserna i artiklarna 6 och 7 skall tillämpas på åtgärden i fråga.
4. Utan hinder av bestämmelserna i punkterna 1-3 får en medlemsstat anta eller bibehålla bestämmelser i anslutning till OPS 1.1105 punkt 6, OPS 1.1110 punkterna 1.3 och 1.4.1, OPS 1.1115 och OPS 1.1125 punkt 2.1 i kapitel Q i bilaga III till dess att gemenskapsbestämmelser har fastställts på grundval av vetenskapliga rön och bästa praxis.
En medlemsstat skall underrätta kommissionen om de bestämmelser som den beslutar att bibehålla.
För nationella bestämmelser som avviker från de bestämmelser i OPS 1 som avses i första stycket och som medlemsstaterna avser att anta efter dagen för tillämpning av bilaga III skall kommissionen inom tre månader efter anmälan från en medlemsstat inleda det förfarande som avses i artikel 12.2 för att besluta om huruvida bestämmelserna är förenliga med säkerhetsmålen i denna förordning och andra regler i gemenskapsrätten och om bestämmelserna får göras tillämpliga.
I så fall skall kommissionen meddela samtliga medlemsstater sitt beslut att godkänna åtgärden och alla skall därvid ha rätt att tillämpa den åtgärden. Tillämpliga bestämmelser i bilaga III får också ändras för att återspegla en sådan åtgärd.
Bestämmelserna i artiklarna 6 och 7 skall tillämpas på åtgärden i fråga."
9. Följande artikel skall införas:
"Artikel 8a
1. Inom … [13] skall Europeiska byrån för luftfartssäkerhet slutföra en vetenskaplig och medicinsk utvärdering av bestämmelserna i kapitel Q och i förekommande fall kapitel O i bilaga III.
2. Utan att det påverkar tillämpningen av artikel 7 i Europaparlamentets och rådets förordning (EG) nr 1592/2002 av den 15 juli 2002 om fastställande av gemensamma bestämmelser på det civila luftfartsområdet och inrättande av en europeisk byrå för luftfartssäkerhet [14] skall Europeiska byrån för luftfartssäkerhet bistå kommissionen med att utarbeta förslag till ändringar av de tillämpliga tekniska bestämmelserna i kapitel Q i bilaga III."
10. Artikel 11.1 skall ersättas med följande:
"1. Enligt det förfarande som avses i artikel 12.2 skall kommissionen göra de ändringar som blivit nödvändiga på grund av vetenskapliga och tekniska framsteg i de gemensamma tekniska krav och administrativa förfaranden som anges i bilaga III."
11. Artikel 12 skall ersättas med följande:
"Artikel 12
1. Kommissionen skall biträdas av luftsäkerhetskommittén, nedan kallad kommittén.
2. När det hänvisas till denna punkt skall artiklarna 5 och 7 i rådets beslut 1999/468/EG [15] tillämpas, med beaktande av bestämmelserna i artikel 8 i det beslutet.
Den tid som fastställs i artikel 5.6 i beslut 1999/468/EG skall vara tre månader.
3. Kommittén skall själv anta sin arbetsordning."
12. Följande artikel skall införas:
"Artikel 12a
När det hänvisas till denna artikel skall förfarandet i fråga om skyddsåtgärder i artikel 6 i beslut 1999/468/EG tillämpas.
Innan kommissionen antar sitt beslut skall den höra kommittén.
Den tid som avses i artikel 6 b i beslut 1999/468/EG skall vara tre månader.
Om en medlemsstat hänskjuter ett beslut som fattats av kommissionen till rådet, får rådet med kvalificerad majoritet fatta ett annat beslut inom tre månader."
13. Texten i bilagan till denna förordning skall läggas till som bilaga III.
Artikel 2
Denna förordning träder i kraft den tjugonde dagen efter det att den har offentliggjorts i Europeiska unionens officiella tidning.
Utan att det påverkar tillämpningen av bestämmelserna i artikel 11 i förordning (EEG) nr 3922/91, skall bilaga III tillämpas från och med … [16].
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Utfärdad i … den …
På Europaparlamentets vägnar
…
Ordförande
På rådets vägnar
…
Ordförande
[1] EGT C 14, 16.1.2001, s. 33.
[2] Europaparlamentets yttrande av den 3 september 2002 (EUT C 272 E, 13.11.2003, s. 103), rådets gemensamma ståndpunkt av den 9 mars 2006 och Europaparlamentets ståndpunkt av den ... (ännu ej offentliggjord i EUT).
[3] EGT L 373, 31.12.1991, s. 4. Förordningen senast ändrad genom Europaparlamentets och rådets förordning (EG) nr 1592/2002 (EGT L 240, 7.9.2002, s. 1).
[4] EGT L 240, 24.8.1992, s. 1.
[5] EGT L 184, 17.7.1999, s. 23.
[6] EGT L 240, 7.9.2002, s. 1. Förordningen senast ändrad genom kommissionens förordning (EG) nr 1701/2003 (EUT L 243, 27.9.2003, s. 5).
[7] EUT L 243, 27.9.2003, s. 6.
[8] EUT L 315, 28.11.2003, s. 1.
[9] Rådets direktiv 2000/79/EG av den 27 november 2000 om genomförande av det europeiska avtal om arbetstidens förläggning för flygpersonal inom civilflyget som har ingåtts mellan Association of European Airlines (AEA), Europeiska transportarbetarfederationen (ETF), European Cockpit Association (ECA), European Regions Airline Association (ERA) och International Air Carrier Association (IACA) (EGT L 302, 1.12.2000, s. 57).
[10] EUT L 143, 30.4.2004, s. 76.
[11] EGT L 184, 17.7.1999, s. 23.
[12] EUT L 315, 28.11.2003, s. 1.
[13] Tre år efter det att denna förordning har trätt i kraft.
[14] EGT L 240, 7.9.2002, s. 1. Förordningen senast ändrad genom kommissionens förordning (EG) nr 1701/2003 (EUT L 243, 27.9.2003, s. 5).
[15] EGT L 184, 17.7.1999, s. 23.
[16] 18 månader efter det att denna förordning har trätt i kraft.
--------------------------------------------------
[pic] | EUROPEISKA GEMENSKAPERNAS KOMMISSION |
Bryssel den 8.2.2006
KOM(2006) 48 slutlig
MEDDELANDE FRÅN KOMMISSIONEN TILL RÅDET, EUROPAPARLAMENTET, EUROPEISKA EKONOMISKA OCH SOCIALA KOMMITTÉN SAMT REGIONKOMMITTÉN
Rapport om hur övergångsordningarna enligt 2003 års anslutningsakt har fungerat under perioden 1 maj 2004–30 april 2006
INNEHÅLLSFÖRTECKNING
1. Rapportens syfte 3
2. Övergångsordningarna 3
3. Samråd med medlemsstaterna och arbetsmarknadens parter 5
4. Statistik över arbetstagnas rörlighet före och efter utvidgningen 6
4.1 Arbetstagarnas rörlighet inom den utvidgade Europeiska unionen 7
4.2 Arbetsmarknadsstatistik för ländernas egna medborgare och EU-medborgare: förvärvsfrekvens 11
4.3. EU 10-arbetskraftens fördelning i EU 15-medlemsstaterna efter bransch och kvalifikationer: komplement eller ersättning? 13
5. Slutsatser och rekommendationer 14
[pic] | EUROPEISKA GEMENSKAPERNAS KOMMISSION |
Bryssel den 27.4.2006
KOM(2006) 192 slutlig
Förslag till
RÅDETS FÖRORDNING
om förlängning av de restriktiva åtgärderna mot Burma/Myanmar och om upphävande av förordning (EG) nr 798/2004
(framlagt av kommissionen)
MOTIVERING
1. Den 28 oktober 1996 införde rådet genom gemensam ståndpunkt 96/635/GUSP vissa restriktiva åtgärder mot Burma/Myanmar, mot bakgrund av det politiska läget i det landet. Dessa åtgärder förlängdes och ändrades därefter genom gemensam ståndpunkt 2000/346/GUSP samt genom gemensam ståndpunkt 2003/297/GUSP, som upphörde att gälla den 29 april 2004. Åtgärderna förlängdes genom gemensam ståndpunkt 2004/423/GUSP, skärptes genom gemensam ståndpunkt 2004/730/GUSP, ändrades genom gemensam ståndpunkt 2005/149/GUSP samt förlängdes och ändrades genom gemensam ståndpunkt 2005/340/GUSP.
2. Vissa av de restriktiva åtgärder som införts mot Burma/Myanmar genomfördes på gemenskapsnivå genom rådets förordning (EG) nr 798/2004.
3. På grund av att rådet hade fortsatt att hysa oro över det politiska läget i Burma/Myanmar och situationen i det landet i fråga om de mänskliga rättigheterna beslutade det genom gemensam ståndpunkt 2006/…/GUSP att bibehålla restriktiva åtgärder mot Burma/Myanmar och att konsolidera och aktualisera texten till den berörda förordningen. 4. Därför bör förordning (EG) nr 798/2004 upphävas och en ny förordning offentliggöras.
Förslag till
RÅDETS FÖRORDNING
om förlängning av de restriktiva åtgärderna mot Burma/Myanmar och om upphävande av förordning (EG) nr 798/2004
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artiklarna 60 och 301,
med beaktande av rådets gemensamma ståndpunkt 2006/…/GUSP om förlängning av restriktiva åtgärder mot Burma/Myanmar[1],
med beaktande av kommissionens förslag[2], och
av följande skäl:
(1) Den 28 oktober 1996 införde rådet, på grund av sin oro över bristen på framsteg i fråga om demokratisering i Burma/Myanmar och de fortsatta kränkningarna av de mänskliga rättigheterna i det landet, genom gemensam ståndpunkt 1996/653/GUSP[3] vissa restriktiva åtgärder mot Burma/Myanmar. Åtgärderna förlängdes och ändrades genom gemensam ståndpunkt 2000/346/GUSP[4] och gemensam ståndpunkt 2003/297/GUSP[5], förlängdes genom gemensam ståndpunkt 2004/423/GUSP[6], skärptes genom gemensam ståndpunkt 2004/730/GUSP[7], ändrades genom gemensam ståndpunkt 2005/149/GUSP[8] samt förlängdes och ändrades genom gemensam ståndpunkt 2005/340/GUSP[9]. Vissa av de restriktiva åtgärder som införts mot Burma/Myanmar genomfördes på gemenskapsnivå genom rådets förordning (EG) nr 798/2004[10].
(2) På grund av det aktuella politiska läget i Burma/Myanmar, vilket exemplifieras av
- de militära myndigheternas underlåtenhet att inleda konkreta diskussioner med den demokratiska rörelsen om en process för att få till stånd nationell försoning, respekt för mänskliga rättigheter och demokrati,
- underlåtenheten att tillåta ett äkta och öppet nationalkonvent,
- underlåtenheten att frige Daw Aung San Suu Kyi och andra medlemmar av National League for Democracy (NLD) samt andra politiska fångar,
- de fortsatta trakasserierna av NLD och andra organiserade politiska rörelser,
- de fortsatta allvarliga kränkningarna av de mänskliga rättigheterna, bland annat underlåtenheten att vidta åtgärder för att göra slut på tvångsarbetet i enlighet med rekommendationerna i rapporten från Internationella arbetsorganisationens högnivågrupp 2001 och senare rekommendationer och förslag från ILO, och
- utvecklingen under den senaste tiden, t.ex. utökade restriktioner för internationella och icke-statliga organisationers verksamhet,
föreskrivs det i gemensam ståndpunkt 2006/…/GUSP att de restriktiva åtgärderna mot militärregimen i Burma/Myanmar, mot dem som drar den största fördelen av dess vanstyre samt mot dem som aktivt obstruerar arbetet med nationell försoning, respekt för mänskliga rättigheter och demokrati skall bibehållas.
(3) De restriktiva åtgärder som föreskrivs i gemensam ståndpunkt 2006/…/GUSP omfattar bland annat ett förbud mot tekniskt stöd, finansiering och finansiellt stöd som har samband med militär verksamhet, ett förbud mot export av utrustning som kan användas för inhemskt förtryck, frysning av penningmedel och ekonomiska resurser tillhörande medlemmar av Burma/Myanmars regering och fysiska eller juridiska personer, enheter eller organ som har anknytning till dessa samt ett förbud mot att göra finansiella lån eller krediter tillgängliga för burmesiska statsägda företag och att förvärva eller utöka en andel i sådana företag.
(4) Dessa åtgärder ligger inom fördragets tillämpningsområde och därför behövs det gemenskapslagstiftning för att genomföra dem för gemenskapens vidkommande, särskilt för att alla medlemsstaters ekonomiska aktörer skall kunna tillämpa dem på ett enhetligt sätt.
(5) Av tydlighetsskäl bör det antas en ny text, som innehåller alla relevanta bestämmelser i deras ändrade lydelse och träder i stället för förordning (EG) nr 798/2004, som bör upphävas.
(6) För att de åtgärder som föreskrivs i denna förordning skall vara verkningsfulla bör förordningen träda i kraft samma dag som den offentliggörs.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
I denna förordning gäller följande definitioner:
(1) tekniskt stöd: allt tekniskt stöd som har samband med reparation, utveckling, tillverkning, montering, testning, underhåll eller någon annan teknisk tjänst och som kan anta sådana former som instruktioner, råd, utbildning, överföring av praktiska kunskaper och färdigheter eller konsulttjänster; tekniskt stöd innefattar muntliga former av stöd.
(2) penningmedel: finansiella tillgångar och ekonomiska förmåner av alla slag, inbegripet men inte begränsat till
a) kontanter, checkar, penningfordringar, växlar, postanvisningar och andra betalningsinstrument,
b) inlåning hos finansinstitut eller andra enheter, kontotillgodohavanden, skuldebrev och skuldförbindelser,
c) börsnoterade och onoterade värdepapper och skuldinstrument, inbegripet aktier och andelar, certifikat för värdepapper, obligationer, växlar, optioner, förlagsbevis och derivatkontrakt, d) räntor, utdelningar eller annan inkomst från tillgångar eller annat värde som härrör från eller skapas genom tillgångar,
e) krediter, kvittningsrätter, garantiförbindelser, fullgörandegarantier eller andra finansiella åtaganden,
f) remburser, fraktsedlar och pantförskrivningar,
g) sådana dokument som utgör bevis på andelar i penningmedel eller andra finansiella resurser.
(3) frysning av penningmedel: förhindrande av varje flyttning, överföring, förändring, användning, tillgång till eller hantering av penningmedel på ett sätt som skulle leda till en förändring av volym, belopp, belägenhet, ägandeförhållanden, innehav, art, bestämmelse eller någon annan förändring som skulle göra det möjligt att utnyttja penningmedlen, inbegripet portföljförvaltning.
(4) ekonomiska resurser: egendom av alla slag, materiell eller immateriell, lös eller fast, som inte utgör penningmedel men som kan användas för att erhålla penningmedel, varor eller tjänster.
(5) frysning av ekonomiska resurser: förhindrande av att dessa resurser på något sätt används för att erhålla penningmedel, varor eller tjänster, inbegripet men inte enbart genom försäljning, uthyrning eller inteckning.
(6) gemenskapens territorium: de till medlemsstaterna hörande territorier på vilka fördraget är tillämpligt på de villkor som fastställs i detta.
Artikel 2
Det skall vara förbjudet
a) att tillhandahålla tekniskt stöd som har samband med militär verksamhet och med tillhandahållande, tillverkning, underhåll eller användning av vapen och vapenrelaterad materiel av alla slag, däri inbegripet vapen och ammunition, militärfordon och militär utrustning, paramilitär utrustning och reservdelar till ovanstående, direkt eller indirekt till alla fysiska och juridiska personer, enheter eller organ i, eller för användning i, Burma/Myanmar,
b) att tillhandahålla finansiering eller finansiellt stöd som har samband med militär verksamhet, särskilt gåvobistånd, lån och exportkreditförsäkring för all försäljning, leverans, överföring eller export av vapen och vapenrelaterad materiel, direkt eller indirekt till alla personer, enheter eller organ i, eller för användning i, Burma/Myanmar,
c) att medvetet och avsiktligt delta i verksamhet vars syfte eller verkan är att kringgå förbudet enligt a eller b.
Artikel 3
Det skall vara förbjudet
a) att sälja, leverera, överföra eller exportera sådan utrustning enligt bilaga I som kan användas för inhemskt förtryck, oavsett om den har sitt ursprung i gemenskapen eller inte, direkt eller indirekt till alla fysiska eller juridiska personer, enheter eller organ i, eller för användning i, Burma/Myanmar,
b) att tillhandahålla tekniskt stöd som har samband med utrustning enligt a direkt eller indirekt till alla fysiska eller juridiska personer, enheter eller organ i, eller för användning i, Burma/Myanmar,
c) att tillhandahålla finansiering eller finansiellt stöd som har samband med utrustning enligt a direkt eller indirekt till alla fysiska eller juridiska personer, enheter eller organ i, eller för användning i, Burma/Myanmar,
d) att medvetet och avsiktligt delta i verksamhet vars syfte eller verkan är att kringgå förbudet enligt a, b eller c.
Artikel 4
1. Genom avvikelse från artiklarna 2 och 3 får de behöriga myndigheter i medlemsstaterna som förtecknas i bilaga II på de villkor som de anser lämpliga ge tillstånd för
a) försäljning, leverans, överföring eller export av icke-dödsbringande militär utrustning som är avsedd endast för humanitärt bruk eller som skydd, eller för Förenta nationernas, Europeiska unionens och gemenskapens program för institutionsuppbyggnad eller för Europeiska unionens och Förenta nationernas krishanteringsinsatser,
b) försäljning, leverans, överföring eller export av sådan utrustning som kan användas för inhemskt förtryck som är avsedd endast för humanitärt bruk eller som skydd, eller för Förenta nationernas, Europeiska unionens och gemenskapens program för institutionsuppbyggnad eller för Europeiska unionens och Förenta nationernas krishanteringsinsatser,
c) försäljning, leverans, överföring eller export av minröjningsutrustning och material som används i minröjningsinsatser,
d) tillhandahållande av finansiering och finansiellt stöd som har samband med sådan utrustning eller med sådana program och insatser,
e) tillhandahållande av tekniskt stöd som har samband med sådan utrustning eller med sådana program och insatser,
2. De tillstånd som avses i punkt 1 får endast beviljas innan den verksamhet som begäran om tillstånd gäller har inletts.
Artikel 5
Artiklarna 2 och 3 skall inte tillämpas på skyddsdräkter, inbegripet skottsäkra västar och militära hjälmar, som tillfälligt exporteras till Burma/Myanmar av Förenta nationernas, Europeiska unionens, gemenskapens eller dess medlemsstaters personal, mediernas företrädare samt bistånds- och utvecklingsarbetare och åtföljande personal och som är avsedda enbart för deras personliga bruk.
Artikel 6
1. Alla penningmedel och ekonomiska resurser som tillhör eller ägs, innehas eller kontrolleras av i bilaga III förtecknade enskilda medlemmar av Burma/Myanmars regering och till dessa knutna fysiska eller juridiska personer, enheter eller organ skall frysas.
2. Inga tillgångar eller ekonomiska resurser får direkt eller indirekt ställas till förfogande för eller göras tillgängliga för fysiska eller juridiska personer, enheter eller organ som förtecknas i bilaga III.
3. Det skall vara förbjudet att medvetet och avsiktligt delta i verksamhet vars syfte eller verkan är att direkt eller indirekt kringgå de åtgärder som avses i punkterna 1 och 2.
Artikel 7
1. De behöriga myndigheter i medlemsstaterna som förtecknas i bilaga II får ge tillstånd till att vissa frysta penningmedel eller ekonomiska resurser frigörs eller att vissa penningmedel eller ekonomiska resurser görs tillgängliga, på sådana villkor som de finner lämpliga, efter det att de har konstaterat att de berörda penningmedlen eller ekonomiska resurserna är
a) nödvändiga för att tillgodose de grundläggande behoven hos de personer som förtecknas i bilaga III och deras beroende familjemedlemmar, inbegripet betalning av livsmedel, hyra eller amorteringar, mediciner och läkarvård, skatter, försäkringspremier och avgifter för samhällstjänster,
b) avsedda endast för betalning av rimliga arvoden och ersättning för utgifter i samband med tillhandahållande av juridiska tjänster,
c) avsedda endast för betalning av avgifter eller serviceavgifter för rutinmässig hantering eller förvaltning av frysta penningmedel eller ekonomiska resurser,
d) nödvändiga för att täcka extraordinära kostnader, förutsatt att den behöriga myndigheten åtminstone två veckor före tillståndsgivningen har anmält till de övriga behöriga myndigheterna och kommissionen på vilka grunder den anser att ett särskilt tillstånd bör beviljas.
Den behöriga myndigheten skall underrätta de behöriga myndigheterna i övriga medlemsstater samt kommissionen om alla tillstånd som beviljats enligt denna punkt.
2. Artikel 6.2 skall inte tillämpas på kreditering av frysta konton med
i) ränta eller övriga intäkter på dessa konton, eller
ii) betalningar i samband med avtal, överenskommelser eller förpliktelser som ingåtts eller uppkommit före den dag från och med vilken dessa konton omfattas av bestämmelserna i förordningarna (EG) nr 1081/2000, (EG) nr 798/2004 eller av den här förordningen, beroende på vilken dag som infaller först, förutsatt att sådan ränta, sådana övriga intäkter och sådana betalningar fortsatt omfattas av artikel 6.1.
Artikel 8
1. Utan att det påverkar de tillämpliga reglerna om rapportering, sekretess och tystnadsplikt skall fysiska och juridiska personer, enheter och organ
a) omedelbart lämna alla uppgifter som underlättar efterlevnaden av denna förordning, till exempel uppgifter om konton och belopp som frysts i enlighet med artikel 6, till de i bilaga II förtecknade behöriga myndigheterna i de medlemsstater där de är bosatta eller belägna och även vidarebefordra dessa uppgifter till kommissionen, direkt eller genom dessa behöriga myndigheter,
b) samarbeta med de behöriga myndigheter som förtecknas i bilaga II vid alla kontroller av dessa uppgifter.
2. Alla ytterligare uppgifter som kommissionen mottar direkt skall göras tillgängliga för den berörda medlemsstatens behöriga myndigheter.
3. Alla uppgifter som lämnas eller mottas enligt denna artikel får användas endast i de syften för vilka de lämnades eller mottogs.
Artikel 9
1. Följande skall vara förbjudet:
a) Beviljande av alla slags lån eller krediter till de burmesiska statsägda företag som förtecknas i bilaga IV, samt förvärv av obligationer, inlåningsbevis, köpoptioner eller förlagsbevis utfärdade av dessa företag.
b) Förvärv eller utökning av en andel i de burmesiska statsägda företag som förtecknas i bilaga IV, inbegripet fullständigt förvärv av dessa företag och förvärv av andelar och värdepapper som motsvarar andelar.
2. Det skall vara förbjudet att medvetet och avsiktligt delta i verksamhet vars syfte eller verkan är att direkt eller indirekt kringgå bestämmelserna i punkt 1.
3. Punkt 1 skall inte påverka genomförandet av handelsavtal om leverans av varor eller tjänster på sedvanliga kommersiella betalningsvillkor, eller vanliga kompletterande överenskommelser i samband med genomförandet av dessa avtal, t.ex. exportkreditförsäkringar.
4. Bestämmelserna i punkt 1 a skall inte påverka genomförandet av en skyldighet i enlighet med kontrakt eller avtal som har ingåtts före den 25 oktober 2004.
5. Förbudet i punkt 1 b skall inte förhindra en utökning av en andel i de burmesiska statsägda företag som förtecknas i bilaga IV, om utökningen är tvingande enligt ett avtal som har ingåtts med det berörda burmesiska statsägda företaget före den 25 oktober 2004. Den berörda behöriga myndigheten enligt förteckningen i bilaga II samt kommissionen skall underrättas före en sådan transaktion. Kommissionen skall underrätta de behöriga myndigheterna i övriga medlemsstater.
Artikel 10
Frysning av penningmedel och ekonomiska resurser eller vägran att tillgängliggöra penningmedel eller ekonomiska resurser, som utförs i god tro att denna åtgärd sker i enlighet med den här förordningen, skall inte medföra ansvar av något slag för den fysiska eller juridiska person eller enhet som vidtar åtgärder, eller för dess ledning eller anställda, såvida det inte kan bevisas att penningmedlen och de ekonomiska resurserna frystes på grund av vårdslöshet.
Artikel 11
Kommissionen och medlemsstaterna skall omedelbart underrätta varandra om de åtgärder som vidtas enligt den här förordningen och lämna varandra alla relevanta upplysningar som de förfogar över med anknytning till den här förordningen, särskilt upplysningar om överträdelser, problem med genomförandet samt domar som avkunnats av nationella domstolar.
Artikel 12
Kommissionen skall ha rätt att
a) ändra bilaga II på grundval av upplysningar som lämnas av medlemsstaterna, och
b) ändra bilagorna III och IV på grundval av beslut som fattas rörande bilagorna I och II till gemensam ståndpunkt 2006/…/GUSP.
Artikel 13
1. Medlemsstaterna skall fastställa regler om påföljder vid överträdelse av bestämmelserna i denna förordning och vidta alla nödvändiga åtgärder för att se till att reglerna tillämpas. Påföljderna skall vara effektiva, proportionella och avskräckande.
2. Medlemsstaterna skall underrätta kommissionen om dessa regler så snart som denna förordning har trätt i kraft och underrätta kommissionen om eventuella senare ändringar.
Artikel 14
Denna förordning skall tillämpas
a) inom gemenskapens territorium, inbegripet dess luftrum,
b) ombord på alla flygplan och fartyg som omfattas av en medlemsstats jurisdiktion,
c) på varje person inom eller utanför gemenskapens territorium, som är medborgare i en medlemsstat,
d) på varje juridisk person, enhet eller organ som har inrättats eller bildats i enlighet med en medlemsstats lagstiftning,
e) på varje juridisk person, enhet eller organ med avseende på varje form av affärsverksamhet som helt eller delvis bedrivs i gemenskapen.
Artikel 15
Förordning (EG) nr 798/2004 skall upphöra att gälla.
Artikel 16
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
[pic] | EUROPEISKA GEMENSKAPERNAS KOMMISSION |
Bryssel den 26.9.2006
KOM(2006) 548 slutlig
2005/0043 (COD)
MEDDELANDE FRÅN KOMMISSIONEN TILL EUROPAPARLAMENTET enligt artikel 251.2 andra stycket i EG-fördraget om
gemensam ståndpunkt antagen av rådet inför antagandet av Europaparlamentets och rådets beslut om Europeiska gemenskapens sjunde ramprogram för verksamhet inom området forskning, teknisk utveckling och demonstration (2007–2013)
2005/0043 (COD)
MEDDELANDE FRÅN KOMMISSIONEN TILL EUROPAPARLAMENTET enligt artikel 251.2 andra stycket i EG-fördraget om
gemensam ståndpunkt antagen av rådet inför antagandet av Europaparlamentets och rådets beslut om Europeiska gemenskapens sjunde ramprogram för verksamhet inom området forskning, teknisk utveckling och demonstration (2007–2013)
1. BAKGRUND
Datum för överlämnande av förslaget till Europaparlamentet och rådet (dokument KOM(2005) 119 slutlig, 2005/0043(COD) och 2005/0044(CNS)): | 13 april 2005 |
Datum för Regionkommitténs yttrande: | 16 november 2005 |
Datum för Europeiska ekonomiska och sociala kommitténs yttrande: | 14 december 2005 |
Datum för Europaparlamentets yttrande efter första behandlingen: | 15 juni 2006 |
Datum för överlämnande av det ändrade förslaget till Europaparlamentet och rådet: | 28 juni 2006 |
Datum för antagande av den gemensamma ståndpunkten: | 25 september 2006 |
2. Kommissionens synpunkter på den gemensamma ståndpunkten
I enlighet med artikel 251 i EG-fördraget innehåller det här meddelandet kommissionens synpunkter på rådets gemensamma ståndpunkt, som den 25 september 2006 antogs med kvalificerad majoritet, om sjunde ramprogrammet för verksamhet inom området forskning och teknisk utveckling, efter det att politisk enighet uppnåtts den 24 juli 2006. Den 24 juli 2006 uppnåddes även politisk enighet om Euratomramprogrammet.
Allmänt sett har den gemensamma ståndpunkten samma struktur och innehåll som kommissionens förslag till ramprogram och överensstämmer generellt med Europaparlamentets yttrande.
Rådet har tagit med en stor del av de ändringsförslag som ingick i yttrandet som Europaparlamentet antog vid den första behandlingen (15 juni 2006) och som kommissionen antog i sitt ändrade förslag.[1]
3. Kommentarer till den gemensamma ståndpunkten
Kommissionen anser att den gemensamma ståndpunkten är en god utgångspunkt för ytterligare förhandlingar om ramprogrammet med målet att nå en överenskommelse vid andra behandlingen.
I fråga om budgeten har rådet (och Europaparlamentet) godkänt det totala belopp på 50 521 miljoner euro som kommissionen föreslog i sitt ändrade förslag[2], efter det att Europaparlamentet, rådet och kommissionen den 17 maj 2006 ingick ett interinstitutionellt avtal om budgetdisciplin och sund ekonomisk förvaltning .[3]
Beträffande uppdelningen av budgeten överensstämmer den gemensamma ståndpunkten i stort med kommissionens ändrade förslag och Europaparlamentets yttrande, förutom i följande:
- I fråga om programmet Samarbete
- Ökade belopp för följande fem teman : Hälsa, Nanovetenskap, nanoteknik, material och ny produktionsteknik, Energi, Miljö samt en liten ökning för Samhällsvetenskap och humaniora.
- Minskade anslag för temat Säkerhets- och rymdforskning.
- I fråga om programmet Kapacitet:
- Större minskning för temat Forskningsinfrastruktur samt minskade anslag för Vetenskapen i samhället.
- Ökade belopp för Forskning till förmån för små och medelstora företag, Forskningspotential samt en liten ökning för Övergripande internationellt samarbete.
Även om det finns en stark koppling mellan de föreslagna verksamheterna och den föreslagna budgeten, kan den krympta budgeten för Infrastruktur och temat Säkerhets- och rymdforskning leda till att de verksamheter som föreslås i den gemensamma ståndpunkten inte förverkligas fullt ut.
Beträffande programmets struktur bibehåller den gemensamma ståndpunkten kommissionens förslag till de olika delarna i programmet, även fokuseringen på teman och flexibiliteten i programmet med beaktande av dess varaktighet på sju år. Kommissionen delar uppfattningen att en sammanhängande utveckling av politiken bör utgöra en separat del av programmet Kapaciteter. Rådet har dock, i likhet med parlamentet, delat upp temat Säkerhets-och rymdforskning i två, och föreslår följaktligen tio teman. Enligt kommissionen kan man uppnå betydande flexibilitet och synergieffekter om man håller ihop de två temana.
Beträffande forskningsinnehållet innehåller den gemensamma ståndpunkten en stor del av de ändringar som Europaparlamentet föreslagit och som kommissionen godkänt och införlivat i sitt ändrade förslag. I sitt ändrade förslag klargjorde kommissionen att beroende på den minskade budgeten, hade den inte tagit med ändringar som skulle innebära att temana fick bredare omfattning, vilket skulle kräva mer resurser. Kommissionen anser att den gemensamma ståndpunkten som helhet respekterar detta. Att ta med ”Exploratory Award Scheme” för små och medelstora företag i temat Kapaciteter överensstämmer inte med den här principen. Kommissionen anser att budgeten enbart bör koncentreras på finansiering av projekt.
Kommissionen stöder förslaget att skärpa texten om små och medelstora företag genom att föreslå konkreta åtgärder i temana, till exempel genom kvantitativ och kvalitativ analys. Enligt kommissionen är det effektivare än artificiella mål som kommissionen inte tog med i det ändrade förslaget.
För parlamentet har de gemensamma teknikinitiativen samt programmen Idéer och Människor varit viktiga frågor.
- I fråga om de gemensamma teknikinitiativen innehåller den gemensamma ståndpunkten ändringarna av kriterierna för identifieringen av dessa initiativ.
- I fråga om programmet Idéer har viktiga förtydliganden infogats i fråga om mandatperioden, förnyelse av det vetenskapliga rådet och dess roll, ledningen och personalfrågor. Även genomförandet av en oberoende genomgång 2010 av Europeiska forskningsrådets struktur och mekanismer, som skall läggas fram för Europaparlamentet och rådet, har infogats.
- I fråga om programmet Människor innehåller en serie ändringar hänvisningar till kopplingar mellan det här programmet och andra delar av ramprogrammet samt andra gemenskapsprogram. Dessa tillägg tydliggör den internationella dimensionen hos den här delen av programmet och innehåller förslag på att skapa lämpliga arbetsvillkor för forskare och instruktioner i fråga om samfinansiering.
Slutligen har kriterierna för stödet till nya forskningsinfrastrukturer gjorts mer detaljerade och vikten av regionala aspekter vid upprättandet erkänns.
I fråga om stamcellsrelalerad forskning godtog kommissionen i sitt ändrade förslag att infoga en artikel om vilka områden som inte skall finansieras inom sjunde ramprogrammet, vilket överensstämde med parlamentets ändringsförslag. Rådet tog även med den här artikeln i sin gemensamma ståndpunkt, och kommissionen bekräftade ännu en gång de metoder som skulle användas (se bilagan).
4. SLUTSATS
Kommissionen anser att den gemensamma ståndpunkten, som antogs med kvalificerad majoritet den 25 september 2006 i mycket hög utsträckning överensstämmer med både Europaparlamentets och kommissionens ståndpunkter. Den beaktar till stor del de ändringsförslag som Europaparlamentet lade fram efter första behandlingen och som kommissionen införlivat i sitt ändrade förslag. Kommissionen ställer sig därför bakom den gemensamma ståndpunkten.
[pic] | EUROPEISKA GEMENSKAPERNAS KOMMISSION |
Bryssel den 12.10.2006
KOM(2006) 564 slutlig
2006/0194 (CNS)
Förslag till
RÅDETS FÖRORDNING om gemenskapens finansiella bidrag till Internationella fonden för Irland (2007-2010)
(framlagt av kommissionen) {SEK(2006) 1227}
MOTIVERING
Internationella fonden för Irland (IFI) inrättades 1986 för att bidra till att genomföra artikel 10 a i det engelsk-irländska avtalet av den 15 november 1985 där det föreskrivs att de två regeringarna skall samarbeta för att främja ekonomisk och social utveckling i de områden i de båda delarna av Irland som har utstått de svåraste lidandena på grund av de närmast föregående årens instabila situation, och att de skall undersöka möjligheterna att få internationellt stöd för detta.
IFI:s mål är att uppmuntra ekonomisk och social utveckling, och att främja kontakt, dialog och försoning mellan nationalister och unionister i hela Irland*.
Efter att Förenta staterna och andra länder redan på ett tidigt stadium lämnat bidrag till dessa strävanden framhöll Europeiska gemenskapen att IFI:s mål låg i linje med de egna målen, vilket resulterade i att även gemenskapen i praktisk handling ville stödja detta initiativ. Gemenskapens bidrag till IFI började betalas ut 1989. EG-stödet utgör nu ca 48 % av de årliga bidragen till fonden och 40 % av de samlade bidragen hittills. Alltsedan början av 1989 har kommissionen företrätts av en observatör vid fondens samtliga styrelsemöten.
Det politiska läget i regionen har förändrats under åren: 1994 proklamerade de mest inflytelserika paramilitära grupperna vapenvila. Genom Belfastavtalet (”långfredagsavtalet”) i april 1998 lades den politiska grunden för en fredsprocess, som inbegrep ett begränsat självstyre med ett nordirländskt parlament (”Assembly”) och en regering (”Executive”) som båda inrättades i slutet av 1999. Det förekommer dock fortfarande en hel del säkerhetsrelaterade incidenter som har samband med religiös tillhörighet, och det psykologiska och fysiska avståndet ökar mellan de största befolkningsgrupperna. Det nordirländska parlamentets verksamhet är för närvarande avbruten, vilket belyser det hot och den osäkerhet som omger fredsprocessen i regionen.
Mot denna bakgrund är ekonomisk och social utveckling till stöd för fred och försoning på gräsrotsnivå en långsiktig process. Som ett instrument för att uppnå detta mål är IFI ett komplement till de insatser som görs genom EU:s program för fred och försoning i Nordirland och de angränsande grevskapen i Irland (”Peace I” 1995–1999, ”Peace II” 2000–2006 och ”Peace III” 2007–2013).
Internationella fonden är dock medveten om att det internationella stödet inte kan fortsätta på samma nivå utan tidsbegränsning, och den gjorde därför en översyn av sina strukturer och prioriteringar 2005 för att anpassa sitt uppdrag till de faktiska förhållandena, och den har antagit en strategi som innebär att fondens verksamhet upphör 2010. Denna strategi går under namnet ”Sharing this Space” och omfattar den sista fasen av fondens verksamhet (2006–2010). Under denna period kommer fonden att koncentrera sig på de områden där behovet är störst och försöka se till att dess arbete får långsiktiga effekter.
I enlighet med förordningen om den nuvarande bidragsrundan**, har Europeiska kommissionen också lagt fram en rapport med en bedömning av IFI:s verksamhet för budgetmyndigheten***. I denna framhålls IFI:s mycket värdefulla och positiva insatser för fred och försoning i regionen och därmed till uppfyllandet av målen. I slutsatserna anges det att kommissionen anser att finansieringen efter 2006 bör beviljas på grundval av de iakttagelser som gjorts i rapporten, vilket skulle kunna ske antingen genom att rådet antar en ny förordning om EG:s bidrag till IFI, eller genom andra lämpliga samarbetsformer mellan kommissionen och IFI.
Mot bakgrund av denna bedömning föreslås det att EU ger 15 miljoner euro i bidrag per år till IFI under en period av ytterligare fyra år. Denna föreslagna nya period kommer således att löpa ut 2010, samtidigt som IFI:s verksamhet upphör.
Den nya rådsförordningen bör också återspegla iakttagelserna i kommissionens rapport, särskilt dem som ger bättre synergieffekter i fråga om mål och samordning med strukturfondernas insatser, i synnerhet det nya Peace-programmet och bestämmelserna om avveckling.
Paketet med förslag som väntar på att antas omfattar följande:
- Förslag till rådets förordning om gemenskapens finansiella bidrag till Internationella fonden för Irland (2007–2010).
- Kommissionens meddelande: Rapport om Internationella fonden för Irland enligt artikel 5 i rådets förordning (EG) nr 177/2005.
2006/0194 (CNS)
Förslag till
RÅDETS FÖRORDNING
om gemenskapens finansiella bidrag till Internationella fonden för Irland (2007-2010)
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 308,
med beaktande av kommissionens förslag[1],
med beaktande av Europaparlamentets yttrande[2], och
av följande skäl:
(1) Internationella fonden för Irland (nedan kallad ”fonden”) inrättades 1986 genom avtalet av den 18 september 1986 mellan Irlands regering och regeringen i Förenade konungariket Storbritannien och Nordirland beträffande Internationella fonden för Irland (nedan kallat ”avtalet”), i syfte att främja ekonomiska och sociala framsteg, uppmuntra till kontakter, dialog och försoning mellan nationalister och unionister över hela Irland och därmed till uppnåendet av ett av de mål som anges i det engelsk-irländska avtalet av den 15 november 1985.
(2) Gemenskapen har sedan 1989 gett finansiellt bidrag till fonden. För perioden 2005–2006 anslogs det, i enlighet med rådets förordning (EG) nr 177/2005 av den 24 januari 2005 om gemenskapens finansiella bidrag till Internationella fonden för Irland (2005–2006)[3], 15 miljoner euro från gemenskapens budget för vart och ett av åren 2005 och 2006. Den förordningen upphör att gälla den 31 december 2006.
(3) Vid de bedömningar som har gjorts i enlighet med artikel 5 i rådets förordning (EG) nr 177/2005 har det bekräftats att det finns ett behov av ytterligare stöd till fondens verksamhet och av bättre synergieffekter i fråga om mål och samordning med strukturfondsinsatserna, i synnerhet med det särskilda program för fred och försoning i Nordirland och de angränsande grevskapen i Irland (nedan kallat ”Peace-programmet”) som inrättats i enlighet med rådets förordning (EG) nr 1260/1999 av den 21 juni 1999 om allmänna bestämmelser för strukturfonderna[4].
(4) Fredsprocessen i Nordirland kräver fortsatt stöd till fonden från gemenskapen även efter den 31 december 2006. Som ett erkännande av de särskilda ansträngningar som gjorts för fredsprocessen har Peace-programmet fått ytterligare stöd från strukturfonderna för perioden 2007–2013, i enlighet med punkt 22 i bilaga II till rådets förordning (EG) nr 1083/2006 av den 11 juli 2006 om allmänna bestämmelser för Europeiska regionala utvecklingsfonden, Europeiska socialfonden och Sammanhållningsfonden samt om upphävande av förordning (EG) nr 1260/1999[5].
(5) Vid sitt möte i Bryssel den 15–16 december 2005 riktade Europeiska rådet en uppmaning till kommissionen om att vidta nödvändiga åtgärder för fortsatt gemenskapsstöd till fonden inför den viktiga slutfasen av dess arbete fram till 2010.
(6) Gemenskapens bidrag till fonden bör utgöras av finansiella bidrag under 2007, 2008, 2009 och 2010, vilket innebär att de avslutas samtidigt med fonden.
(7) Vid fördelningen av gemenskapens bidrag bör fonden prioritera projekt som involverar människor från båda sidor av gränsen eller från båda befolkningsgrupperna och på ett sådant sätt att de kompletterar de insatser som finansieras genom Peace-programmet under perioden 2007–2010.
(8) I enlighet med avtalet deltar samtliga bidragsgivare till fonden som observatörer i de möten som hålls i styrelsen för Internationella fonden för Irland.
(9) Det är av avgörande betydelse att det finns en nära samordning mellan fondens verksamhet och de insatser som finansieras genom gemenskapens strukturfonder enligt artikel 159 i fördraget, särskilt Peace-programmet.
(10) Stödet från fonden bör betraktas som effektivt endast om det leder till hållbara ekonomiska och sociala förbättringar, och om det inte ersätter annan offentlig eller privat finansiering.
(11) Det bör göras en översyn av bestämmelserna om avveckling av fonden före den 1 juli 2008.
(12) Ett finansiellt referensbelopp enligt punkt 38 i det interinstitutionella avtalet av den 17 maj 2006 mellan Europaparlamentet, rådet och kommissionen om budgetdisciplin och sund ekonomisk förvaltning[6] har införts i denna förordning för hela den tid som programmet pågår, utan att detta påverkar budgetmyndighetens befogenheter enligt fördraget.
(13) Gemenskapens bidrag till fonden bör uppgå till 15 miljoner euro för vart och ett av åren 2007, 2008, 2009 och 2010, uttryckt i löpande penningvärde.
(14) Detta stöd kommer att bidra till att stärka solidariteten mellan medlemsstaterna och mellan folken.
(15) Fördraget innehåller inte några andra befogenheter för att anta denna förordning än de som anges i artikel 308.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
Det finansiella referensbeloppet för Internationella fonden för Irland (nedan kallad ”fonden”) för perioden 2007–2010 skall vara 60 miljoner euro.
De årliga anslagen skall beviljas av budgetmyndigheten enligt riktlinjerna i finansieringsramen.
Artikel 2
Fonden skall använda bidraget i enlighet med avtalet av den 18 september 1986 mellan Irlands regering och regeringen i Förenade konungariket Storbritannien och Nordirland beträffande Internationella fonden för Irland (nedan kallat ”avtalet”).
Vid fördelningen av bidraget skall fonden prioritera projekt som genomförs över gränsen eller mellan befolkningsgrupperna, på ett sådant sätt att de kompletterar de insatser som finansieras genom strukturfonderna, särskilt Peace-programmets verksamhet i Nordirland och de angränsande grevskapen i Irland.
Bidraget skall användas på ett sådant sätt att det leder till hållbar ekonomisk och social förbättring i de berörda områdena. Det får inte användas för att ersätta annan offentlig eller privat finansiering.
Artikel 3
Kommissionen skall företräda gemenskapen som observatör vid mötena i fondens styrelse (nedan kallad ”styrelsen”).
Fonden skall företrädas genom en observatör vid de möten som Peace-programmets och andra strukturfondsprograms övervakningskommittéer håller.
Artikel 4
Kommissionen skall tillsammans med fondens styrelse fastställa lämpliga förfaranden för att främja samordning på alla nivåer mellan fonden och de förvaltningsmyndigheter och genomförandeorgan som inrättats för de berörda strukturfondsinsatserna, särskilt inom ramen för Peace-programmet.
Artikel 5
Kommissionen skall i samarbete med fondens styrelse fastställa lämpliga förfaranden för offentliggörande och information i syfte att sprida kunskap om gemenskapens bidrag till de projekt som finansieras av fonden.
Artikel 6
Senast den 30 juni 2008 skall fonden till kommissionen överlämna sin strategi för att avveckla fondens verksamhet, inklusive
a) en handlingsplan med förväntade utbetalningar och förväntat avvecklingsdatum,
b) principer för återtagande av medel,
c) hantering av eventuella resterande belopp och ränta vid fondens avveckling.
Senare utbetalningar till fonden är beroende av kommissionens godkännande av avvecklingsstrategin. Om strategin inte har lagts fram senast den 30 juni 2008 skall utbetalningarna till fonden stoppas tills strategin har mottagits.
Artikel 7
1. Kommissionen skall förvalta bidragen.
Om inte annat följer av punkt 2 skall det årliga bidraget överföras genom delutbetalningar enligt följande:
a) Ett första förskott på 40 % skall betalas ut efter att kommissionen har mottagit ett åtagande som undertecknats av fondens styrelseordförande, och av vilket det framgår att fonden skall uppfylla villkoren för beviljande av det bidrag som fastställs i denna förordning.
b) Ett andra förskott på 40 % skall betalas ut sex månader senare.
c) En slutlig utbetalning på 20 % skall göras efter att kommissionen har mottagit och godkänt fondens årliga verksamhetsrapport och reviderade räkenskaper för året i fråga.
2. Innan en delutbetalning görs skall kommissionen göra en bedömning av fondens finansiella behov på grundval av fondens kassabehållning vid tidpunkten för varje planerad utbetalning. Om bedömningen är att fondens finansiella behov inte motiverar en av delutbetalningarna skall denna utbetalning skjutas upp. Kommissionen skall se över detta beslut på grundval av ny information från fonden och fortsätta utbetalningarna så snart som dessa anses vara motiverade.
Artikel 8
Ett bidrag från fonden får betalas ut till en insats som tar emot eller som skall ta emot finansiellt bistånd från strukturfonderna endast om summan av det finansiella biståndet plus 40 % av bidraget från fonden uppgår till högst 75 % av de totala stödberättigande kostnaderna.
Artikel 9
En slutrapport skall överlämnas till kommissionen sex månader före det datum för fondens avveckling som förutses i strategin för avveckling och som avses i artikel 6.1 a eller sex månader efter kommissionens sista utbetalning, beroende på vilket som infaller först, och den skall omfatta all nödvändig information som kan möjliggöra för kommissionen att utvärdera genomförandet av biståndet och måluppfyllelsen.
Artikel 10
Bidraget för det sista året skall betalas ut efter den analys av fondens finansiella behov som avses i artikel 7.2 och förutsatt att fondens verksamhet bedrivs i överensstämmelse med den strategi för avveckling som föreskrivs i artikel 6.
Artikel 11
Slutdatum för stödberättigande utgifter skall vara den 31 december 2013.
Artikel 12
Denna förordning träder i kraft den 1 januari 2007.
Den löper ut den 31 december 2010.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
[pic] | EUROPEISKA GEMENSKAPERNAS KOMMISSION |
Bryssel den 9.10.2006
KOM(2006) 579 slutlig
2006/0184 (CNS)
Förslag till
RÅDETS BESLUT
om makroekonomiskt stöd till Republiken Moldavien
(framlagt av kommissionen) {SEK(2006) 1258}
MOTIVERING
BAKGRUND |
110 | Motiv och syfte Kommissionen föreslår att Moldavien skall ges makroekonomiskt stöd på maximalt 45 miljoner euro i form av ett bidrag i syfte att stödja betalningsbalansen och bygga upp valutareserven. Det föreslagna stödet kommer att hjälpa Moldavien att klara de ekonomiska påfrestningar som genomförandet av landets ekonomiska program innebär. Det kommer också att underlätta och uppmuntra myndigheternas insatser för att genomföra reformer inom ramen för handlingsplanen för den europeiska grannskapspolitiken för EU-Moldavien och strategidokumentet för ökad tillväxt och fattigdomsminskning. Det föreslagna makroekonomiska stödet kommer att vara av engångskaraktär, tidsbegränsat och komplettera stödet från Bretton Woods-institutioner, bilaterala givare och Parisklubben. Det kommer dessutom att ges på villkor att framsteg görs, framför allt i genomförandet av den IMF-stödda överenskommelsen om mekanismen för ökad tillväxt och fattigdomsminskning. Stödet kommer i ett skede när förbindelserna mellan EU och Moldavien går in i en ny och djupare fas inom ramen för den europeiska grannskapspolitiken. |
120 | Allmän bakgrund I inledningen av övergången till marknadsekonomi genomförde Moldavien flera reformer av första generationen. I slutet av 90-talet och början av 2000-talet minskade dock reformtakten och regeringens administrativa påverkan på ekonomin ökade. Mot den bakgrunden avbröts policybaserade lån från Bretton Woods-institutionerna. Två makroekonomiska EU-stöd till Moldavien, ett lån på 15 miljoner euro som det fattades beslut om år 2000 och ett bidrag på samma belopp som det beslutades om 2002[1], kunde därför inte genomföras. Under den perioden ökade Moldaviens BNP med 7 % per år. Tillväxten har drivits på av inhemsk efterfrågan som eldats på av starkt stigande antal överföringar som ökat till mer än 30 % av BNP. Från år 2000 till 2005 mer än fördubblades Moldaviens BNP per capita (räknat i dollar). Det hindrar inte att landets BNP är den överlägset lägsta i Europa på 812 dollar. Moldavien är det enda land i Europa som Världsbanken klassificerar som låginkomstland. Under 2004-2005 kom strukturreformer åter upp på den politiska dagordningen i Moldavien, vilket framförallt tog sig uttryck i att regeringen antog strategidokumentet för ökad tillväxt och fattigdomsminskning. Regeringens reformambitioner har fått ytterligare näring av EU-ambitionerna, som bekräftades genom antagandet i februari 2005 av handlingsplanen för den europeiska grannskapspolitiken för EU-Moldavien. Under större delen av 2005 förde regeringen en ekonomisk politik som skulle illustrera den förnyade stabiliteten och reformbeslutsamheten. Mot bakgrund av de resultat som i slutet av 2005 uppnåtts, återupptog IMF diskussionerna om ett nytt program som skulle kunna få stöd genom ett finansieringsavtal med fonden. I februari 2006 uppnåddes en överenskommelse om villkoren för programmet och i maj 2006 godkände IMF:s styrelse ett treårigt finansieringsavtal inom ramen för mekanismen för fattigdomsminskning och ökad tillväxt. Godkännandet av avtalet följdes av en överenskommelse med Moldaviens officiella fordringsägare i Parisklubben om en omstrukturering av ackumulerade skulder och löpande betalningar som skall betalas under programperioden på de så kallade Houstonvillkoren. Ett av målen för arrangemanget var att hjälpa regeringen att normalisera Moldaviens förhållande till de officiella långivarna. Programmet för ökad tillväxt och fattigdomsminskning är utformat för att bibehålla makroekonomisk stabilitet och på så sätt stödja tillväxt och fattigdomsminskning, inte minst mot bakgrund av ett fortsatt starkt inflöde av överföringar och betydligt högre priser på importerad energi. Enligt programmet måste myndigheterna begränsa budgetunderskottet till 0,5 % av BNP och centralbanken har som mål att till slutet av 2008 öka valutareserven till motsvarande tre månaders import. De prioriterade åtgärderna för strukturpolitiken kommer främst att ske på områdena avreglering av utrikeshandeln, styrning av företag, reformering av banksektorn och skatteförvaltning. När programmet antogs antog man att de föreslagna åtgärderna skulle leda till en BNP-tillväxt på 6 % under 2006 och 5 % perioden 2007-2008, en gradvis minskning av inflationen till cirka 7 % i slutet av 2008 och ett underskott i bytesbalansen på omkring 5 % av BNP. Programmet skall dock genomföras under synnerligen svåra förhållanden. Beroende på enorma oljeprishöjningar försämrades Moldaviens handels- och bytesbalans kraftigt redan 2005. Sedan början av 2006 har Moldavien drabbats av ytterligare chocker som drabbat betalningsbalansen. Till exempel beslöt det ryska gasmonopolet Gazprom i januari 2006 att öka gaspriserna från 80 dollar per tusen kubikmeter till 110 dollar, och till 160 dollar i juli och Moldaviens export av vin och alkohol till Ryssland förbjöds. Sammantaget gör det utsikterna för att uppnå målen i PRGF-programmet mycket dystra. Moldaviens försvagade utrikeshandel kommer också att försvåra för regeringen att uppnå sina mål på medellång sikt i fråga om tillväxt och fattigdomsminskning som ingår i regeringens strategidokument för ökad tillväxt och fattigdomsminskning, och målen i handlingsplanen för den europeiska grannskapspolitiken för EU och Moldavien. Den ekonomiska utvecklingen i Moldavien kommer först och främst att kräva vissa ändringar av programmet för ökad tillväxt och fattigdomsminskning samt ytterligare finansiering av engångskaraktär förutom den finansiering som för närvarande finns. EU har vid flera tillfällen bistått Moldavien med makroekonomiskt stöd i syfte att lindra de chocker betalningsbalansen utsatts för. Kommissionen anser att dagens situation motiverar att ytterligare resurser förs över till samma instrument. Det makroekonomiska stödet från EU skulle bidra till Moldaviens externa finansieringsbehov under 2007 och 2008. Det kan också motiveras av det fördjupade samarbetet mellan EU och Moldavien inom ramen för den europeiska grannskapspolitiken. Sedan grannskapspolitiken lanserades 2004 är Moldavien ett av EU:s partnerländer. Tillsammans med Ukraina är Moldavien också det enda östeuropeiska grannskapsland som för närvarande genomför handlingsplanen för den europeiska grannskapspolitiken. Grannskapspolitiken har som mål att utveckla ett allt djupare förhållande mellan EU och partnerländerna, som går längre än det hittillsvarande samarbetet och som omfattar ett intensivare politiskt samarbete, till exempel inom utrikes- och säkerhetspolitik. Vidare syftar den till att främja den ekonomiska utvecklingen och fattigdomsminskningen. |
130 | Gällande bestämmelser Inga. |
140 | Förenlighet med Europeiska unionens politik och mål på andra områden Sedan grannskapspolitiken inleddes har relationerna mellan EU och Moldavien fördjupats. Gemenskapens stöd genom det makroekonomiska stödinstrumentet skulle bidra till att stärka de bilaterala relationerna med Moldavien. Enligt planerna kommer det europeiska grannskaps- och partnerskapsinstrumentet att göras tillgängligt för Moldavien 2007 och framåt. Det medger stöd även i form av budgetstöd. Förberedelserna av program för sektoriellt och/eller allmänt budgetstöd som gynnar Moldavien förväntas inledas så snart som grannskaps- och partnerskapsinstrumentet träder i kraft. Inga utbetalningar inom ramen för budgetstödet till det instrumentet väntas inom den närmaste framtiden. Det instrument för budgetstöd inom grannskaps- och partnerskapsinstrumentet som är avsett att stödja strukturpolitiken på medellång till lång sikt är inte särskilt välavpassat till Moldaviens aktuella problem, som till stor del på chocker som påverkar den kortsiktiga betalningsbalansen. Finansiering genom instrumentet för makroekonomiskt stöd förväntas bli tillgänglig i god tid före ett eventuellt budgetstöd inom ramen för grannskaps- och partnerskapsinstrumentet. Det makroekonomiska stödet, som ett kortsiktigt instrument, kommer att inriktas på Moldaviens akuta externa finansieringsbehov som beror på en kraftig försämring av det externa ekonomiska klimatet. Under övergångsperioden kommer det makroekonomiska stödet också att stödja de strukturreformer som diskuteras i handlingsplanen för EU och Moldavien och i strategidokumentet för ökad tillväxt och fattigdomsminskning. |
SAMRÅD MED BERÖRDA PARTER OCH KONSEKVENSANALYS |
Samråd med berörda parter |
219 | I maj 2006 begärde Moldaviens finansminister Mihail Pop ekonomiskt stöd från EG. Kommissionens berörda avdelningar har varit i kontakt med IMF, Världsbanken och bilaterala givare under förberedelserna av detta förslag från kommissionen för att diskutera vilka stödbehov som finns. Under arbetet med förslaget har kommissionen också rådfrågat Ekonomiska och finansiella kommittén. Efter det att rådets beslut har antagits kommer kommissionens avdelningar att förhandla fram ett samförståndsavtal med Moldaviens myndigheter och en bidragsöverenskommelse för att fastställa närmare bestämmelser för genomförandet. |
Extern experthjälp |
229 | Någon extern experthjälp har inte behövts. |
230 | Konsekvensanalys Eftersom det makroekonomiska stödet är ett policybaserat instrument lämpar det sig särskilt väl för att stödja Moldaviens myndigheters satsning på att förbättra de offentliga finansernas hållbarhet på kort till medellång sikt. Makroekonomiskt stöd kommer att få omedelbara konsekvenser för Moldaviens betalningsbalans och valutareserver och kommer att på så sätt bidra till att lindra de ekonomiska påfrestningarna förknippade med genomförandet av myndigheternas ekonomiska program. Stödet från EG kommer också att underlätta för myndigheterna att genomföra de åtgärder på kort och medellång sikt som anges i handlingsplanen för den europeiska grannskapspolitiken för EU-Moldavien och strategidokumentet för ökad tillväxt och fattigdomsminskning. |
RÄTTSLIGA ASPEKTER |
305 | Sammanfattning av den föreslagna åtgärden Kommissionen skall ge Moldavien makroekonomiskt stöd i form av ett bidrag på högst 45 miljoner euro. Stödet kommer att betalas ut i tre delutbetalningar under en tvåårsperiod. Programmets genomförandeperiod kan komma att utökas med ett år. Stödet förvaltas av kommissionen som tillsammans med myndigheterna skall fastställa de särskilda ekonomisk-politiska och finansiella villkoren knutna till bidragsutbetalningarna. Man kommer att ta hänsyn till särskilda bestämmelser för att förhindra bedrägerier och oegentligheter i enlighet med budgetförordningen. |
310 | Rättslig grund Artikel 308 i fördraget. |
329 | Subsidiaritetsprincipen Förslaget avser ett område där gemenskapen är ensam behörig. Subsidiaritetsprincipen är därför inte tillämplig. |
Proportionalitetsprincipen Förslaget är förenligt med proportionalitetsprincipen av följande skäl: |
331 | Stödet uppgår grovt räknat till en tredjedel av Moldaviens finansieringsbehov för åren 2007-2008, som täcks av stödet. Eftersom Moldavien får stöd av bilaterala givare och långivare samt internationella givare i allmänhet anses detta vara en lämplig fördelning av bördorna för gemenskapen. Stödet kommer att vara fullständigt förenligt med de makroekonomiska mål som finns angivna i Moldaviens dokument över landets ekonomiska politik, till exempel avsiktsförklaringen och avtalet om ekonomiska och finansiella frågor i avtalet om ökad tillväxt och fattigdomsbekämpning med IMF, godkänt i maj 2006. Det kommer också att vara förenligt med de långsiktiga mål som diskuterades i strategidokumentet för ökad tillväxt och fattigdomsminskning i maj 2004 och med handlingsplanen för grannskapspolitiken EU och Moldavien som antogs i februari 2005. Vad gäller de särskilda villkoren som skall knytas till utbetalningen av bidraget kommer kommissionen att koncentrera sig på ett begränsat antal områden, och i synnerhet förvaltning av offentliga medel. Kommissionen kan också överväga att rikta stödet mot viss sektorspolitik av särskilt intresse och som ringats in som sådan i handlingsplanen för grannskapspolitiken för EU och Moldavien. |
Val av regleringsform |
341 | Föreslagen regleringsform: annan. |
342 | Övriga regleringsformer skulle vara olämpliga av följande skäl: I avsaknad av en ramförordning för den makroekonomiska stödordningen är särskilda beslut för ändamålet i rådet enligt artikel 308 i fördraget det enda tillgängliga rättsliga instrumentet för detta stöd. |
BUDGETKONSEKVENSER |
401 | Stödet skulle finansieras genom åtagandebemyndiganden under 2007 under budgetrubrik 01 03 02 (makroekonomiskt stöd), under förutsättning att EG-budgeten för 2007 godkänns, med utbetalningar under 2007 och 2008. |
ÖVRIGA UPPLYSNINGAR |
Översyn/ändring/tidsbegränsning |
533 | Förslaget innehåller en bestämmelse om tidsbegränsning. |
1. 2006/0184 (CNS)
Förslag till
RÅDETS BESLUT
om makroekonomiskt stöd till Republiken Moldavien
EUROPEISKA UNIONENS RÅD HAR BESLUTAT FÖLJANDE
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 308,
med beaktande av kommissionens förslag,[2]
med beaktande av Europaparlamentets yttrande,[3]
efter samråd med Ekonomiska och finansiella kommittén, och
av följande skäl:
2. Myndigheterna i Moldavien arbetar för ekonomisk stabilitet och strukturreformer med stöd av Internationella valutafonden (IMF) genom en treårig åtgärd inom ramen för mekanismen för fattigdomsminskning och ökad tillväxt som godkändes den 5 maj 2006. Därefter godkände fordringsägarna i Parisklubben den 12 maj 2006 en omstrukturering av Moldaviens bilaterala offentliga skulder enligt Houstonvillkoren.
3. I maj 2004 antog de moldaviska myndigheterna ett strategidokumentet för ökad tillväxt och fattigdomsminskning, som innehöll prioriteringarna på medellång sikt för regeringens åtgärder.
4. Moldavein, å ena sidan, och Europeiska gemenskapen och dess medlemsstater, å andra sidan, har undertecknat ett partnerskaps- och samarbetsavtal, som trädde i kraft den 1 juli 1998.
5. Relationerna mellan Moldavien och Europeiska unionen utvecklas inom ramen för den europeiska grannskapspolitiken, som förväntas leda till fördjupad ekonomisk integration. EU och Moldavien har överenskommit om en handlingsplan för den europeiska grannskapspolitiken som innehåller prioriteringar på kort och medellång sikt i relationerna mellan EU och Moldavien och berörda politikområden.
6. Finansieringsbehovet är omfattande i Moldavien beroende på en grav försämring av landets externa situation.
7. De moldaviska myndigheterna har begärt förmånligt finansiellt stöd från de internationella finansinstituten, gemenskapen och andra bilaterala givare. Utöver den finansiering som IMF och Världsbanken tillhandahåller finns det ett avsevärt behov av ytterligare finansiering som måste täckas för att landet skall klara av betalningsbalansen, kunna stärka valutareserven och uppnå de ekonomisk-politiska målen för myndigheternas reformåtgärder.
8. Moldavien är berättigat till mycket fördelaktiga lån och bidrag från Världsbanken och IMF.
9. Under dessa omständigheter bör gemenskapens makroekonomiska stöd till Moldavien ske i form av ett bidrag, som en lämplig åtgärd för att hjälpa landet i dess kritiska läge.
10. För att säkra ett effektivt skydd av gemenskapens ekonomiska intressen knutna till det aktuella makroekonomiska stödet måste man sörja för att Moldavien vidtar lämpliga åtgärder för att förhindra och bekämpa bedrägerier, korruption och andra oegentligheter i samband med detta stöd, samt att kommissionen och revisionsrätten genomför kontroller.
11. Budgetmyndighetens befogenheter påverkas inte av att detta stöd i form av bidrag frigörs.
12. Detta makroekonomiska stöd bör förvaltas av kommissionen i samråd med Ekonomiska och finansiella kommittén.
13. Fördraget innehåller inte några andra befogenheter för att anta detta beslut, än de som anges i artikel 308.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
14. Gemenskapen skall ge Moldavien ett makroekonomiskt stöd i form av ett bidrag på upp till 45 miljoner euro i syfte att stödja Moldaviens betalningsbalans och, på så vis, lindra de ekonomiska påfrestningar genomförandet av regeringens ekonomiska program medför.
15. Gemenskapens ekonomiska stöd skall förvaltas av kommissionen i nära samråd med Ekonomiska och finansiella kommittén och med beaktande av bestämmelserna i de avtal och överenskommelser som ingåtts mellan IMF och Moldavien.
16. Gemenskapens ekonomiska stöd skall vara tillgängligt i två år från och med den första dagen efter att detta beslut träder i kraft. Om omständigheterna så kräver kan emellertid kommissionen, efter samråd med Ekonomiska och finansiella kommittén, besluta att förlänga tillgänglighetsperioden med högst ett år.
Artikel 2
17. Kommissionen är bemyndigad att, efter samråd med Ekonomiska och finansiella kommittén, enas med Moldaviens myndigheter om vilken ekonomisk politik och vilka finansiella villkor som skall knytas till stödet och detta skall formuleras i ett samförståndsavtal och en bidragsöverenskommelse. Villkoren skall vara förenliga med de avtal och överenskommelser som avses i artikel 1.2.
18. Under det faktiska genomförandet av gemenskapsstödet skall kommissionen övervaka att Moldavien har sunda finansiella flöden, administrativa förfaranden samt interna och externa kontrollmekanismer som är relevanta för detta makroekonomiska stöd från gemenskapen.
19. Kommissionen skall regelbundet, i samarbete med Ekonomiska och finansiella kommittén och samordnat med IMF, kontrollera att Moldaviens ekonomiska politik överensstämmer med syftena med detta stöd, samt att överenskommelserna om ekonomisk politik och finansiella villkor följs på tillfredsställande sätt.
Artikel 3
20. Kommissionen skall tillhandahålla Moldavien stödet i tre delutbetalningar.
21. Den första delutbetalningen skall ske efter ett tillfredsställande genomförande av det IMF-stödda ekonomiska programmet inom ramen för mekanismen för fattigdomsminskning och ökad tillväxt och handlingsplanen för den europeiska grannskapspolitiken för EU och Moldavien.
22. Den andra och eventuella ytterligare delutbetalningar skall ske efter ett tillfredsställande genomförande av det IMF-stödda ekonomiska programmet inom ramen för mekanismen för fattigdomsminskning och ökad tillväxt och handlingsplanen för den europeiska grannskapspolitiken för EU och Moldavien, samt andra eventuella åtgärder som överenskommits med kommissionen i enlighet med artikel 2.1, dock tidigast ett kvartal efter den förra delutbetalningen.
23. Medlen skall utbetalas till Moldaviens centralbank. Slutmottagare av medlen är Moldaviens finansministerium.
Artikel 4
Detta stöd skall genomföras i enlighet med budgetförordningen för Europeiska gemenskapernas allmänna budget samt dess genomförandebestämmelser. I synnerhet gäller att det samförståndsavtal och den bidragsöverenskommelse som ingås med Moldaviens myndigheter skall innehålla lämpliga åtgärder som Moldavien skall vidta för att förhindra och bekämpa bedrägerier, korruption och andra oegentligheter i samband med detta stöd. Det skall också innehålla bestämmelser om kontroller som skall utföras av kommissionen, inklusive Europeiska byrån för bedrägeribekämpning (OLAF), med rätt att utföra inspektioner och kontroller på plats samt om revisionsrättens rätt att utföra revision, där så krävs på platsen.
Artikel 5
Kommissionen skall minst en gång om året senast den 31 augusti överlämna en rapport till Europaparlamentet och rådet som skall innehålla en utvärdering av genomförandet av detta beslut under föregående år.
Artikel 6
Detta beslut får verkan samma dag som det offentliggörs i Europeiska unionens officiella tidning .
[pic] | EUROPEISKA GEMENSKAPERNAS KOMMISSION |
Bryssel den 25.10.2006
KOM(2006) 622 slutlig
2006/0198 (ACC)
Förslag till
RÅDETS FÖRORDNING
om handel med vissa stålprodukter mellan Europeiska gemenskapen och Ukraina
(framlagt av kommissionen)
MOTIVERING
BAKGRUND |
110 | Motiv och syfte I Europeiska gemenskapens avtal om partnerskap och samarbete med Ukraina fastställs att handel med vissa stålprodukter skall omfattas av ett avtal mellan parterna. |
120 | Allmän bakgrund Det nuvarande avtalet löper ut den 31 december 2006. Båda parter vill ingå ett nytt avtal för 2007 och följande år, men det nya avtalet kommer inte att träda i kraft den 1 januari 2007. I avvaktan på att avtalet träder i kraft måste därför autonoma åtgärder som fastställer kvoter från och med den 1 januari 2007 vidtas. |
130 | Gällande bestämmelser Rådets beslut 2005/638/EG om ingående av avtalet (EUT L 232, 8.9.2005, s. 42) och rådets förordning (EG) nr 1440/2005 (EUT L 232, 8.9.2005, s. 1) om tillämpningen av detta avtal. |
141 | Förenlighet med Europeiska unionens politik och mål på andra områden Ej tillämpligt. |
SAMRÅD MED BERÖRDA PARTER OCH KONSEKVENSANALYS |
Samråd med berörda parter |
219 | Parterna har konsulterats om ett förslag som hänger samman med detta förslag. Denna förordning innebär en fortsatt tillämpning av ett system som redan tillämpats sedan flera år tillbaka. |
Extern experthjälp |
229 | Någon extern experthjälp har inte behövts. |
230 | Konsekvensanalys Ej tillämpligt. |
RÄTTSLIGA ASPEKTER |
305 | Sammanfattning av den föreslagna åtgärden I denna rådsförordning fastställs kvantitativa begränsningar som skall gälla från och med den 1 januari 2007 tills den nya förordningen träder i kraft. |
310 | Rättslig grund Artikel 133 i fördraget om upprättandet av Europeiska gemenskapen. |
329 | Subsidiaritetsprincipen Förslaget avser ett område där gemenskapen är ensam behörig. Subsidiaritetsprincipen är därför inte tillämplig. |
Proportionalitetsprincipen Förslaget är förenligt med proportionalitetsprincipen av följande skäl: |
331 | Importen av stålprodukter som omfattas av denna förordning är underkastad ett system med kvoter och importtillstånd. Importörer i EU ansöker om det importtillstånd som krävs hos en medlemsstats behöriga myndighet. Den behöriga myndigheten kontrollerar att de handlingar som den sökande lämnat in följer gällande bestämmelser, kontrollerar elektroniskt i en central databas att de kvantiteter som ansökan avser finns tillgängliga och utfärdar därefter importtillståndet. Den praktiska tillämpningen av systemet är så utformad att antalet inblandade parter begränsas till ett minimum. Systemet är följaktligen ganska smidigt, eftersom antalet nivåer är begränsat och det inte kräver kommissionens medverkan. |
332 | Sedan flera år tillbaka har internationella avtal med samma föremål och operativa regler ingåtts. Det faktum att ingen av de berörda parterna har begärt någon ändring kan tolkas som en bekräftelse på att aktörerna och de nationella myndigheterna anser att systemet är förhållandevis lätt att hantera. |
Val av regleringsform |
341 | Föreslagen regleringsform: förordning. |
342 | Övriga regleringsformer skulle vara olämpliga av följande skäl: Kvantitativa begränsningar kan bara fastställas genom en förordning. |
BUDGETKONSEKVENSER |
409 | Förslaget påverkar inte gemenskapens budget. |
1. 2006/0198 (ACC)
Förslag till
RÅDETS FÖRORDNING
om handel med vissa stålprodukter mellan Europeiska gemenskapen och Ukraina
EUROPEISKA UNIONENS RÅD HAR ANTAGIT DENNA FÖRORDNING
med beaktande av fördraget om upprättandet av Europeiska gemenskapen, särskilt artikel 133,
med beaktande av kommissionens förslag, och
av följande skäl:
(1) Enligt artikel 22.1 i avtalet om partnerskap och samarbete mellan Europeiska gemenskaperna och deras medlemsstater, å ena sidan, och Ukraina, å andra sidan[1], skall handel med vissa stålprodukter regleras genom ett särskilt avtal om kvantitativa arrangemang.
(2) Det nuvarande bilaterala avtalet om handel med vissa stålprodukter mellan Europeiska gemenskapen och Ukrainas regering, som undertecknades den 29 juli 2005[2], löper ut den 31 december 2006.
(3) Preliminära diskussioner mellan parterna tyder på att båda har för avsikt att ingå ett nytt avtal för 2007 och följande år.
(4) I avvaktan på att det nya avtalet undertecknas och träder i kraft bör kvantitativa begränsningar fastställas för 2007.
(5) Eftersom omständigheterna idag är desamma som de som rådde när de kvantitativa begränsningarna för 2006 fastställdes, är det lämpligt att behålla de kvantitativa begränsningarna för 2007 på samma nivå som de låg 2006.
(6) Det är nödvändigt att genom så liknande bestämmelser som möjligt sörja för att denna ordning kan administreras inom gemenskapen på ett sådant sätt som underlättar genomförandet av det nya avtalet.
(7) Det är nödvändigt att se till att de berörda produkternas ursprung kontrolleras och att lämpliga metoder för administrativt samarbete införs för detta ändamål.
(8) Produkter som placeras i en frizon eller som importeras enligt förfarandena för tullager, temporär import eller aktiv förädling (suspensionssystemet) bör inte avräknas mot de begränsningar som fastställts för produkterna i fråga.
(9) För en effektiv tillämpning av denna förordning bör det införas ett krav på en EG-importlicens för de berörda produkternas övergång till fri omsättning i gemenskapen.
(10) För att säkerställa att de kvantitativa begränsningarna inte överskrids är det nödvändigt att införa ett förfarande som innebär att de behöriga myndigheterna i medlemsstaterna inte utfärdar importlicenser förrän kommissionen har bekräftat att det fortfarande finns utrymme inom den kvantitativa begränsningen i fråga.
HÄRIGENOM FÖRESKRIVS FÖLJANDE.
Artikel 1
1. Denna förordning skall tillämpas från och med den 1 januari 2007 till och med den 31 december 2007 på import till gemenskapen av stålprodukter enligt förteckningen i bilaga I med ursprung i Ukraina.
2. Stålprodukterna skall klassificeras i de produktgrupper som anges i bilaga I.
3. Klassificeringen av produkterna i bilaga I skall baseras på den kombinerade nomenklatur (KN) som fastställts genom rådets förordning (EEG) nr 2658/87[3].
4. Ursprunget för de produkter som avses i punkt 1 skall bestämmas enligt de bestämmelser som gäller i gemenskapen.
Artikel 2
1. Import till gemenskapen av stålprodukter enligt förteckningen i bilaga I med ursprung i Ukraina skall omfattas av de kvantitativa begränsningar som fastställs i bilaga V. För övergång till fri omsättning i gemenskapen av produkter enligt förteckningen i bilaga I med ursprung i Ukraina skall krävas att det uppvisas ett ursprungscertifikat enligt bilaga II och en importlicens som utfärdats av medlemsstaternas myndigheter i enlighet med artikel 4.
2. För att säkra att de kvantiteter för vilka importlicenser utfärdas inte vid något tillfälle överstiger de sammanlagda kvantitativa begränsningarna för varje produktgrupp skall de behöriga myndigheter som anges i bilaga IV utfärda importlicenser först efter det att kommissionen har bekräftat att det fortfarande finns tillgängliga kvantiteter inom de för leverantörslandet gällande kvantitativa begränsningarna för den stålproduktgrupp som berörs av en eller flera importörers ansökningar till de behöriga myndigheterna.
3. Beviljad import skall avräknas mot de kvantitativa begränsningar som anges i bilaga V. Avsändningen av produkterna skall anses ha ägt rum den dag då de lastades på det transportmedel som användes för exporten.
Artikel 3
1. De kvantitativa begränsningar som anges i bilaga V skall inte gälla för produkter som placeras i en frizon eller ett frilager eller som importeras enligt förfarandena för tullager, temporär import eller aktiv förädling (suspensionssystemet).
2. Om de produkter som avses i punkt 1 senare övergår till fri omsättning, i oförändrat skick eller efter bearbetning eller behandling, skall artikel 2.2 tillämpas och de produkter som övergår till fri omsättning skall avräknas mot den relevanta kvantitativa begränsningen i bilaga V.
Artikel 4
1. Vid tillämpning av artikel 2.2 skall de behöriga myndigheterna i medlemsstaterna – angivna i bilaga IV – innan de utfärdar importlicenser, till kommissionen anmäla de kvantiteter för vilka de har mottagit ansökningar om importlicenser, underbyggda med exportlicenser i original. Kommissionen skall omgående, i den ordning medlemsstaternas anmälningar tas emot (”först till kvarn”-principen), meddela huruvida de begärda kvantiteterna är tillgängliga för import.
2. De ansökningar som omfattas av anmälningarna till kommissionen skall vara giltiga om de i varje enskilt fall klart och tydligt anger exportlandet, det berörda produktnumret, den kvantitet som skall importeras, exportlicensens nummer, kvotåret och den medlemsstat där produkterna avses övergå till fri omsättning.
3. Kommissionen skall, så långt det är möjligt, för myndigheterna bekräfta hela den kvantitet som anges i de anmälda ansökningarna för varje produktgrupp.
4. De behöriga myndigheterna skall så snart de får kännedom om kvantiteter som inte utnyttjats under en importlicens giltighetstid anmäla dessa kvantiteter till kommissionen. Sådana outnyttjade kvantiteter skall automatiskt överföras till de återstående kvantiteterna av gemenskapens sammanlagda kvantitativa begränsning för varje berörd produktgrupp.
5. De anmälningar som avses i punkterna 1–4 skall sändas på elektronisk väg via det integrerade nät som upprättats för detta ändamål, såvida det inte av tvingande tekniska skäl är nödvändigt att tillfälligt använda andra kommunikationssätt.
6. Importlicenserna eller motsvarande dokument skall utfärdas i enlighet med artiklarna 12-16.
7. Medlemsstaternas behöriga myndigheter skall underrätta kommissionen om redan utfärdade importlicenser eller motsvarande dokument upphävs i de fall då de motsvarande exportlicenserna har återkallats eller upphävts av de behöriga myndigheterna i Ukraina. Om kommissionen eller en medlemsstats behöriga myndigheter har underrättats av de behöriga myndigheterna i Ukraina om återkallandet eller upphävandet av en exportlicens efter det att de berörda produkterna har importerats till gemenskapen, skall kvantiteterna i fråga dock avräknas mot den relevanta kvantitativa begränsning som anges i bilaga V.
Artikel 5
1. Om kommissionen har indikationer på att produkter enligt förteckningen i bilaga I med ursprung i Ukraina har omlastats eller omdirigerats eller på annat sätt importerats till gemenskapen på ett sätt som utgör kringgående av de kvantitativa begränsningar som avses i artikel 2 och om den konstaterar att anpassningar måste göras, skall den begära att samråd inleds så att en överenskommelse kan nås om en motsvarande anpassning av de berörda kvantitativa begränsningarna.
2. I avvaktan på resultatet av det samråd som avses i punkt 1 får kommissionen begära att Ukraina vidtar nödvändiga försiktighetsåtgärder för att säkra att de anpassningar av de kvantitativa begränsningarna som parterna kommer överens om vid samrådet kan genomföras.
3. Om gemenskapen och Ukraina inte når en tillfredsställande lösning och om kommissionen konstaterar att klara bevis för kringgående föreligger, skall kommissionen från de kvantitativa begränsningarna dra av en motsvarande kvantitet produkter med ursprung i Ukraina.
Artikel 6
1. En exportlicens – utfärdad av de behöriga myndigheterna i Ukraina – skall krävas för alla sändningar av stålprodukter som omfattas av de kvantitativa begränsningarna i bilaga V, upp till nivån för dessa begränsningar.
2. Originalet av exportlicensen skall uppvisas av importören för att den importlicens som avses i artikel 12 skall kunna utfärdas.
Artikel 7
1. Exportlicensen för produkter som omfattas av kvantitativa begränsningar skall överensstämma med förlagan i bilaga II och skall intyga bland annat att den berörda mängden varor har avräknats mot den kvantitativa begränsning som fastställts för den berörda produktgruppen.
2. Varje exportlicens skall avse endast en av de produktgrupper som anges i bilaga I.
Artikel 8
Export skall avräknas mot de kvantitativa begränsningar som anges i bilaga V och avsändas i den mening som avses i artikel 2.3.
Artikel 9
1. Den exportlicens som avses i artikel 6 får inbegripa kopior, vilka skall vara vederbörligen märkta som sådana. Exportlicensen, ursprungscertifikatet och kopiorna av dessa skall vara avfattade på engelska.
2. Om de dokument som avses i punkt 1 fylls i för hand skall uppgifterna textas med bläck.
3. Exportlicenser eller motsvarande dokument skall ha måtten 210 × 297 mm. Det papper som används skall vara vitt skrivpapper, limbehandlat, fritt från mekanisk massa och med en vikt av minst 25 g/m². Varje del skall ha en tryckt guillocherad bakgrund som gör all förfalskning på mekanisk eller kemisk väg synlig.
4. Endast originalet skall godtas av gemenskapens behöriga myndigheter såsom giltigt för import i enlighet med bestämmelserna i denna förordning.
5. Varje exportlicens eller motsvarande dokument skall genom tryck eller på annat sätt förses med ett standardiserat löpnummer som möjliggör identifiering av dokumentet.
6. Löpnumret skall vara sammansatt på följande sätt:
– Två bokstäver som anger exportlandet enligt följande: UA = Ukraina
– Två bokstäver som anger avsedd bestämmelsemedlemsstat enligt följande:
BE = Belgien
BG = Bulgarien
CZ = Tjeckien
DK = Danmark
DE = Tyskland
EE = Estland
EL = Grekland
ES = Spanien
FR = Frankrike
IE = Irland
IT = Italien
CY = Cypern
LV = Lettland
LT = Litauen
LU = Luxemburg
HU = Ungern
MT = Malta
NL = Nederländerna
AT = Österrike
PL = Polen
PT = Portugal
RO = Rumänien
SI = Slovenien
SK = Slovakien
FI = Finland
SE = Sverige
UK = Förenade kungariket
– Ett ensiffrigt nummer som anger kvotåret i fråga och som utgörs av den sista siffran i det årtalet, t.ex. ”4” för 2004.
– Ett tvåsiffrigt nummer som anger det utfärdande kontoret i exportlandet.
– Ett femsiffrigt nummer som löper i följd från 00 001 till 99 999 och som tilldelas bestämmelsemedlemsstaten i fråga.
Artikel 10
Exportlicenser får utfärdas efter avsändandet av de produkter de avser. I sådana fall skall de vara försedda med påskriften ”issued retrospectively”.
Artikel 11
Om en exportlicens stulits, förlorats eller förstörts, får exportören hos den behöriga myndighet som utfärdat dokumentet ansöka om ett duplikat, som skall utfärdas på grundval av de exporthandlingar som exportören förfogar över.
Ett sålunda utfärdat duplikat av en licens skall ha påskriften ”duplicate”. Det skall ha samma datum som den ursprungliga licensen.
Artikel 12
1. Om kommissionen, i enlighet med artikel 4, har bekräftat att den begärda mängden finns tillgänglig inom den kvantitativa begränsningen i fråga, skall medlemsstaternas behöriga myndigheter utfärda en importlicens inom fem arbetsdagar efter det att importören har uppvisat motsvarande exportlicens i original. Exportlicensen måste uppvisas senast den 31 mars året efter det år då de varor som omfattas av licensen avsändes. Importlicenser skall utfärdas av de behöriga myndigheterna i vilken som helst av medlemsstaterna, oavsett vilken medlemsstat som anges på exportlicensen, om kommissionen i enlighet med artikel 4 har bekräftat att den begärda mängden finns tillgänglig inom den kvantitativa begränsningen i fråga.
2. Importlicenserna skall vara giltiga i fyra månader från och med den dag de utfärdades. En medlemsstats behöriga myndigheter får, efter en väl motiverad begäran från importören, förlänga giltighetstiden med ytterligare högst fyra månader.
3. Importlicenserna skall utformas enligt förlagan i bilaga III och de skall vara giltiga i hela gemenskapens tullområde.
4. Den deklaration eller ansökan som importören lämnar in för att få importlicensen skall innehålla följande uppgifter:
a) Exportörens fullständiga namn och adress.
b) Importörens fullständiga namn och adress.
c) En exakt beskrivning av varorna och numret eller numren i Taric.
d) Varornas ursprungsland.
e) Avsändningsland.
f) Korrekt produktgrupp för och kvantiteten av de produkter det är fråga om.
g) Nettovikt för varje Taric-nummer.
h) Produkternas värde cif vid gemenskapens gräns för varje Taric-nummer.
i) Uppgift om huruvida de berörda produkterna är andrasorteringsprodukter eller av bristfällig kvalitet.
j) I tillämpliga fall, betalnings- och leveransdatum och en kopia av konossementet och av köpeavtalet.
k) Exportlicensens datum och nummer.
l) Interna koder för administrativa ändamål.
m) Datum samt importörens underskrift.
5. Importörerna skall inte vara skyldiga att importera hela den kvantitet som omfattas av en importlicens i en och samma sändning.
Artikel 13
Giltigheten av importlicenser som utfärdats av medlemsstaternas myndigheter skall vara beroende av giltigheten av och de kvantiteter som anges i de exportlicenser som utfärdats av de behöriga myndigheterna i Ukraina och som legat till grund för utfärdandet av importlicenserna.
Artikel 14
Importlicenser eller motsvarande dokument skall utfärdas av medlemsstaternas behöriga myndigheter i enlighet med artikel 2.2 till varje importör i gemenskapen utan åtskillnad, oavsett var i gemenskapen denne är etablerad, och utan att det påverkar tillämpningen av övriga krav som ställs enligt gällande bestämmelser.
Artikel 15
1. Om kommissionen konstaterar att de sammanlagda kvantiteter som omfattas av exportlicenser som utfärdats av Ukraina för en viss produktgrupp överstiger den kvantitativa begränsning som fastställts för den produktgruppen, skall de behöriga myndigheter som utfärdar licenser i medlemsstaterna genast underrättas så att inga ytterligare importlicenser utfärdas. I sådana fall skall kommissionen genast inleda samråd.
2. En medlemsstats behöriga myndigheter skall neka att utfärda importlicenser för produkter med ursprung i Ukraina som inte omfattas av exportlicenser utfärdade i enlighet med bestämmelserna i artiklarna 6–11.
Artikel 16
1. De formulär som medlemsstaternas behöriga myndigheter skall använda för att utfärda de importlicenser som avses i artikel 12 skall överensstämma med förlagan till importlicens i bilaga III.
2. Importlicensformulär och utdrag ur dessa skall upprättas i två exemplar: det ena skall vara märkt ”Innehavarens exemplar" och ha nummer 1 och utfärdas till den som ansöker om importlicensen, det andra skall vara märkt ”Utfärdande myndighets exemplar” och ha nummer 2 och behållas av den myndighet som utfärdar licensen. De behöriga myndigheterna får för administrativa ändamål lägga till ytterligare kopior av formulär nr 2.
3. Formulären skall tryckas på vitt skrivpapper, fritt från mekanisk massa och med en vikt på mellan 55 och 65 g/m². De skall ha måtten 210 × 297 mm. Radavståndet skall vara 4,24 mm (en sjättedels tum). Formulärens utformning skall noga följas. Båda sidor av exemplar nr 1, som utgör själva licensen, skall dessutom ha en röd, tryckt guillocherad bakgrund som gör all förfalskning på mekanisk eller kemisk väg synlig.
4. Medlemsstaterna skall ansvara för tryckningen av formulären. Formulären får också tryckas av tryckerier som godkänts av den medlemsstat där de är etablerade. I det senare fallet skall det på varje formulär finnas en hänvisning till detta godkännande. Varje formulär skall vara försett med tryckeriets namn och adress eller ett märke som gör det möjligt att identifiera tryckeriet.
5. Vid utfärdandet skall importlicenserna eller utdragen av dessa ges ett utfärdandenummer som fastställs av de behöriga myndigheterna i medlemsstaten. Importlicensens nummer skall anmälas till kommissionen på elektronisk väg inom det integrerade nät som upprättats enligt artikel 4.
6. Licenser och utdrag skall fyllas i på det officiella språket eller ett av de officiella språken i den utfärdande medlemsstaten.
7. I fält 10 skall de behöriga myndigheterna ange tillämplig stålproduktgrupp.
8. De myndigheter som utfärdar licenserna och handhar avräkningarna skall sätta sin stämpel på dokumenten. Den utfärdande myndighetens stämpel får dock ersättas med ett relieftryck kombinerat med bokstäver eller siffror som anbringas på licensen genom perforering eller tryckning. De utfärdande myndigheterna skall vid registrering av den tilldelade kvantiteten använda en metod som omöjliggör förfalskning, så att det inte är möjligt att lägga till siffror eller hänvisningar.
9. På baksidan av exemplar nr 1 och nr 2 skall det finnas ett fält i vilket kvantiteter kan anges, antingen av tullmyndigheterna när importformaliteterna fullgörs eller av de behöriga förvaltningsmyndigheterna när ett utdrag utfärdas. Om utrymmet för avräkningar på licensen eller utdraget av denna är otillräckligt, får de behöriga myndigheterna använda tilläggsblad med fält som motsvarar fälten på baksidan av exemplar nr 1 och 2 av licensen eller utdraget. De myndigheter som svarar för avräkningen skall placera sin stämpel på sådant sätt att ena halvan är på licensen eller utdraget av denna och andra halvan på tilläggsbladet. Om det finns mer än ett tilläggsblad skall ytterligare en stämpel placeras på samma sätt tvärs över varje blad och det föregående bladet.
10. Importlicenser och utdrag som utfärdats, uppgifter som fyllts i och påskrifter som gjorts av myndigheterna i en medlemsstat skall ha samma rättsliga verkan i var och en av de andra medlemsstaterna som handlingar som utfärdats, uppgifter som fyllts i och påskrifter som gjorts av myndigheterna i dessa medlemsstater.
11. Medlemsstaternas behöriga myndigheter får när det är nödvändigt kräva att innehållet i licenserna eller utdragen översätts till det officiella språket eller ett av de officiella språken i den berörda medlemsstaten.
Artikel 17
Denna förordning träder i kraft samma dag som den offentliggörs i Europeiska unionens officiella tidning.
Denna förordning är till alla delar bindande och direkt tillämplig i alla medlemsstater.
Sammanfattande information om statligt stöd som beviljats enligt kommissionens förordning (EG) nr 1/2004 av den 23 december 2003 om tillämpningen av artiklarna 87 och 88 i EG-fördraget på statligt stöd till små och medelstora företag som är verksamma inom produktion, bearbetning och saluföring av jordbruksprodukter
(2006/C 2/03)
Stöd nr : XA 37/04
Medlemsstat : Italien
Region : Venetien
Namnet på stödordningen eller namnet på det företag som tar emot det enskilda stödet : Stöd till investeringar i samband med bearbetning och saluföring av jordbruksprodukter
Rättslig grund : Legge Regionale 12 Dicembre 2003, n. 40 Titolo VI Capo III artt. 24, 25, 26, 27 e 28 %quot%Nuove norme per gli interventi in agricoltura%quot% e successive modifiche ed integrazioni. Il testo coordinato della legge è pubblicato sul Bollettino Ufficiale della Regione del Veneto n. 40 del 13.4.2004
Stödordningens beräknade utgifter per år eller totalt belopp som beviljats företaget som enskilt stöd : Det årliga stödbeloppet fastställs genom den finansieringslag (Legge finanziaria) som varje år antas av regionrådet (Consiglio regionale). Man kan utgå från att ett belopp på 2000000 EUR kommer att ställas till förfogande varje år. Denna siffra är endast vägledande
Högsta tillåtna stödnivå : 40 % av de stödberättigande kostnaderna
Datum för genomförande : 1 september 2004
Stödordningens eller det enskilda stödets varaktighet : 30 juni 2007
Stödets syfte 1) Sysselsättning
2) Sektorsutveckling
3) Miljöskydd
Artikel 7 i förordning 1/2004 av den 23 december 2003
Stödberättigande kostnader: miljöskydd och avlägsnande av förorenande biprodukter från bearbetningsverksamhet; ombyggnation, modernisering och rationalisering av anläggningar för lagring, hantering, beredning, bearbetning och saluföring av jordbruksprodukter; förvärv av anläggningar, maskiner och redskap för att modernisera arbetsprocesser och produkter; inköp av datautrustning och –program till styrning av produktionsprocessen; förbättring av arbetsmiljön och anpassning till säkerhetsföreskrifter; inköp av företag, anläggningar och tillhörande utrustning, med undantag av jordarealer; förbättring av de hygieniska förhållandena på företagen; anpassning av företagen i syfte att införa system för kontroll och styrning av produkternas kvalitet och spårbarhet
Sektor(er) av ekonomin som berörs : Stödordningen omfattar bearbetning och/eller saluföring av de jordbruksprodukter som ingår i bilaga I till fördraget och berör samtliga produktionssektorer
Den beviljande myndighetens namn och adress Regione Veneto
Giunta Regionale
Direzione politiche agroalimentari e per le imprese
Via Torino 110, I-30174 Mestre (VE)
Webbplats : http://www.consiglioveneto.it/leggi/2003/03lr0040.html
Stöd nr : XA 40/05
Medlemsstat : Spanien
Region : Kastilien-León
Namnet på stödordningen : Stöd för att främja bevattnade grödor i den självstyrande regionen Kastilien-León
Rättslig grund :
Orden AYG …/2005, de … junio, de la Consejería de Agricultura y Ganadería, por la que se establece un plan de dinamización de los cultivos de regadío en la Comunidad Autónoma de Castilla y León.
Denna stödordning beviljas enligt det undantag som fastställs genom kommissionens förordning (EG) 1/2004 av den 23 december 2003 och följer bestämmelserna i artiklarna 7, 13 och 14 i denna förordning vad gäller investeringar i bearbetning och saluföring, stöd för att uppmuntra produktion och saluföring av kvalitetsprodukter från jordbruket och tillhandahållande av tekniskt stöd inom jordbrukssektorn
Stödordningens beräknade utgifter per år : Stödet för 2005 beräknas till 3500000 EUR
Högsta stödnivå - Artikel 7 i förordning 1/2004. Den högsta stödnivån kommer att vara 50 % av de stödberättigande investeringarna.
- Artikel 13 i förordning 1/2004. Det högsta totala stödet per stödmottagare är 100000 EUR för en period på tre år.
- Artikel 14 i förordning 1/2004. Stödet per stödmottagare får inte överskrida det största av följande belopp: 100000 EUR under tre år eller 50 % av de stödberättigande kostnaderna
Datum för genomförande : Stödordningen träder i kraft i juni 2005
Stödordningens eller det enskilda stödets varaktighet : Stödordningen skall vara giltig fram till och med den 31 december 2006
Stödets syfte Allmänt syfte
Att främja utvecklingen av bevattnade grödor i den självstyrande regionen Kastilien-León.
Sekundärt syfte
- Stimulera investeringar i bearbetning och saluföring av bevattnade grödor i de områden i regionen som är särskilt lämpliga för odling av grödorna i fråga. - Främja uppmuntra produktion och saluföring av kvalitetsprodukter.
- Tillhandahålla tekniskt stöd inom sektorn för bevattnade grödor genom genomförande av revisioner, förvaltningsanalyser, genomförbarhetsanalyser, investeringsanalyser och marknadsstudier.
- Berörda artiklar
- Stödordningen följer bestämmelserna i följande artiklar i förordning 1/2004:
- Artikel 7 om investeringar i bearbetning och saluföring.
- Artikel 13 om stöd för att uppmuntra produktion och saluföring av kvalitetsprodukter från jordbruket.
- Artikel 14 om tillhandahållande av tekniskt stöd inom jordbrukssektorn.
- Även artiklarna 17–20 i kapitel 3 i förordningen – allmänna bestämmelser och slutbestämmelser – har beaktats.
- Stödberättigande kostnader
- Artikel 7 i förordning 1/2004. Investeringar i bearbetning och saluföring av bevattnade grödor
- Kostnader för uppförande och förvärv av fast egendom, dock inte förvärv av mark.
- Kostnader för förvärv av nya maskiner och ny utrustning, inklusive datorprogram upp till produktens marknadsvärde.
- Allmänna kostnader, exempelvis för arvoden till arkitekter, ingenjörer, konsulter, värderingsmän och revisorer samt kostnader för genomförbarhetsstudier och förvärv av patent och licenser.
- Artikel 13 i förordning 1/2004. Stöd för att uppmuntra produktion och saluföring av kvalitetsprodukter från jordbruket.
- Kostnader som hänför sig till införandet av system som skall främja och förbättra produktkvaliteten. Till dessa kostnader kan man också lägga följande kostnader: kostnader för förstudier för ansökningar om godkännande av kvalitetsmärkning; kostnader som hänför sig till införandet av kvalitetssäkringssystemet; kostnader för externa konsulter; kostnader för certifiering; kostnader för utbildning av personalen om tillämpningen av dessa system.
- Artikel 14 i förordning 1/2004. Tillhandahållande av tekniskt stöd inom jordbrukssektorn.
- Kostnader som hänför sig till genomförande av revisioner, förvaltningsanalyser, genomförbarhetsanalyser, investeringsanalyser och marknadsstudier
Berörd sektor : Jordbrukssektorn i allmänhet
Den beviljande myndighetens namn och adress :
Stödet skall beviljas av Kastilien-Leóns regering, och administreras av Jordbruks- och boskapsministeriets generaldirektorat för industrialisering och modernisering av jordbruket.
C/ Rigoberto Cortejoso, 14 – E-47014-Valladolid
Webbplats : Stödordningens fullständiga text offentliggörs på Kastilien-Leóns regerings webbplats http://www.jcyl.es/agrocomercializacion
Övriga upplysningar : Förvaltningen av stödet skall ske enligt förordningen och måste uppfylla artikel 18 i förordningen vad gäller kumulering
Stöd nr : XA 55/05
Medlemsstat : Polen
Region : Provinsen Opolskie (NTS – 2.16)
Stödsystemets titel eller namn på det företag som erhåller individuellt stöd : Przedsiębiorstwo Produkcyjno-Handlowe %quot%Ferma-Pol%quot% Sp. z o. o. w Zalesiu, PL-46-146 Domaszowice (individuellt stöd)
Rättslig grund : Ustawa z dnia 27 kwietnia 2001 r. Prawo ochrony środowiska (Dz.U. nr 62, poz. 627, z późn. zm.) — art. 405 oraz art. 411 ust. 10
Stödordningens beräknade utgifter per år inom ramen för stödsystemet, eller sammanlagt individuellt stöd som tilldelats företaget : Stödet tilldelas i form av ett mjukt lån på 500000 PLN (nominellt värde). Lånet betalas ut till januari 2006, och återbetalas från januari 2006 till november 2010. Lånets bruttovärde uppgår till 42770,54 PLN.
Högsta stödnivå : Bruttostödnivån är 6,66 %
Genomförandedatum : Efter godkännande i form av en anmälan tillsammans med ett identifieringsnummer som visar att kommissionen har erhållit denna sammanfattande information om det tilldelade individuella stödet
Stödordningens eller det enskilda stödets varaktighet : Ungefär från juli 2005 till november 2010
Stödets syfte :
Det individuella stödet betalas ut för investeringar i ett centrum för djuruppfödning i syfte att upprätthålla skyddsnivån för miljön och förbättra de hygieniska förhållandena och djurens välbefinnande. Investeringen kommer att användas för att ta bort farligt takmaterial som innehåller asbest och ersätta det med ett asbestfritt tak.
Denna insats krävs främst på grund av ett beslut av byggnadsinspektionen i distriktet Namysłowski av den 2 juli 2004 i vilket %quot%FERMA-POL%quot% i Zalesie uppmanades att avlägsna alla asbesthaltiga material från sina anläggningar. I beslutet hävdades det att skador på eternitskivor kan leda till att asbestfibrer kommer ut i luften och därmed utgöra ett hot mot människors hälsa och miljön, inbegripet för tamdjur.
Exponering för asbest medför risk för sjukdomar i luftvägarna, t.ex. asbestos, lungcancer, skador i lungsäckarna osv. Detta har belagts genom experiment som utfördes på 1970-talet. 1977 sammanställde Europeiska unionens sakkunniga en rapport om de risker för folkhälsan som uppstår genom miljöexponering för asbestdamm, och bekräftade ämnets patogena effekter.
Investeringen omfattas även av det program för att avskaffa asbest och produkter som innehåller asbest i Polen, som antogs av polska ministerrådet den 14 maj 2002, och som bland annat syftar till att befria Polen från asbest och asbesthaltiga produkter som har använts i många år.
Stödet kommer att tilldelas i enlighet med artikel 4 i förordning (EG) nr 1/2004 för investering i en anläggning för djuruppfödning. De stödberättigande kostnaderna omfattar investeringskostnader för att förbättra anläggningen
Berörd(a) sektor(er) : Stödet betalas ut till företag som bedriver jordbruksverksamhet inom sektorn djuruppfödning
Den beviljande myndighetens namn och adress : Stödet kommer att tilldelas av nationella fonden för miljöskydd och vattenhushållning, ul. Konstruktorska 3A, PL-02-673 Warszawa, via Bank Ochrony Środowiska S.A. (Banken för miljöskydd), Al. Jana Pawła II 12, PL-00-950 Warszawa
Webbplats : http://www.bosbank.pl/i.php?i=421
Övriga upplysningar - Bruttostödet (bruttostödnivån) har beräknats i enlighet med definitionen i artikel 2.5 i kommissionens förordning (EG) nr 1/2004 av den 23 december 2003 om tillämpningen av artiklarna 87 och 88 i EG-fördraget på statligt stöd till små och medelstora företag som är verksamma inom produktion, bearbetning och saluföring av jordbruksprodukter. Det utgör därför en procentandel av de stödberättigande kostnaderna.
- Bruttostödsekvivalenten för det mjuka lånet har beräknats i enlighet med den metod som avses i punkt 3 i bilaga I till Riktlinjer för statligt stöd för regionala ändamål (EGT C 74, 10.3.1998, s. 9), men med en skillnad: inkomstskatt har inte tagits med i beräkningen. Bruttostödsekvivalenten uppgår till 42770,54 PLN.
- De stödberättigande kostnaderna uppgår till 642183,67 PLN.
- Bruttostöd = 42770,54 PLN/642183,67 PLN = 6,66 %
Stödnummer : XA 59/05
Medlemsstat : Förenade kungariket
Region : England
Stödordningens namn, eller namnet på det företaget som får enskilt stöd : Jordbruksprogrammet 2005–06 för England (Farming Activities Programme (England) 2005–06)
Rättslig grund : Det finns ingen särskild lagstiftning för stödordningen i fråga. Avsnitt 1 i jordbrukslagen från 1986 (Agriculture Act, section 1) är den rättsliga grunden för regeringens rådgivning i jordbruksfrågor
Årliga utgifter under stödordningen : 1000000 GBP
Högsta stödnivå : Stödnivån är 100 %
Stödordningen gäller från och med : Det första mötet kommer att äga rum tidigast den 12 september 2005
Stödordningens eller det enskilda stödets varaktighet : Stödordningen kommer hela tiden att vara öppen för nya deltagare. Verksamhet inom ramen för stödordningen kommer att pågå under perioden 12 september 2005– 31 mars 2006. Programmet avslutas den 31 mars 2005
Stödets syfte :
Utveckling av en viss sektor. Programmet inriktas på yrkesverksamma jordbrukare. Syftet är att med hjälp av konferenser, studiecirklar och seminarier sätta in jordbrukare i aktuella frågor som kan påverka deras företag, t.ex. nyheterna i den gemensamma jordbrukspolitiken, jordbruk i känsliga avrinningsområden och de nya stödordningarna för miljöhänsyn (Environmental Stewardship Schemes). Detta kommer att höja kompetensen inom sektorn.
Stöd kommer att beviljas i enlighet med artikel 14 i förordning 1/2004, och berättigande kostnader är kostnader för arrangemang av utbildningsprogram
Berörda sektorer : Stödordningen gäller företag som framställer någon form av jordbruksprodukter
Den beviljande myndighetens namn och adress Department for Environment, Food %amp% Rural Affairs
Farm Advice Unit
Rural Development Service
Area 4A, Ergon House
Horseferry Road
London
SW1P 2JR
United Kingdom
Webbplats : www.defra.gov.uk/farm/state-aid/setup/exist-exempt.htm. Klicka på Farming Activities Programme (England) 2005–06, eller gå direkt till http://defraweb/farm/state-aid/setup/schemes/farmingactivities-0506.pdf
Stöd nr: : XA 60/05
Medlemsstat : Italien
Region : Sardinien
Stödordningens namn : Lag nr 1329/65 (%quot%Sabatini-lagen%quot%): stöd för inköp eller leasing av nya maskiner och ny utrustning inom jordbruket
Rättslig grund :
Legge 28 novembre 1965 n. 1329.
Legge regionale 29 novembre 2002 n. 22.
Deliberazione della Giunta Regionale n. 27/7 del 21.6.2005 relativa alle Direttive di attuazione dei benefici di cui alla Legge 1329/65.
Decreto dell'Assessore dell'Agricoltura n. 801/2005 del 4 agosto 2005.
Stödordningens beräknade utgifter per år : 5472000 EUR
Högsta tillåtna stödnivå :
Räntebidrag som uppgår till nettoskillnaden mellan den europeiska referensräntan och den ränta som fastställs för bidraget den dag som det beviljas.
För företag i mindre gynnade områden (artiklarna 18-20 i förordning 1257/1999) får bruttonivån uppgå till högst 50 % av de stödberättigande kostnaderna.
För företag i övriga områden får denna bruttonivå uppgå till högst 40 % av de stödberättigande kostnaderna.
För unga jordbrukare, inom fem år efter den första etableringen, får stödnivån i mindre gynnade områden uppgå till högst 60 % av de stödberättigande kostnaderna; i övriga områden är den övre gränsen 50 %
Genomförandeperiod : Från och med meddelandet om stödet
Stödordningens varaktighet : 31.12.2006
Stödets syfte - lägre produktionskostnader,
- bättre eller omlagd produktion,
- högre kvalitet,
- bevarad eller bättre miljö, bättre hygien och djurskydd,
- diversifiering av jordbruksverksamheten,
Stödet beviljas i enlighet med artikel 4 i förordning (EG) nr 1/2004 av den 23 december 2003, offentliggjord i EUT L den 3 januari 2004
Berörd(a) sektorer : Små och medelstora företag inom jordbruksproduktionen
Den beviljande myndighetens namn och adress Regione Autonoma della Sardegna
Assessorato dell'Agricoltura e Riforma Agro-Pastorale
Via Mario Siddi n. 4, I-09126 Cagliari
Webbplats : www.regione.sardegna.it
Stödnummer : XA 61/05
Medlemsstat : Förenade kungariket
Region : England
Stödordningens namn, eller namnet på det företag som får enskilt stöd : Rådgivning till jordbruksföretag – vilka möjligheter har du? (Farm Business Advice Service – Knowing Your Options)
Rättslig grund : Det finns ingen särskild lagstiftning för tjänsten i fråga. Avsnitt 1 i jordbrukslagen från 1986 (Agriculture Act, section 1) är den rättsliga grunden för regeringens rådgivning i jordbruksfrågor
Utgifter för stödordningen 2005/06: 3500000 GBP
2006/07: 4500000 GBP
Högsta stödnivå : Stödnivån är 100 %
Stödordningen gäller från och med : 26 september 2005
Stödordningens eller det enskilda stödets varaktighet : Stödordningen löper ut den 31 mars 2007. Stöd kommer att betalas ut till och med den 30 april 2007
Stödets syfte : Utveckling av en viss sektor. Syftet med tjänsten är att ge råd och utbildning som kan hjälpa jordbrukare att förstå hur det samlade gårdsstödet påverkar deras verksamhet. Tjänsten ska uppmuntra jordbrukare att överväga omorganisering och diversifiering av verksamheten, samarbete samt alternativa försörjningsmöjligheter om jordbruksverksamheten avvecklas. Berättigande kostnader är sålunda konsultarvoden och utbildningskostnader för jordbrukare och jordbruksanställda enligt artikel 14 i förordning (EG) nr 1/2004
Berörda sektorer : Stödordningen gäller alla företag som framställer jordbruksprodukter och är registrerade för det samlade gårdsstödet i England. Rådgivningen kan gälla produktionen, men även diversifiering till bearbetning och försäljning. Alla undersektorer omfattas
Den beviljande myndighetens namn och adress Department for Environment, Food and Rural Affairs:
Rural Development Service
Ergon House
Horseferry Road
London
SW1P 2AL
United Kingdom
Webbplats : www.defra.gov.uk/farm/state-aid/setup/exist-exempt.htm. Klicka på Farm Business Advice Service – Knowing Your Options, eller gå direkt till www.defra.gov.uk/farm/state-aid/setup/schemes/farmbusinessadvice.pdf
Övrig information :
Den nya tjänsten kommer att starta den 26 september 2005. Den ska erbjuda jordbruksföretag gratis rådgivning för att hjälpa dem att se vilka möjligheter som det samlade gårdsstödet – i kraft sedan den 1 januari 2005 – erbjuder. Tjänsten ersätter den tredagarstjänst som avslutades den 31 mars 2005 (Farm Business Advice Service, stödnummer XA 7/04).
Rent praktiskt kommer tjänsten att tillhandahållas över hela England av tre företag som har valts ut efter upphandling i enlighet med artikel 14.5 i förordning (EG) nr 1/2004
Stöd nr : XA 62/05
Medlemsstat : Nederländerna
Region : Provinserna Limburg, Noord-Brabant, Utrecht, Gelderland och Overijssel
Stödordningens namn Limburg:
Algemene subsidieverordening 2004; Subsidieregels Project Verplaatsing Intensieve Veehouderijen Noord- en Midden-Limburg; Beleidsregels Project Verplaatsing Intensieve Veehouderijen Noord- en Midden-Limburg
Noord-Brabant:
Verordening subsidies kwaliteits- en structuurverbetering Landelijk Gebied provincie Noord-Brabant 2001; Subsidieregeling Verplaatsingskosten Veehouderij 2005
Utrecht:
Subsidieverordening verplaatsing intensieve veehouderij provincie Utrecht 2005
Gelderland:
Subsidieregeling Verplaatsing intensieve veehouderijen Gelderland
Overijssel:
Uitvoeringsbesluit Subsidies Overijssel; Beleidsregel Verplaatsing intensieve veehouderijen Overijssel 2005
Rättslig grund : Artikel 105 juncto artikel 145 Provinciewet, alsmede artikel 158 Provinciewet
| 2005 | 2006 | 2007 | 2008-2012 | Totalt |
Limburg | 0 | 0,225 | 3,415 | 3,96 | 7,7 |
Noord-Brabant | 12,5 | 13 | 13 | 2 | 40,5 |
Utrecht | 0 | 0 | 0 | 1,6 | 1,6 |
Gelderland | 1 | 1 | 3 | 8 | 13 |
Overijssel | 0 | 1,17 | 0 | 5,73 | 6,9 |
Ministerie van LNV | 1,5 | 18,23 | 2,25 | 71,22 | 93,2 |
Preliminära årliga utgifter enligt bestämmelserna, i miljoner EUR Högsta stödnivå 1. 100 % av priset på de anläggningsbyggnader (grundat på taxeringsvärdet) där den intensiva djuruppfödning som skall utlokaliseras äger rum. Taxeringsvärdet relateras till de utgifter som behövs för att inrätta eller förvärva en motsvarande produktionskapacitet med samma tekniska och funktionella livslängd.
2. 25 EUR per kvadratmeter markyta i den rivna anläggningsbyggnaden. Detta avser en kompensation för rivningskostnader för de anläggningsbyggnader som avses i punkt 1.
3. 100 % av priset för den mark (grundat på taxeringsvärdet) på vilken de anläggningsbyggnader står i vilka intensiv djuruppfödning genomfördes. Taxeringsvärdet relateras till markvärdet efter utlokalisering av den intensiva djuruppfödningen och rivning av anläggningsbyggnaderna. Detta motsvarar odlingsmarkens värde.
4. De faktiska kostnaderna för rådgivning, planering och undersökning i samband med nyetableringen, med ett tak på 1000 EUR per utlokaliserad NGE, men maximalt 100000 EUR sammanlagt. NGE (Nederlandse Grootte Eenheid – nederländsk enhet för beståndsstorlek) är en enhet som utgående från antalet djur per art och antalet hektar visar den ekonomiska omfattningen av ett jordbruksföretag eller en enskild produktionsanläggning inom företaget, så som det hanteras av det ekonomiska jordbruksinstitutet (Landbouw Economisch Instituut).
5. 25 EUR per kvadratmeter markyta för icke-användbara anläggningsbyggnader på platsen för nyetableringen som rivits av denna anledning. Detta utgör en kompensation för rivningskostnaderna
Datum för genomförande : Genomförandet inleds efter det offentliggörande i Europeiska unionens officiella tidning som avses i artikel 19 första stycket i kommissionens förordning (EG) nr 1/2004
Varaktighet : Från september 2005 till och med september 2012
Stödets syfte : Utlokalisering – i allmänhetens intresse – av anläggningsbyggnader för intensiv djuruppfödning. Stödet avser utlokalisering av intensiva djurhållningsföretag med goda ekonomiska förutsättningar (små och medelstora företag) som är belägna i extensifieringsområden. Extensifieringsområden är geografiskt avgränsade delar av de omstruktureringsområden som avses i Reconstructiewet, där bosättning och natur prioriteras och där utvidgning, återetablering och nyetablering av intensiv djurhållning inte är möjlig.
Berörd(a) sektor(er): :
Stödet är avsett för intensiva djuruppfödningsföretag (små och medelstora företag) i extensifieringsområden.
Stödet tilldelas inom ramen för bestämmelserna i artikel 6 första och andra stycket i kommissionens förordning (EG) nr 1/2004.
Den beviljande myndighetens namn och adress: Provincie Limburg
Limburglaan 10
Postbus 5700
6202 MA Maastricht
Nederland
Provincie Noord-Brabant
Brabantlaan 1
Postbus 90151
5200 MC 's-Hertogenbosch
Nederland
Provincie Utrecht
Pythagoraslaan 101
Postbus 80300
3508 TH Utrecht
Nederland
Provincie Gelderland
Markt 11
Postbus 9090
6800 GX Arnhem
Nederland
Provincie Overijssel
Luttenbergstraat 2
Postbus 10078
8000 GB Zwolle
Nederland
Webbplats :
www.limburg.nl
www.brabant.nl
www.provincie-utrecht.nl
www.gelderland.nl
www.overijssel.nl
Stöd nr : XA 64/05
Medlemsstat : Spanien
Region : Murcia
Benämning på stödordningen eller namn på det företag som mottar ett individuellt stöd : Stöd under 2005 till företag som genomför projekt som syftar till ökad användning av förnybar energi
Rättslig grund : Orden de 28 de julio de 2005, de la Consejería de Industria y Medio Ambiente, de modificación de la Orden de 20 de enero de 2005 de la Consejería de Economía, Industria e Innovación, publicada en el BORM no 23 de 29 de enero de 2005, por la que se regulan las bases y la convocatoria de ayudas a empresas y a familias e instituciones sin fines de lucro, con destino a la ejecución y explotación de proyectos de instalaciones de aprovechamiento de recursos energéticos renovables, para el ejercicio 2005
Planerade årliga utgifter inom stödordningen eller totalt belopp för individuellt stöd som beviljats företaget : För företag: 400000 EUR
Högsta stödnivå : 40 % brutto av de totala stödberättigande kostnaderna
Genomförandetid : Från och med den dag då stödordningen offentliggörs i regionen Murcias officiella tidning
Varaktighet för stödordningen eller det individuella stödet : Till och med december 2005
Syfte - Under 2005 kan små och medelstora företag i regionen Murcia få stöd för projekt som syftar till ökad användning av förnybar energi.
- Under 2005 kan även små och medelstora företag i regionen Murcia som är verksamma inom produktion, bearbetning och saluföring av jordbruksprodukter få stöd för ökad användning av förnybar energi. Det ursprungliga beslutet om den här typen av stöd fattades genom det ovan nämnda dekretet av den 20 januari 2005 (Orden de 20 de enero de 2005 de la Consejería de Economía, Industria e Innovación) som offentliggjordes i regionen Murcias officiella tidning nr 23 av den 29 januari 2005 (i enlighet med förordning 70/2001).
- Stöden beviljas i enlighet med artikel 4 i kommissionens förordning (EG) nr 1/2004, och de stödberättigande kostnaderna är följande:
1. Kostnader som avser fasta tillgångar (uppförande av byggnader; utrustning; montering och installation) som är nödvändiga för att nå de uppsatta målen.
2. Följande kostnader är inte stödberättigande:
a) Moms på köp av varor eller tjänster, andra typer av skatter.
b) IT-utrustning som inte uttryckligen används för de ändamål som anges i ansökan.
c) Investeringar i begagnad utrustning.
d) Förvärv eller arrende av mark.
e) Projekteringskostnader.
f) Kostnader som inte specificeras på ett entydigt sätt eller som inte direkt avser användning av förnybar energi.
g) Investeringar i anläggningar där förnybar energi skall användas
Berörda sektorer : Bearbetning och saluföring av jordbruksprodukter
Den beviljande myndighetens namn och adress Comunidad Autónoma de la Región de Murcia
Consejería de Industria y Medio Ambiente
C/San Lorenzo, no 6
E-30071 Murcia
Webbplats :
www.carm.es (Consejería de Industria y Medio Ambiente/ Ayudas y subvenciones:
http://www.carm.es/ceii/subv_detalle_ini.asp?S=TODOS)
Stödnummer : XA 66/05
Medlemsstat : Förenade kungariket
Region : Wales
Stödordningens namn : Projekt om vattenmiljövänligt jordbruk i känsliga avrinningsområden i Wales (Wales Catchment Sensitive Farming Project)
Rättslig grund : Agriculture Act 1986 (Section 1(1)(C) to be read in conjunction with Government of Wales Act 1998 (Sections 40 and 85))
2005: | 5200 GBP |
2006: | 382480 GBP |
2007: | 209180 GBP |
Totalt: | 596860 GBP |
Årliga utgifter under stödordningen Högsta stödnivå 1. Tekniskt bistånd – stöd beviljas upp till 100 %.
2. Investeringsstöd som kan kopplas till en förbättring av miljön – stöd beviljas upp till 60 %
Stödordningen gäller från och med : Den 26 september 2005
Stödordningens varaktighet : Stöd får beviljas till och med den 31 mars 2007. Sista utbetalningsdag är den 30 juni 2007.
Stödets syfte Miljöskydd.
I syfte att skydda vattenmiljön kommer Wales nationalförsamling att inrätta och driva ett projekt för främjande av vattenmiljövänligt jordbruk i känsliga avrinningsområden. Projektet kommer att drivas i två områden med 80 gårdar.
Konsulter kommer att anlitas för att kartlägga föroreningsrisker och gällande krav på skadebegränsning. För den del av stödet som beviljas i enlighet med artikel 14 i förordning 1/2004 kommer konsultarvoden att räknas som berättigande kostnader.
Stöd kan också beviljas till strukturella investeringar som förbättrar vattenmiljön. Sådant stöd beviljas i enlighet med artikel 4 i förordning 1/2004, och följande kommer att räknas som berättigande kostnader:
- Byggnation, förvärv eller förbättring av fast egendom.
- Inköp eller leasing av nya maskiner och utrustning, inklusive datorprogram, upp till tillgångens marknadsvärde. Övriga kostnader i samband med leasingavtal (skatt, uthyrarens påslag, räntekostnader, fasta kostnader, försäkring, m.m.) är inte stödberättigande.
Bara utgifter som leder till väsentligt minskad föroreningsrisk är stödberättigande. Begagnade maskiner är inte stödberättigande
Berörda sektorer :
Syftet med stödordningen är att minska jordbrukets effekter på vattenmiljön. Alla lönsamma jordbruk (oavsett företagsform) i projektområdena kan få stöd.
Det ena området är ett höglänt område där djurhållning (främst nöt och får) är vanligast. Det andra området är ett låglänt område där mjölkproduktion och djurhållning (nöt och får) dominerar.
Den beviljande myndighetens namn och adress National Assembly for Wales
Cathays Park (CP2)
Cardiff CF10 3NQ
United Kingdom
Webbplats :
www.defra.gov.uk/farm/state-aid/setup/exist-exempt.htm. Klicka på Wales Catchment Sensitive Farming Project, eller gå direkt till
http://defraweb/farm/state-aid/setup/schemes/walescatchment.pdf (på engelska) eller http://defraweb/farm/state-aid/setup/schemes/walescatchment-welsh.pdf (på walesiska).
Övrig information Stephen Anderson
Agricultural State Aid Team Leader
Defra
8E9 Millbank
17 Smith Square
London
SW1P 3JR
United Kingdom
Stöd nr : XA 68/05
Medlemsstat : Nederländerna
Region : Ej tillämpligt
Namnet på stödordningen eller namnet på det företag som tar emot det enskilda stödet : Stöd från Hoofdbedrijfschap Agrarische Groothandel för grossisthandel inom den nederländska frukt- och grönsakssektorn
Rättslig grund : Heffingsverordening groenten en fruit 2004, Verordening heffing groenten en fruit 2005 alsmede hun jaarlijkse rechtsopvolgers, welke heffingsverordeningen hun wettelijke basis vinden in artikel 126 van de Wet op de bedrijfsorganisatie
Stödordningens beräknade utgifter per år eller totalt belopp som beviljats företaget som enskilt stöd : Hoofdbedrijfschap Agrarische Groothandel har anslagit 100000 EUR för tekniskt stöd till grossistföretag inom den nederländska frukt- och grönsakssektorn
Högsta stödnivå : 100000 EUR
Datum för genomförande : Efter det nationella godkännandet av avgiftsförordningen (se %quot%Rättslig grund%quot%), dvs. efter det att den tidsfrist på tio arbetsdagar som föreskrivs i förordning (EG) nr 1/2004 har löpt ut
Stödordningens eller det enskilda stödets varaktighet : Med tanke på det fortlöpande behovet av aktuella kunskaper kommer det tekniska stödet att ha obegränsad varaktighet
Stödets syfte : Stödet är riktat till grossistföretag inom frukt- och grönsakssektorn och är avsett att öka deras konkurrenskraft genom att se till att de får tillgång till allmängiltiga kunskaper och information som företagen själva är för små för att skaffa sig. Det är fråga om ett tekniskt stöd i enlighet med artikel 14 i förordning (EG) nr 1/2004
Berörd(a) sektor(er) : Stödordningen är tillämplig på grossistföretag inom frukt- och grönsakssektorn och följaktligen på saluföring av jordbruksprodukter, i synnerhet frukt och grönsaker, utan åtskillnad i fråga om produkternas ursprung
Den beviljande myndighetens namn och adress : Hoofdbedrijfschap Agrarische Groothandel; adres: Postbus 1012, 1430 BA Aalsmeer, Nederland
Webbadress: : www.hbag.nl och www.hbaggroenten.nl
--------------------------------------------------
Sammanfattande information om statliga stöd som beviljas i enlighet med kommissionens förordning (EG) nr 1/2004 av den 23 december 2003 om tillämpningen av artiklarna 87 och 88 i EG-fördraget på statligt stöd till små och medelstora företag som är verksamma inom produktion, bearbetning och saluföring av jordbruksprodukter
(2006/C 16/04)
Stöd nr : XA 57/05
Medlemsstat : Finland
Region : Finländska fastlandet, region utanför mål 1-området
Namn på stödordningen : Stöd till utbildningsprojekt
Rättslig grund : Valtioneuvoston asetus maaseudun kehittämisestä (609/2000, myöhemmin tehtyine muutoksineen), 52 pykälän 2 momentin 4 kohta
Stödordningens beräknade utgifter per år : Under 2006 beräknas 1,9 miljoner EUR beviljas för utbildningsprojekt
Högsta stödnivå :
För ett utbildningsprojekt kan stöd beviljas till högst 90 % av de stödberättigande kostnaderna, dock högst 100000 EUR per stödmottagare över en treårsperiod. Vid beräkning av stödet anses mottagaren vara den person som tar emot det tekniska stödet.
Stödet beviljas i form av bidrag
Datum för genomförande : Från och med den 1.1.2006
Stödordningens eller det enskilda stödets varaktighet : Stöd till utbildningsprojekt beviljas under 2006
Stödets syfte : Att genom stöd till utbildning förbättra jordbrukares och jordbruksanställdas kompetens och yrkeskvalifikationer. Stödet beviljas på grundval av artikel 14 kommissionens förordning (EG) nr 1/2004. Vid beviljandet av stödet följs punkt 14 i gemenskapens riktlinjer för statligt stöd till jordbrukssektorn
Berörda sektorer : Jordbruk
Den beviljande myndighetens namn och adress Södra Österbottens TE-central
Huhtalantie 2
FIN-60220 Seinäjoki
Tavastlands TE-central
Rauhankatu 10
FIN-15110 Lahtis
Sydöstra Finlands TE-central
Salpausselänkatu 22, PB 1041
FIN-45101 Kouvola
Mellersta Finlands TE-central
Cygnaeuksenkatu 1, PL 44
FIN-40101 Jyväskylä
Birkalands TE-central
Kauppakatu 4, PB 467
FIN-33101 Tammerfors
Österbottens TE-central
Hovrättsesplanaden 19 A, PB 131
FIN-65101 Vasa
Norra Österbottens TE-central
Viestikatu 1, PB 86
FIN-90101 Uleåborg
Satakunta TE-central
Pohjoisranta 11 E, PB 266
FIN-28100 Björneborg
Nylands TE-central
Magistratsporten 2, PB 15
FIN-00241 Helsingfors
Egentliga Finlands TE-central
Bangårdsgatan 36, PB 592
FIN-20101 Åbo
Webbplats : www.mmm.fi/tuet/valtiontuet/ryhmapoikkeusasetus
--------------------------------------------------
Republiken Libanons uppfyllande av vissa administrativa samarbetsformaliteter för att bevisa produktens ursprung
(Meddeland enligt artikel 11 i kommissionens förordning (EG) nr 565/2002)
(2006/C 34/03)
I enlighet med artikel 11 i förordning (EG) nr 565/2002 [1] meddelar kommissionen härmed importörer och berörda administrationer att Republiken Libanon till kommissionen har översänt avtryck av de stämplar som används av de libanesiska myndigheterna, och namn och adress till de libanesiska myndigheter som ansvarar för att utfärda och ta emot ansökningar om kontroller i efterhand av ursprungscertifikat. Dessa krav uppfylldes den 13 oktober 2005.
[1] EUT L 86, 3.4.2002, s. 11. Förordningen senast ändrad genom förordning (EG) nr 537/2004 (EUT L 86, 24.3.2004, s. 9).
--------------------------------------------------
Förlängning och ändring av bestämmelserna om allmän trafikplikt för regelbunden lufttrafik på flyglinjer i Grekland i enlighet med rådets förordning (EEG) nr 2408/92
(2006/C 46/06)
(Text av betydelse för EES)
1. Grekland har beslutat att från och med den 1 april 2006 förlänga och delvis ändra de bestämmelser om allmän trafikplikt för regelbunden lufttrafik på flyglinjer inom Grekland som införts i enlighet med artikel 4.1 a i rådets förordning (EEG) nr 2408/92 av den 23 juli 1992 om EG-lufttrafikföretags tillträde till flyglinjer inom gemenskapen och som offentliggjorts i Europeiska gemenskapernas officiella tidning C 164 av den 10 juli 2002.
2. Ändringarna av den allmänna trafikplikten omfattar följande:
A) När det gäller minsta antal flygningar och minsta antal tillgängliga platser per vecka på följande linjer:
- Aten – Karpathos
- Aten – Sitia
- Thessaloniki – Kerkira (Korfu)
Aten – Karpathos
Tre flygningar tur och retur per vecka, med sammanlagt 150 platser per vecka i båda riktningarna under vinterhalvåret.
Sju flygningar tur och retur per vecka, med sammanlagt 350 platser per vecka i båda riktningarna under sommarhalvåret.
Aten – Sitia
Tre flygningar tur och retur per vecka, med sammanlagt 90 platser per vecka i båda riktningarna under vinterhalvåret.
Fyra flygningar tur och retur per vecka, med sammanlagt 120 platser per vecka i båda riktningarna under sommarhalvåret.
Thessaloniki – Kerkira (Korfu)
Tre flygningar tur och retur per vecka, med sammanlagt 180 platser per vecka i båda riktningarna under vinterhalvåret.
Fyra flygningar tur och retur per vecka, med sammanlagt 240 platser per vecka i båda riktningarna under sommarhalvåret.
B) När det gäller priset:
Priset för en enkel biljett i ekonomiklass får inte överstiga följande:
—Mellan Aten och Kithira: | 40 EUR |
—Mellan Aten och Naxos: | 54 EUR |
—Mellan Aten och Paros: | 53 EUR |
—Mellan Aten och Karpathos: | 64 EUR |
—Mellan Aten och Sitia: | 62 EUR |
—Mellan Aten och Skiathos: | 45 EUR |
—Mellan Thessaloniki och Korfu: | 60 EUR |
—Mellan Rhodos och Kos: | 38 EUR |
—Mellan Rhodos och Astypalea: | 44 EUR |
—Mellan Rhodos och Leros: | 44 EUR |
—Mellan Kos och Astypalea: | 44 EUR |
—Mellan Kos och Leros: | 38 EUR |
—Mellan Astypalea och Leros: | 38 EUR |
—Mellan Kerkira och Aktio: | 33 EUR |
—Mellan Kerkira och Kefalinia: | 33 EUR |
—Mellan Kerkira och Zakynthos: | 44 EUR |
—Mellan Aktio och Kefalinia: | 28 EUR |
—Mellan Aktio och Zakynthos: | 33 EUR |
—Mellan Kefalinia och Zakynthos: | 26 EUR |
3. Viktiga upplysningar:
Om inget lufttrafikföretag senast den 1 mars 2006 har meddelat Civil Aviation Department, Directorate for Air Operations sin avsikt att från och med den 1 april 2006 bedriva regelbunden trafik på en eller flera av de ovannämnda flyglinjerna, utan att begära ekonomisk ersättning, har Grekland beslutat att, enligt det förfarande som föreskrivs i artikel 4.1 d i förordning (EEG) nr 2408/92, begränsa tillträdet till en eller flera av flyglinjerna till endast ett trafikföretag under tre år och efter anbudsinfordran bevilja rätten att bedriva trafik på flyglinjerna från och med den 1 april 2006.
På de tre ovannämnda flyglinjerna ersätter skyldigheterna och priserna dem som fastställs i Europeiska gemenskapernas officiella tidning C 239 av den 25 augusti 2001.
I övriga avseenden skall den allmänna trafikplikt som offentliggjordes i Europeiska gemenskapernas officiella tidning C 239 av den 25 augusti 2001 fortsätta att gälla.
--------------------------------------------------
Kommissionens meddelande inom ramen för genomförandet av Rådets direktiv 89/686/EEG av den 21 december 1989 om tillnärmning av medlemsstaternas lagstiftning om personlig skyddsutrustning
(2006/C 91/03)
(Text av betydelse för EES)
(Offentliggörande av titlar på och hänvisningar till harmoniserade standarder inom ramen för direktivet)
ESO [1] | Titel på och hänvisning till standarden (samt referensdokument) | Första offentliggörandet EGT | Hänvisning till den ersatta standarden | Datum då standarden upphör att gälla Anm. 1 |
CEN | EN 132:1998 Andningsskydd – Definitioner | 4.6.1999 | EN 132:1990 | Datum passerat ( 30.6.1999) |
CEN | EN 133:2001 Andningsskydd – Klassifikation | 10.8.2002 | EN 133:1990 | Datum passerat ( 10.8.2002) |
CEN | EN 134:1998 Andningsskydd – Terminologi för komponenter och detaljer | 13.6.1998 | EN 134:1990 | Datum passerat ( 31.7.1998) |
CEN | EN 135:1998 Andningsskydd – Ordlista | 4.6.1999 | EN 135:1990 | Datum passerat ( 30.6.1999) |
CEN | EN 136:1998 Andningsskydd – Helmasker – Fordringar, provning, märkning | 13.6.1998 | EN 136:1989 EN 136-10:1992 | Datum passerat ( 31.7.1998) |
EN 136:1998/AC:1999 | | | |
CEN | EN 137:1993 Andningsskydd – Bärbar tryckluftsapparat med öppet system – Fordringar, provning, märkning | 23.12.1993 | EN 137:1986 | Datum passerat ( 23.12.1993) |
EN 137:1993/AC:1993 | | | |
CEN | EN 138:1994 Andningsskydd – Sugslangsapparat för helmask, halvmask eller bitmunstycke – Fordringar, provning, märkning | 16.12.1994 | — | |
CEN | EN 140:1998 Andningsskydd – Halv- och kvartsmasker – Fordringar, provning, märkning | 6.11.1998 | EN 140:1989 | Datum passerat ( 31.3.1999) |
EN 140:1998/AC:1999 | | | |
CEN | EN 142:2002 Andningsskydd – Bitmunstycksenheter – Fordringar, provning, märkning | 10.4.2003 | EN 142:1989 | Datum passerat ( 10.4.2003) |
CEN | EN 143:2000 Andningsskydd – Partikelfilter – Fordringar, provning, märkning | 24.1.2001 | EN 143:1990 | Datum passerat ( 24.1.2001) |
Varning! När det gäller partikelfilter, vars filtereffekt helt eller delvis baseras på elektrostatiskt laddade fiberfiltermaterial, gäller detta offentliggörande inte punkt 8.7.2.4 sista meningen, punkt 8.7.3.4 sista meningen och punkt 10 i standarden, för vilka offentliggörandet inte innebär något antagande om överensstämmelse med de grundläggande hälso- och säkerhetskraven i direktiv 89/686/EEG. Denna varning skall också beaktas vid tillämpningen av följande harmoniserade standarder: EN 149:2001, EN 405:2001, EN 1827:1999, EN 12083:1998, EN 12941:1998, EN 12941:1998+A1:2003, EN 12942:1998, EN 12942:1998+A1:2002, EN 13274-7:2002. |
CEN | EN 144-1:2000 Andningsskydd – Gasflaskventiler – Del 1: Flaskhalsgängor | 24.1.2001 | EN 144-1:1991 | Datum passerat ( 24.1.2001) |
EN 144-1:2000/A1:2003 | 21.2.2004 | Anmärkning 3 | Datum passerat ( 31.10.2003) |
EN 144-1:2000/A2:2005 | 6.10.2005 | Anmärkning 3 | Datum passerat ( 31.12.2005) |
CEN | EN 144-2:1998 Andningsskydd – Gasflaskventiler – Del 2: Utlopp | 4.6.1999 | — | |
CEN | EN 144-3:2003 Andningsskydd – Gasflaskventiler – Del 3: Utlopp för dykgaserna Nitrox-blandningar och syrgas | 21.2.2004 | — | |
CEN | EN 145:1997 Andningsskydd – Bärbar andningsapparat med slutet system för komprimerad oxygen eller komprimerad oxygen/nitrogen – Fordringar, provning, märkning | 19.2.1998 | EN 145:1988 EN 145-2:1992 | Datum passerat ( 28.2.1998) |
EN 145:1997/A1:2000 | 24.1.2001 | Anmärkning 3 | Datum passerat ( 24.1.2001) |
CEN | EN 148-1:1999 Andningsskydd – Gängor för ansiktsmasker – Del 1: Anslutning med standardgänga | 4.6.1999 | EN 148-1:1987 | Datum passerat ( 31.8.1999) |
CEN | EN 148-2:1999 Andningsskydd – Gängor för ansiktsmasker – Anslutning med centrumgänga | 4.6.1999 | EN 148-2:1987 | Datum passerat ( 31.8.1999) |
CEN | EN 148-3:1999 Andningsskydd – Gängor för ansiktsmasker – Del 3: Anslutning med gänga M45x3 | 4.6.1999 | EN 148-3:1992 | Datum passerat ( 31.8.1999) |
CEN | EN 149:2001 Andningsskydd – Filtrerande halvmasker mot partiklar – Fordringar, provning, märkning | 21.12.2001 | EN 149:1991 | Datum passerat ( 21.12.2001) |
CEN | EN 165:2005 Ögonskydd – Terminologi | Detta är det första offentliggörandet | EN 165:1995 | 31.5.2006 |
CEN | EN 166:2001 Ögonskydd – Fordringar och specifikationer | 10.8.2002 | EN 166:1995 | Datum passerat ( 10.8.2002) |
CEN | EN 167:2001 Ögonskydd – Optiska provningsmetoder | 10.8.2002 | EN 167:1995 | Datum passerat ( 10.8.2002) |
CEN | EN 168:2001 Ögonskydd – Icke-optiska provningsmetoder | 10.8.2002 | EN 168:1995 | Datum passerat ( 10.8.2002) |
CEN | EN 169:2002 Ögonskydd – Filter vid svetsning och besläktade förfaranden – Fordringar på transmittans | 28.8.2003 | EN 169:1992 | Datum passerat ( 28.8.2003) |
CEN | EN 170:2002 Ögonskydd – Filter mot ultraviolett strålning – Fordringar på transmittans | 28.8.2003 | EN 170:1992 | Datum passerat ( 28.8.2003) |
CEN | EN 171:2002 Ögonskydd – Filter mot infraröd strålning – Fordringar på transmittans | 10.4.2003 | EN 171:1992 | Datum passerat ( 10.4.2003) |
CEN | EN 172:1994 Ögonskydd – Solglasögon för yrkesarbete | 15.5.1996 | — | |
EN 172:1994/A1:2000 | 4.7.2000 | Anmärkning 3 | Datum passerat ( 31.10.2000) |
EN 172:1994/A2:2001 | 10.8.2002 | Anmärkning 3 | Datum passerat ( 10.8.2005) |
CEN | EN 174:2001 Ögonskydd – Skidglasögon för utförsåkning | 21.12.2001 | EN 174:1996 | Datum passerat ( 21.12.2001) |
CEN | EN 175:1997 Personligt skydd – Ögon- och ansiktsskydd vid svetsning och likartatarbete | 19.2.1998 | — | |
CEN | EN 207:1998 Ögonskydd – Filter mot laserstrålning | 21.11.1998 | EN 207:1993 | Datum passerat ( 31.3.1999) |
EN 207:1998/A1:2002 | 28.8.2003 | Anmärkning 3 | Datum passerat ( 28.8.2003) |
CEN | EN 208:1998 Ögonskydd – Filter för användning under justering av lasrar och lasersystem | 21.11.1998 | EN 208:1993 | Datum passerat ( 31.3.1999) |
EN 208:1998/A1:2002 | 28.8.2003 | Anmärkning 3 | Datum passerat ( 28.8.2003) |
CEN | EN 250:2000 Andningsskydd – Bärbar tryckluftsapparat med öppet system för dykning – Fordringar, provning, märkning | 8.6.2000 | EN 250:1993 | Datum passerat ( 19.7.2000) |
CEN | EN 269:1994 Andningsskydd – Fläktassisterad sugslangsapparat med huva – Fordringar, provning, märkning | 16.12.1994 | — | |
CEN | EN 340:2003 Skyddskläder – Allmänna fordringar | 6.10.2005 | EN 340:1993 | Datum passerat ( 6.10.2005) |
CEN | EN 341:1992 Personlig fallskyddsutrustning – Nedfirningsdon | 23.12.1993 | — | |
EN 341:1992/A1:1996 | 6.11.1998 | Anmärkning 3 | Datum passerat ( 6.11.1998) |
EN 341:1992/AC:1993 | | | |
CEN | EN 342:2004 Skyddskläder – Hela dräkter och plagg till skydd mot kyla | 6.10.2005 | — | |
CEN | EN 343:2003 Skyddskläder – Skydd mot dåligt väder | 21.2.2004 | — | |
CEN | EN 348:1992 Skyddskläder – Provningsmetod: Bestämning av materials motstånd vid påverkan av små stänk av smält metall | 23.12.1993 | — | |
EN 348:1992/AC:1993 | | | |
CEN | EN 352-1:2002 Hörselskydd – Allmänna fordringar – Del 1: Kåpor | 28.8.2003 | EN 352-1:1993 | Datum passerat ( 28.8.2003) |
CEN | EN 352-2:2002 Hörselskydd – Allmänna fordringar – Del 2: Proppar | 28.8.2003 | EN 352-2:1993 | Datum passerat ( 28.8.2003) |
CEN | EN 352-3:2002 Hörselskydd – Allmänna fordringar – Del 3: Kåpor monterade på industrihjälm | 28.8.2003 | EN 352-3:1996 | Datum passerat ( 28.8.2003) |
CEN | EN 352-4:2001 Hörselskydd – Fordringar och provning – Del 4: Nivåberoende kåpor | 10.8.2002 | — | |
EN 352-4:2001/A1:2005 | Detta är det första offentliggörandet | Anmärkning 3 | 30.4.2006 |
CEN | EN 352-5:2002 Hörselskydd – Fordringar och provning – Del 5: Kåpor med aktiv bullerdämpning | 28.8.2003 | — | |
CEN | EN 352-6:2002 Hörselskydd – Fordringar och provning – Del 6: Kåpor med elektrisk ljudingång | 28.8.2003 | — | |
CEN | EN 352-7:2002 Hörselskydd – Fordringar och provning – Del 7: Nivåberoende proppar | 28.8.2003 | — | |
CEN | EN 353-1:2002 Personlig fallskyddsutrustning – Del 1: Styrt glidlås på fast förankringslina eller skena | 28.8.2003 | EN 353-1:1992 | Datum passerat ( 28.8.2003) |
CEN | EN 353-2:2002 Personlig fallskyddutrustning – Styrt glidlås på flexibel förankringslina | 28.8.2003 | EN 353-2:1992 | Datum passerat ( 28.8.2003) |
CEN | EN 354:2002 Personlig fallskyddsutrustning – Kopplingslinor | 28.8.2003 | EN 354:1992 | Datum passerat ( 28.8.2003) |
CEN | EN 355:2002 Personlig fallskyddsutrustning – Falldämpare | 28.8.2003 | EN 355:1992 | Datum passerat ( 28.8.2003) |
CEN | EN 358:1999 Personlig skyddsutrustning med stödjande och fallhindrande funktion – Stödbälten och fallhindrande kopplingslinor för stödutrustning | 21.12.2001 | EN 358:1992 | Datum passerat ( 21.12.2001) |
CEN | EN 360:2002 Personlig fallskyddsutrustning – Säkerhetsblock | 28.8.2003 | EN 360:1992 | Datum passerat ( 28.8.2003) |
CEN | EN 361:2002 Personlig fallskyddsutrustning – Helselar | 28.8.2003 | EN 361:1992 | Datum passerat ( 28.8.2003) |
CEN | EN 362:2004 Personlig fallskyddsutrustning – Kopplingsanordningar | 6.10.2005 | EN 362:1992 | Datum passerat ( 6.10.2005) |
CEN | EN 363:2002 Personlig fallskyddsutrustning – Fallskyddssystem | 28.8.2003 | EN 363:1992 | Datum passerat ( 28.8.2003) |
CEN | EN 364:1992 Personlig fallskyddsutrustning – Provningsmetoder | 23.12.1993 | — | |
EN 364:1992/AC:1993 | | | |
CEN | EN 365:2004 Personlig fallskyddsutrustning – Allmänna fordringar för bruksanvisningar, användning, underhåll, periodisk kontroll, reparation, märkning och förpackning | 6.10.2005 | EN 365:1992 | Datum passerat ( 6.10.2005) |
CEN | EN 367:1992 Skyddskläder – Skydd mot hetta och flamma – Metod för bestämningav värmegenomgång vid påverkan av flamma | 23.12.1993 | — | |
EN 367:1992/AC:1992 | | | |
CEN | EN 373:1993 Skyddskläder – Bedömning av motstånd hos material vid stänk av smält metall | 23.12.1993 | — | |
CEN | EN 374-1:2003 Skyddshandskar mot kemikalier och mikroorganismer – Del 1: Terminologi och fordringar på prestanda | 6.10.2005 | EN 374-1:1994 | Datum passerat ( 6.10.2005) |
CEN | EN 374-2:2003 Skyddshandskar mot kemikalier och mikroorganismer – Del 2: Bestämning av motstånd mot penetration | 6.10.2005 | EN 374-2:1994 | Datum passerat ( 6.10.2005) |
CEN | EN 374-3:2003 Skyddshandskar mot kemikalier och mikroorganismer – Del 3: Bestämning av motstånd mot permeation av kemikalier | 6.10.2005 | EN 374-3:1994 | Datum passerat ( 6.10.2005) |
CEN | EN 379:2003 Ögonskydd – Automatiska svetsfilter | 6.10.2005 | EN 379:1994 | Datum passerat ( 6.10.2005) |
CEN | EN 381-1:1993 Skyddskläder för användare av handhållna kedjesågar – Del 1: Provningsutrustning för provning av motstånd mot genomsågning med kedjesåg | 23.12.1993 | — | |
CEN | EN 381-2:1995 Sågningsskydd – Del 2: Provningsmetoder för benskydd | 12.1.1996 | — | |
CEN | EN 381-3:1996 Sågningsskydd – Del 3: Provningsmetoder för skyddskodon | 10.10.1996 | — | |
CEN | EN 381-4:1999 Sågningsskydd – Del 4: Provningsmetoder för handskar till skydd mot kedjesåg | 16.3.2000 | — | |
CEN | EN 381-5:1995 Sågningsskydd – Del 5: Fordringar för benskydd | 12.1.1996 | — | |
CEN | EN 381-7:1999 Sågningsskydd – Del 7: Fordringar för handskar till skydd mot kedjesåg | 16.3.2000 | — | |
CEN | EN 381-8:1997 Skyddskläder för användare av handhållna kedjesågar – Del 8: Provningsmetoder för damasker till skydd mot kedjesåg | 18.10.1997 | — | |
CEN | EN 381-9:1997 Skyddskläder för användare av handhållna kedjesågar – Del 9: Fordringar för damasker till skydd mot kedjesåg | 18.10.1997 | — | |
CEN | EN 381-10:2002 Sågningsskydd – Del 10: Provningsmetoder för skydd för överkroppen | 28.8.2003 | — | |
CEN | EN 381-11:2002 Sågningsskydd – Del 11: Fordringar för skydd för överkroppen | 28.8.2003 | — | |
CEN | EN 388:2003 Skyddshandskar mot mekaniska risker | 6.10.2005 | EN 388:1994 | Datum passerat ( 6.10.2005) |
CEN | EN 393:1993 Flytvästar – Flytplagg – 50 N | 16.12.1994 | — | |
EN 393:1993/A1:1998 | 6.11.1998 | Anmärkning 3 | Datum passerat ( 6.11.1998) |
EN 393:1993/AC:1995 | | | |
CEN | EN 394:1993 Flytvästar – Tilläggsutrustning | 16.12.1994 | — | |
CEN | EN 395:1993 Flytvästar – Räddningsvästar – 100 N | 16.12.1994 | — | |
EN 395:1993/A1:1998 | 6.11.1998 | Anmärkning 3 | Datum passerat ( 6.11.1998) |
EN 395:1993/AC:1995 | | | |
CEN | EN 396:1993 Flytvästar – Räddningsvästar – 150 N | 16.12.1994 | — | |
EN 396:1993/A1:1998 | 6.11.1998 | Anmärkning 3 | Datum passerat ( 6.11.1998) |
EN 396:1993/AC:1995 | | | |
CEN | EN 397:1995 Industrihjälmar | 12.1.1996 | — | |
EN 397:1995/A1:2000 | 24.1.2001 | Anmärkning 3 | Datum passerat ( 24.1.2001) |
CEN | EN 399:1993 Flytvästar – Räddningsvästar – 275 N | 16.12.1994 | — | |
EN 399:1993/A1:1998 | 6.11.1998 | Anmärkning 3 | Datum passerat ( 6.11.1998) |
EN 399:1993/AC:1995 | | | |
CEN | EN 402:2003 Andningsskydd, flyktutrustning – Bärbar tryckluftsapparat med öppet system med helmask eller bitmunstycksenhet – Fordringar, provning, märkning | 21.2.2004 | EN 402:1993 | Datum passerat ( 21.2.2004) |
CEN | EN 403:2004 Andningsskydd – Flyktfilterskydd med huva vid brand – Fordringar, provning, märkning | 6.10.2005 | EN 403:1993 | Datum passerat ( 6.10.2005) |
CEN | EN 404:2005 Andningsskydd – Flyktfilter – Fordringar, provning, märkning | 6.10.2005 | EN 404:1993 | Datum passerat ( 2.12.2005) |
CEN | EN 405:2001 Andningsskydd – Filtrerande halvmasker med ventiler mot gaser eller gaser och partiklar – Fordringar, provning, märkning | 10.8.2002 | EN 405:1992 | Datum passerat ( 10.8.2002) |
CEN | EN 407:2004 Skyddshandskar mot termiska risker (hetta och/eller brand) | 6.10.2005 | EN 407:1994 | Datum passerat ( 6.10.2005) |
CEN | EN 420:2003 Allmänna fordringar för handskar Anmärkning 4 | 2.12.2005 | EN 420:1994 | Datum passerat ( 2.12.2005) |
CEN | EN 421:1994 Skyddshandskar mot joniserande strålning och radioaktiv förorening | 16.12.1994 | — | |
CEN | EN 443:1997 Skyddshjälmar för brandmän | 19.2.1998 | — | |
CEN | EN 458:2004 Hörselskydd – Rekommendationer för val, användning, skötsel och underhåll – Vägledande dokument | 6.10.2005 | EN 458:1993 | Datum passerat ( 6.10.2005) |
CEN | EN 463:1994 Skyddskläder – Skydd mot kemikalier i vätskeform – Provningsmetod: Bestämning av motstånd mot penetration av en vätskestråle (vätskestrålprovning) | 16.12.1994 | — | |
CEN | EN 464:1994 Skyddskläder – Skydd mot kemikalier i vätske- och gasform, inklusive vätskeaerosoler och fasta partiklar – Provningsmetod: Bestämning av täthet hos gastäta dräkter (trycktäthetsprovning) | 16.12.1994 | — | |
CEN | EN 468:1994 Skyddskläder – Skydd mot kemikalier i vätskeform – Provningsmetod: Bestämning av motstånd mot penetration av stänk(stänkprovning) | 16.12.1994 | — | |
CEN | EN 468:1994 Skyddskläder – Skydd mot kemikalier i vätskeform – Provningsmetod: Bestämning av motstånd mot penetration av stänk(stänkprovning) | Detta är det första offentliggörandet | EN 469:1995 | 30.6.2005 |
CEN | EN 470-1:1995 Skyddskläder för användning vid svetsarbete ellerlikartat arbete – Del 1: Allmänna fordringar | 12.1.1996 | — | |
EN 470-1:1995/A1:1998 | 13.6.1998 | Anmärkning 3 | Datum passerat ( 31.8.1998) |
CEN | EN 471:2003 Skyddskläder med god synbarhet (Varselklädsel) för yrkesbruk | 6.10.2005 | EN 471:1994 | Datum passerat ( 6.10.2005) |
CEN | EN 510:1993 Specifikation för skyddskläder som används där risk föreligger att fastna i rörliga delar | 16.12.1994 | — | |
CEN | EN 511:1994 Skyddshandskar mot kyla | 16.3.2000 | — | |
CEN | EN 530:1994 Nötningshållfasthet hos material för skyddskläder – Provningsmetoder | 30.8.1995 | — | |
EN 530:1994/AC:1995 | | | |
CEN | EN 531:1995 Skyddskläder för industriarbetare som exponeras för hetta (med undantag för brandmansdräkter och svetsarbetskläder) | 6.11.1998 | — | |
EN 531:1995/A1:1998 | 4.6.1999 | Anmärkning 3 | Datum passerat ( 4.6.1999) |
CEN | EN 533:1997 Skyddskläder – Skydd mot hetta och flamma – Material och materialkombinationer för begränsad flamspridning | 14.6.1997 | — | |
CEN | EN 564:1997 Klätterutrustning – Repsnöre – Säkerhetskrav och provningsmetoder | 10.8.2002 | — | |
CEN | EN 565:1997 Klätterutrustning – Band – Säkerhetskrav och provningsmetoder | 10.8.2002 | — | |
CEN | EN 566:1997 Klätterutrustning – Slingor – Säkerhetskrav och provningsmetoder | 10.8.2002 | — | |
CEN | EN 567:1997 Klätterutrustning – Repklämmor – Säkerhetskrav och provningsmetoder | 10.8.2002 | — | |
CEN | EN 568:1997 Klätterutrustning – Issäkringar – Säkerhetskrav och provningsmetoder | 14.6.1997 | — | |
CEN | EN 569:1997 Klätterutrustning – Bultar – Säkerhetskrav och provningsmetoder | 10.8.2002 | — | |
CEN | EN 659:2003 Skyddshandskar för brandmän | 21.2.2004 | EN 659:1996 | Datum passerat ( 21.2.2004) |
CEN | EN 702:1994 Skyddskläder – Skydd mot hetta och flamma – Provningsmetod: Bestämning av kontaktvärmegenomgång genom skyddsklädereller deras material | 12.1.1996 | — | |
CEN | EN 795:1996 Fallskydd – Förankringsutrustning – Fordringar och provning | 12.2.2000 | — | |
Anmärkning: Detta offentliggörande gäller inte klass A ("structural anchors"), C ("anchor devices employing horizontal flexible lines") eller D ("anchor devices employing horizontal rigid anchor rails") som omnämns i punkterna 3.13.1, 3.13.3, 3.13.4, 4.3.1, 4.3.3, 4.3.4, 5.2.1, 5.2.2, 5.2.4, 5.2.5, 5.3.2 (vad gäller klass A 1) 5.3.3, 5.3.4, 5.3.5, 6 (vad gäller klass A, C och D), bilaga A (stycke A.2, A.3, A.5 och A.6), bilaga B, bilaga ZA (vad gäller klass A, C och D). Dessa kan inte förutsättas överensstämma med bestämmelserna i direktiv 89/686/EEG. |
| EN 795:1996/A1:2000 | 24.1.2001 | Anmärkning 3 | Datum passerat ( 30.4.2001) |
CEN | EN 812:1997 Stötskyddsmössor | 19.2.1998 | — | |
EN 812:1997/A1:2001 | 10.8.2002 | Anmärkning 3 | Datum passerat ( 10.8.2002) |
CEN | EN 813:1997 Personlig skyddsutrustning med fallhindrande funktion – Sittselar | 14.6.1997 | — | |
CEN | EN 863:1995 Skyddskläder – Mekaniska egenskaper – Provningsmetod: Motstånd mot punktering | 15.5.1996 | — | |
CEN | EN 892:2004 Utrustning för bergsklättring – Dynamiska klätterrep – Säkerhetskrav och provningsmetoder | 6.10.2005 | EN 892:1996 | Datum passerat ( 6.10.2005) |
CEN | EN 893:1999 Klätterutrustning – Isbroddar – Säkerhetskrav och provningsmetoder | 10.8.2002 | — | |
CEN | EN 943-1:2002 Skyddskläder för användning mot kemikalier i vätske- och gasform inklusive vätskeaerosoler och fasta partiklar – Del 1: Fordringar på prestanda för ventilerade och ej ventilerade "gastäta" (Typ 1) och "ej gastäta" (Typ 2) skyddskläder | 28.8.2003 | — | |
CEN | EN 943-2:2002 Skyddskläder mot kemikalier i vätske- och gasform inklusive vätskeaerosoler och fasta partiklar – Del 2: Funktionskrav för gastäta (Typ 1) skyddsdräkter för insatsstyrkor | 10.8.2002 | — | |
CEN | EN 958:1996 Klätterutrustning – Falldämpande system för användning vid klättring på klätterstigar (via ferrata) – Säkerhetskrav ochprovningsmetoder | 14.6.1997 | — | |
CEN | EN 960:1994 Skyddshjälmar – Modellhuvud för provning | 15.5.1996 | — | |
EN 960:1994/A1:1998 | 6.11.1998 | Anmärkning 3 | Datum passerat ( 6.11.1998) |
CEN | EN 966:1996 Luftsporthjälmar | 10.10.1996 | — | |
EN 966:1996/A1:2000 | 4.7.2000 | Anmärkning 3 | Datum passerat ( 30.9.2000) |
CEN | EN 1073-1:1998 Skyddskläder – Skydd mot hetta och flamma – Provningsmetod: Bestämning av kontaktvärmegenomgång genom skyddsklädereller deras material | 6.11.1998 | — | |
CEN | EN 1073-2:2002 Skyddskläder mot radioaktiva föroreningar – Del 2: Fordringar och provningsmetoder för icke ventilerade skyddskläder mot radioaktiva föreningar i partikelform | 28.8.2003 | — | |
CEN | EN 1077:1996 Skidhjälmar | 10.10.1996 | — | |
CEN | EN 1078:1997 Hjälmar för cyklister, skateboard- och rullskridskoåkare | 14.6.1997 | — | |
EN 1078:1997/A1:2005 | Detta är det första offentliggörandet | Anmärkning 3 | 30.6.2006 |
CEN | EN 1080:1997 Småbarnshjälmar | 14.6.1997 | — | |
EN 1080:1997/A1:2002 | 28.8.2003 | Anmärkning 3 | Datum passerat ( 28.8.2003) |
EN 1080:1997/A2:2005 | Detta är det första offentliggörandet | Anmärkning 3 | 30.6.2006 |
CEN | EN 1082-1:1996 Skyddskläder – Handskar och armskydd mot skär och stick av handhållna knivar – Del 1: Brynjehandskar och armskydd | 14.6.1997 | — | |
CEN | EN 1082-2:2000 Skyddskläder – Handskar och armskydd mot skär och stick av handhållna knivar – Del 2: Handskar och armskydd av andra material än ringbrynjor | 21.12.2001 | — | |
CEN | EN 1082-3:2000 Skyddskläder – Handskar och armskydd mot skär och stick av handhållna knivar – Del 3: Stöt- och skärprovning av tyg, läder och andra material | 21.12.2001 | — | |
CEN | EN 1095:1998 Säkerhetsselar och säkerhetslinor för fritidsbåtar – Säkerhetskrav och provningsmetoder | 6.11.1998 | — | |
CEN | EN 1146:2005 Andningsskydd, flyktutrustning – Bärbar tryckluftsapparat med öppet system, med huva för utrymning – Fordringar, provning, märkning | Detta är det första offentliggörandet | EN 1146:1997 | 30.4.2006 |
CEN | EN 1149-1:1995 Skyddskläder – Elektrostatiska egenskaper – Del 1: Ytresistivitet (Provningsmetoder och fordringar) | 10.10.1996 | — | |
CEN | EN 1149-2:1997 Skyddskläder – Elektrostatiska egenskaper – Del 2: Provningsmetod för mätning av elektrisk resistans genom ett material (vertikal resistans) | 19.2.1998 | — | |
CEN | EN 1149-3:2004 Skyddskläder – Elektrostatiska egenskaper – Del 3: Provningsmetoder för mätning av avklingningstid | 6.10.2005 | — | |
CEN | EN 1150:1999 Skyddskläder – Kläder med god synbarhet för icke yrkesmässigt bruk – Provningsmetoder och fordringar | 4.6.1999 | — | |
CEN | EN 1384:1996 Ridhjälmar | 14.6.1997 | — | |
EN 1384:1996/A1:2001 | 10.8.2002 | Anmärkning 3 | Datum passerat ( 10.8.2002) |
CEN | EN 1385:1997 Kanothjälmar | 13.6.1998 | — | |
EN 1385:1997/A1:2005 | 6.10.2005 | Anmärkning 3 | Datum passerat ( 6.10.2005) |
CEN | EN 1486:1996 Skyddskläder för brandmän – Provningsmetoder och fordringar för värmereflekterande kläder för speciell brandbekämpning | 3.12.1996 | — | |
CEN | EN 1621-1:1997 Skyddskläder mot mekaniska stötar för motorcyklister – Del 1: Fordringar och provningsmetoder för stötskydd | 13.6.1998 | — | |
CEN | EN 1621-2:2003 Skyddskläder mot mekanisk påverkan för motorcyklister – Del 2: Ryggskydd – Krav och provningsmetoder | 6.10.2005 | — | |
CEN | EN 1731:1997 Ögon- och ansiktsskydd av nättyp, för industrielleller icke-industriell användning mot mekaniska och/eller värmerisker | 14.6.1997 | — | |
EN 1731:1997/A1:1997 | 13.6.1998 | Anmärkning 3 | Datum passerat ( 30.6.1998) |
CEN | EN 1809:1997 Dykutrustning – Avvägningsvästar – Funktions- ochsäkerhetskrav, provningsmetoder | 13.6.1998 | — | |
CEN | EN 1827:1999 Andningsskydd – Halvmasker utan inandningsventiler och med separata filter mot gaser eller gaser och partiklar eller enbar partiklar – Fordringar, provning, märkning | 24.2.2001 | — | |
CEN | EN 1836:2005 Ögonskydd – Solglasögon och solskyddsfilter för allmänt bruk samt filter för direkt iakttagelse av solen | 2.12.2005 | EN 1836:1997 | Datum passerat ( 31.3.2006) |
CEN | EN 1868:1997 Personlig fallskyddsutrustning – Ordlista | 18.10.1997 | — | |
CEN | EN 1891:1998 Personlig fallskyddsutrustning – Statiska kärnmantelrep | 6.11.1998 | — | |
CEN | EN 1938:1998 Ögonskydd – Skyddsglasögon för motorcykel- och mopedförare | 4.6.1999 | — | |
CEN | EN ISO 4869-2:1995 Akustik – Hörselskydd – Del 2: Uppskattning av effekt A-vägd ljudtrycksnivå vid användning av hörselskydd (ISO 4869-2:1994) | 15.5.1996 | — | |
CEN | EN ISO 4869-4:2000 Akustik – Hörselskydd – Del 4: Mätning av effektiv ljudtrycksnivå för nivåberoende hörselskydd med ljudåtergivningssystem (ISO/TR 4869-4:1998) | 6.10.2005 | — | |
CEN | EN ISO 6529:2001 Skyddskläder – Skydd mot kemikalier – Bestämning av motstånd mot penetration av vätskor och gaser hos material för skyddskläder (ISO 6529:2001) | 6.10.2005 | EN 369:1993 | Datum passerat ( 6.10.2005) |
CEN | EN ISO 6530:2005 Skyddskläder – Skydd mot kemikalier i vätskeform – Provningsmetod för bestämning av motstånd mot penetration av vätskor hos material för skyddskläder (ISO 6530:2005) | 6.10.2005 | EN 368:1992 | Datum passerat ( 6.10.2005) |
CEN | EN ISO 6942:2002 Skyddskläder – Skydd mot hetta och brand – Provningsmetod: Utvärdering av material och materialkombinationer som exponeras för en källa med strålningsvärme (ISO 6942:2002) | 28.8.2003 | EN 366:1993 | Datum passerat ( 28.8.2003) |
CEN | EN ISO 10256:2003 Huvud- och ansiktsskydd för ishockeyspelare (ISO 10256:2003) | 6.10.2005 | EN 967:1996 | Datum passerat ( 6.10.2005) |
CEN | EN ISO 10819:1996 Vibration och stöt – Hand-armvibrationer – Metod att mäta och bedöma vibrationsöverföring hos handskar till handflatan (ISO 10819:1996) | 3.12.1996 | — | |
CEN | EN 12083:1998 Andningsskydd – Filter ej monterade på mask – Partikelfilter, gasfilter och kombinerade filter – Fordringar, provning, märkning | 4.7.2000 | — | |
EN 12083:1998/AC:2000 | | | |
CEN | EN 12270:1998 Klätterutrustning – Kilar – Säkerhetskrav och provningsmetoder | 16.3.2000 | — | |
CEN | EN 12275:1998 Klätterutrustning – Kabinhakar – Säkerhetskrav och provningsmetoder | 16.3.2000 | — | |
CEN | EN 12276:1998 Klätterutrustning – Fläns – Säkerhetskrav och provningsmetoder | 24.2.2001 | — | |
EN 12276:1998/AC:2000 | | | |
CEN | EN 12277:1998 Klätterutrustning – Säkerhetsselar – Säkerhetskrav och provningsmetoder | 6.11.1998 | — | |
CEN | EN 12278:1998 Klätterutrustning – Block – Säkerhetskrav och provningsmetoder | 6.11.1998 | — | |
CEN | EN 12477:2001 Skyddshandskar för svetsare | 10.8.2002 | — | |
EN 12477:2001/A1:2005 | 6.10.2005 | Anmärkning 3 | Datum passerat ( 31.12.2005) |
CEN | EN 12492:2000 Klätterutrustning – Klätterhjälmar – Säkerhetskrav och provningsmetoder | 21.12.2001 | — | |
EN 12492:2000/A1:2002 | 28.8.2003 | Anmärkning 3 | Datum passerat ( 28.8.2003) |
CEN | EN 12568:1998 Fot- och benskydd – Fordringar och provningsmetoder för skyddståhättor samt spiktrampsskydd av metall | 6.11.1998 | — | |
CEN | EN 12628:1999 Dykutrustning – Kombinerade flyt- och räddningsanordningar – Funktions- och säkerhetskrav, provningsmetoder | 4.7.2000 | — | |
EN 12628:1999/AC:2000 | | | |
CEN | EN 12941:1998 Andningsskydd – Fläktassisterade filterskydd med hjälp eller huva – Fordringar, provning, märkning | 4.6.1999 | EN 146:1991 | Datum passerat ( 4.6.1999) |
EN 12941:1998/A1:2003 | 6.10.2005 | Anmärkning 3 | Datum passerat ( 6.10.2005) |
CEN | EN 12942:1998 Andningsskydd – Fläktassisterade filterskydd med helmasker, halvmasker eller kvartsmasker – Fordringar, provning, märkning | 4.6.1999 | EN 147:1991 | Datum passerat ( 4.6.1999) |
EN 12942:1998/A1:2002 | 28.8.2003 | Anmärkning 3 | Datum passerat ( 28.8.2003) |
CEN | EN 13034:2005 Skyddskläder för kemikalier i vätskeform – Funktionskrav för kemisk skyddsdräkt med begränsad skyddsfunktion mot kemikalier i vätskeform (typ 6 utrustning) | 6.10.2005 | — | |
CEN | EN 13061:2001 Skyddskläder – Benskydd för fotbollsspelare – Fordringar och provningsmetoder | 10.8.2002 | — | |
CEN | EN 13087-1:2000 Skyddshjälmar – Provningsmetoder – Del 1: Provningsbetingelser och konditionering | 10.8.2002 | — | |
EN 13087-1:2000/A1:2001 | 10.8.2002 | Anmärkning 3 | Datum passerat ( 10.8.2002) |
CEN | EN 13087-2:2000 Skyddshjälmar – Provningsmetoder – Del 2: Stötdämpande förmåga | 10.8.2002 | — | |
EN 13087-2:2000/A1:2001 | 10.8.2002 | Anmärkning 3 | Datum passerat ( 10.8.2002 |
CEN | EN 13087-3:2000 Skyddshjälmar – Provningsmetoder – Del 3: Motstånd mot penetration | 10.8.2002 | — | |
EN 13087-3:2000/A1:2001 | 10.8.2002 | Anmärkning 3 | Datum passerat ( 10.8.2002) |
CEN | EN 13087-4:2000 Skyddshjälmar – Provningsmetoder – Del 4: Fastspänningens effektivitet | 21.12.2001 | — | |
CEN | EN 13087-5:2000 Skyddshjälmar – Provningsmetoder – Del 5: Hakbandets hållfasthet | 24.2.2001 | — | |
CEN | EN 13087-6:2000 Skyddshjälmar – Provningsmetoder – Del 6: Synfält | 10.8.2002 | — | |
EN 13087-6:2000/A1:2001 | 10.8.2002 | Anmärkning 3 | Datum passerat ( 10.8.2002) |
CEN | EN 13087-7:2000 Skyddshjälmar – Provningsmetoder – Del 7: Flamhärdighet | 10.8.2002 | — | |
EN 13087-7:2000/A1:2001 | 10.8.2002 | Anmärkning 3 | Datum passerat ( 10.8.2002) |
CEN | EN 13087-8:2000 Skyddshjälmar – Provningsmetoder – Del 8: Elektriska egenskaper | 21.12.2001 | — | |
EN 13087-8:2000/A1:2005 | 6.10.2005 | Anmärkning 3 | Datum passerat ( 6.10.2005) |
CEN | EN 13087-10:2000 Skyddshjälmar – Provningsmetoder – Del 10: Motstånd mot strålningsvärme | 21.12.2001 | — | |
CEN | EN 13138-1:2003 Flythjälpmedel för att lära sig simma – Del 1: Flythjälpmedel att ha på sig – Säkerhetskrav och provningsmetoder | 6.10.2005 | — | |
CEN | EN 13158:2000 Skyddsutrustning – Skyddsjacka, kropps- och axelskydd för ryttare – Krav och provningsmetoder | 24.2.2001 | — | |
CEN | EN 13178:2000 Ögonskydd – Ögon- och ansiktsskydd för snöskoteråkare | 21.12.2001 | — | |
CEN | EN 13274-1:2001 Andningsskydd – Testmetoder – Del 1: Bestämning av inläckage och totalt inläckage | 21.12.2001 | — | |
CEN | EN 13274-2:2001 Andningsskydd – Testmetoder – Del 2: Praktisk provning | 21.12.2001 | — | |
CEN | EN 13274-3:2001 Andningsskydd – Testmetoder – Del 3: Bestämning av andningsmotstånd | 10.8.2002 | — | |
CEN | EN 13274-4:2001 Andningsskydd – Testmetoder – Del 4: Flamtester | 10.8.2002 | — | |
CEN | EN 13274-5:2001 Andningsskydd – Testmetoder – Del 5: Klimatvillkor | 21.12.2001 | — | |
CEN | EN 13274-6:2001 Andningsskydd – Testmetoder – Del 6: Bestämning av koldioxidhalten i inandningsluft | 10.8.2002 | — | |
CEN | EN 13274-7:2002 Andningsskydd – Testmetoder – Del 7: Bestämning av aerosolpenetration genom partikelfilter | 28.8.2003 | — | |
CEN | EN 13274-8:2002 Andningsskydd – Testmetoder – Del 8: Bestämning av igensättning med damm på partikelfilter | 28.8.2003 | — | |
CEN | EN 13277-1:2000 Skyddsutrustning för kampsporter – Del 1: Allmänna krav och provningsmetoder | 24.2.2001 | — | |
CEN | EN 13277-2:2000 Skyddsutrustning för kampsporter – Del 2: Tilläggskrav och provningsmetoder för vrist-, knä- och underarmsskydd | 24.2.2001 | — | |
CEN | EN 13277-3:2000 Skyddsutrustning för kampsporter – Del 3: Tilläggskrav och provningsmetoder för bålskydd | 24.2.2001 | — | |
CEN | EN 13277-4:2001 Skyddsutrustning för kampsporter – Del 4: Tilläggskrav och provningsmetoder för huvudskydd | 10.8.2002 | — | |
CEN | EN 13277-5:2002 Skyddsutrustning för kampsporter – Del 5: Tilläggskrav och provningsmetoder för genital- och kroppsskydd | 10.8.2002 | — | |
CEN | EN 13277-6:2003 Personlig skyddsutrustning för kampsporter – Del 6: Tilläggskrav och provningsmetoder för bröstskydd för kvinnor | 21.2.2004 | — | |
CEN | EN 13287:2004 Personlig skyddsutrustning – Skodon – Provningsmetod för bestämning av halkskydd | 6.10.2005 | — | |
CEN | EN 13356:2001 Personreflexer med god synbarhet för icke yrkesmässigt bruk – Provningsmetoder och fordringar | 21.12.2001 | — | |
CEN | EN 13484:2001 Rodelhjälmar | 10.8.2002 | — | |
CEN | EN 13546:2002 Krav och testmetoder för hand-, arm-, bröst-, buk-, ben-, fot- och underlivsskydd för landhockeymålvakter samt benskydd för utespelare | 28.8.2003 | — | |
CEN | EN 13567:2002 Kroppsskydd – Hand-, arm-, buk-, ben-, underlivs- och ansiktsskydd för fäktare – Fordringar och testmetoder | 28.8.2003 | — | | CEN | EN 13594:2002 Krav och testmetoder på skyddsutrustning och dess beständighet mot mekanisk påverkan för professionella motorcyklister – Skyddshandskar | 28.8.2003 | — | |
CEN | EN 13595-1:2002 Skyddskläder för professionella motorcyklister – Jacka, byxor och hel eller delad dräkt – Del 1: Allmänna krav | 28.8.2003 | — | |
CEN | EN 13595-2:2002 Skyddskläder för professionella motorcyklister – Jacka, byxor och hel eller delad dräkt – Del 2: Provningsmetoder för slitmotstånd | 28.8.2003 | — | |
CEN | EN 13595-3:2002 Skyddskläder för professionella motorcyklister – Jacka, byxor och hel eller delad dräkt – Del 3: Provningsmetoder för bestämning av sprickmotstånd | 28.8.2003 | — | |
CEN | EN 13595-4:2002 Skyddskläder för professionella motorcyklister – Jacka, byxor och hel eller delad dräkt – Del 4: Provningsmetoder för skärmotstånd | 28.8.2003 | — | |
CEN | EN 13634:2002 Krav och testmetoder för fotskydd för professionella motorcyklister | 28.8.2003 | — | |
CEN | EN 13781:2001 Skyddshjälmar för passagerare och förare av terrängskotrar och bobsleighs | 10.8.2002 | — | |
CEN | EN 13794:2002 Andningsskydd – Bärbar flyktapparat med slutet system – Fordringar, provning, märkning | 28.8.2003 | EN 1061:1996 EN 400:1993 EN 401:1993 | Datum passerat ( 28.8.2003) |
CEN | EN 13819-1:2002 Hörselskydd – Provning – Del 1: Fysikaliska provningsmetoder | 28.8.2003 | — | |
CEN | EN 13819-2:2002 Hörselskydd – Provning – Del 2: Akustiska provningsmetoder | 28.8.2003 | — | |
CEN | EN 13911:2004 Skyddskläder för brandmän – Fordringar och provningsmetoder för huvor för brandmän | 6.10.2005 | — | |
CEN | EN 13949:2003 Andningsskydd – Bärbar Nitroxapparat med öppet system för dykning – Fordringar, provning, märkning | 21.2.2004 | — | |
CEN | EN ISO 13982-1:2004 Skyddskläder för användning mot fasta partiklar – Del 1: Fodringar på prestanda för skyddskläder mot kemikalier som ger skydd för hela kroppen mot luftburna fasta partiklar (Skyddskläder Typ 5) (ISO 13982-1:2004) | 6.10.2005 | — | |
CEN | EN ISO 13982-2:2004 Skyddskläder för användning mot fasta partiklar – Del 2: Provningsmetod för bestämning av inläckage i dräkter av aerosoler av fina partiklar (ISO 13982-2:2004) | 6.10.2005 | — | |
CEN | EN ISO 13995:2000 Skyddskläder – Mekaniska egenskaper – Provningsmetod för bestämning av motstånd mot punktering och dynamisk rivstyrka hos material (ISO 13995:2000) | 6.10.2005 | — | |
CEN | EN ISO 13997:1999 Skyddskläder – Mekaniska egenskaper – Bestämning av motstånd mot skärning med vassa föremål (ISO 13997:1999) | 4.7.2000 | — | |
EN ISO 13997:1999/AC:2000 | | | |
CEN | EN ISO 13998:2003 Skyddskläder – Förkläden, byxor och västar till skydd mot skär och stick av handhållna knivar (ISO 13998:2003) | 28.8.2003 | EN 412:1993 | Datum passerat ( 28.8.2003) |
CEN | EN 14021:2003 Förarskydd mot stensprut vid motorcykelåkning i terräng – Krav och provningsmetoder | 6.10.2005 | — | |
CEN | EN 14052:2005 Industrihjälmar med hög skyddsförmåga | Detta är det första offentliggörandet | — | |
CEN | EN 14058:2004 Skyddskläder – Plagg till skydd i kalla miljöer | 6.10.2005 | — | |
CEN | EN 14120:2003 Kroppsskydd – Handleds-, hand-, knä- och armbågsskydd för rullskridskoåkare – Krav och provningsmetoder | 21.2.2004 | — | |
CEN | EN 14126:2003 Skyddskläder – Funktionskrav och provningsmetoder för skyddskläder mot smittsamma ämnen | 6.10.2005 | — | |
CEN | EN 14143:2003 Andningsskydd – Bärbar andningsapparat för dykning med slutet/halvslutet gasregleringssystem | 6.10.2005 | — | |
CEN | EN 14225-1:2005 Dykardräkter – Del 1: Våtdräkter – Krav och provningsmetoder | 6.10.2005 | — | |
CEN | EN 14225-2:2005 Dykardräkter – Del 2: Torrdräkter – Krav och provningsmetoder | 6.10.2005 | — | |
CEN | EN 14225-3:2005 Dykardräkter – Del 3: Aktivt uppvärmda eller kylda dräkter – Krav och provningsmetoder | 6.10.2005 | — | |
CEN | EN 14225-4:2005 Dykardräkter – Del 4: Enatmosfärsdräkter – Fordringar och provningsmetoder | 6.10.2005 | — | |
CEN | EN 14325:2004 Skyddskläder mot kemikalier – Provningsmetoder och klassificering av egenskaper hos material, sömmar, skarvar och förbindningar hos skyddskläder mot kemikalier | 6.10.2005 | — | |
CEN | EN 14328:2005 Skyddskläder – Handskar och armskydd till skydd mot maskindrivna knivar – Krav och provningsmetoder | 6.10.2005 | — | |
CEN | EN 14360:2004 Skyddskläder mot dåligt väder – Provningsmetod för regntäthet hos beklädnader – Påverken av högt fallande regndroppar | 6.10.2005 | — | |
CEN | EN 14387:2004 Andningsskydd – Gasfilter och kombinationsfilter – Fordringar, provning, märkning | 6.10.2005 | EN 141:2000 EN 371:1992 EN 372:1992 | Datum passerat ( 6.10.2005) |
CEN | EN 14404:2004 Skyddskläder – Knäskydd för arbete i knästående ställning | 6.10.2005 | — | |
CEN | EN 14435:2004 Andningsskydd – Bärbar tryckluftsapparat med öppet system och halvmask – Fordringar, provning, märkning | 6.10.2005 | — | |
CEN | EN 14458:2004 Ögonskydd – Ansiktsskärmar och visir på skyddshjälm för användning av personal inom räddnings- och ambulanstjänst | 6.10.2005 | — | |
CEN | EN ISO 14460:1999 Skyddskläder för förare av tävlingsbilar – Skydd mot hetta och flamma – Funktionskrav och provningsmetoder (ISO 14460:1999) | 16.3.2000 | — | |
EN ISO 14460:1999/A1:2002 | 10.8.2002 | Anmärkning 3 | Datum passerat ( 30.9.2002) |
EN ISO 14460:1999/AC:1999 | | | |
CEN | EN 14529:2005 Andninsskydd – Bärbar tryckluftsapparat med öppet system för halvmask inkluderande överstrycksventil avsedd enbart för flykt – Fordringar, provning, märkning | Detta är det första offentliggörandet | — | |
CEN | EN 14572:2005 Stötskyddsmössor | 6.10.2005 | — | |
CEN | EN 14593-1:2005 Andningsskydd – Tryckluftsapparat med behovsstyrt flöde – Del 1: Apparat med helmask – Fordringar, provning, märkning | 6.10.2005 | EN 139:1994 | Datum passerat ( 2.12.2005) |
CEN | EN 14593-2:2005 Andningsskydd – Tryckluftsapparat med behovsstyrt flöde – Del 2: Apparat med halvmask med övertryck – Fordringar, provning, märkning | 6.10.2005 | EN 139:1994 | Datum passerat ( 2.12.2005) |
EN 14593-2:2005/AC:2005 | | | |
CEN | EN 14594:2005 Andningsskydd – Tryckluftsapparat med kontinuerligt flöde – Fordringar, provning, märkning | 6.10.2005 | EN 271:1995 EN 12419:1999 EN 139:1994 EN 1835:1999 EN 270:1994 | Datum passerat ( 2.12.2005) |
EN 14594:2005/AC:2005 | | | |
CEN | EN 14605:2005 Skyddskläder mot kemikalier i vätskeform – Funktionskrav för skyddskläder mot kemikalier, med vätsketäta (typ 3) eller stänktäta (typ 4) anslutningar mellan olika delar av beklädnanden samt beklädnad begränsad till delar av kroppen | 6.10.2005 | EN 467:1995 EN 466:1995 EN 465:1995 | Datum passerat ( 6.10.2005) |
CEN | EN ISO 14877:2002 Skyddskläder vid blästring med kornigt slipmedel (ISO 14877:2002) | 28.8.2003 | — | |
CEN | EN ISO 15025:2002 Skyddskläder – Skydd mot hetta och flamma – Provningsmetod för begränsad flamspridning (ISO 15025:2000) | 28.8.2003 | EN 532:1994 | Datum passerat ( 28.8.2003) |
CEN | EN ISO 15027-1:2002 Sjöräddningsdräkter – Del 1: Räddningsdräkter för arbete, fordringar för säkerhet (ISO 15027-1:2002) | 10.4.2003 | — | |
CEN | EN ISO 15027-2:2002 Sjöräddningsdräkter – Del 2: Räddningsdräkter för nödläge, fordringar för säkerhet (ISO 15027-2:2002) | 10.4.2003 | — | |
CEN | EN ISO 15027-3:2002 Sjöräddningsdräkter – Del 3: Provningsmetoder (ISO 15027-3:2002) | 10.4.2003 | — | |
CEN | EN ISO 15831:2004 Beklädnad – Fysiologisk inverkan – Mätning av värmeisolering med hjälp av en termisk docka (ISO 15831:2004) | 6.10.2005 | — | |
CEN | EN ISO 17249:2004 Skyddsskor till skydd mot kedjesåg (ISO 17249:2004) | 6.10.2005 | — | |
CEN | EN ISO 20344:2004 Personlig skyddsutrustning – Provningsmetoder för skodon (ISO 20344:2004) | 6.10.2005 | EN 344:1992 EN 344-2:1996 | Datum passerat ( 6.10.2005) |
CEN | EN ISO 20345:2004 Personlig skyddsutrustning – Skyddsskor (ISO 20345:2004) | 6.10.2005 | EN 345:1992 EN 345-2:1996 | Datum passerat ( 6.10.2005) |
CEN | EN ISO 20346:2004 Personlig skyddsutrustning – Lätta skyddsskor (ISO 20346:2004) | 6.10.2005 | EN 346-2:1996 EN 346:1992 | Datum passerat ( 6.10.2005) |
CEN | EN ISO 20347:2004 Personlig skyddsutrustning – Yrkesskor (ISO 20347:2004) | 6.10.2005 | EN 347:1992 EN 347-2:1996 | Datum passerat ( 6.10.2005) |
CEN | EN 24869-1:1992 Akustik – Hörselskydd – Del 1: Subjektiv metod för mätning av ljuddämpning (ISO 4869-1:1990) | 16.12.1994 | — | |
CEN | EN 24869-3:1993 Akustik – Hörselskydd – Del 3: Förenklad metod för mätning av ljuddämpning (ISO/TR 4869-3:1989) | 16.12.1994 | — | |
CENELEC | EN 50237:1997 Arbete med spänning – Isolerande handskar med skydd mot yttre påverkan | 4.6.1999 | — | |
CENELEC | EN 50286:1999 Elektriskt isolerande skyddskläder för lågspänning | 16.3.2000 | — | |
CENELEC | EN 50321:1999 Elektriskt isolerande fotbeklädnad för användning i lågspänningsanläggningar | 16.3.2000 | — | |
CENELEC | EN 50365:2002 Elektriskt isolerande hjälmar för användning i lågspänningsinstallationer | 10.4.2003 | — | |
CENELEC | EN 60743:2001 Arbete med spänning – Terminologi (IEC 60743:2001) | 10.4.2003 | EN 60743:1996 Anmärkning 2.1 | Datum passerat ( 1.12.2004) |
CENELEC | EN 60895:2003 Arbete med spänning – Elektriskt ledande kläder (IEC 60895:2002 (Ändrad)) | 6.10.2005 | EN 60895:1996 Anmärkning 2.1 | 1.7.2006 |
CENELEC | EN 60903:2003 Utrustning för arbete under spänning – Isolerande handskar (IEC 60903:2002 (Ändrad)) | 6.10.2005 | EN 60903:1992 och dess tillägg + EN 50237:1997 Anmärkning 2.1 | 1.7.2006 |
CENELEC | EN 60984:1992 Utrustning för arbete under spänning – Isolerande armskydd (IEC 60984:1990 (Ändrad)) | 4.6.1999 | — | |
EN 60984:1992/A1:2002 (IEC 60984:1990/A1:2002) | 10.4.2003 | Anmärkning 3 | Datum passerat ( 6.10.2005) |
EN 60984:1992/A11:1997 | 4.6.1999 | Anmärkning 3 | Datum passerat ( 4.6.1999) |
Anmärkning 1 Det datum då den ersatta standarden upphör att gälla är i allmänhet det datum då den upphävs av det europeiska standardiseringsorganet. Användare av dessa standarder bör dock vara medvetna om att det i vissa undantagsfall kan vara ett annat datum.
Anmärkning 2.1 Den nya (eller ändrade) standarden har samma tillämpningsområde som den standard den ersätter. Vid angivet datum upphör den ersatta standarden att ge presumtion om överensstämmelse med de väsentliga kraven i direktivet.
Anmärkning 3 Om tillägg förekommer innefattar hänvisningen såväl standarden EN CCCCC:YYYY som eventuella tidigare tillägg och det nya, angivna, tillägget. Den ersatta standarden (kolumn 3) består därför av EN CCCCC:YYYY med eventuella tidigare tillägg, men utan det nya, angivna, tillägget. Vid angivet datum upphör den ersatta standarden att gälla.
Anmärkning 4 BHSR 1.2.1.1 får förutsättas överensstämma med EN 420:2003 när det gäller halten av Cr(VI) i handskmaterialen, så länge som provningsmetodens detektionsgräns för Cr(VI) är 3 mg/kg eller lägre.
ANMÄRKNING:
- Närmare upplysningar om standarderna kan erhållas från de europeiska och nationella standardiseringsorgan som anges i bilagan till Europaparlamentets och rådets direktiv 98/34/EG [2], ändrat genom direktiv 98/48/EG [3].
- Offentliggörandet av hänvisningarna i Europeiska unionens officiella tidning innebär inte att de aktuella standarderna är tillgängliga på alla gemenskapsspråken.
- Denna förteckning ersätter alla tidigare förteckningar som har publicerats i Europeiska unionens officiella tidning. Kommissionen skall fortlöpande uppdatera denna förteckning.
Mer information återfinns på Europa-servern på Internet:
http://europa.eu.int/comm/enterprise/newapproach/standardization/harmstds/
[1] ESO: Europeiskt standardiseringsorgan:
- CEN: rue de Stassart 36, B-1050 Bryssel, Tfn (32-2) 550 08 11; fax (32-2) 550 08 19 (http://www.cenorm.be)
- CENELEC: rue de Stassart 35, B-1050 Bryssel, Tfn (32-2) 519 68 71; fax (32-2) 519 69 19 (http://www.cenelec.org)
- ETSI: 650, route des Lucioles, F-06921 Sophia Antipolis, Tfn (33) 492 94 42 00; fax (33) 493 65 47 16 (http://www.etsi.org)
[2] EGT L 204, 21.7.1998, s. 37
[3] EGT L 217, 5.8.1998, s. 18.
--------------------------------------------------
Statligt stöd – Belgien
Statligt stöd C 46/2005 (f.d. NN 9/2004 %amp% N 55/2005) – Inter Ferry Boats
(Text av betydelse för EES)
(2006/C 159/02)
Uppmaning enligt artikel 88.2 i EG-fördraget att inkomma med synpunkter
Genom den skrivelse av den 7 december 2005 som återges på det giltiga språket på de sidor som följer på denna sammanfattning, underrättade kommissionen Belgien om sitt beslut att inleda det förfarande som anges i artikel 88.2 i EG-fördraget avseende ovannämnda stöd.
Kommissionen uppmanar berörda parter att inom en månad från dagen för detta offentliggörande inkomma med sina synpunkter på stödet/åtgärderna i fråga. Synpunkterna skall sändas till följande adress:
Europeiska gemenskapernas kommission
Generaldirektoratet för energi och transport
Direktorat A – Allmänna frågor och resursförvaltning
DM 28, kontor 6/100
B-1049 Bryssel
Fax: (32-2) 296 41 04
Synpunkterna kommer att meddelas Belgien. Den berörda part som inkommer med synpunkter kan skriftligen begära konfidentiell behandling av sin identitet, med angivande av skälen för begäran.
SAMMANFATTNING
1. FÖRFARANDE
Ej anmält ärende.
2. BESKRIVNING AV DEN ÅTGÄRD AVSEENDE VILKEN KOMMISSIONEN INLEDER FÖRFARANDET
nationell rättslig grund : beslut i SNCB:s styrelse.
myndighet i medlemsstaten som beviljar stödet : Société nationale des chemins de fer belge (SNCB)
stödform : Beviljande av en tidsfrist för betalning av 63 miljoner euro, beviljande av ett förskott som kan återkrävas på 5 miljoner euro, beviljande av en kredit på 15 miljoner euro för kapitalökning, en ytterligare kapitalökning på 5 miljoner euro i form av andelar i företaget TRW.
varaktighet : ej fastställd
mottagare : Société InterFerryBoats SA
syfte/ändamål : Stöd till omstrukturering
budget, ursprung för de medel som används för finansiering av stödet samt stödbeloppet (per år) : Beviljande av en tidsfrist för betalning av 63 miljoner euro, beviljande av ett förskott som kan återkrävas på 5 miljoner euro, beviljande av en kredit på 15 miljoner euro, omvandling till en nettofordran av 63 miljoner euro och ett lån på 15 miljoner euro för kapitalökning, en ytterligare kapitalökning på 5 miljoner euro i form av andelar i företaget TRW.
3. BEDÖMNING AV ÅTGÄRDEN
SNCB:s beslut att bevilja företaget IFB ett omstruktureringsstöd fattades den 7 april 2003 och kan tillskrivas belgiska staten, eftersom meddelandet om omstruktureringsplanen som lämnats till belgiska staten och tidningsartiklar låter förstå att belgiska staten påverkat SNCB:s beslut. Å andra sidan tvivlar kommissionen på att det tysta medgivandet att skjuta upp SNCB:s betalningar till IFB mellan 2001och den 19 september 2002 kan tillskrivas staten.
SNCB agerade inte som en fordringsägare (när det gällde tidsfristen för betalningarna) eller en investerare som kände till marknaden (när det gäller övriga åtgärder), och räntan på det investerade kapitalet ligger under den som skulle ha kunnat godtas av en sådan investerare.
Likviditetsstöden kan inte deklareras som undsättningsstöd eftersom varaktigheten är längre än tolv månader.
För att stöden skall kunna anses förenliga med den gemensamma marknaden i egenskap av omstruktureringsstöd, skall företaget vara stödberättigande i enlighet med riktlinjerna för omstruktureringar och stödet skall uppfylla fem villkor:
(1) Omstruktureringsplanen skall göra det möjligt att inom en rimlig tid återge företaget dess ekonomiska hållbarhet på lång sikt.
(2) Åtgärder bör vidtas för att i möjligaste mån motverka negativa effekter som stödet får för konkurrenterna.
(3) Stödet bör begränsas till det absoluta minimum som krävs för att möjliggöra omstruktureringen och företaget skall själv bidra till omstruktureringen.
(4) Kommissionen skall ges möjlighet att konstatera att omstruktureringen förlöper väl i form av regelbundna och detaljerade rapporter.
(5) Stöd till omstrukturering skall inte beviljas mer än en gång.
Kommissionen kan i det här skedet inte utesluta att företaget IFB fick en del av stödet mindre än tre år efter att företaget startades. Kommissionen uttrycker därför sina tvivel på att IFB är ett företag som kan berättiga till omstruktureringsstöd.
Kommissionens granskning visade att villkoren 1, 4 och 5 är uppfyllda. Å andra sidan hyser kommissionen tvivel om att de åtgärder som har vidtagits för i möjligaste mån motverka negativa effekter som stödet får för konkurrenterna är tillräckliga, och om IFB:s eget bidrag är tillräckligt.
När det gäller att motverka negativa effekter för konkurrenterna: De belgiska myndigheterna förklarar att IFB vidtog två åtgärder för att i möjligaste mån motverka negativa effekter som stödet får för konkurrenterna:
- De upphörde med sin verksamhet i Frankrike
- De stängde terminalen i Bressoux i Belgien och sålde aktierna i terminalerna i Bryssel och Zeebrugge i Belgien.
Dessa två åtgärder innebar att man sänkte omsättningen från 62 miljoner euro 2002 till 58 miljoner euro 2003. Eftersom det emellertid rör sig om insatser som inriktades på icke vinstgivande delar av verksamheten ställer sig kommissionen tveksam till om den kan beakta åtgärderna.
För att ta reda på om dessa två åtgärder var tillräckliga för att i möjligaste mån motverka negativa effekter som stödet får för konkurrenterna är det lämpligt att erinra om de viktigaste aspekterna av utvecklingen på de två marknader där IFB är aktivt, nämligen logistikmarknaden och lossning och lastning av varor. Vidare är det lämpligt att analysera om de åtgärder som har föreslagit verkligen i möjligaste mån motverkar negativa effekter som stödet får för konkurrenterna.
a) Marknaden för logistik och stödet till IFB
Marknaden för logistik genomgår för närvarande en djupgående förändring på grund av att marknaden för järnvägstransporter har öppnats och järnvägs- och postföretag har kommit in på marknaden, med ett stort antal mindre aktörer och flera stora, specialiserade företag med integrerade tjänster.
Kommissionen noterar att de åtgärder som har föreslagits inte rör marknaden för logistik. IFB:s andel av den marknaden ökade avsevärt under 2004 i jämförelse med 2003. Belgien har inte lagt fram något som helst åtagande, inte ens tillfälligt, som skulle begränsa IFB:s insatser på den marknaden.
Kommissionen anser att avsaknaden av förslag till åtgärder på logistikmarknaden, liksom det faktum att marknaden håller på att förändras och att IFB har ökat sin omsättning avsevärt leder till tvivel på om Belgien i möjligaste mån har motverkat negativa effekter som stödet får för konkurrenterna när det gäller IFB:s logistikverksamhet.
b) Marknaden för lossning och lastning av varor och stödet till IFB
De två åtgärder som har föreslagits gäller marknaden för lossning och lastning av varor. IFB har nästan helt upphört med verksamheten i Frankrike och har vidare stängt en terminal i Belgien och sålt sitt aktieinnehav i två andra terminaler.
Den enda marknad där detta kan få negativa konsekvenser på konkurrensen är alltså den belgiska. IFB har mindre än 7 % av denna.
För att begränsa de negativa effekter stödet kan få på den belgiska marknaden stängde IFB en terminal och sålde sitt aktieinnehav i två andra. Kommissionen noterar emellertid både att det var den minsta av terminalerna som stängdes och att stängningen främst var avsedd att minska IFB:s förluster, och att IFB efter kapitalökningen på nytt kommer att använda de två terminaler som det sålde, för företaget TRW, från vilket SNCB kommer att överföra 47 % av aktieinnehavet till IFB, har ett avsevärt aktieinnehav i terminalerna i Bruxelles och Zeebrugge.
Vidare utnyttjar TRW flera andra terminaler i Belgien. Följaktligen kommer kapitalökningen i form av aktieinnehav i TRW att innebära att IFB:s andel av den belgiska marknaden växer.
Vidare noterar kommissionen att IFB är minoritetsägare av aktierna i ett stort antal belgiska terminaler.
Följaktligen tvivlar kommissionen på att de åtgärder som IFB har föreslagit för att i möjligaste mån motverka negativa effekter som stödet får för konkurrenterna faktiskt är tillräckliga.
När det gäller IFB:s eget bidrag: Enligt den belgiska regeringens uppgifter tycks IFB inte ha bidragit med egna medel till omstruktureringen. Ett sådant bidrag krävs enligt riktlinjerna från 1999 och 2004. Kommissionen tvivlar följaktligen på att IFB:s eget bidrag är tillräckligt.
SJÄLVA SKRIVELSEN
"1. PROCÉDURE
1.1. Cas NN 9/2004
1. Par lettre du 12 août 2003, enregistrée à la Commission européenne le 20 août 2003 (TREN/A(03)27718), les autorités belges ont notifié certains accords entre la Société Nationale des Chemins de Fer Belges (SNCB) et sa filiale Inter Ferry Boats (IFB) au titre de l'article 88 paragraphe 3 du traité CE. D'après cette notification, il s'agit de mesures de sauvetage pour IFB de la part de la SNCB.
2. Le 13 octobre 2003 (D(03)17546), la Direction générale de l'énergie et des transports a invité les autorités belges à fournir à la Commission des renseignements complémentaires. Une réunion bilatérale à ce sujet avec les autorités belges a eu lieu le 12 décembre 2003. Lors de cette réunion, un plan de restructuration pour IFB, élaboré par McKinsey, a été présenté.
3. Les autorités belges ont répondu à la lettre de la Commission par courrier du 7 janvier 2004, enregistrée à la Commission le 13 janvier 2004 (TREN/A(04)10708). De ce courrier, il ressort que les mesures de sauvetage notifiées ont partiellement été mises en œuvre. Par conséquent, le cas a été enregistré sous le numéro NN 9/2004. Une deuxième réunion a eu lieu le 30 avril 2004. Les autorités belges ont envoyé des documents supplémentaires, demandés par la Commission lors de cette réunion, par lettre du 15 juin 2004, enregistrée à la Commission le 21 juin 2004 (TREN/A(04)23691).
4. Par lettre du 26 janvier 2005 (D(05)100339), la Direction générale de l'énergie et des transports a invité les autorités belges à fournir des renseignements complémentaires quant au développement de la société IFB, et notamment de sa restructuration.
5. Par lettre du 25 mars 2005, enregistrée à la Commission le 30 mars 2005 (TREN/A(05)7712), les autorités belges ont transmis à la Commission les renseignements complémentaires demandés par la lettre du 26 janvier 2005.
1.2. Cas N 55/2005
6. Par lettre du 28 janvier 2005 (SG(2005)A1133), les autorités belges ont notifié à la Commission l'intention de la SNCB de procéder à une augmentation de capital de la société IFB,. Les autorités belges considèrent que cela n'est pas une aide d'État, mais ont notifié cette intention pour des raisons de sécurité juridique. La Commission a enregistré ce cas comme un nouveau dossier "aide d'État notifié" sous le numéro N 55/2005.
7. Par lettre du 29 mars 2005 (D(05)106199), la Direction générale de l'énergie et des transports a invité les autorités belges à fournir des renseignements complémentaires quant aux mesures de restructuration de la société IFB.
8. Par lettre du 28 avril 2005, enregistrée à la Commission le 3 mai 2005 (SG(2005)A(05)4155), les autorités belges ont transmis à la Commission les renseignements complémentaires demandés par la lettre du 29 mars 2005.
9. Par lettre du 31 mai 2005 (D(05)111096), la Direction générale de l'énergie et des transports a invité les autorités belges à fournir des renseignements complémentaires quant aux informations transmises le 28 avril 2005.
10. Par lettre du 30 juin 2005, enregistrée à la Commission le 1 juillet 2005 (TREN/A(05)16598), les autorités belges ont transmis à la Commission les renseignements complémentaires demandés par la lettre du 31 mai 2005.
11. Le 16 septembre 2005, une réunion de travail a eu lieu entre la Commission et les autorités belges. Lors de cette réunion, la Commission a demandé aux autorités belges de transmettre des informations complémentaires. Par courriel du 21 octobre 2005, enregistré à la Commission le 24 octobre 2005 (TREN/A(05)27067), les autorités belges ont transmis ces informations.
2. DESCRIPTION DÉTAILLÉE DES MESURES DE SAUVETAGE ET DE RESTRUCTURATION
2.1. Les parties du contrat cadre concernant le sauvetage et la restructuration d'IFB
2.1.1. IFB
2.1.1.1. Description de la société
12. Inter Ferry Boats ("IFB") est une société anonyme de droit belge. La SNCB détient 89,03 % du capital social. Les autres actionnaires sont CNC Transports, une filiale à 93,8 % de la SNCF (7,41 %), ICF (2,08 %), et EWS (English Welsh and Scottish Railway — 1,22 %). IFB compte aujourd'hui 245 employés.
13. La société IFB a été créée le 1er avril 1998 par la fusion des trois sociétés suivantes: Ferry Boats Ltd., Interferry Ltd. et le département "rail" de Edmond Depaire Ltd. Avant la création d'IFB, Ferry Boats Ltd a été une entreprise contrôlée de manière conjointe par les chemins de fer britannique et les chemins de fer belge. Interferrry Ltd et Edmond Depaire Ltd ont été contrôlés par les chemins de fer belge. Il ne ressort pas clairement des documents fournis par la Belgique si IFB continue la personnalité juridique d'une des trois sociétés.
14. La société Ferry Boats Ltd. a été créée en 1923 sous le nom "Société Belgo-Anglaise des Ferry-Boats". La société Interferry a été créée en 1967 sous le nom d' "Intercontainer", et la société Edmond Depaire en 1906 comme une société privé de transport des containers.
15. IFB poursuit surtout deux types d'activités:
- Le secteur d'activité "IFB Logistics", qui commercialise les activités d'expédition d'IFB et;
- Le secteur d'activité "IFB Terminals", qui exploite des terminaux continentaux.
À ces activités, il faut ajouter les participations et filiales qu'IFB détient ou détenait en Belgique et à l'étranger.
a) L'activité IFB Logistics
16. L'activité "IFB Logistics" concerne la commercialisation par IFB, ainsi que par les sociétés dans lesquelles elle détient une participation, de:
- Activités d'expédition (y compris des services complémentaires de "transport engineering"), et
- Activités logistiques.
17. Les activités d'expédition sont les activités principales d'"IFB Logistics". Elles consistent à offrir aux clients des solutions de transport aussi complètes que possible. Pour les activités d'expédition, le transport ferroviaire, qu'il soit conventionnel ou combiné, représente pour IFB le mode de transport principal, mais IFB offre aussi le transport par voie navigable et le transport routier. Pour IFB, le transport ferroviaire est surtout un transport de "courte" ou de "moyenne" distance (de 100 à 500 km, avec IFB se présentant surtout comme partenaire des armateurs pour le développement du "carrier haulage", qui est une activité complémentaire à celle des opérateurs ferroviaires, qui se concentrent plutôt sur les transports de "longue distance").
18. Les marchandises expédiées par IFB sont des produits en vrac, des conteneurs et des produits divers (general cargo). Le tableau suivant montre le volume de fret transporté par IFB en 2003 et 2004 par rail conventionnel, rail intermodal et voies navigables. Le transport routier n'est utilisé par IFB que pour l'acheminement des unités de transport vers ou leur évacuation depuis des terminaux ferroviaires et ce uniquement dans les cas où le client a demandé une prestation porte-à-porte ou de/vers un terminal maritime.
19. Les principaux clients d'IFB Logistics sont les sociétés de fret maritime […] [1] [2] et […] ainsi que les sociétés […] [3], […], […] [4] et […]. Les produits transportés sont notamment des produits chimiques, le charbon, et les granulâts. Le tableau suivant montre les volumes transportés par IFB en 2003 et 2004.
Année | Rail conventionnel [5] | Rail intermodal | Voie navigable |
2003 | 0,672 millions de tonnes | 423583 TEU [6] | 0,385 millions de tonnes |
2004 | 1,995 millions de tonnes | 481556 TEU | 1,023 millions de tonnes |
20. Les activités d'expédition comprennent également des services complémentaires de "transport engineering", tels le stockage en magasin, la distribution, les transbordements,…, qui y sont intimement liés.
21. Dans le cadre de son système d'organisation, l'activité d'agence pour compte d'expéditeurs/transporteurs ferroviaires tiers est également rattachée à IFB Logistics. IFB est active en tant qu'agent logistique en Belgique pour un certain nombre d'entreprises étrangères.
22. Le marché de l'expédition et des activités logistiques a connu une croissance importante pendant les dernières années, qui est liée à la globalisation croissante de l'industrie, la tendance vers la sous-traitance et une spécialisation de plus en plus poussée des entreprises de production (just in time production).
23. Les barrières à l'entrée sur le marché sont réduites, et le marché connaît à la fois la présence d'un nombre importants de petits acteurs spécialisés et de grands acteurs intégrés (DHL, UPS, …). Suite à l'ouverture des marchés du transport ferroviaire et des services postaux, des entreprises ferroviaires (Deutsche Bahn, SNCB) et des entreprises postales (Deutsche Post) ont fait leur entrée sur ce marché.
24. La combinaison de la croissance du marché, de l'entrée de nouveaux acteurs importants et de la libéralisation du transport ferroviaire fait de ce marché un marché en pleine mutation et mouvement.
b) IFB Terminals
25. IFB Terminals exploite des terminaux ferroviaires (transbordement d'Unités de Transport Intermodal (UTI) du/vers le chemin de fer) continentaux.
26. L'activité principale des terminaux continentaux ("dry ports") concerne le chargement de conteneurs maritimes de camions sur des wagons. Au total, IFB exploite six terminaux continentaux avec connexion au réseau ferroviaire en Belgique, dont quatre sont situés dans le port d'Anvers et trois autres à l'intérieur de la Belgique.
27. Les terminaux continentaux dans le port d'Anvers sont "Mainhub", "Cirkeldyck", "Zomerweg" et "Schijnpoort". Le gouvernement belge souligne que ces quatre terminaux se trouvent dans une situation spécifique, car ils sont situés au port d'Anvers, au cœur même de l'activité maritime à laquelle ils sont indissociablement liés. Les UTI traités dans ces terminaux sont principalement des conteneurs maritimes qui sont d'abord déchargés des navires vers des camions dans un terminal maritime, qui n'est pas exploité par IFB. Ce n'est que par la suite que ces conteneurs sont déchargés des camions vers des wagons de chemin de fer dans un terminal continental exploité par IFB. Pour l'exportation maritime, l'ordre inverse est suivi. En 2004, les quatre terminaux continentaux d'IFB situés dans le port d'Anvers ont traité un volume de 0,4 millions TEU.
28. IFB exploite deux terminaux continentaux qui ne sont pas situés dans le port d'Anvers, à savoir le terminal de Muizen (situé près de Malines, terminal route-rail) et le terminal de Rénory (situé près de Liège, trafic route-rail-barge). Un troisième terminal, celui de Bressoux, a été fermé en 2003.
29. Le marché des terminaux est un marché plus stable que le marché de la logistique. Le nombre des terminaux exploités en Belgique reste constant. Cependant, le nombre de containeurs transportés est en augmentation, suite à la croissance de trafic dans le port d'Anvers et aux efforts de transporter d'avantage de biens par le transport combiné.
c) Les participations d'IFB
30. IFB détient ou détenait des participations dans des sociétés exploitant des terminaux maritimes et continentaux ainsi que dans des sociétés de transport. Au total, IFB détient ou détenait une trentaine de participations.
31. Participations dans les terminaux maritimes et continentaux à Dunkerque. IFB a réalisé des investissements importants dans le port de Dunkerque, où elle détenait des participations majoritaires dans Acimar (terminal pour produits d'acier, filiale à 100 % de NFTI-ou), NFTI-ou (terminal de conteneurs maritimes, participation de 60 % en 2003, réduite à 30 % depuis), Dry Port Dunkerque (DPD, un terminal ferroviaire, participation de 90 % restée inchangée depuis 2003), Short Sea Terminal Dunkirk (SSTD, chargement et déchargement de semi-remorques, participation de 50 % en 2003, réduite à 0 % depuis), et IFB France (société de holding et de services aux sociétés liées sises à Dunkerque, participation de 100 %, vendue entièrement à NFTI-ou depuis).
32. IFB France a été renommée Administration Gestion Entreprise Portuaires (AGEP). IFB a cédé la totalité de ses parts dans cette société à la société NFTI-ou.
33. En décembre 2002, une procédure de redressement judiciaire a été entamée concernant Acimar. Acimar n'exerce plus d'activités depuis le 1er septembre 2003. La totalité des actions qu'IFB possédait dans Acimar a été cédée à AGEP (voir ci-dessous).
34. IFB a réduit sa participation dans NFTI-ou, qui détient AGEP et, via AGEP, Acimar, de 60 % à 30 %. IFB a révoqué tout patronage de NFTI-ou, en dénonçant sa lettre de confort. Ainsi, IFB s'est libérée de toute obligation de se porter garante pour NFTI-ou, cette obligation étant reportée intégralement sur l'actionnaire majoritaire, le Port Autonome de Dunkerque, qui détient 70 % des parts de NFTI-ou. IFB cherche maintenant à se défaire de sa participation minoritaire dans NFTI-ou.
35. IFB avait une participation de 90 % dans DPD. En juin 2003, IFB a dénoncé sa lettre de confort; ensuite, IFB a vendu les infrastructures et des équipements de DPD au Port Autonome de Dunkerque et dissout la société DPD en juin 2004. La liquidation s'est terminée à l'été 2005.
36. IFB a vendu sa participation dans SSTD en avril 2005.
37. En conclusion, IFB a vendu toutes ses participations dans le port de Dunkerque, à l'exception de sa participation minoritaire dans NFTI-ou, pour laquelle il est à la recherche d'un acquéreur.
38. Participation dans des terminaux en Belgique. En Belgique, IFB détenait des participations dans des terminaux à Zeebrugge, Bruxelles, Mouscron, Athus, Liège et Charleroi.
39. À Zeebrugge, IFB et Hesse-Noord Natie avaient créé le groupement d'intérêt économique OCHZ, dont IFB et Hesse-Noord Natie étaient les copropriétaires à 50 %. En septembre 2004, IFB s'est retiré de OCHZ et a vendu ses droits à OCHZ.
40. À Bruxelles, IFB possédait des intérêts dans un terminal à conteneurs tri-modal, situé dans le port de Bruxelles, par le biais des sociétés Brussels Port Invest (BPI) et Brussels Terminal Intermodal (BTI). BTI a entre-temps été dissoute et mise en liquidation. Quant à BPI, IFB a cédé sa participation à une autre société étrangère au groupe SNCB.
41. À Mouscron, IFB détient une participation de 16,76 % dans la SA Dryport Mouscron Lille (DPM Li). Cette société a des capitaux propres de 530000 EUR, et a réalisé en 2004 un résultat net de 76000 EUR.
42. À Athus, IFB détient une participation de 24,89 % dans la SA Terminal Athus (Terminal Athus). Cette société a des capitaux propres de 1,7 millions EUR, et a réalisé en 2002 un résultat net de 61000 EUR (pas de données plus récentes).
43. À Liège, IFB détient une participation de 45,12 % dans Liège Logistics Intermodal. La Commission ne dispose pas de plus d'informations sur cette participation.
44. À Charleroi, IFB détient une participation de 14,28 % dans la SA Charleroi Dry Port (Charleroi DP). Cette société a des capitaux propres de 36000 EUR, et a réalisé en 2002 un résultat net de 899 EUR (pas de données plus récentes).
45. En conclusion, IFB détient aujourd'hui des participations minoritaires dans quatre terminaux en Belgique, à savoir les terminaux Mouscron, Liège, Athus, Charleroi. En plus, IFB détient une participation dans la société qui exploite ces terminaux, qui est la société TRW, à la hauteur de 0,9 %. La SNCB détient dans TRW une participation directe de 47 %.
46. En revanche, IFB a vendu ses participations dans les terminaux de Zeebrugge et Bruxelles.
47. Participations dans des entreprises de transport. IFB possède ou possédait les participations suivantes dans des sociétés de transport:
- CNC Ferry Boats intermodal, Belgique, 50 % (capitaux propres: 61000 EUR, résultat net 2004: pas connu), et sa filiale à 100 %, Rail Web. Cette société a été dissoute le 31 mars 2005.
- Affrètements Van Reeth, Belgique, 100 % (capitaux propres: 412000 EUR; résultat net en 2002: 150000 EUR).
- SA Unilog, Belgique, 55 % (capitaux propres: 1,9 millions EUR, résultat net 2004: 21000 EUR).
- SA Unilog, Royaume uni, 100 % (pas d'informations supplémentaires).
- SA Rail Infra Logistics, Belgique, 99,93 % (capitaux propres: 500000 EUR; résultat net 2004: 55000 EUR).
- ACTS België, Belgique, 12,5 % (pas d'informations supplémentaires). Cette société a été dissoute le 29 mars 2005.
- RKE, Belgique, 61,46 % (capitaux propres: 2,6 millions EUR, résultat net 2004: 250000 EUR).
- Coil Terminal, indirectement par RKE, car RKE détient une participation de 50 % dans Coil Terminal.
- CARRE (pas d'informations supplémentaires). Pour cette société, des négociations de vente sont en cours.
- GIE Cigogne Shuttle, Belgique (pas d'informations supplémentaires). Pour cette société, IFB prévoit le retrait d'IFB de la société.
- Haeger Schmidt International, Allemagne, 100 % (capitaux propres: 2,1 millions EUR, résultat net 2004: pas connu).
- Compagnie nouvelle des conteneurs Transports Nationaux et Internationaux, France, 2 % (pas d'informations supplémentaires).
- GIE NEN (pas d'informations supplémentaires). Ce GIE est en voie de dissolution.
- ACTS Belgique, 13 % (pas d'informations supplémentaires). Cette société a été dissoute le 5 novembre 2003.
- TRW, Belgique, 0,89 %.
48. Participation dans Haeger and Schmidt International. A travers sa filiale à 100 % Haeger and Schmidt International, IFB détient des participations dans les sociétés Best Logistics (Pologne), A van Reeth (France), KREAS et SITRA. Haeger et Schmidt réalise un chiffre d'affaires annuelles de EUR 50 millions, principalement par le transport fluvial.
49. Aperçu d'ensemble. L'organigramme suivant reprend toutes les participations d'IFB dans un aperçu d'ensemble. La systématique est la suivante:
Première colonne: les participations dans les sociétés actives exploitant des terminaux;
Deuxième colonne: les participations dans les sociétés actives dans le domaine du transport;
troisième colonne: les participations dans les sociétés prestataires de services;
quatrième colonne: les participations dans les sociétés (allemandes) actives dans le domaine du transport fluvial (barge);
+++++ TIFF +++++
2.1.1.2. Définition des marchés concernés et parts de marchés de IFB
50. La Commission a statué dans le passé sur la définition des marchés pertinents pour les activités d'expédition et les activités logistiques dans ses décisions COMP/M.3603 "UPS/Menlo" et COMP/M.3496 "TNT FORWARDING HOLDING/WILSON LOGISTICS"; elle a retenu comme marché de produit pertinent:
- Pour les activités d'expédition ou freight forwarding: "the organisation of transportation items (possibly including ancillary activities such as customs clearance, warehousing, ground services, etc.) on behalf of customers according to their needs."
- Pour les activités de logistique ou general logistic services: "the part of the supply chain process that plans, implements and controls the efficient, effective flow and storage of goods, services and related information from the point of origin to the point of consumption in order to meet customers' requirements."
51. Ces marchés ont été définis comme des marchés nationaux, malgré une tendance vers plus d'internationalisation.
52. Selon les informations transmises par le gouvernement belge, la part de marché d'IFB Logistics sur ces deux marchés est comprise entre 2 % et 5 %, ce qui s'expliquerait par la partie relativement faible des biens qui sont transportés par le transport combiné et le transport ferroviaire.
53. Cette estimation paraît crédible, si l'on compare le chiffre d'affaires d'IFB, qui a été de EUR […] millions en 2003, aux chiffres d'affaires des autres acteurs belges sur ce marché, qui ont eu en 2003 les chiffres d'affaires suivants en Belgique:
Entreprise | Chiffre d'affaires |
Hesse-Noordnatie | 485 millions EUR |
Danzas | 176 millions EUR |
Ziegler | 129 millions EUR |
Schenker | 156 millions EUR |
54. En ce qui concerne le marché des terminaux, il y a lieu d'opérer une distinction entre les terminaux continentaux et les terminaux maritimes.
55. En ce qui concerne les terminaux continentaux, la Commission a pris position sur la définition des marchés pertinents dans ses décisions COMP M 2632 "DEUTSCHE BAHN/ECT INTERNAIONAL/UNITED DEPOTS" et IV/M 1651 "MAERSK/SEA LAND" et IV/M.831 "PO/Nedlloyd".
56. Dans la décision COMP M 2632, la Commission a défini le marché de produit en cause comme le marché "für das Erbringen von Umschlagdienstleistungen im Containergüter-Hinterlandverkehr per Binnenschiff zwischen ARA-Häfen und deutschem Niederrhein/Ruhrgebiet", le marché géographique étant "die Containerterminals entlang des Niederrheins von Nijmeggen bis Köln". En d'autres mots, tous les terminaux du bas Rhin seraient le marché pertinent. Dans les décisions IV M 1651 et IV M 831, le marché géographique d'un port est défini comme suit: "Ports or groups of ports serve a particular hinterland or are used for transshipment to smaller ports. The geographic area they generally serve determines the geographic scope related to their services." Il s'en suit que le marché de produit est le marché du transbordement du fret, et que son étendue géographique couvre le hinterland d'un port donné.
57. Pour le cas d'espèce, on arrive donc à la conclusion que le marché de produit en cause peut être défini comme le marché des services de transbordement d'UTI du/vers le transport terrestre (route — chemin de fer — barge). Le marché géographique pertinent est au minimum la région d'Anvers et ses environs, éventuellement même la région des ports ARA.
58. Á part les terminaux continentaux d'IFB, les terminaux au moins trimodaux de Hesse-Noordnatie (Noordzeeterminal, Europaterminal) et P O Ports (Seaport terminal) offrent les services de transbordement d'UTI du/vers le transport terrestre (route — chemin de fer — barge). Ces terminaux sont bien plus importants en volumes d'UTI traités que les terminaux d'IFB. En 2004, Hesse-Noordnatie a traité 4,9 millions TEU, P O Ports 0,7 millions TEU, tandis qu'IFB a traité 0,4 millions TEU. Le part de marché d'IFB est donc d'environ 6,7 %.
59. Les deux terminaux maritimes dans lesquels IFB détient des participations n'ont que des parts de marchés marginales en Belgique et en France. IFB ne détient pas de participations dans des terminaux dans d'autres pays.
2.1.2. La SNCB
60. La SNCB a été créée par la loi belge du 23 juillet 1926 créant la Société Nationale des Chemins de Fer Belges [7]. Depuis le 14 octobre 1992 [8], elle est une entreprise publique autonome et société anonyme de droit public [9]. Ainsi, la SNCB est soumise aux dispositions légales et réglementaires de droit commercial national qui sont applicables aux sociétés anonymes pour tout ce qui n'est pas expressément prévu par ou en vertu du titre premier de la loi du 21 mars 1991 portant réforme de certaines entreprises publiques économiques, précitée, ou en vertu d'une loi spécifique quelconque.
61. L'État belge a réformé la structure de la SNCB au 1er janvier 2005. Elle a été transformée en trois sociétés distinctes, à savoir:
- la SNCB Holding: une société "de type holding" qui détiendra des participations dans les deux autres sociétés;
- Infrabel, le gestionnaire de l'infrastructure ferroviaire;
- la nouvelle SNCB, l'entreprise ferroviaire.
62. L'objet social de la SNCB est défini à l'art. 1bis de la loi du 23 juillet 1926, précité, inséré par la loi du 1er août 1966 [10] et modifié par l'art. 155 de la loi du 21 mars 1991, précité, comme suit:
"(1) La société a pour objet le transport de voyageurs et de marchandises par chemin de fer."
"(2) La société peut, par elle-même ou par voie de participations à des organismes existants ou a créer, belges, étrangers ou internationaux, faire toutes opérations commerciales, industrielles ou financières se rapportant directement ou indirectement, en tout ou en partie, à son objet social ou qui seraient susceptibles d'en faciliter ou d'en favoriser la réalisation ou le développement."
"(3) Est notamment considéré comme susceptible de favoriser la réalisation de l'objet social, le fait de fabriquer et de vendre des biens ou des services ayant trait directement ou indirectement à l'activité ferroviaire."
63. Cet article a toujours été interprété de manière extensive par la jurisprudence et la doctrine belge. Selon les autorités belges, les activités d'IFB sont clairement couvertes par lui.
64. Les organes de gestion de la SNCB sont le Conseil d'administration, le Comité de direction et l'Administrateur délégué. Le Conseil d'administration est composé de 10 membres, y compris l'Administrateur délégué. Les administrateurs sont nommés par le Roi, par arrêté délibéré en Conseil des Ministres. Ils sont choisis, après une procédure ouverte, en fonction de la complémentarité de leurs compétences telle que l'analyse financière et comptable, les aspects juridiques, la connaissance du secteur du transport, l'expertise en matière de mobilité, la stratégie du personnel et les relations sociales. Une fois nommés, les membres du Conseil d'administration exercent leur mandat de manière indépendante, et ne doivent pas obéir aux instructions de quiconque.
65. Les membres du Comité de direction, à l'exception de l'Administrateur délégué, nommé par le Roi, sont nommés par le Conseil d'administration, qui en détermine aussi le nombre. Le Comité de direction forme un collège.
2.2 Les difficultés financières rencontrées par IFB
66. Au cours des exercices 2001 et 2002, IFB a enregistré des pertes considérables: Selon les comptes annuels de 2002 d'IFB, les pertes cumulées au 31 décembre 2002 s'élevaient à EUR 137 millions (dont EUR 25 millions reporté de 2001), ce qui avait pour résultat des fonds propres négatifs de EUR 84 millions. A la fin de l'exercice 2001, ses fonds propres s'étaient encore élevés à EUR 28 millions.
67. Toujours selon les comptes annuels de 2002, les pertes opérationnelles de l'exercice 2002, c'est-à-dire la différence entre les dépenses courantes et les revenues courantes, s'élevaient à 13,4 millions d'EUR. Il y a lieu d'analyser d'abord les raisons pour les difficultés financières, et de décrire ensuite la réaction de l'encadrement d'IFB et de la SNCB, ainsi que la réaction des créanciers privés d'IFB.
2.2.1. Les raisons pour les difficultés financières
68. La principale raison pour les difficultés financières d'IFB a été les difficultés financières rencontrées par ses participations en France dans le port de Dunkerque, qui ont obligé IFB à faire d'importantes provisions dans ses comptes annuels de 2001 et 2002.
69. De plus, les activités "IFB Logistics" et "IFB Terminals" réalisaient de légères pertes en 2001 et 2002.
2.2.2. La réaction de l'encadrement d'IFB et de la SNCB
70. Depuis 2000, IFB n'avait plus payé toutes les factures que la SNCB lui avait envoyées pour les prestations de service de train. En 2001 et surtout en 2002, IFB a continué cette pratique. La SNCB semble avoir toléré cette pratique. Ainsi, IFB se trouvait fin janvier 2003 avec des factures impayées de la SNCB d'une valeur totale de EUR 63 millions.
71. En réaction aux difficultés financières rencontrées par IFB, tant le conseil d'administration d'IFB que son actionnaire principal, la SNCB, sont devenus de plus en plus convaincus que la survie du groupe IFB à long terme impliquait une modification structurelle du plan de la gestion de l'entreprise.
72. Le 19 septembre 2002, l'administrateur délégué d'IFB a chargé deux réviseurs de rédiger un rapport spécial afin d'évaluer la situation financière de l'entreprise. Le 24 décembre 2002, l'Assemblée Générale extraordinaire des Actionnaires ("AGE") d'IFB a pris connaissance du fait que la SNCB, suite à la réunion du Conseil d'administration qui a eu lieu le 20 décembre 2002, était disposée à souscrire une augmentation de capital à raison de maximum EUR 80 millions afin de redresser la situation financière d'IFB, dont EUR 20 millions pour répondre aux besoins d'IFB en liquidités. Les deux conseils d'administration de la SNCB et d'IFB ont donc donné leur accord de principe à deux augmentations de capital — de EUR 60 millions en convertissant des créances de la SNCB sur IFB en capital et de EUR 20 millions en mettant à la disposition d'IFB des moyens en liquide — à souscrire par la SNCB afin d'assurer la continuité de l'activité d'IFB.
73. IFB et la SNCB ont conclu le 7 avril 2003 un "contrat cadre concernant la restructuration d'IFB" afin de mettre en œuvre ces augmentations de capital. Ce contrat, qui est un contrat de droit privé, prévoit deux volets: un volet "mesures de sauvetage" et un volet "mesures de restructuration".
74. Vu ces circonstances, le Conseil d'administration d'IFB, après concertation avec son actionnaire principal, la SNCB, a décidé de convoquer une AGE, comme prévu à l'article 633 du Code belge des Sociétés en cas de pertes au moins égales à la moitié du capital social. Lors de cette assemblée, réunie le 20 mai 2003, les actionnaires d'IFB ont pris connaissance du rapport spécial du conseil d'administration d'IFB, dans lequel le contrat cadre entre la SNCB et IFB a été décrit et dans lequel il a été proposé de poursuivre les activités d'IFB moyennant la mise en œuvre d'une restructuration. Sur cette base, les actionnaires d'IFB ont marqué leur accord avec la poursuite des activités d'IFB.
2.2.3. La réaction des créanciers privés d'IFB
75. IFB a obtenu de la part des banques d'affaires privées des prêts et des garanties bancaires. Selon les informations transmises par le gouvernement belge, les difficultés financières rencontrées par IFB n'a eu le moindre impact sur les relations entre IFB et les banques: Ces banques ont tous maintenu les conditions contractuellement prévues, sans exiger des garanties complémentaires à celles d'usage ou autres cautions ou sûretés. Toujours selon le gouvernement belge, elles ont toutes été disposées à accorder de nouveaux prêts à des conditions concurrentielles.
76. Au 31 décembre 2004, IFB avait les contrats de prêt suivants auprès des banques privées:
Objet du prêt | Banque | Année | Taux | Montant (en EUR) | Situation au 31.12.2004 (en EUR) |
[…] | […] | 1997 | [entre 2 et 6 %] | 328334,97 | […] |
[…] | […] | 1999 | [entre 2 et 6 %] | 1264930,18 | […] |
[…] | […] | 1999 | [entre 2 et 6 %] | 1611307,91 | […] |
[…] | […] | 2001 | [entre 2 et 6 %] | 4945476,00 | […] |
[…] | […] | 2003 | [entre 2 et 6 %] | 2000000,00 | […] |
Total | | | | 10150049,06 | 5550066,03 |
77. Le dernier contrat de prêt a été conclu en juillet 2003, donc après la conclusion de l'accord cadre entre IFB et la SNCB et après que les banques ont appris les difficultés financières d'IFB.
78. Les garanties bancaires dont disposait IFB au 31 décembre 2004 ont été les suivants:
Bénéficiaire de la garantie bancaire | Montant (en EUR) |
Service public Fédéral FINANCES Garantie Douanes et Accises | 2401220,64 |
Service public Fédéral FINANCES Garantie Différend fiscal | 1772817,63 |
Service Public Fédéral MOBILITE ET TRANSPORT Garantie Commissionnaire de transport | 111552,12 |
Autres garanties | 44767,12 |
79. Les lignes de crédit afférentes à ces garanties ont toutes été maintenues, sans modification des conditions contractuellement prévues.
2.3. Les dispositions principales du "contrat cadre entre la SNCB et IFB concernant la restructuration d'IFB"
80. Afin d'assurer la continuité d'IFB, la SNCB et IFB ont conclu le contrat cadre mentionné ci-dessus qui stipule que l'exécution des mesures proposées se fera en deux phases: dans une première phase, une série de mesures de sauvetage seront prises à l'égard d'IFB jusqu'au moment où un plan de restructuration pourra être mis en œuvre pour IFB; dans une deuxième phase, des mesures seraient élaborées dans le cadre d'un plan de restructuration touchant IFB, les mesures de sauvetage pouvant à cette occasion être converties en capital.
81. Dans le préambule du contrat, la SNCB confirme son intention de "donner son approbation à une augmentation de capital d'IFB à souscrire par la SNCB à concurrence d'environ 60 millions EUR en convertissant les créances de la SNCB sur IFB et en mettant à la disposition d'IFB un montant supplémentaire de 20 millions EUR, dont 5 millions EUR seraient libérés immédiatement."
82. L'article 2 du contrat cadre entre la SNCB et IFB prévoit deux volets, à savoir un volet "mesures de sauvetage" et un volet "mesures de restructuration".
2.3.1. Modalités et conditions d'octroi des mesures de sauvetage
83. Le premier volet de l'article 2 prévoit trois mesures de sauvetage:
(1) l'octroi d'une avance récupérable de EUR 5 millions;
(2) l'octroi d'une facilité de crédit d'un maximum de EUR 15 millions et
(3) l'octroi d'un délai de paiement provisoire portant sur les dettes d'IFB.
84. L'article 3 du contrat cadre stipule que le taux d'intérêt sur l'avance récupérable et les sommes prélevées sur la facilité de crédit sera au moins égal au taux d'intérêt de référence appliqué par la Commission européenne pour l'aide d'État [11]. Il prévoit aussi que les intérêts sont capitalisés. Leur paiement aura lieu au même moment que le paiement des créances dues.
85. L'avance et la facilité de crédit sont mises à disposition à titre provisoire afin de répondre aux besoins financiers urgents d'IFB et seront converties en capital dans le cadre du plan de restructuration à établir.
86. En ce qui concerne en particulier l'octroi d'une facilité de crédit d'un maximum de EUR 15 millions, IFB pourra imputer les créances de la SNCB vis-à-vis d'IFB facturées à partir du 1er janvier 2003 à l'exception d'une facture du 31 janvier 2003 d'un montant de EUR 8 millions.
87. L'octroi d'un délai de paiement provisoire porte sur toutes les dettes d'IFB qui étaient facturées au 31 décembre 2002, y compris la facture du 31 janvier 2003 d'un montant de EUR 8 millions, ainsi que les dettes dont le montant était certain et liquide au 31 décembre 2002, mais qui ne sont en général pas facturées. Le total des montants dus à la SNCB s'élevait à EUR 63 millions. En plus, le montant en question doit être augmenté d'un intérêt de retard conventionnel, fixé à [entre 1 et 2] pro mille par décade indivisible [12], ou d'un taux d'intérêt légal applicable. Les intérêts sont capitalisés, et seront payé au moment du paiement de la créance principale.
88. Les intérêts dus par IFB à la SNCB pour les dettes et la facilité de crédit étaient de 2,2 millions EUR en 2002, de 3, 9 millions EUR en 2003 et de 4,7 millions EUR en 2004. Le contrat cadre prévoit que le paiement des intérêts a lieu en même temps que le paiement des créances.
89. IFB a aussi renoncé, vis-à-vis de la SNCB, à la prescription de ses dettes. L'ensemble de ces mesures, à l'exception de l'avance récupérable, a été mis en œuvre dès la signature du contrat cadre, à savoir le 7 avril 2003. En ce qui concerne le délai de paiement, il avait de facto déjà été accordé avant la conclusion du contrat cadre, et formalisé par le contrat cadre.
2.3.2. Modalités et conditions d'octroi des mesures de restructuration
90. En ce qui concerne le deuxième volet de l'article 2 du contrat cadre, il prévoit que les "mesures de restructuration" seront développées par les conseils d'administration de la SNCB et de IFB et ensuite soumis à l'État belge pour approbation.
91. L'article 4 du contrat cadre, intitulé "modalités d'octroi du volet 'mesures de restructuration", est rédigé comme suit:
"Les Parties confirment leur intention de mettre à exécution les mesures suivantes pour autant qu'elles soient conformes à un plan de restructuration approuvé par leurs deux Conseils d'administration, par l'État belge et si nécessaire par la CE, et sous réserve d'approbation par les actionnaires d'IFB:
- La conversion en capital d l'avance récupérable d'un montant de 5 millions EUR
- La conversion en capital de la partie de facilité de crédit prélevée pour un montant maximum de 15 millions EUR […]
- La conversion en capital des dettes de […] 63 millions EUR
- Eventuellement et à condition que les deux parties soient d'accord à ce sujet, une augmentation de capital supplémentaire […]"
92. Le gouvernement belge a informé la Commission dans les réunions du 12 décembre 2003 et du 16 septembre 2005 ainsi que dans ses lettres du 13 janvier 2004, du 28 janvier 2005, du 25 mars 2005 et du 30 juin 2005 sur les détails prévus pour les mesures de restructuration, qui comprennent des mesures ad hoc entamées par IFB vis-à-vis de ses filiales exploitant des terminaux en France, un plan de restructuration pour la société IFB, ainsi qu'une augmentation de capital.
93. À ce jour, aucune de ces mesures n'a été mise en œuvre.
2.3.2.1. Les mesures ad hoc entamées par IFB vis-à-vis de ses filiales exploitant des terminaux en France
94. Comme expliqué ci-dessous, IFB a poursuivi une stratégie de désinvestissement pour ses filiales françaises. Cette politique est quasiment achevée (cf. ci-dessus la description des participations); elle a été accompagnée d'une dénonciation des lettres de confort.
2.3.2.2. Le plan de restructuration
95. IFB et la SNCB ont élaboré avec le consultant McKinsey un plan de restructuration pour IFB, qui garantit la viabilité économique à longue terme d'IFB. Ce plan de restructuration prévoit deux parties:
- Restructuration de l'activité "IFB Logistics";
- Restructuration de l'activité "IFB Terminals".
96. La mise en œuvre du plan de restructuration a commencé dès 2003, et sera achevée en 2005. Le plan de restructuration prévoyait qu'IFB réalisera des bénéfices opérationnels de 0,5 millions d'EUR en 2003 et de 0,8 millions d'EUR en 2004, après avoir réalisé des pertes opérationnelles de 13,4 millions d'EUR en 2002.: Le tableau suivant montre la répartition des bénéfices et des pertes entre les différentes activités prévue pour les années 2002 à 2004:
| 2002 | 2003 | 2004 |
Filiales | […] | […] | […] |
IFB Terminals | […] | […] | […] |
IFB Logistics | […] | […] | […] |
Total | - 13,4 | 0,5 | 0,8 |
97. Les résultats réalisés en 2003 étaient inférieurs aux prévisions, le résultat d'exploitation étant de — 2,9 millions d'euros. Cela était dû notamment aux pertes des filiales (pertes de […] millions d'euros au lieu d'un bénéfice de […] millions d'euros) et aux faibles bénéfices d'IFB Logistics (bénéfice de […] millions d'euros au lieu d'un bénéfice escompté de […] millions d'euros).
98. Les résultats réalisés en 2004 étaient supérieurs aux prévisions, le résultat d'exploitation étant un bénéfice de 5,7 millions d'euros. IFB Logistics y contribuait pour […] millions d'euros, IFB Terminals pour […] millions d'euros, et les filiales pour […] millions d'euros.
99. Le plan de restructuration prévoit aussi la nécessité de nouveaux investissements d'une hauteur de […] millions d'EUR. Il y a lieu de présenter de plus près les mesures de restructuration prévues dans les différents secteurs d'activités et le besoin pour de nouveaux investissements.
a) Restructuration de l'activité logistique
100. En ce qui concerne l'activité "IFB Logistics", le plan de restructuration prévoyait un bénéfice opérationnel de […] millions d'EUR en 2003, après des pertes de […] millions d'EUR en 2002. Pour y arriver, le plan prévoyait un total de neuf mesures qui devaient permettre de réaliser des économies de […] millions d'EUR. Suite à la réduction du volume du transport conventionnel, qui devrait entraîner des pertes de […] millions d'EUR, l'amélioration totale serait donc de […] millions d'EUR. Les neuf mesures repris dans le tableau suivant:
Mesures | Bénéfice |
1.Effet de la réduction de la charge salariale | […] millions |
2.Consultance et outsourcing | […] millions |
3.Réductions de valeur et amortissement exceptionnel | […] millions |
4.Cessation des branches non rentables du North European Network | […] millions |
5.Perte de volume de trafic conventionnel | […] millions |
6.Reprise de provisions entretien wagons | […] millions |
7.Croissance de l'intermodal | […] millions |
8.Révision du contrat Railbarge (augmentation des prix et reengineering produit) | […] millions |
9.Augmentation des commissions des représentations (agent) | […] millions |
10.Réduction des frais généraux | […] millions |
101. Pour l'essentiel, les mesures de restructuration consistaient donc dans une augmentation des prix, liée à un nouveau design des produits, des reprises des provisions et des amortissements exceptionnels, une réduction des coûts salariaux et frais généraux, ainsi qu' une cessation d'activités non rentables.
102. Dans l'activité "IFB Logistics", il a donc été prévu que la restructuration s'achèverait entre mi-2003 et mi-2004.
b) Restructuration de l'activité terminal
103. La restructuration de l'activité "IFB Terminal", en revanche, devrait prendre trois ans. Il a été prévu que cette activité réduirait ses pertes opérationnelles de […] millions d'EUR en 2002 à […] millions d'EUR en 2003 et […] millions d'EUR en 2004, avant de conclure l'année 2005 avec un bénéfice opérationnel de […] millions d'EUR. Pour y arriver, le plan de restructuration prévoyait les 8 mesures suivantes:
Mesures | Bénéfice |
1.Mainhub:Réduction du personnelAdaptations informatiquesRéduction des amortissements et reprise des provisionsAugmentation du nombre des manipulations | […] millions |
2.CirkeldijckRéduction des opérations du terrainVente des actifsLocation du terminalRéduction du volumeRéduction du personnel | […] millions |
3.ZomerwegTransfer RailbargeAugmentation volumeExpansionsInvestissements | […] millions |
4.Dry port MuizenRéduction de coûts de personnel grâce au nouveau système de surveillanceAugmentation de volume | […] millions |
5.SchijnpoortAugmentation de volumeRéduction de coût d'exploitation | […] millions |
6.RenoryVente d'un stackerArrêt de la solidarité financière d'IFB | […] millions |
7.Bressoux: Fermeture du terminal | […] millions |
104. Les mesures les plus importantes concernent donc les terminaux Mainhub, Cirkeldijck et Zomerweg. Ils seront expliqués plus en détail dans les paragraphes qui suivent.
105. Mainhub. Le Mainhub fera, dès le deuxième semestre 2003 jusqu'à fin 2005, l'objet d'une réorganisation intégrale, qui permettra, grâce notamment à des adaptations informatiques importantes, une réduction du personnel combinée avec une augmentation du nombre des manipulations. Cela permettra une meilleure utilisation de la capacité du terminal, qui n'a été utilisé qu'à la hauteur de […] % en 2002.
106. Cirkeldijck. Dans le terminal Cirkeldijck, IFB renforcera sa coopération avec Hesse NoordNatie (HNN). HNN reprendra les opérations de terrain, tandis que IFB maintient le planning et le chargement du transport ferroviaire. […].
107. Zomerweg. Le terminal Zomerweg sera transformé de terminal bimodal en terminal trimodal, avec le transfert de tout le trafic Railbarge vers ce terminal. Dans ce contexte, le terrain et le quai seront élargis, le terrain, l'entrée et les chemins seront adaptés, et des investissements en matériel seront nécessaires.
c) Besoin d'investissement
108. La restructuration de Mainhub ainsi que la restructuration de Zomerweg impliquent la nécessité de nouveaux investissements d'une hauteur de […] millions d'EUR chacun. En même temps, la vente de la grue portique du terminal Cirkeldijck permettra de réduire ce besoin à […] millions d'EUR au total.
2.3.2.3. L'augmentation du capital
109. Par lettre du 28 janvier 2005, le gouvernement belge a informé la Commission que l'encadrement d'IFB ainsi que l'encadrement de la SNCB estiment qu'il est nécessaire d'accompagner le plan de restructuration d'une augmentation de capital d'IFB, comme l'avait prévu le contrat cadre. Le montant nécessaire, légèrement revu à la hausse par rapport aux prévisions du contrat cadre, serait de 96,5 millions EUR.
110. L'augmentation de capital se déroulera comme suit: d'abord, les dettes d'IFB vis-à-vis de la SNCB, qui s'élèvent à 78 millions EUR, et les intérêts dus sur ces dettes, qui s'élèveront à 13,5 millions EUR à la fin de l'année 2005, seront converties en capital. L'origine de ces dettes sont les mesures de sauvetage 1 et 2, donc le délai de paiement ainsi que la facilité de crédit. Ensuite, la SNCB apportera le reste, c'est-à-dire 5 millions EUR, en nature. La procédure correspond donc à la procédure prévue à l'article 4 du contrat cadre.
111. L'apport en nature consiste dans la participation de la SNCB dans la société TRW. Cette participation s'élève, comme expliqué ci-dessus, à 47 %, IFB détenant déjà une participation de 0,9 % dans la société. TRW exploite des terminaux à Anvers, Zeebrugge, Oostende, Charleroi, Liège, Bruxelles, Etge, Genk et Muizen, et offre des trains de fret pour 11 pays de l'UE.
112. Le montant de l'augmentation de capital est plus élevé que ce qui avait été prévu lors de la conclusion du contrat cadre entre IFB et la SNCB, qui prévoyait une augmentation de capital de 80 millions EUR, mais moins élevé que la proposition du consultant McKinsey, qui dans le plan de restructuration tablait sur une augmentation de capital de 120 millions EUR.
113. Le gouvernement belge estime que cette augmentation de capital laisserait à IFB, après réduction du capital pour résorber les pertes reportées, des capitaux propres de 23,9 millions EUR, ce qui présenterait une structure de capital saine avec un rapport entre le financement par fonds propres et les dettes adapté aux activités d'IFB.
114. Le taux de solvabilité, c'est-à-dire le ratio capitaux propres/passif, d'IFB avant et après l'augmentation du capital est illustré par la table suivante:
| Situation au 30.06.2005 | Augmentation proposée | Situation après l'augmentation |
Capitaux propres | - 72,6 | 96,5 | 23,9 |
Provisions et impôts différés | 14,3 | | 14,3 |
Dettes | 125,6 | - 91,5 | 34,1 |
Total du passif | 67,3 | | 72,3 |
Taux de solvabilité | | | 33 % [13] |
115. L'augmentation du capital est prévue pour le deuxième semestre 2005, après approbation par la Commission européenne et le Conseil d'Administration de la SNCB.
116. Contrairement à ce qui était prévu à l'article 4 du contrat cadre, le plan pour l'augmentation du capital n'a pas été soumis au gouvernement belge pour approbation. Le gouvernement belge estime qu'une telle approbation n'est pas nécessaire, car il s'agit d'une décision purement commerciale de la SNCB, que cette dernière peut prendre sans approbation par l'État.
2.4. Développement financier d'IFB depuis la conclusion du contrat cadre
117. La situation économique et financière d'IFB s'est améliorée substantiellement depuis la conclusion du contrat cadre en avril 2003. Ainsi, le résultat d'exploitation a connu une évolution positive de — 47,36 millions EUR en 2002 à 5,74 millions EUR en 2004. Le résultat de l'exercice avant impôts s'est amélioré de — 109,76 millions EUR en 2002 à 13,21 millions EUR en 2004.
118. Le tableau suivant donne un aperçu du développement des principaux indicateurs économiques et financiers d'IFB:
Tableau: Situation économique et financière d'IFB (en 000 EUR).
| 31.12.2002 (audité) | 30.09.2003 | 31.12.2003 (audité) | 30.09.2004 | 31.12.2004 (audité) |
Ventes et prestations | 65377 | 43184 | 59091 | 61369 | 85751 |
Dont chiffre d'affaires | 63669 | 42445 | 58079 | 59903 | 83343 |
Coût des ventes et des prestations | 112734 | 43781 | 62051 | 58759 | 80011 |
Résultat d'exploitation | (47357) | (1336) | (2960) | 2610 | 5740 |
Résultat financier | (3034) | — | (4458) | (3247) | (3303) |
Résultat exceptionnel | (59369) | — | 7342 | 6754 | 10773 |
Résultat de l'exercice avant impôt | (109760) | (1200) | (76) | 6117 | 13210 |
Cash Flow | | (101) | | | |
Capitaux propres | (84068) | (85277) | (83941) | (77775) | (74850) |
119. L'amélioration de la situation économique et financière est due d'un côté à la réalisation du plan de restructuration, de l'autre à la poursuite de la stratégie de désinvestissement en ce qui concerne les participations.
120. Dans le premier semestre 2005, IFB a continué à enregistrer des bénéfices: le résultat d'exploitation était de 1,6 millions EUR, le résultat avant impôt de 2,2 millions EUR.
2.4.1. La mise en œuvre du plan de restructuration
121. Pour la mise en œuvre du plan de restructuration, il faut distinguer entre les mesures qui affectent l'ensemble des activités d'IFB, et les mesures spécifiques à IFB Logistics et IFB Terminals.
2.4.1.1. Mesures qui affectent l'ensemble des activités d'IFB
122. La conclusion d'une nouvelle convention de travail au niveau de l'entreprise et la modification du règlement de travail ont permis d'atteindre un taux d'activité plus élevé (le nombre de jours à prester par an a augmenté) à des coûts inférieurs (la rémunération pour le travail de week-end et celle pour le travail d'équipe a été réduite). Les services administratifs et commerciaux ont été centralisés à Berchem, ce qui a permis de fermer l'établissement à Gand et de réduire la capacité de celui de Zeebruges.
123. Ces mesures ont contribué à limiter le personnel nécessaire et à baisser les frais généraux.
2.4.1.2. Mesures spécifiques à IFB Terminals
124. En plus des mesures prévues par le plan de restructuration deux mesures ont été prises: Pour le terminal de Cirkeldijck, le prix de manutention a été revu à la hausse. En général, les trafics ont été analysés et, par la suite, réorientés en concertation avec les clients.
125. L'ensemble des mesures, ainsi que la croissance des volumes manutentionnés, ont permis à IFB Terminals de re-devenir rentable dès 2004, avec un bénéfice avant impôts de […] EUR, après des pertes avant impôts de […] millions EUR en 2003. L'objectif fixé par le plan de restructuration a donc été plus que respecté (pour rappel: le plan de restructuration prévoyait des pertes de […] EUR.)
2.4.1.3. Mesures spécifiques à IFB Logistics
126. En plus des mesures prévues par le plan de restructuration, IFB Logistics a réalisé une analyse profonde de ses produits ferroviaires, qui a révélé l'existence de produits non rentables, qu'IFB a arrêté de produire depuis.
127. Pour d'autres produits, cette analyse a démontré la nécessité d'améliorations sur le plan technique. Ces améliorations ont été faites, notamment pour le secteur du transport intermodal des conteneurs.
128. L'ensemble des mesures a permis à IFB Logistics de re-devenir rentable dès 2003, avec un bénéfice avant impôts de […] EUR. En 2004, le résultat a encore été amélioré à […] millions EUR. IFB Logistics n'a donc pas pu atteindre l'objectif fixé par le plan de restructuration pour 2003 ([…] millions EUR), mais a pu l'atteindre en 2004 (l'objectif était de […] millions EUR).
2.5. Budget
129. Le montant prévisionnel total des mesures de sauvetage s'élève à maximum EUR 78 millions [14].
130. Le montant total de l'augmentation de capital prévu s'élève à 96,5 millions EUR, dont 78 millions EUR résulteront de la conversion des dettes existantes (63 millions) et des mesures de sauvetage (15 millions) en capital, et 13,5 millions EUR de la conversion des intérêts capitalisés en capital. 5 millions EUR supplémentaires seront apportés par la SNCB en nature, par le transfert de la participation de la SNCB dans TRW à IFB.
2.6. Mise à disposition des ressources financières et durée
131. Dans ses lettres du 28 janvier 2005 et du 25 mars 2005, le gouvernement belge explique que les mesures 2 (facilité de crédit de 15 millions d'euro) et 3 (délai de payement pour les dettes existantes de 63 millions d'euro) du volet "mesures de sauvetage" ont été mises en œuvre par la SNCB et IFB à partir du 7 avril 2003. En revanche, IFB n'a pas eu besoin de l'avance récupérable prévue par la mesure 1.
132. Le contrat cadre prévoit que, sauf conversion en capital dans le cadre d'un éventuel plan de restructuration approuvé ou de toute autre mesure comparable convenue, les sommes majorées des intérêts sont remboursables douze mois après avoir été effectivement mises à la disposition d'IFB par la SNCB. L'encadrement d'IFB et de la SNCB ayant convenu du principe d'une augmentation de capital, ils considèrent que le contrat de prêt a été tacitement prolongé jusqu'à ce que l'augmentation du capital ait lieu. IFB continue en attendant d'accumuler les intérêts prévus par le contrat cadre, à savoir un intérêt de retard conventionnel, fixé à [entre 1 et 2] pro mille par décade indivisible [15], ou un taux d'intérêt légal applicable. Le taux moyen des intérêts est de [entre 3,6 et 7,2] %. La totalité des intérêts devra être payée au moment du paiement de la créance, ou sera convertie en capital social.
133. L'augmentation de capital est prévue pour le deuxième semestre 2005, après son approbation par la Commission.
3. APPRÉCIATION
3.1. Evaluation du caractère d'aide des mesures de sauvetage et de restructuration
134. Selon l'article 87, paragraphe 1, du traité, "sont incompatibles avec le marché commun, dans la mesure où elles affectent les échanges entre Etats membres, les aides accordées par les Etats ou au moyen de ressources de l'État sous quelque forme que ce soit qui faussent ou menacent de fausser la concurrence en favorisant certaines entreprises ou certaines productions".
3.1.1. Accordée par l'État ou au moyen de ressources de l'État
135. Il se pose donc d'abord la question de savoir si le soutien financier de la SNCB à IFB a été "accordées par les Etats ou au moyen de ressources de l'État". Selon la jurisprudence Stardust Marine de la CJCE [16], ce critère est rempli si d'une part il s'agit de ressources d'Etat et si d'autre part l'octroi de ceux-ci est imputable à l'État en question, à savoir la Belgique.
3.1.1.1. Ressources d'État
136. En ce qui concerne l'aspect "fonds publics", la Commission constate que la SNCB est qualifiable d'entreprise publique au sens de l'article 2 de la Directive de la Commission 2000/52/CE [17]: l'État belge détient 100 % du capital souscrit de la SNCB, et le Conseil d'administration, ainsi que l'administrateur délégué, sont nommés par le Roi, par arrêté délibéré en Conseil des Ministres. Ainsi, et le critère a) et le critère c) à l'alinéa 2 de l'article 2 de la Directive sont remplis.
137. Dans ce contexte, "… il convient de rappeler qu'il découle déjà de la jurisprudence de la Cour que l'article 87, paragraphe 1, CE englobe tous les moyens pécuniaires que les autorités publiques peuvent effectivement utiliser pour soutenir des entreprises, sans qu'il soit pertinent que ces moyens appartiennent ou non de manière permanente au patrimoine de l'État. En conséquence, même si les sommes correspondant à la mesure en cause ne sont pas de façon permanente en possession du Trésor public, le fait qu'elles restent constamment sous contrôle public, et donc à la disposition des autorités nationales compétentes, suffit pour qu'elles soient qualifiées de ressources d'État. " [18]
138. En conséquence, la Commission estime que les sommes mises à la disposition d'IFB sont à qualifier de ressources d'État.
3.1.1.2. Imputabilité
3.1.1.3. En ce qui concerne le critère de l'imputabilité des mesures à l'État concerné, l'arrêt Stardust Marine stipule que "…le seul fait qu'une entreprise publique soit sous contrôle étatique ne suffit pas pour imputer des mesures prises par celle-ci, telles que les mesures de soutien financier en cause, à l'État. Il est encore nécessaire d'examiner si les autorités publiques doivent être considérées comme ayant été impliquées, d'une manière ou d'une autre, dans l'adoption de ces mesures. …. [19]"
139. Il ressort donc de la jurisprudence de la Cour que le critère de l'imputabilité à l'État doit faire l'objet d'un examen au cas par cas par la Commission. La Cour admet qu'en règle générale, "… il sera très difficile pour un tiers, précisément à cause des relations privilégiées existant entre l'État et une entreprise publique, de démontrer dans un cas concret que des mesures d'aide prises par une telle entreprise ont effectivement été adoptées sur instruction des autorités publiques. A cet égard, il ne saurait être exigé qu'il soit démontré, sur le fondement d'une instruction précise, que les autorités publiques ont incité concrètement l'entreprise publique à prendre les mesures d'aide en cause" [20]. Pour ces motifs, selon la même jurisprudence, "…il y a lieu d'admettre que l'imputabilité à l'État d'une mesure d'aide prise par une entreprise peut être déduite d'un ensemble d'indices résultant des circonstances de l'espèce et du contexte dans lequel cette mesure est intervenue."
140. Dans le cas d'espèce, il faut distinguer, en ce qui concerne l'imputabilité, entre la période avant la conclusion du contrat cadre le 7 avril 2003 et la période après.
141. En ce qui concerne la période avant la conclusion du contrat cadre, il se pose la question de savoir si la décision de la SNCB de ne pas demander le paiement des sommes pour les prestations de service de transport à partir de 2000 est imputable à l'État belge.
142. La Commission ne dispose d'aucune information sur la question de savoir comment et pourquoi la SNCB a décidé de ne pas demander le paiement de ses factures dues. Puisque le non paiement des factures semble avoir été systématique dans la période fin 2000 jusque début 2003, la Commission a cependant des doutes qu'une telle décision aurait pu être prise par l'encadrement moyen de l'entreprise. Il semble que les auditeurs de l'entreprise ont dû le constater et alerter l'encadrement supérieur, et éventuellement aussi le commissaire du gouvernement en charge de la SNCB. La Commission exprime donc à ce stade des doutes si la décision de la SNCB de ne plus demander le paiement de ses factures à IFB à partir de fin 2000 a été imputable à l'État belge, et invite les autorités belges à lui fournir tout élément utile pour établir comment cette décision a été prise.
143. En ce qui concerne la période après la conclusion du contrat cadre, l'analyse du dossier par la Commission a relevé trois indices concrets pour une imputabilité des mesures de sauvetage et de restructuration en faveur d'IFB à l'État belge:
- La soumission du plan de restructuration à l'approbation par l'État belge
- Les articles de presse démontrant une forte influence du gouvernement belge sur la SNCB pendant l'année 2003
- L'ampleur, le contenu et les conditions du contrat cadre
a) L'approbation par les autorités publiques
144. Dans ses arrêts Van der Kooy [21], Italie/Commission [22] et Commission/France [23], la Cour a déduit l'imputabilité de l'aide du fait que l'octroi de l'aide ait été sujet à l'approbation par les autorités publiques. Dans l'arrêt Van der Kooy, cet élément suffit à lui seul pour établir l'imputabilité; dans les arrêts Italie/Commission et Commission/France, l'approbation est combinée avec d'autres éléments qui montrent l'influence des pouvoirs publics [24]. La récente décision Space Park Development GmbH, qui a été la première décision de la Commission appliquant l'arrêt Stardust Marine, a déduit l'imputabilité d'une aide également du fait que le prêt en question devait recevoir l'agrément des autorités du Land de Brême [25]. Par conséquent, la soumission d'une mesure à l'État membre pour approbation constitue un indice pour l'imputabilité.
145. Dans le présent dossier, l'article 2 du contrat cadre oblige les Conseils d'administration de la SNCB et d'IFB de soumettre le plan de restructuration pour approbation par l'État belge. Cela constitue un indice supplémentaire de l'imputabilité des décisions de la SNCB dans le présent cas à l'État belge.
146. Le gouvernement belge a informé la Commission entre-temps que, à la différence de ce qui a été prévu dans le contrat cadre, la SNCB et IFB n'ont pas soumis le plan de restructuration à l'approbation du gouvernement belge, car cela aurait violé l'autonomie commerciale de la SNCB.
147. La Commission considère que cela n'a pas pour conséquence de rendre cet indice d'imputabilité inopérant: il paraît exclu que les deux parties au contrat, la SNCB et IFB, aient inclus une telle clause dans le contrat, s'il n'y avait pas une prise d'influence du gouvernement belge dans ce sens. Dès lors, le fait que le gouvernement belge n'ait pas insisté à être formellement consulté sur la mise en œuvre de la restructuration ne suffit pas pour exclure une prise d'influence informelle de la part du gouvernement belge lors de la préparation du contrat cadre, qui contient déjà les grandes lignes du sauvetage et de la restructuration.. En tout état de cause, le fait que l'État belge ait omis d'utiliser des moyens de contrôle dont il disposait ne signifie pas que la mesure ne lui soit pas imputable.
b) Articles de presse
148. Des indices pour une intervention du gouvernement belge dans la présente affaire se trouvent aussi dans des articles de presse [26]. Ainsi, un article paru dans La libre Belgique du 19 Mai 2003 [27] cite la cellule presse de la SNCB, qui explique que la Belgique n'avait pas encore notifié les mesures de sauvetage à la Commission le 19 mai 2003, tandis que le contrat cadre avait été signé le 7 avril 2003, par le fait que "le pouvoir fédéral a[vait] son mot à dire ". Dans un article paru en mars 2003 dans www.cheminots.be, Karel Vinck, à l'époque administrateur délégué de la SNCB, est cité à propos des dossiers ABX et IFB comme suit: "Il réclame une marge de manœuvre suffisante pour le management de la société". Cela laisse sous-entendre que l'encadrement de la SNCB considérait que l'État intervenait trop dans ces affaires.
c) Ampleur, contenu, conditions du contrat cadre
149. De manière plus générale, la Commission rappelle que, selon le point 56 de l'arrêt Stardust Marine, précité, "tout autre indice indiquant, dans le cas concret, une implication des autorités publiques ou l'improbabilité d'une absence d'implication dans l'adoption d'une mesure, eu égard également à l'ampleur de celle-ci, à son contenu ou aux conditions qu'elle comporte" doit être pris en compte pour établir l'imputabilité d'une mesure à l'État membre en question. S'agissant en l'espèce d'importantes mesures de restructuration, qui devaient être conditionnées par l'approbation des autorités belges, la Commission considère que l'ampleur, le contenu et les conditions du contrat cadre constituent dans ce cas concret des indices supplémentaires d'imputabilité.
d) Conclusion
150. Par conséquent, la Commission considère, à ce stade, que le soutien financier est imputable à l'État belge en ce qui concerne la période après la conclusion du contrat cadre. Il faut donc analyser si l'aide a conféré un avantage au bénéficiaire, ou si, au contraire, la Belgique a agi comme l'aurait fait un investisseur avisé en économie de marché.
3.1.2. Soutien financier favorisant certaines entreprises
151. S'il s'avère que la décision de la SNCB de ne plus demander le paiement de ses factures à IFB à partir de fin 2000 est imputable à la Belgique, il faudrait analyser si ce soutien aurait était accordé par un investisseur privé en économie de marché.
152. La décision de la SNCB de signer le contrat cadre avec IFB étant imputable à la Belgique, il faut ensuite analyser si la SNCB, en accordant à IFB d'abord un financement de sauvetage et ensuite à un financement de la restructuration, a favorisé IFB par rapport à d'autres entreprises. Tel n'est pas le cas si la SNCB a agi, vis-à-vis d'IFB, comme l'aurait fait un investisseur avisé/un créditeur avisé en économie de marché. Pour effectuer cette deuxième appréciation, il y a lieu de distinguer entre les mesures de sauvetage et les mesures de restructuration.
3.1.2.1. Le non-paiement des factures de la SNCB par IFB entre 2000 et 2003
153. En ce qui concerne le non-paiement des factures de la SNCB par IFB, il faut vérifier si un créancier avisé aurait accepté, à la place de la SNCB, qu'IFB ne paye pas ses factures, ou si un créancier avisé aurait entamé, à la place de la SNCB, une procédure en justice, pour obtenir le paiement de ses factures.
154. À ce titre, il y a d'abord lieu de relever qu'il est une pratique commerciale courante d'accorder à un client qui connaît des problèmes de liquidités momentanés, mais qui est pour le reste en bonne santé économique, un délai de paiement tacite pour ses factures, en attendant le paiement plutôt que de l'assigner tout de suite en justice.
155. Il semble que les difficultés financières de l'entreprise ne sont devenues apparentes que dans le courant de l'année 2002 (voir description de la situation financière ci-dessus). Le fait qu'IFB ait obtenu un prêt de plus de 4 millions EUR de la part de la banque commerciale […] en 2001 à un taux de marché, et que les fonds propres d'IFB étaient de 28 millions EUR à la fin de l'année 2001 pointent aussi dans cette direction.
156. Cependant, la Commission ne peut pas exclure à ce stade que la SNCB en tant que société mère d'IFB aurait du se rendre compte des problèmes d'IFB plus en amont, durant l'année 2001.
157. C'est donc au plus tôt à partir de 2001 qu'un investisseur privé aurait agi de manière plus prudente. Il est difficile de dire à partir de quand un créancier privé aurait cherché à obtenir un remboursement de ses créances ou des sécurités additionnelles; à ce stade, la Commission considère que ce moment était venu au plus tard le 19 septembre 2002, quand l'administrateur délégué d'IFB a chargé deux réviseurs de rédiger un rapport spécial sur la situation financière d'IFB.
158. Ce processus a mené au développement du contrat cadre, qui prévoit explicitement des mesures de sauvetage et de restructuration. En continuant à fournir à IFB des prestations de transport par chemin de fer, la SNCB a accordé au plus tôt courant 2001 et au plus tard depuis le 19 septembre 2002 des avantages économiques à IFB, qui doivent être considéré comme des aides d'État. En ne poursuivant pas IFB devant la justice afin d'obtenir le paiement des factures datant de 2000 et de 2001 au plus tard à partir de ce moment, la SNCB a aussi accordé un avantage à IFB en ce qui concerne le non-paiement de ces factures.
159. La SNCB a donc accordé de facto une aide à IFB au plus tôt depuis 2001, au plus tard depuis le 19 septembre 2002; cette aide n'a été que formalisée par le contrat cadre.
3.1.2.2. Les mesures de sauvetage
160. Les mesures de sauvetage ont été décrites ci-dessus dans la partie 2. Pour rappel, il s'agissait de:
- l'octroi d'un délai de paiement pour des dettes de 63 millions d'euros;
- l'octroi d'une facilité de crédit de 15 millions d'euros;
- l'octroi d'une avance récupérable de 5 millions d'euros.
161. Parmi ces mesures, il y a lieu de distinguer entre les actions que la SNCB a prises en tant que créancier d'IFB, à savoir l'octroi du délai de paiement pour les dettes déjà existantes de 63 millions d'euros, et les actions que la SNCB a pris en tant qu'investisseur en IFB, à savoir l'octroi d'une nouvelle facilité de crédit de 15 millions EUR et l'octroi d'une nouvelle avance récupérable de 5 millions EUR.
162. Comme l'explique l'avocat général Poiares Maduro, "le critère du créancier privé ne doit pas être confondu avec celui […] de l'investisseur privé. Tandis que l'investisseur prétend réaliser un bénéfice en intervenant auprès des entreprises concernées, le créancier cherche à obtenir le paiement des sommes qui lui sont dues par un débiteur connaissant des difficultés financières. […] Dans ce cas, le critère décisif n'est donc pas de savoir s'il existe un avantage économique, mais de savoir si cet avantage correspond à un traitement plus favorable que celui qui serait accordé, dans des conditions similaires, par un créancier privé à son entreprise débitrice" [28].
163. Il y a donc lieu d'analyser dans la suite d'abord si la Belgique a agi comme un créancier avisé en économie de marché en ce qui concerne l'octroi du délai de paiement, et ensuite si la Belgique a agi comme l'aurait fait un investisseur avisé en économie de marché en ce qui concerne l'octroi de la facilité de crédit et de l'avance récupérable.
a) La SNCB a-t-elle agi comme l'aurait fait un créancier avisé en économie de marché en accordant le délai de paiement ?
164. Selon le Tribunal, il faut comparer le comportement de l'État à celui d'"un créancier privé cherchant à obtenir le paiement des sommes qui lui sont dues par un débiteur connaissant des difficultés financières" [29]. La décision à laquelle le créancier SNCB était confronté dans le cas d'espèce était donc de déterminer si un créancier avisé aurait préféré mettre IFB en faillite plutôt que de lui accorder un délai de paiement.
165. Le contrat cadre a été signé le 7 avril 2003, mais des délais de paiement pouvant constituer des aides d'État avaient été accordés dès 2001. Il faut placer l'analyse sous l'angle des faits connus de la SNCB à ce moment [30].
166. Pour l'année 2002, IFB avait enregistré des pertes d'exploitation d'EUR 47,4 millions, dont 34 millions étaient des dépréciations spécifiques déjà constatées au niveau des charges d'exploitation, et des pertes exceptionnelles de EUR 59,369 millions. Les pertes exceptionnelles étaient surtout dues à des moins-values dans un certain nombre de filiales, principalement françaises. A cause de ces pertes, IFB avait des fonds propres négatifs de EUR 84,07 millions à la fin de l'exercice 2002.
167. Dans l'hypothèse d'une faillite, la SNCB, qui détenait 89,03 % du capital social de l'IFB, n'aurait eu éventuellement accès aux résultats de la liquidation qu'après satisfaction des créanciers. De plus, ses créances découlant des factures non payées n'auraient probablement été satisfaites qu'en partie.
168. C'est d'ailleurs pour cela que, dans ses comptes annuels de 2002, la SNCB avait mis la valeur des ces titres et créances à zéro, [31] au motif que, "compte tenu de la situation financière de ce groupe [i.e. IFB] et dans l'attente d'une finalisation du plan de restructuration de ce groupe au sein du secteur fret de la SNCB, les créances commerciales et les commandes en cours que la SNCB possède [doivent être] comptabilisées comme douteuses." [32].
169. La SNCB était de loin le créancier le plus important d'IFB à ce moment: selon les comptes annuels d'IFB de 2003, IFB avait des dettes auprès des établissements de crédit de 12 millions d'euros, et des dettes vis-à-vis ses fournisseurs, donc principalement vis-à-vis de la SNCB, de 108 millions d'euros.
170. Dans l'hypothèse d'une faillite, la SNCB aurait aussi dû réintégrer 50 employés, qui avaient été détachés à IFB, au sein de l'entreprise. Dans un contexte où la SNCB essaie de réduire le nombre de ses employés, cela aurait constitué un désavantage supplémentaire pour la SNCB.
171. En conclusion, la mise en faillite d'IFB aurait engendré des coûts supplémentaires pour la SNCB, sans qu'elle ait la certitude de voir ses créances honorées.
172. Cependant, il se pose la question de savoir si l'alternative, à savoir l'octroi du délai de paiement, accompagnée du paiement des intérêts moratoires au taux légal ou au taux de marché (selon les dettes, cf. description ci-dessus), d'un engagement de ne pas invoquer la prescription des créances et de nouveaux investissements, permettait à la SNCB de raisonnablement s'attendre à ce qu'IFB une rentabilité suffisante pour rémunérer ses nouveaux investissements à un niveau acceptable pour un investisseur privé en économie de marché et pour améliorer les perspectives de satisfaction des créances antérieures à moyen ou longue terme.
173. En avril 2003, au moment de la conclusion du contrat cadre, IFB avait commencé sa restructuration, qui impliquait d'un côté une restructuration en profondeur des opérations d'IFB lui-même, d'un autre côté une stratégie de désinvestissement pour endiguer les pertes opérationnelles des filiales françaises, comme décrit ci-dessus dans la partie 2.3.2.
174. En ce qui concerne les chances pour un retour à la rentabilité économique d'IFB, force est de constater que les difficultés financières étaient notamment dues à sa stratégie d'expansion en France, et seulement dans une moindre mesure à des problèmes structurels de IFB Logistics et IFB Terminals..
175. Cependant, le contrat cadre prévoit que le délai de paiement soit accompagné d'une facilité de crédit de 15 millions EUR et d'une avance récupérable de 5 millions EUR. Afin de pouvoir raisonnablement s'attendre aux paiements des créances, la SNCB devait donc investir de capital frais. Dès lors, un investisseur privé n'aurait accordé un délai de paiement que si son investissement additionnel de 20 millions de capital frais constituait un investissement avec un rendement acceptable.
176. Le délai de paiement doit donc être analysé ensemble avec les décisions d'investissement prises par la SNCB dans le contrat cadre, car les mesures forment un ensemble au sens de la jurisprudence BP Chemicals [33].
b) La SNCB a-t-elle agi comme l'aurait fait un investisseur avisé en économie de marché en accordant l'octroi d'une facilité de crédit et l'octroi d'une avance récupérable?
177. En ce qui concerne l'octroi de la facilité de crédit de 15 millions d'EUR, et l'octroi de l'avance récupérable de 5 millions d'EUR, la SNCB n'agissant pas en tant qu'investisseur n'était pas un créancier d'IFB, mais avait le libre choix d'investir cet argent dans IFB ou bien ailleurs, et était donc un investisseur.
178. Il convient donc d'analyser si la SNCB a agi comme l'aurait fait un investisseur avisé en économie de marché. Selon la jurisprudence de la Cour, il y a lieu d'apprécier si, dans des circonstances similaires, un investisseur privé d' une taille qui puisse être comparée à celle de la SNCB aurait pu être amené à procéder aux apports de capitaux de cette importance [34].
179. La Cour a précisé que si le comportement de l' investisseur privé, auquel doit être comparée l'intervention de l'investisseur public poursuivant des objectifs de politique économique, n'est pas nécessairement celui de l'investisseur ordinaire plaçant des capitaux en vue de leur rentabilisation à plus ou moins court terme, il doit, au moins, être celui d' un holding privé ou d' un groupe privé d' entreprises poursuivant une politique structurelle, globale ou sectorielle, et guidé par des perspectives de rentabilité à plus long terme [35]. Le Tribunal a défini de manière plus précise la méthode d'évaluation à suivre par la Commission. Il a précisé que la Commission est obligée "de faire une analyse complète de tous les éléments pertinents de l'opération litigieuse et de son contexte" afin de savoir si l'État a agi comme l'aurait fait un investisseur avisé en économie de marché [36].
180. Il faut donc établir, dans le cas d'espèce, la rentabilité de l'intervention de la SNCB, ce qui suppose de regarder si l'investissement dans IFB devait dégager une marge bénéficiaire normale.
181. La SNCB a, à travers les mesures de sauvetage, décidé de mobiliser en avril 2003 20 millions d'EUR dans la société IFB, sous forme de prêt (facilité de crédit de 15 millions d'euros et avance récupérable de 5 millions d'euros).
182. Le contrat cadre, qui accordait les mesures de sauvetage, a été conclu le 7 avril 2003. En ce qui concerne l'investissement de 20 millions d'EUR fait à ce moment au titre de mesure de sauvetage, leur analyse doit donc être placée sous l'angle des faits connus de la SNCB à ce moment [37].
183. Généralement, pour déterminer si un taux d'intérêt pour un prêt correspond aux conditions normales du marché, la Commission établit une comparaison avec la valeur, à la même date, du taux de référence fixé pour l'État membre considéré [38]. Les prêts en espèces étant rémunérés au taux de marché et en partie même à un taux supérieur au taux de marché, il semble de prime abord ne pas y avoir un élément d'aide. Cependant, il faut constater qu'IFB était, au moment de l'octroi des prêts, une entreprise confrontée à de très graves difficultés financières. Il semble invraisemblable qu'il aurait pu obtenir, sur le marché de capital, un prêt à des conditions comparables à celles offertes par la SNCB. Une banque aurait donc très probablement demandé un taux de rémunération supérieur au taux demandé par la SNCB ou aurait même refuser d'octroyer un prêt à IFB. D'ailleurs, la décision de la SNCB d'accorder un délai de paiement sur ses créances existantes est un indice de la difficulté que devait rencontrer IFB à se refinancer ailleurs.
184. Les autorités belges considèrent que le fait qu'IFB ait obtenu en juillet 2003, donc après la conclusion du contrat cadre, un prêt sur 2 millions EUR de la part de la banque ING démontre que les banques privées ne demandaient pas une rémunération supérieure au taux de marché.
185. Cet argument n'est pas convaincant, pour deux raisons. D'abord, le montant de 2 millions EUR est très faible comparé aux engagements de la SNCB, qui prévoyaient des investissements de 20 millions EUR ainsi que la possibilité de convertir les créances de 63 millions EUR en capital. Ensuite, ING n'a accordé ce prêt qu'après que la SNCB s'était engagée de garantir la survie d'IFB, en signant le contrat cadre.
186. Dès lors, force est de constater que la SNCB, en accordant les prêts à un taux inférieur au taux qui aurait été adéquat pour la situation financière d'IFB, n'a pas agi comme l'aurait fait un investisseur avisé en économie de marché.
187. Le gouvernement belge considère pour sa part que la SNCB a agi comme l'aurait fait toute société mère, dont une filiale est en difficulté, sans préciser davantage cet argument. La Commission observe à cet égard que la Belgique n'a pas démontré cet argument et en particulier, n'a pas démontré que le nouvel investissement était nécessaire pour pouvoir espérer en retirer un montant supérieur à l'ensemble de ses créances existantes et nouvelles.
c) Conclusion en ce qui concerne les mesures de sauvetage
188. En conclusion, la Commission considère, à ce stade, que la SNCB n'a pas agi comme l'aurait fait un investisseur avisé en économie de marché en ce qui concerne l'octroi de la facilité de crédit de 15 millions d'euros et en ce qui concerne l'octroi de l'avance récupérable de 5 millions d'euros. Puisque l'octroi du délai de paiement n'était raisonnable pour un créancier privé que si l'investissement l'était aussi, il s'ensuit que la SNCB n'a pas non plus agi comme l'aurait fait un créancier avisé en économie de marché en ce qui concerne l'octroi d'un délai de paiement pour IFB.
3.1.2.3. Les mesures de restructuration
189. Les mesures de restructuration ont été décrites ci-dessus dans la partie 2. Pour rappel, il s'agissait de:
- La conversion des dettes de 63 millions d'euros pour lesquelles un délai de paiement a été octroyé en capital social.
- La conversion de la facilité de crédit de 15 millions d'euros en capital social.
- La conversion des intérêts sur le délai de paiement capitalisés de 11 millions d'euros en capital social.
- La conversion des intérêts sur l'avance récupérable capitalisés de 2,5 millions d'euros en capital social.
- L'injection de 5 millions d'euros par l'apport en nature de la participation de la SNCB dans TRW.
190. En total, l'augmentation de capital sera donc de 96,5 millions d'euros. IFB ayant en ce moment des fonds propres négatifs de 72,6 millions d'euros, l'augmentation de capital lui laissera des capitaux propres de 23,8 millions d'euros.
191. Parmi ces mesures, il y a lieu de distinguer entre les actions que la SNCB a pris en tant que créancier d'IFB, à savoir la conversion des dettes existantes de 63 millions d'euros et des intérêts liés de 11 millions d'euros en capital social, et les actions que la SNCB a pris en tant qu'investisseur en IFB, à savoir la conversion de la facilité de crédit de 15 millions EUR et des intérêts liés de 2,5 millions d'euros en capital social et l'injection de capital frais de 5 millions EUR.
192. En ce qui concerne la conversion de la facilité de crédit de 15 millions en capital social, il pourrait être objecté qu'au moment de la conversion, la SNCB n'était plus un investisseur, mais un créancier. Cela ignore cependant le fait qu'il était prévu dans le contrat cadre de convertir éventuellement la facilité de crédit en capital social (voir description dans la partie 2), et que la facilité de crédit n'était qu'une mesure temporaire. Dès lors, il faut considérer que la conversion de la facilité de crédit en capital social doit être comparée à un investissement.
a) La SNCB a-t-elle agi comme l'aurait fait un créancier avisé en économie de marché en convertissant ses créances de 63 millions d'euros et les intérêts liés de 11 millions d'euros en capital social?
193. En convertissant ses créances de 63 millions d'euros et les intérêts liés de 11 millions d'euros en capital social, la SNCB renonce au paiement de ses dettes. En contrepartie, elle aura droit aux dividendes qu'IFB payera à ses propriétaires, et acquiert des parts sociales.
194. Comme démontré ci-dessus, il y a lieu de considérer, à ce stade, qu'un créancier privé avisé n'aurait pas accordé le délai de paiement accordé par la SNCB, mais il aurait mis IFB en faillite et aurait essayer d'obtenir le paiement des créances dans le cadre de la procédure collective.
195. Dès lors, un créancier privé avisé n'aurait pas non plus converti ses créances en capital social d'une entreprise qui ne pouvait survivre que s'il injectait en même du capital frais. La SNCB n'a donc pas agi comme l'aurait fait un créancier privé en économie de marché en convertissant ses créances en capital social.
b) La SNCB a-t-elle agi comme l'aurait fait un investisseur avisé en économie de marché en convertissant la facilité de crédit de 15 millions d'euros et les intérêts liés de 2,5 millions d'euros en capital social, et en injectant des capitaux frais de 5 millions d'euros?
196. Il convient d'analyser si la SNCB a agi comme l'aurait fait un investisseur avisé en économie de marché en ce qui concerne la conversion en capital social de la facilité de crédit de 15 millions d'euros et des intérêts liés de 2,5 millions d'euros ainsi que l'augmentation de capital d'IFB à l'hauteur de 5 millions d'EUR.
197. Selon la jurisprudence de la Cour, il y a lieu d'apprécier si, dans des circonstances similaires, un investisseur privé d' une taille qui puisse être comparée à celle de la SNCB aurait pu être amené à procéder aux apports de capitaux de cette importance [39].
198. La Cour a précisé que si le comportement de l' investisseur privé, auquel doit être comparée l'intervention de l'investisseur public poursuivant des objectifs de politique économique, n'est pas nécessairement celui de l'investisseur ordinaire plaçant des capitaux en vue de leur rentabilisation à plus ou moins court terme, il doit, au moins, être celui d' un holding privé ou d' un groupe privé d' entreprises poursuivant une politique structurelle, globale ou sectorielle, et guidé par des perspectives de rentabilité à plus long terme [40]. Le Tribunal a défini de manière plus précise la méthode d'évaluation à suivre par la Commission. Il a précisé que la Commission est obligée "de faire une analyse complète de tous les éléments pertinents de l'opération litigieuse et de son contexte" afin de savoir si l'État a agi comme l'aurait fait un investisseur avisé en économie de marché [41].
199. Il faut donc établir, dans le cas d'espèce, la rentabilité de l'intervention de la SNCB, ce qui suppose de démontrer que l'investissement dans IFB dégagera une marge bénéficiaire normale.
200. Par sa décision de convertir la facilité de crédit de 15 millions d'euros et les intérêts liés de 2,5 millions d'euros, qui était une mesure temporelle de sauvetage, en une augmentation de capital, la SNCB pérennisera cet investissement.
201. En décidant d'ajouter à cette augmentation de capital la somme de 5 millions d'EUR, elle a décidé de faire un investissement supplémentaire de 5 millions d'EUR.
202. La conversion de la facilité de crédit de 15 millions d'euros et des intérêts liés de 2,5 millions d'euros en capital social et le principe de l'augmentation de capital additionnel de 5 millions d'euros ont été décidés au printemps 2005; leur analyse doit donc être placée sous l'angle des faits connus de la SNCB à ce moment [42].
203. Ces deux mesures doivent être comparées à la décision d'un investisseur privé de participer à une augmentation de capital d'IFB.
204. La Commission note d'abord l'absence d'un investisseur privé, qui aurait participé, avec la SNCB, à l'augmentation de capital d'IFB.
205. Le gouvernement belge considère que la SNCB a agi comme l'aurait fait un investisseur avisé en économie de marché. Pour démontrer cela, il donne l'exemple suivant: Si la SNCB avait recapitalisé IFB au 1er janvier 2004 par conversion des dettes d'IFB vis-à-vis de la SNCB (de l'ordre de 79 millions EUR à ce moment) et d'un apport supplémentaire de l'ordre de 21 millions EUR, IFB aurait disposé de fonds propres en début d'exercice d'environ 16 millions EUR. En outre, elle aurait réalisé un bénéfice d'exploitation de 5,74 millions EUR (rendement de 36 % sur fonds propres) et un bénéfice courant avant impôts de plus de 7,18 millions EUR (45 % sur fonds propres). La marge opérationnelle bénéficiaire sur le chiffre d'affaires aurait alors été de l'ordre de 7 % en 2004. Le résultat de 2004 étant fortement influencé par l'utilisation et la reprise de certaines provisions faites en 2001 et 2002 pour les pertes attendues des filiales françaises, le gouvernement belge propose de neutraliser ces événements extraordinaires, ce qui laisse une marge opérationnelle bénéficiaire sur le chiffre d'affaire de 2,9 % pour 2004. Le gouvernement belge n'a pas transmis d'estimation pour les bénéfices d'IFB pour les années suivantes.
206. La Commission considère que le développement d'IFB depuis 2003 témoigne certes de la viabilité économique d'IFB. Cependant, le test de l'investisseur privé en économie de marché vise non seulement la viabilité économique d'une entreprise, mais la rentabilité de celle-ci. Selon la Cour, "il convient d'apprécier si, dans des circonstances similaires, un associé privé se basant sur les possibilités de rentabilités prévisibles, abstraction faite de toute considération de caractère social ou de politique régionale ou sectorielle, aurait procédé à un tel apport de capital" [43]. Cette possibilité de rentabilité doit, "au moins, être celui d' un holding privé ou d' un groupe privé d' entreprises poursuivant une politique structurelle, globale ou sectorielle, et guidé par des perspectives de rentabilité à plus long terme" [44].
207. La rémunération normale s'apprécie en tenant compte notamment de la rentabilité moyenne des concurrents. A cet égard, le gouvernement belge a informé la Commission que le chiffre d'affaires et la rentabilité des concurrents d'IFB était la suivante (en millions EUR):
| Chiffres d'affaires 2003 | Bénéfice en 2003 | Bénéfice en 2003 en % | Chiffres d'affaires 2004 | Bénéfice en 2004 | Bénéfice en 2004 en % |
CEMAT | 164,1 | 1,4 | 0,9 | 176,6 | 3,9 | 2,2 |
CNC | 193,5 | - 17,0 | - 8,8 | 164,4 | - 20,6 | - 12,5 |
HUPAC | 195,2 | 5,7 | 2,9 | 225,6 | 6,0 | 2,7 |
ICF | 276,5 | 0,5 | 0,2 | 261,1 | - 3,7 | - 1,4 |
Kombiverkehr | 289,2 | 0,8 | 0,3 | n/a | n/a | n/a |
Novatrans | 109,0 | - 7,1 | - 6,5 | 102,5 | - 5,5 | - 5,4 |
208. Il faut noter que ce tableau ne donne pas le rendement pour les grands concurrents Hesse-Noordnatie, Danzas, Ziegler, et Schenker, et que la plupart des entreprises citées par le gouvernement belge ont réalisé des pertes en 2004.
209. Les chiffres fournis par le gouvernement belge ne peuvent donc pas être utilisés pour apprécier si le rendement d'IFB est un rendement normal. En absence d'un chiffre de comparaison adéquate, la Commission constate qu'un rendement de 2,9 % est un rendement très faible, car il correspond à peu près au rendement des obligations gouvernementales. Cependant, un investissement dans IFB présente un risque nettement supérieur au risque des obligations gouvernementales.
210. Dès lors, la Commission considère que le rendement d'un investissement dans IFB ne serait pas suffisant pour convaincre un investisseur avisé en économie de marché de procéder à un tel investissement. Un investisseur avisé n'aurait donc pas procédé aux investissements que la SNCB a faits dans IFB.
c) Conclusion en ce qui concerne les mesures de restructuration
211. La Commission considère donc, à ce stade, que la SNCB n'a pas agi comme l'aurait fait un créancier privé en économie de marché, en convertissant les dettes de 63 millions d'euros et les intérêts liés de 11 millions d'euros en capital social. Elle considère que la SNCB n'a pas non plus agi comme l'aurait fait un investisseur avisé en économie de marché en ce qui concerne la conversion de la facilité de crédit de 15 millions d'euros et les intérêts liés de 2,5 millions d'euros en capital social et en ce qui concerne l'injection de 5 millions d'euros dans IFB.
3.1.3. Distorsion de concurrence et affectation des échanges entre les Etats membres
212. La Commission doit analyser la situation du marché concerné et les parts de marché des bénéficiaires sur ce marché, ainsi que l'impact que le soutien financier aura sur la situation de concurrence [45].
213. En l'espèce, le soutien financier a été accordé à une entreprise active sur des marchés ouverts à la concurrence, qui est en situation de concurrence avec d'autres acteurs de plusieurs Etats membres, comme démontré ci-dessus dans la partie "description". Le soutien financier fausse ou menace de fausser donc la concurrence, et menace d'affecter ou affecte les échanges entre les États membres.
3.1.4. Conclusion: présence d'une aide d'État
214. En conclusion, la Commission considère, à ce stade, que la SNCB n'a pas agi comme l'aurait fait un créancier avisé en économie de marché en ce qui concerne le délai de paiement et la conversion des créances de 63 millions d'euros dues et non payées le 31 janvier 2003, et qu'elle n'a pas agi comme l'aurait fait un investisseur avisé en économie de marché en ce qui concerne l'octroi d'une facilité de crédit de 15 millions d'euros, l'octroi d'une avance récupérable de 5 millions d'euros, la conversion de la facilité de crédit de 15 millions d'euros en capital social ainsi qu'en ce qui concerne l'injection de capitaux frais de 5 millions EUR.
3.2. Compatibilité de l'aide
215. L'art. 87 §3 lit. c du traité CE prévoit que "peuvent être considérés comme compatibles avec le marché commun les aides destinées à faciliter le développement de certaines activités ou de certaines régions économiques, quand elles n'altèrent pas les conditions des échanges dans une mesure contraire à l'intérêt commun."
216. L'aide accordée par la Belgique à travers la SNCB pourrait être compatible avec le marché commun en vertu de l'article 87 § 3 c, tel qu'interprété par la Commission dans ses lignes directrices communautaires concernant les aides d'État au sauvetage et à la restructuration d'entreprises en difficulté (ci-après: les lignes directrices) [46].
217. Afin de pouvoir bénéficier d'aides au sauvetage et d'aides à la restructuration, une entreprise doit d'abord être éligible pour l'application des lignes directrices. Pour être éligible, une entreprise ne doit pas être une entreprise nouvellement créée, et doit être une entreprise en difficulté.
218. Pas d'entreprise nouvellement créée. Le point 12 des lignes directrices de 2004 précisent à ce propos, reprenant et précisant les lignes directrices de 1999, point 7:
Aux fins des présentes lignes directrices, une entreprise nouvellement créée ne peut bénéficier d'aides au sauvetage ou à la restructuration, même si sa position financière initiale est précaire. Tel est notamment le cas lorsqu'une nouvelle entreprise naît de la liquidation d'une entreprise préexistante ou de la reprise de ses seuls actifs. Une entreprise est en principe considérée comme nouvellement créée pendant les premières trois années qui suivent son entrée en activité dans le domaine concerné.
219. Il se pose donc d'abord la question de savoir si IFB est une entreprise nouvellement créée. Comme décrit ci-dessus dans la partie 2, IFB a été créée le 1er avril 1998, par la fusion de trois autres sociétés, qui avaient été créées en 1906, 1923 et 1967 respectivement.
220. Comme expliqué ci-dessus dans la partie 3.1.2.1, le premier avantage octroyé par la SNCB à IFB était l'octroi tacite d'un délai de paiement pour les services prestés par la SNCB, mais non payé par IFB, à partir de l'année 2001 au plus tôt.
221. L'entreprise IFB a été créée le 1er avril 1998 par la fusion de trois sociétés préexistantes. A ce stade, il n'est pas clair si l'entreprise continue la personnalité juridique d'une de ces trois sociétés. Si telle était le cas, IFB serait clairement une entreprise de plus de trois ans en 2001.
222. Si IFB ne continuait pas la personnalité juridique d'une de ces sociétés, mais était une entreprise nouvellement créée le 1er avril 1998, il dépasserait l'age de trois ans le 1er avril 2001. Dans cette hypothèse, elle ne serait éligible pour des aides à la restructuration qu'à partir du 1er avril 2001.
223. La Commission exprime donc des doutes si IFB est une entreprise éligible aux aides à la restructuration, et invite les autorités belges de lui fournir tout renseignement utile afin de vérifier si IFB, vu ces considérations, est une entreprise éligible pour les aides à la restructuration.
224. Entreprise en difficulté. Il n'existe pas de définition communautaire de l'entreprise en difficulté. Les lignes directrices considèrent dans leur paragraphe 5 (version de 1999) respectivement 10 (version de 2004) qu'une société à responsabilité limitée, comme l'est IFB, qui est une société par actions, est en tout cas considérée comme en difficulté lorsque plus de la moitié de son capital souscrit a disparu et que plus du quart de ce capital a été perdu au cours des douze derniers mois. Les comptes annuels de 2002 montrent un capital souscrit de EUR 48 millions et des pertes courantes avant impôts de 50 millions EUR. Par conséquent, le capital social avait disparu quant la SNCB avait décidé en avril 2003 d'accorder des aides au sauvetage. Plus de la moitié du capital souscrit ayant disparu à ce moment, dont plus d'un quart dans les douze derniers mois, IFB est une entreprise en difficulté au sens des lignes directrices.
225. Les lignes directrices sont donc applicables. Il y a lieu d'analyser si les aides accordées par la SNCB à IFB les ont respectées. A cet égard, il y a lieu d'abord d'analyser si au moins une partie des aides ont été des aides au sauvetage compatibles avec les lignes directrices.
3.2.1. Compatibilité en tant qu'aides au sauvetage
226. Seules les mesures consistant en une aide de trésorerie pourraient être compatibles en tant qu'aides au sauvetage. Dans le présent cas, les aides de trésorerie sont l'accord d'un délai de paiement tacite au plus tôt en 2001, au plus tard le 19 septembre 2002, devenu délai de paiement exprès dès le 7 avril 2003, la facilité de crédit et l'avance récupérable.
227. Il se pose d'abord la question de savoir qu'elle version des lignes directrices est applicable. La dernière version de ces lignes directrices est entrée en vigueur le 10 octobre 2004. Elle dispose dans son point 7 "date d'application et durée":
102. La Commission appliquera les présentes lignes directrices à partir du 10 octobre 2004 et jusqu'au 9 octobre 2009.
103. Les notifications enregistrées par la Commission avant le 10 octobre 2004 seront examinées au regard des critères en vigueur au moment de la notification.
104. La Commission examinera la compatibilité avec le marché commun de toute aide au sauvetage ou à la restructuration octroyée sans son autorisation et donc en violation de l'article 88, paragraphe 3, du traité sur la base des présentes lignes directrices si l'aide, ou une partie de celle-ci, a été octroyée après leur publication au Journal officiel de l'Union européenne. Dans tous les autres cas elle fera l'examen sur la base des lignes directrices applicables au moment de l'octroi de l'aide.
228. Les aides de trésorerie ont été octroyées au plus tôt en 2001, ou courant 2002 et dans leur ensemble le 7 avril 2003, sans notification préalable à la Commission et donc en violation de l'article 88 § 3 du traité CE. L'appréciation de leur compatibilité en tant qu'aides au sauvetage, en faisant abstraction des autres mesures à considérer comme des aides à la restructuration, se fera donc sur base des lignes directrices de 1999.
229. Le paragraphe 23 des lignes directrices de 1999, qui sont d'application pour les aides au sauvetage que la SNCB a accordées à IFB éventuellement en 2001, certainement en 2002 et 2003, définit les cinq conditions pour qu'une aide au sauvetage puisse être compatible avec le marché commun. Ces cinq conditions sont les suivantes:
a) consister en des aides de trésorerie prenant la forme de garanties de crédits ou de crédits. Dans les deux cas de figures, le crédit doit être soumis à un taux au moins comparable aux taux observés pour des prêts à des entreprises saines et notamment aux taux de référence adoptés par la Commission;
b) être liées à des crédits dont la durée de remboursement qui suit le dernier versement à l'entreprise des sommes prêtées ne dépasse pas douze mois; le remboursement du prêt lié à l'aide au sauvetage peut éventuellement être couvert par l'aide à la restructuration qui serait autorisée ultérieurement par la Commission;
c) être justifiées par des raisons sociales aiguës et ne pas avoir des effets graves de débordement ("spillover") négatif dans d'autres États membres;
d) être accompagnées, lors de leur notification, d'un engagement de l'État membre de transmettre à la Commission, dans un délai de six mois à compter de l'autorisation de l'aide au sauvetage, soit un plan de restructuration, soit un plan de liquidation, soit la preuve que le prêt a été intégralement remboursé et/ou qu'il a été mis fin à la garantie;
e) se borner dans leur montant à ce qui est nécessaire pour l'exploitation de l'entreprise (par exemple, la couverture des charges salariales ou des approvisionnements courants) pendant la période pour laquelle l'aide est autorisée.
3.2.1.1. Aide consistant en une aide de trésorerie
230. Pour rappel, les mesures de sauvetage consistent en un délai de paiement pour des créances d'une valeur totale de 63 millions EUR, en une avance récupérable de 5 millions EUR, qui a été accordée, mais non pas utilisée par IFB, et en une facilité de crédit de 15 millions EUR.
231. Par conséquent, l'aide consiste en une aide de trésorerie, qui se compose d'un délai de paiement, d'une avance récupérable et d'une facilité de crédit.
3.2.1.2. Aide liée à des crédits dont la durée de remboursement qui suit le dernier versement à l'entreprise ne dépasse pas douze mois
232. La durée de remboursement prévue par le contrat cadre est de douze mois. Néanmoins, le gouvernement belge a informé la Commission que la durée a été tacitement prolongée entre les parties jusqu'au moment de l'augmentation de capital.
233. De plus, l'avantage résultant du délai de paiement a déjà été octroyé au plus tôt courant l'année 2001, au plus tard le 19 décembre 2002. La Commission considère donc que ce critère n'est pas rempli, et que les aides de trésorerie ne peuvent pas être autorisées comme des aides au sauvetage.
3.2.1.3. Conclusion
234. En conclusion, la Commission considère, à ce stade, que les aides de trésorerie que la SNCB a accordées à IFB ne sont pas compatibles avec le marché commun en vertu de l'article 87 § 3 c du traité en tant qu'aides au sauvetage. Elles pourraient néanmoins être compatibles avec le marché commun en tant qu'aides à la restructuration.
3.2.2. Compatibilité des aides à la restructuration
235. Il se pose de nouveau la question de savoir quelle version des lignes directrices est applicable. Pour rappel, la dernière version de ces lignes directrices est entrée en vigueur le 10 octobre 2004. Elle dispose dans son point 7 "date d'application et durée":
102. La Commission appliquera les présentes lignes directrices à partir du 10 octobre 2004 et jusqu'au 9 octobre 2009.
103. Les notifications enregistrées par la Commission avant le 10 octobre 2004 seront examinées au regard des critères en vigueur au moment de la notification.
104. La Commission examinera la compatibilité avec le marché commun de toute aide au sauvetage ou à la restructuration octroyée sans son autorisation et donc en violation de l'article 88, paragraphe 3, du traité sur la base des présentes lignes directrices si l'aide, ou une partie de celle-ci, a été octroyée après leur publication au Journal officiel de l'Union européenne. Dans tous les autres cas elle fera l'examen sur la base des lignes directrices applicables au moment de l'octroi de l'aide.
236. Les aides de trésorerie ont été octroyées en partie au plus tôt courant l'année 2001, au plus tard le 19 septembre 2002, et dans leur ensemble le 7 avril 2003, sans notification préalable à la Commission et donc en violation de l'article 88 § 3 du traité CE. Leur conversion en capital était prévue depuis la conclusion du contrat cadre le 7 avril 2003, mais n'a pas eu lieu jusqu'à ce jour.
237. Puisque la SNCB a mis en œuvre l'aide de trésorerie sans accord préalable de la Commission, il faut appliquer le point 104 des lignes directrices de 2004 pour déterminer les lignes directrices applicables au présent cas. L'aide de trésorerie a été accordé en partie au plus tôt courant l'année 2001, au plus tard le 19 septembre 2002, et pour le reste le 7 avril 2003, et donc avant la publication des lignes directrices de 2004 au Journal officiel. Si l'aide était limitée aux aides de trésorerie, il faudrait donc appliquer les lignes directrices de 1999, car l'octroi de l'aide aurait eu lieu avant la publication des lignes directrices de 2004.
238. Cependant, la conversion des créances en capital constitue une mesure ultérieure, qui modifie la nature des avantages antérieurement consentis à IFB. A cet égard, le contrat-cadre fait état de l'intention des parties de procéder à cette conversion, mais sous réserve notamment de l'approbation du plan de restructuration par les deux Conseils d'administration et par l'État belge, ainsi que de l'approbation par les actionnaires d'IFB. A ce stade, il n'est donc pas démontré que la mesure a été définitivement octroyée avant la publication des lignes directrices de 2004, en ce sens que l'autorité compétente s'est engagée par un acte juridiquement contraignant à accorder l'aide avant cette date [47]. Si tel n'était pas le cas, et considérant que la conversion des créances en capital n'a pas été notifiée avant le 10 octobre 2004, les lignes directrices de 2004 seraient applicables.
239. Les autorités belges ont notifié à la Commission, par lettre du 28 janvier 2005, que la SNCB devrait accorder un nouveau avantage de 5 millions EUR sous forme d'une augmentation de capital par apport en nature en 2005 ou 2006. Dans un tel cas, une aide aurait été notifiée après le 10 octobre 2004. En vertu du point 103 des lignes directrices de 2004, il faudrait alors appliquer les lignes directrices de 2004 à cette nouvelle notification.
240. La Commission est tenue de statuer sur l'ensemble des mesures qui lui ont été notifiées; elle base donc son appréciation juridique sur les lignes directrices de 2004. Cependant, elle attire l'attention du gouvernement belge et des parties tiers intéressées sur le fait que si la SNCB décide de ne pas accorder de nouveau avantage à IFB, et si la preuve était apportée que la SNCB s'était engagée à convertir ses créances en capital avant la publication des lignes directrices de 2004, la Commission devrait examiner dans sa décision finale les aides accordées par la SNCB à IFB sur la base des lignes directrices de 1999. Les doutes exprimés ci-dessous sur la base du texte de 2004 valent aussi, mutatis mutandis, pour le texte de 1999.
241. Le point 3.2.2 des lignes directrices de 2004 énonce les conditions pour l'autorisation d'une aide à la restructuration. Les conditions sont les suivantes:
- Le plan de restructuration doit permettre de rétablir dans un délai raisonnable la viabilité à long terme de l'entreprise
- Des mesures doivent être prises pour atténuer, autant que possible, les conséquences défavorables de l'aide pour les concurrents.
- L'aide doit être limitée au strict minimum nécessaire pour permettre la restructuration.
- La Commission doit être mise en mesure de s'assurer du bon déroulement du plan de restructuration, au travers de rapports réguliers et détaillés.
- Les aides à la restructuration ne doivent être accordées qu'une seule fois.
3.2.2.1. Plan de restructuration
242. L'octroi des aides à la restructuration est conditionné par la mise en œuvre d'un plan de restructuration, qui doit permettre de rétablir dans un délai raisonnable la viabilité à long terme de l'entreprise, sur la base d'hypothèses réalistes concernant les conditions d'exploitation future.
243. Les paragraphes 32 à 34 des lignes directrices précisent les conditions minimales pour l'acceptation d'un plan de restructuration par la Commission. Le plan de restructuration doit notamment contenir les éléments suivants:
- Une étude de marché.
- Une description des circonstances ayant entraîné les difficultés de l'entreprise, permettant d'évaluer si les mesures proposées dans le plan sont adaptées pour permettre le retour à la viabilité de l'entreprise.
- Une description des changements prévus pour que l'entreprise puisse, une fois la restructuration achevée, couvrir tous ses coûts, y compris les coûts d'amortissement et les charges financières, et affronter la concurrence en ne comptant plus que sur ses seules forces.
244. Le gouvernement belge a présenté un plan de restructuration pour IFB en décembre 2003, et détaillé ce plan dans la suite, qui contient ces éléments et dont les détails sont décrits dont la partie 2 de la présente décision.
245. Ce plan contient une analyse des marchés de la logistique et du transbordement du fret, ainsi que la position d'IFB sur ce marché. Il décrit les raisons pour les difficultés d'IFB, qui ont leur racine notamment dans une politique d'expansion en France, qui a été mal menée, et dans une mauvaise gestion des activités "IFB Terminals" et "IFB Logistics".
246. Finalement, ce plan décrit les changements prévus pour que l'entreprise puisse, une fois la restructuration achevée, couvrir tous ses coûts en ne comptant que sur ses seules forces. Les changements prévus sont notamment la cessation des filiales françaises, ainsi qu'une restructuration des activités "IFB Logistics" et "IFB Terminals". Ces restructurations impliquent notamment une concentration sur les offres rentables, une nouvelle convention collective, et une réorganisation des terminaux.
247. La mise en œuvre de ce plan de restructuration a été terminée, avec succès, en 2005.
3.2.2.2. Viabilité économique de l'entreprise
248. Le plan de restructuration contient les mesures prévues par IFB pour retrouver sa viabilité économique. Comme décrit ci-dessus, IFB n'a pas su atteindre ses objectifs financiers en 2003. Cependant, dès l'exercice 2004, il a pu atteindre les objectifs fixés par le plan de restructuration, et a même réalisé un bénéfice supérieur à ce qui était prévu. Ce bon développement s'est poursuivi en 2005.
249. IFB a réussi à augmenter sensiblement le volume de fret transporté depuis le début du programme de restructuration (voir description ci-dessus dans la partie 2). Cela explique aussi la croissance de son chiffre d'affaires, de 58 millions d'euros en 2003 à 83 millions d'euros en 2004.
250. L'entreprise IFB a donc su démontrer sa viabilité économique à la fois dans son plan de restructuration, présenté en 2003, et dans ses résultats réalisés depuis lors.
3.2.2.3. Mesures pour atténuer, autant que possible, les conséquences défavorables de l'aide pour les concurrents
251. Des mesures compensatoires doivent être prises pour atténuer, autant que possible, les conséquences défavorables de l'aide pour les concurrents. A défaut, l'aide d'État devrait être considérée comme contraire à l'intérêt commun, et donc incompatible avec le marché commun.
252. Les autorités belges expliquent que, afin d'atténuer, autant que possible, les conséquences défavorables de l'aide pour les concurrents, IFB a pris deux mesures:
- Le retrait de ses activités de transbordement en France.
- La fermeture du terminal de Bressoux en Belgique et la vente des participations dans les terminaux à Bruxelles et à Zeebrugge en Belgique.
253. Ces deux mesures ont eu pour conséquence une baisse de son chiffre d'affaires de 62 millions d'euros en 2002 à 58 millions d'euros en 2003. Cependant, son chiffre d'affaires en 2004 a déjà été supérieur au chiffre d'affaires de 2002, avec 83 millions d'euros.
254. La Commission attire cependant l'attention de la Belgique sur le point 40 des lignes directrices de 2004, qui dispose:
Les radiations comptables et la fermeture d'activités déficitaires qui seraient en tout état de cause nécessaires pour rétablir la viabilité ne seront pas considérées comme une réduction de la capacité ou de la présence sur le marché aux fins de l'appréciation des contreparties.
255. D'après les informations que le gouvernement belge a transmis à la Commission, il semble que le retrait du marché français, ainsi que la fermeture des terminaux en Belgique, concernaient des activités déficitaires.
256. Afin de savoir si ces deux mesures sont suffisantes pour atténuer, autant que possible, les conséquences défavorables de l'aide pour les concurrents, il convient de rappeler les principaux développements des deux marchés sur lesquels IFB est actif, à savoir le marché de la logistique et le marché du transbordement du fret. Ensuite, il convient d'analyser si les mesures proposées atténuent autant que possible les conséquences défavorables de l'aide pour les concurrents.
a) Le marché de la logistique et les aides pour IFB
257. Comme expliqué dans la partie 2 de cette décision, le marché de la logistique est un marché en plein mutation, due à l'ouverture des marchés du transport ferroviaire et à l'entrée sur le marché des entreprises ferroviaires et postales, avec à la fois un grand nombre de petits acteurs spécialisés et de grands acteurs intégrés.
258. La Commission note que les mesures proposées ne concernent pas le marché de la logistique. Comme le montre le tableau du paragraphe 16 de la présente décision, IFB a su augmenter son volume sur ce marché de manière importante en 2004 (par rapport à 2003). La Belgique n'a présenté aucun engagement qui aurait limité, pendant la période de la restructuration, la présence d'IFB sur ce marché.
259. La Commission considère dès lors que l'absence de mesures proposées pour le marché de la logistique, ainsi que les faits que le marché est en plein mutation et qu'IFB a su augmenter son volume de manière importante, créent des doutes si la Belgique a limité, autant que possible, les conséquences défavorables pour la concurrence en ce qui concerne les activités de logistique d'IFB.
b) Le marché du transbordement de fret et les aides pour IFB
260. Les deux mesures proposées concernent le marché du transbordement de fret. IFB a quasiment arrêté ses activités en France, et a clôturé un terminal en Belgique et a vendu ses participations dans deux autres terminaux.
261. Le seul marché pour lequel l'aide peut avoir des conséquences négatives pour la concurrence est donc le marché belge. Sur ce marché, IFB a moins de 7 % des parts de marchés (cf. description des marchés dans la partie 2 de cette décision).
262. Afin de limiter les effets négatifs de l'aide sur le marché belge, IFB a clôturé un terminal, et a vendu ses participations dans deux autres. La Commission note cependant d'un côté que la fermeture concernait le plus petit des terminaux, et que la fermeture servait en premier lieu à réduire les pertes d'IFB Terminals, et de l'autre côté qu'IFB exploitera de nouveau les deux terminaux qu'il a vendu après l'augmentation de capital, car la société TRW, dont la SNCB apportera 47 % des parts sociales à IFB, détient des participations importantes dans les terminaux de Bruxelles et de Zeebrugge.
263. Ensuite, la Commission note qu'IFB possède des participations minoritaires dans un nombre importants de terminaux belges.
264. Par conséquent, la Commission a des doutes sur la question de savoir si les mesures proposées par IFB pour limiter, autant que possible, les effets négatifs de l'aide pour la concurrence sur le marché du transbordement du fret sont suffisantes.
3.2.2.4. Limitation de l'aide au strict minimum et contribution du bénéficiaire
265. Afin de démonter que l'aide est limitée au strict minimum, le gouvernement belge explique que l'augmentation du capital se limite à restaurer le capital social d'IFB, qui était devenu négatif suite aux pertes enregistrées en 2001 et 2002, à une hauteur qui lui permet de retrouver la viabilité économique. Comme expliqué ci-dessus dans la partie 2, le taux de solvabilité, c'est-à-dire le ratio fonds propres/passif, d'IFB sera de 33 % après l'augmentation de capital.
266. La Belgique a communiqué à la Commission les taux de solvabilité des principaux concurrents d'IFB. Ils sont les suivants:
Sociétés de terminaux | |
ABP Ports | 59,60 |
Hesse-Noord Natie | 58,19 |
Katoennatie Terminals | 54,97 |
Schelde Container Terminal Noord | 53,33 |
Sea-Ro-Terminal | 43,75 |
RSC | 74,24 |
Moyenne | 57,35 |
| |
Sociétés de Transport | |
DHL Freight (route) | 34,60 |
ECS European Containers (route) | 14,27 |
Gefco Benelux (rail) | 39,92 |
Henri Essers (route) | 15,71 |
Rhinecontainer (barge) | 18,63 |
TRW (rail) | 20,74 |
Ziegler (route) | 20,42 |
Moyenne | 23,47 |
| |
Sociétés aux activités mixtes | |
Gosselin | 38,92 |
Hupac | 34,90 |
Moyenne | 36,91 |
| |
Moyenne générale | 39,24 |
267. La Commission prend note de la circonstance que le taux de solvabilité envisagé pour IFB est inférieur à celui des sociétés de terminaux et aussi, bien que dans une moindre mesure, à celui des sociétés ayant des activités mixtes. Cependant, ce taux est supérieur à la moyenne des taux enregistrés dans les sociétés de transport. Il est vrai également que l'augmentation du capital est inférieure de 20 millions EUR à ce que le consultant McKinsey avait préconisé dans le plan de restructuration. Toutefois, à ce stade, la Commission ne dispose pas d'éléments suffisants pour conclure de manière définitive que l'aide a été limitée au strict minimum.
268. La Commission attire l'attention du gouvernement belge sur les dispositions des points 42 et suivants des lignes directrices de 2004, qui prévoient:
Les bénéficiaires de l'aide doivent contribuer de manière importante au plan de restructuration sur leurs propres ressources, y compris par la vente d'actifs qui ne sont pas indispensables à la survie de l'entreprise, ou par un financement extérieur obtenu aux conditions du marché. Cette contribution est un signe indiquant que les marchés croient à la faisabilité du retour à la viabilité. Elle doit être réelle, c'est-à-dire effective, à l'exclusion de tous bénéfices potentiels, tels que du cash flow, et doit être la plus élevée possible.
La Commission considèrera normalement que les contributions suivantes à la restructuration seront appropriées: au moins 25 % dans le cas des petites entreprises, au moins 40 % pour les entreprises de taille moyenne et au moins 50 % pour les grandes entreprises. Dans des circonstances exceptionnelles et dans des situations de difficulté particulière qui doivent être démontrées par l'État membre, la Commission pourra accepter une contribution propre réelle moins élevée.
Pour limiter l'effet de distorsion de la concurrence, le montant de l'aide ou la forme sous laquelle elle est accordée, doit être de nature à éviter que l'entreprise ne dispose de liquidités excédentaires qu'elle pourrait consacrer à des activités agressives susceptibles de provoquer des distorsions sur le marché qui ne seraient pas liées au processus de restructuration. À cet effet, la Commission examinera le niveau du passif de l'entreprise après sa restructuration, y compris après tout report ou réduction de ses dettes, en particulier dans le cadre de son maintien en activité à la suite d'une procédure collective de droit national relative à son insolvabilité. L'aide ne doit en aucune façon servir à financer de nouveaux investissements qui ne sont pas indispensables au retour à la viabilité de l'entreprise.
269. La Commission note que d'après le plan de restructuration, IFB ne semble pas faire de contribution propre à sa restructuration. Dès lors, la Commission a des doutes si IFB contribue, comme l'exige les lignes directrices de 2004, à son aide à la restructuration de manière suffisante.
3.2.2.5. Rapport annuel et "one time, last time"
270. Le gouvernement belge a accepté de fournir à la Commission un rapport annuel pour permettre à la Commission d'évaluer si le plan de restructuration est mis en oeuvre selon les engagements pris par les autorités belges.
271. Finalement, il y a lieu de vérifier si l'aide à la restructuration a respecté le principe "One time, last time". D'après les informations fournies par les autorités belges, IFB n'a pas bénéficié d'une aide à la restructuration auparavant. La Commission n'a pas encore pris de décision par rapport à IFB auparavant. Elle considère donc que le critère "one time, last time" a été respecté.
3.3. Conclusion
272. La Commission considère, à ce stade, que l'octroi d'un délai de paiement pour les dettes existantes de 63 millions d'euros et leur conversion, ainsi que la conversion des intérêts y liés de 11 millions d'euros, en capital social constituent une aide d'État, car la SNCB n'a pas agi comme l'aurait fait un investisseur privé en économie de marché.
273. De même, l'octroi d'une avance récupérable de 5 millions d'euros et l'octroi d'une facilité de crédit de 15 millions d'euros, la conversion de la facilité de crédit de 15 millions et des intérêts y liés de 2,5 millions d'euros en capital social, ainsi que l'apport en nature de 5 millions d'euros de nouveau capital social constituent des aides d'État.
274. Dans la mesure où ces aides constituent des aides de trésorerie, elles ne peuvent pas être déclarées compatibles avec le marché commun en tant qu'aides à la restructuration, car elles ont été octroyées pour une période qui dépasse 12 mois.
275. La Commission a des doutes sur la question de savoir si l'ensemble des aides peut être déclarées compatibles avec le marché commun en tant qu'aides à la restructuration.
276. Ses doutes portent sur l'imputabilité d'une partie de l'aide à l'État belge, le caractère suffisant des mesures prises pour atténuer, autant que possible, les conséquences défavorables de l'aide pour les concurrents, ainsi que sur la limitation de l'aide au strict minimum et sur la suffisance de la contribution propre de l'entreprise IFB aux aides à la restructuration.
4. DÉCISION
La Commission a décidé de considérer, à ce stade, que les mesures de sauvetage et les mesures de restructuration en faveur d'IFB constituent des aide d'État au sens de l'article 87 (1) du traité CE.
Elle émet des doutes sur la question de savoir si ces aides peuvent être déclarées compatibles avec le marché commun en vertu des lignes directrices pour les aides à la restructuration et ouvre donc pour cette partie du dossier la procédure prévue à l'article 88 § 2 du traité CE.
Compte tenu des considérations qui précédent, la Commission invite la Belgique, dans le cadre de la procédure de l'article 88, paragraphe 2, du traité CE, à présenter ses observations et à fournir toute information utile pour l'évaluation de l'aide dans un délai d'un mois à compter de la date de réception de la présente. Elle invite vos autorités à transmettre immédiatement une copie de cette lettre au bénéficiaire potentiel de l'aide.
La Commission rappelle à la Belgique l'effet suspensif de l'article 88, paragraphe 3, du traité CE et se réfère à l'article 14 du règlement (CE) no 659/1999 du Conseil qui prévoit que toute aide illégale pourra faire l'objet d'une récupération auprès de son bénéficiaire.
Par la présente, la Commission avise la Belgique qu'elle informera les intéressés par la publication de la présente lettre et d'un résumé de celle-ci au Journal officiel de l'Union européenne. Elle informera également les intéressés dans les pays de l'AELE signataires de l'accord EEE par la publication d'une communication dans le supplément EEE du Journal officiel, ainsi que l'autorité de surveillance de l'AELE en leur envoyant une copie de la présente. Tous les intéressés susmentionnés seront invités à présenter leurs observations dans un délai d'un mois à compter de la date de cette publication."
"1. PROCEDURE
1.1. Zaak NN 9/2004
1. Bij schrijven van 12 augustus 2003, geregistreerd bij de Europese Commissie op 20 augustus 2003 (TREN/A(03)27718), hebben de Belgische autoriteiten enkele door de Nationale Maatschappij der Belgische Spoorwegen (NMBS) en haar dochtermaatschappij Inter Ferry Boats (IFB) gesloten overeenkomsten aangemeld krachtens artikel 88, lid 3, van het EG-Verdrag. Deze aanmelding behelst reddingsmaatregelen die de NMBS heeft genomen ten gunste van IFB.
2. Op 13 oktober 2003 (D(03)17546) heeft het directoraat-generaal Energie en vervoer de Belgische autoriteiten verzocht de Commissie aanvullende inlichtingen te verstrekken. In verband hiermee heeft op 12 december 2003 een bilaterale ontmoeting met de Belgische autoriteiten plaatsgevonden. Tijdens deze ontmoeting werd een door McKinsey opgesteld herstructureringsplan voor IFB gepresenteerd.
3. De Belgische autoriteiten hebben de brief van de Commissie beantwoord met het schrijven van 7 januari 2004, dat op 13 januari 2004 (TREN/A(04)10708) bij de Commissie is geregistreerd. Uit genoemd schrijven blijkt dat de aangemelde reddingsmaatregelen reeds gedeeltelijk zijn uitgevoerd. Derhalve is de zaak geregistreerd onder nummer NN 9/2004. Op 30 april 2004 heeft nogmaals een vergadering plaatsgevonden. De Belgische autoriteiten hebben bij schrijven van 15 juni 2004, dat bij de Commissie op 21 juni 2004 is geregistreerd (TREN/A(04)23691), de aanvullende documenten toegestuurd waarom de Commissie tijdens deze vergadering had verzocht.
4. Bij schrijven van 26 januari 2005 (D(05)100339) heeft het directoraat-generaal Energie en vervoer de Belgische autoriteiten verzocht aanvullende inlichtingen te verstrekken betreffende de ontwikkeling van IFB, en met name haar herstructurering.
5. Bij schrijven van 25 maart 2005, dat bij de Commissie is geregistreerd op 30 maart 2005 (TREN/A(05)7712), hebben de Belgische autoriteiten de Commissie de aanvullende inlichtingen toegestuurd waarom zij in haar schrijven van 26 januari 2005 had verzocht.
1.2. Zaak N 55/2005
6. Bij schrijven van 28 januari 2005 (SG(2005)A1133) hebben de Belgische autoriteiten bij de Commissie het voornemen van de NMBS om het kapitaal van IFB te verhogen, aangemeld. De Belgische autoriteiten zijn van mening dat het niet om staatssteun gaat, maar hebben dit voornemen aangemeld om redenen van rechtszekerheid. De Commissie heeft deze zaak als een nieuw dossier "aangemelde staatssteunmaatregel" geregistreerd onder nummer N 55/2005.
7. Bij schrijven van 29 maart 2005 (D(05)106199) heeft het directoraat-generaal Energie en vervoer de Belgische autoriteiten verzocht aanvullende inlichtingen te verstrekken over de herstructureringsmaatregelen van IFB.
8. Bij schrijven van 28 april 2005, geregistreerd bij de Commissie op 3 mei 2005 (SG(2005)A(05)4155), hebben de Belgische autoriteiten de Commissie de aanvullende inlichtingen toegezonden waarom in de brief van 29 maart 2005 was verzocht.
9. Bij brief van 31 mei 2005 (D(05)111096) heeft het directoraat-generaal Energie en vervoer de Belgische autoriteiten verzocht aanvullende inlichtingen te verstrekken betreffende de op 28 april 2005 toegezonden informatie.
10. Bij schrijven van 30 juni 2005, dat bij de Commissie is geregistreerd op 1 juli 2005 (TREN/A(05)16598), hebben de Belgische autoriteiten de Commissie de aanvullende inlichtingen toegezonden waarom in de brief van 31 maart 2005 was verzocht.
11. Op 16 september 2005 heeft een werkvergadering plaatsgevonden tussen de Commissie en de Belgische autoriteiten. Tijdens deze vergadering heeft de Commissie de Belgische autoriteiten verzocht aanvullende inlichtingen te verstrekken. De Belgische autoriteiten hebben deze inlichtingen toegezonden per e-mail van 21 oktober 2005, die bij de Commissie is geregistreerd op 24 oktober 2005 (TREN/A(05)27067).
2. GEDETAILLEERDE BESCHRIJVING VAN DE REDDINGS- EN HERSTRUCTURERINGSMAATREGELEN
2.1. De partijen in de kaderovereenkomst betreffende de redding en herstructurering van IFB
2.1.1. IFB
2.1.1.1. Beschrijving van IFB
12. Inter Ferry Boats (IFB) is een naamloze vennootschap volgens Belgisch recht. De NMBS bezit 89,03 % van het maatschappelijk kapitaal. De overige aandeelhouders zijn CNC Transports, voor 93,8 % een dochtermaatschappij van de NMBS (7,41 %), ICF (2,08 %) en EWS (English Welsh and Scottish Railway — 1,22 %). IFB telt momenteel 245 werknemers.
13. IFB werd op 1 april 1998 opgericht door de fusie van de volgende drie bedrijven: Ferry Boats Ltd., Interferry Ltd. en de spoordivisie van Edmond Depaire Ltd. Vóór de oprichting van IFB was Ferry Boats Ltd. een onderneming die onder de gezamenlijke zeggenschap stond van de Britse spoorwegen en de Belgische spoorwegen. Interferry Ltd. en Edmond Depaire Ltd. vielen onder de zeggenschap van de Belgische spoorwegen. Uit de door België verstrekte documenten blijkt niet duidelijk of IFB de rechtspersoonlijkheid van een van de drie ondernemingen heeft voortgezet.
14. Ferry Boats Ltd. werd in 1923 opgericht onder de naam "Société Belgo-Anglaise des Ferry-Boats". Interferry is in 1967 opgericht onder de naam "Intercontainer" en de onderneming Edmond Depaire in 1906 opgericht als een particuliere onderneming voor het vervoer van containers.
15. De activiteiten van IFB zijn geconcentreerd in twee sectoren:
- de activiteitensector "IFB Logistics", voor het commerciële beheer van de expeditieactiviteiten van IFB, en
- de activiteitensector "IFB Terminals", die de inlandterminals exploiteert.
Aan deze activiteiten moeten de participaties en de dochtermaatschappijen worden toegevoegd die IFB heeft of had in België en in het buitenland.
a) De activiteit IFB Logistics
16. De activiteit "IFB Logistics" betreft het commerciële beheer door IFB, alsmede door de ondernemingen waarin zij een participatie heeft, van:
- expeditieactiviteiten (inclusief aanvullende "transport engineering"-diensten) en
- logistieke diensten.
17. De expeditieactiviteiten zijn de belangrijkste activiteiten van "IFB Logistics". Deze activiteiten bestaan erin aan de cliënten zo volledig mogelijke vervoersoplossingen aan te bieden. Wat de expeditieactiviteiten betreft, vertegenwoordigt het spoorvervoer, ongeacht of het gaat om conventioneel dan wel om gecombineerd vervoer, voor IFB de belangrijkste wijze van vervoer, maar IFB biedt ook vervoer over de binnenwateren en over de weg aan. Voor IFB is het spoorvervoer vooral vervoer over "korte" of "middellange" afstand (100 à 500 km, waarbij IFB vooral optreedt als partner van de reders voor de ontwikkeling van "carrier haulage", een activiteit welke die van de spoorwegexploitanten (die zich veeleer concentreren op langeafstandsvervoer) aanvult.
18. De door IFB verzonden goederen zijn bulkproducten, containers en diverse producten (general cargo). In onderstaande tabel wordt de hoeveelheid vracht aangegeven die door IFB in 2003 en 2004 over het conventionele spoor, het intermodale spoor en over de binnenwateren is vervoerd. Uitsluitend in gevallen waarin de cliënt heeft verzocht om dienstverlening van deur tot deur of van/naar een zeeterminal, maakt IFB gebruik van het vervoer over de weg om transporteenheden naar of vanuit spoorwegterminals te vervoeren.
19. De belangrijkste cliënten van IFB Logistics zijn de zeevrachtbedrijven […] [48] [49] en […], alsmede […] [50], […], […] [51] en […]. De producten die worden vervoerd zijn met name chemische producten, steenkool en granulaat. In onderstaande tabel zijn de door IFB in 2003 en 2004 vervoerde volumes aangegeven.
Jaar | Conventioneel spoor [52] | Intermodaal spoor | Binnenvaart |
2003 | 0,672 miljoen ton | 423583 TEU [53] | 0,385 miljoen ton |
2004 | 1,995 miljoen ton | 481556 TEU | 1,023 miljoen ton |
20. De expeditieactiviteiten omvatten ook aanvullende "transport engineering"-diensten, zoals opslag, distributie, overslag, …, die er nauw mee samenhangen.
21. In het kader van haar organisatie valt ook de activiteit van agent voor rekening van derde spoorwegexpediteurs/vervoerders onder IFB Logistics. IFB is als logistiek agent in België actief voor een aantal buitenlandse ondernemingen.
22. De markt voor expeditieactiviteiten en logistieke activiteiten heeft de voorbije jaren een aanzienlijke groei gekend, die samenhangt met de toenemende mondialisering van het bedrijfsleven, de trend naar uitbesteding en een steeds verdergaande specialisatie van de productieondernemingen (just in time production).
23. De belemmeringen voor de toegang tot de markt zijn afgenomen en op de markt zijn zowel tal van kleine gespecialiseerde actoren als grote geïntegreerde actoren (DHL, UPS, …) aanwezig. Als gevolg van de liberalisering van de spoorwegmarkt en van de markt voor postdiensten hebben spoorwegondernemingen (Deutsche Bahn, NMBS) en postondernemingen (Deutsche Post) hun intrede gedaan op die markt.
24. De combinatie van marktgroei, toetreding van belangrijke nieuwkomers en liberalisering van het spoorvervoer heeft gemaakt dat deze markt volop aan het veranderen en bewegen is.
b) IFB Terminals
25. IFB Terminals exploiteert inlandterminals (overladen van intermodale transporteenheden (ITU) van/naar het spoor).
26. De voornaamste activiteit van de inlandterminals ("dry ports") bestaat in het overladen van zeecontainers van vrachtwagens op spoorwagons. IFB exploiteert in totaal zes inlandterminals die zijn aangesloten op het Belgische spoorwegnet en waarvan er zich vier in de haven van Antwerpen en drie in het Belgische achterland bevinden.
27. De inlandterminals in de haven van Antwerpen zijn "Mainhub", "Cirkeldijck", "Zomerweg" en "Schijnpoort". De Belgische regering onderstreept dat deze vier terminals zich in een bijzondere situatie bevinden, aangezien zij gelegen zijn in de haven van Antwerpen, in het centrum van de zeevaartactiviteiten waarmee zij onlosmakelijk zijn verbonden. De ITU die in deze terminals worden behandeld, zijn hoofdzakelijk zeecontainers, die eerst van schepen naar vrachtwagens worden overgeslagen in een niet door IFB geëxploiteerde zeeterminal. Pas nadien worden deze containers van de vrachtwagens naar treinwagons overgeslagen in een door IFB geëxploiteerde inlandterminal. In geval van export over zee is de volgorde omgekeerd. In 2004 hebben de vier inlandterminals van IFB in de haven van Antwerpen 0,4 miljoen TEU behandeld.
28. IFB exploiteert twee inlandterminals die zich niet in de haven van Antwerpen bevinden, namelijk de terminal van Muizen (in de buurt van Mechelen, terminal weg-spoor) en de terminal van Rénory (in de buurt van Luik, verkeer weg-spoor-binnenschip). Een derde terminal, die van Bressoux, is in 2003 gesloten.
29. De markt voor terminals is een stabielere markt dan die voor logistiek. Het aantal in België geëxploiteerde terminals blijft constant. Het aantal vervoerde containers neemt echter toe ten gevolge van de groei van het verkeer in de haven van Antwerpen en de inspanningen om meer goederen via het gecombineerde vervoer te transporteren.
c) De participaties van IFB
30. IFB heeft of had participaties in ondernemingen die zee- en inlandterminals exploiteren, alsmede in vervoersondernemingen. IFB heeft of had in totaal een dertigtal participaties.
31. Participaties in de zee- en inlandterminals in Duinkerke. IFB heeft belangrijke investeringen gedaan in de haven van Duinkerke, waar zij meerderheidsparticipaties bezat in Acimar (terminal voor staalproducten, volle dochtermaatschappij van NFTI-ou) en NFTI-ou (terminal voor zeecontainers, participatie van 60 % in 2003, sindsdien verminderd tot 30 %), Dry Port Dunkerque (DPD, een spoorwegterminal, sinds 2003 ongewijzigd gebleven participatie van 90 %), Short Sea Terminal Dunkirk (SSTD, laden en lossen van opleggers, participatie van 50 % in 2003, sindsdien tot 0 % teruggebracht), en IFB France (holdingmaatschappij en onderneming voor dienstverlening aan in Duinkerke gevestigde verbonden ondernemingen, participatie van 100 %, sindsdien volledig verkocht aan NFTI-ou).
32. IFB France is omgedoopt tot Administration Gestion Entreprise Portuaires (AGEP). IFB heeft de totaliteit van haar aandelen in deze ondernemingen overgedragen aan NFTI-ou.
33. In december 2002 is een insolventieprocedure ingeleid tegen Acimar. Acimar is niet meer actief sinds 1 september 2003. Alle aandelen die IFB in Acimar bezat, zijn overgedragen aan AGEP (zie hierna).
34. IFB heeft haar participatie in NFTI-ou, die AGEP en, via AGEP, Acimar in haar bezit heeft, van 60 % teruggebracht tot 30 %. IFB heeft haar patronaat (door een moedermaatschappij tegenover derden aangegane verbintenis dat zij zal instaan voor de nakoming van de verplichtingen van haar dochtermaatschappij) ingetrokken door de opzegging van haar "comfort letter" (patronaatsverklaring). IFB is aldus bevrijd van elke verplichting om als garant voor NFTI-ou op te treden, aangezien deze verplichting volledig werd overgedragen aan de meerderheidsaandeelhouder, de Port Autonome de Dunkerque, die 70 % van de aandelen van NFTI-ou bezit. IFB tracht nu haar minderheidsparticipatie in NFTI-ou van de hand te doen.
35. IFB had een participatie van 90 % in DPD. In juni 2003 heeft IFB haar patronaatsverklaring opgezegd; vervolgens heeft IFB de infrastructuur en de apparatuur van DPD aan de Port Autonome de Dunkerque verkocht en DPD in juni 2004 ontbonden. De liquidatie werd afgesloten in de zomer van 2005.
36. IFB heeft haar participatie in SSTD verkocht in april 2005.
37. IFB heeft bijgevolg al haar participaties in de haven van Duinkerke verkocht, met uitzondering van haar minderheidsparticipatie in NFTI-ou, waarvoor zij een koper zoekt.
38. Participatie in terminals in België. In België had IFB participaties in de terminals van Zeebrugge, Brussel, Moeskroen, Athus, Luik en Charleroi.
39. In Zeebrugge hadden IFB en Hesse-Noord Natie het economische samenwerkingsverband OCHZ opgericht, waarvan IFB en Hesse-Noord Natie elk voor de helft mede-eigenaar waren. In september 2004 is IFB uit OCHZ gestapt en heeft zij haar rechten aan OCHZ verkocht.
40. In Brussel had IFB via Brussels Port Invest (BPI) en Brussels Terminal Intermodal (BTI) belangen in een trimodale containerterminal in de haven van Brussel. BTI is intussen ontbonden en aan een liquidatieprocedure onderworpen. Haar participatie in BPI heeft IFB overgedragen aan een andere onderneming buiten de NMBS-groep.
41. In Moeskroen heeft IFB een participatie van 16,76 % in de onderneming SA Dryport Mouscron Lille (DPM Li). Deze onderneming beschikt over een eigen kapitaal van 530000 euro en heeft in 2004 een nettoresultaat van 76000 euro gerealiseerd.
42. In Athus heeft IFB een participatie van 24,89 % in de onderneming SA Terminal Athus (Terminal Athus). Deze onderneming heeft een eigen kapitaal van 1,7 miljoen euro en heeft in 2002 een nettoresultaat van 61000 euro behaald (er zijn geen recentere gegevens beschikbaar).
43. In Luik heeft IFB een participatie van 45,12 % in Liège Logistics Intermodal. De Commissie beschikt niet over meer informatie over deze participatie.
44. In Charleroi heeft IFB een participatie van 14,28 % in de onderneming SA Charleroi Dry Port (Charleroi DP). Deze onderneming heeft een eigen kapitaal van 36000 euro en heeft in 2002 een nettoresultaat van 899 euro gerealiseerd (er zijn geen recentere gegevens beschikbaar).
45. IFB heeft op dit ogenblik bijgevolg minderheidsparticipaties in vier terminals in België, namelijk de terminals van Moeskroen, Luik, Athus en Charleroi. IFB heeft bovendien een participatie van 0,9 % in de onderneming die deze terminals exploiteert, namelijk TRW. De NMBS heeft een directe participatie van 47 % in TRW.
46. IFB heeft daarentegen haar participaties in de terminals van Zeebrugge en Brussel verkocht.
47. Participaties in vervoersondernemingen. IFB heeft of had de volgende participaties in vervoersondernemingen:
- CNC Ferry Boats intermodal, België, 50 % (eigen kapitaal: 61000 euro, nettoresultaat 2004: niet bekend) en haar volle dochtermaatschappij Rail Web. Rail Web is op 31 maart 2005 ontbonden.
- Affrètements Van Reeth, België, 100 % (eigen kapitaal: 412000 euro; nettoresultaat in 2002: 150000 euro).
- SA Unilog, België, 55 % (eigen kapitaal: 1,9 miljoen euro, nettoresultaat in 2004: 21000 euro).
- SA Unilog, Verenigd Koninkrijk, 100 % (geen andere informatie beschikbaar).
- SA Rail Infra Logistics, België, 99,93 % (eigen kapitaal: 500000 euro; nettoresultaat in 2004: 55000 euro).
- ACTS België, 12,5 % (geen andere informatie beschikbaar). Deze onderneming is op 29 maart 2005 ontbonden.
- RKE, België, 61,46 % (eigen kapitaal: 2,6 miljoen euro, nettoresultaat in 2004: 250000 euro).
- Coil Terminal, onrechtstreeks via RKE, aangezien RKE een participatie van 50 % heeft in Coil Terminal.
- CARRE (geen andere informatie beschikbaar). Er zijn onderhandelingen over de verkoop van CARRE aan de gang.
- GIE Cigogne Shuttle, België (geen andere informatie beschikbaar). IFB denkt eraan om uit deze onderneming te stappen.
- Haeger Schmidt International, Duitsland, 100 % (eigen kapitaal: 2,1 miljoen euro, nettoresultaat in 2004: niet bekend)
- Compagnie nouvelle des conteneurs Transports Nationaux et Internationaux, Frankrijk, 2 % (geen andere informatie beschikbaar).
- GIE NEN (geen andere informatie beschikbaar). GIE wordt ontbonden.
- ACTS Belgique, 13 % (geen andere informatie beschikbaar). Deze onderneming is op 5 november 2003 ontbonden.
- TRW, België, 0,89 %.
48. Participatie in Haeger and Schmidt International. Via haar volle dochtermaatschappij, Haeger and Schmidt International, heeft IFB participaties in Best Logistics (Polen), A. van Reeth (Frankrijk), KREAS en SITRA. Haeger and Schmidt heeft een jaaromzet van 50 miljoen euro, hoofdzakelijk door de binnenvaart.
49. Overzicht. In onderstaand schema wordt een algemeen overzicht gegeven van alle participaties van IFB. Het overzicht is als volgt opgebouwd:
eerste kolom: de participaties in ondernemingen die terminals exploiteren;
tweede kolom: de participaties in vervoersondernemingen;
derde kolom: de participaties in ondernemingen die diensten verrichten;
vierde kolom: de participaties in (Duitse) ondernemingen die actief zijn op het gebied van de binnenvaart (binnenschepen).
+++++ TIFF +++++
2.1.1.2. Definitie van de relevante markten en marktaandelen van IFB
50. De Commissie heeft in het verleden in haar beschikkingen COMP/M.3603 "UPS/Menlo" en COMP/M.3496 "TNT FORWARDING HOLDING/WILSON LOGISTICS" uitspraak gedaan over de definitie van de relevante markten voor expeditieactiviteiten en logistieke activiteiten; als relevante productmarkt heeft zij aangemerkt:
- voor de expeditieactiviteiten of freight forwarding: "the organisation of transportation items (possibly including ancillary activities such as customs clearance, warehousing, ground services, etc.) on behalf of customers according to their needs."
- voor de logistieke activiteiten of general logistic services: "the part of the supply chain process that plans, implements and controls the efficient, effective flow and storage of goods, services and related information from the point of origin to the point of consumption in order to meet customers' requirements."
51. Deze markten zijn, ondanks een trend naar een sterkere internationalisering, als nationaal aangemerkt.
52. Volgens de door de Belgische regering verstrekte informatie ligt het marktaandeel van IFB Logistics op deze beide markten tussen 2 % en 5 %, wat zou kunnen worden verklaard door het betrekkelijk kleine deel van de goederen dat via gecombineerd vervoer en via het spoor wordt getransporteerd.
53. Deze raming lijkt betrouwbaar, wanneer de omzet van IFB, die in 2003 […] euro bedroeg, wordt vergeleken met de omzet van de andere Belgische actoren op die markt, die in 2003 in België de volgende omzet hebben gerealiseerd:
Onderneming | Omzet |
Hesse-Noordnatie | 485 miljoen euro |
Danzas | 176 miljoen euro |
Ziegler | 129 miljoen euro |
Schenker | 156 miljoen euro |
54. Wat de markt voor terminals betreft, moet een onderscheid worden gemaakt tussen inlandterminals en zeeterminals.
55. De Commissie heeft in verband met de inlandterminals een standpunt over de definitie van de relevante markten ingenomen in haar beschikkingen COMP M 2632 "DEUTSCHE BAHN/ECT INTERNATIONAL/UNITED DEPOTS", IV/M 1651 "MAERSK/SEA LAND" en IV/M.831 "PT/Nedlloyd".
56. In haar beschikking COMP M 2632 heeft de Commissie de relevante productmarkt gedefinieerd als de markt "für das Erbringen von Umschlagdienstleistungen im Containergüter-Hinterlandverkehr per Binnenschiff zwischen ARA-Häfen und deutschem Niederrhein/Ruhrgebiet", en de geografische markt als "die Containerterminals entlang des Niederrheins von Nijmeggen bis Köln". Alle terminals van de Benedenrijn zouden met andere woorden de relevante markt zijn. In de beschikkingen IV M 1651 en IV M 831 wordt de geografische markt van een haven als volgt gedefinieerd: "Ports or groups of ports serve a particular hinterland or are used for transshipment to smaller ports. The geographic area they generally serve determines the geographic scope related to their services". Hieruit volgt dat de productmarkt de markt voor de overslag van vracht is en het geografische gebied dat erdoor wordt bestreken het achterland van een bepaalde haven.
57. In het onderhavige geval moet derhalve worden geconcludeerd dat de relevante productmarkt kan worden gedefinieerd als de markt voor diensten op het gebied van de overslag van ITU van/naar het vervoer over land (weg — spoorweg — binnenschip). De relevante geografische markt is op zijn minst de regio Antwerpen en omgeving, eventueel zelfs de regio van de ARA-havens.
58. Behalve de inlandterminals van IFB bieden ook de op zijn minst trimodale terminals van Hesse-Noordnatie (Noordzeeterminal, Europaterminal) en P O Ports (Seaport terminal) diensten op het gebied van de overslag van ITU van/naar het vervoer over land (weg — spoorweg — binnenschip) aan. Deze terminals zijn, wat het volume behandelde ITU betreft, heel wat belangrijker dan de terminals van IFB. In 2004 heeft Hesse-Noordnatie 4,9 miljoen TEU behandeld en P O Ports 0,7 miljoen TEU, terwijl IFB 0,4 miljoen TEU heeft behandeld. Het marktaandeel van IFB bedraagt derhalve ongeveer 6,7 %.
59. De twee zeeterminals waarin IFB participaties heeft, hebben in België en Frankrijk slechts marginale marktaandelen. IFB heeft geen participaties in terminals in andere landen.
2.1.2. De NMBS
60. De NMBS is opgericht bij de Belgische wet van 23 juli 1926 tot oprichting van de Nationale Maatschappij der Belgische Buurtspoorwegen [54]. Sinds 14 oktober 1992 [55] is de NMBS een autonoom overheidsbedrijf en een naamloze vennootschap van publiek recht [56]. De NMBS valt bijgevolg onder de voor naamloze vennootschappen geldende wettelijke en bestuursrechtelijke bepalingen van het handelsrecht voor alle aspecten die niet uitdrukkelijk zijn geregeld bij of krachtens titel I van de wet van 21 maart 1991 houdende hervorming van sommige economische overheidsbedrijven dan wel door of krachtens een specifieke wet.
61. De Belgische staat heeft de structuur van de NMBS op 1 januari 2005 hervormd. Zij is omgevormd tot drie afzonderlijke vennootschappen, namelijk:
- NMBS Holding: een vennootschap "van het type holding" die participaties in de twee andere vennootschappen zal hebben,
- Infrabel, de infrastructuurbeheerder,
- Nieuwe NMBS, de spoorwegmaatschappij.
62. Het maatschappelijk doel van de NMBS staat omschreven in artikel 1bis van voornoemde wet van 23 juli 1926, dat in de wet van 1 augustus 1966 [57] is ingevoegd en bij artikel 155 van voornoemde wet van 21 maart 1991 als volgt is gewijzigd:
"(1) De maatschappij heeft tot doel het vervoer van reizigers en goederen per spoor."
"(2) De maatschappij kan, op eigen gezag, of door middel van deelneming in bestaande of op te richten Belgische, vreemde of internationale organismen, alle commerciële, industriële of financiële handelingen verrichten, die rechtstreeks of onrechtstreeks, geheel of ten dele in verband staan met haar maatschappelijk doel, dan wel de verwezenlijking of de uitbreiding van dat doel kunnen vergemakkelijken of bevorderen."
"(3) Het feit dat er goederen of diensten worden gefabriceerd en verkocht, die rechtstreeks of onrechtstreeks op de spoorwegactiviteiten betrekking hebben, is inzonderheid van aard de verwezenlijking of de uitbreiding van het maatschappelijk doel te bevorderen."
63. Dit artikel is door de Belgische jurisprudentie en rechtsleer steeds ruimer geïnterpreteerd. Volgens de Belgische autoriteiten vallen de activiteiten van IFB duidelijk onder dit artikel.
64. De beheersorganen van de NMBS zijn de raad van bestuur, het directiecomité en de gedelegeerd bestuurder. De raad van bestuur is samengesteld uit tien leden, met inbegrip van de gedelegeerd bestuurder. De bestuurders worden door de koning benoemd bij een besluit vastgesteld na overleg in de Ministerraad. Zij worden gekozen overeenkomstig de complementariteit van hun competentie inzake financiële en boekhoudkundige analyse, juridische aspecten, hun kennis van de vervoerssector, hun deskundigheid inzake mobiliteit, personeelsstrategie en sociale relaties. Nadat zij zijn benoemd oefenen de leden van de raad van bestuur hun mandaat op onafhankelijke wijze uit en aanvaarden zij van niemand instructies.
65. De leden van het directiecomité worden met uitzondering van de gedelegeerd bestuurder benoemd door de raad van bestuur, die ook het aantal leden bepaalt. Het directiecomité vormt een college.
2.2 De financiële moeilijkheden van IFB
66. Over de jaren 2001 en 2002 heeft IFB aanzienlijke verliezen geboekt: volgens de jaarrekeningen van IFB betreffende 2002 bedroeg het gecumuleerde verlies op 31 december 2002 137 miljoen euro (waarvan 25 miljoen euro overgedragen van 2001), met als resultaat negatieve eigen middelen ten belope van 84 miljoen euro. Aan het einde van het boekjaar 2001 bedroegen deze eigen middelen nog 28 miljoen euro.
67. Steeds volgens de jaarrekeningen van 2002 bedroegen de operationele verliezen in het boekjaar 2002, d.w.z. het verschil tussen de lopende uitgaven en de lopende ontvangsten, 13,4 miljoen euro. Eerst dienen de oorzaken van de financiële moeilijkheden te worden onderzocht en vervolgens moet de reactie van het management van IFB en van de NMBS, alsmede die van de particuliere schuldeisers van IFB worden beschreven.
2.2.1. De oorzaken van de financiële moeilijkheden
68. De financiële moeilijkheden waarmee IFB werd geconfronteerd bij haar participaties in Frankrijk in de haven van Duinkerke en die haar ertoe hebben verplicht belangrijke voorzieningen in haar jaarrekeningen van 2001 en 2002 op te nemen, zijn de belangrijkste oorzaak van de financiële moeilijkheden van IFB.
69. Bovendien leden de activiteiten "IFB Logistics" en "IFB Terminals" in 2001 en 2002 lichte verliezen.
2.2.2. De reactie van het management van IFB en van de NMBS
70. Sinds 2000 had IFB niet meer alle facturen betaald die de NMBS haar voor treindiensten had toegezonden. In 2001, en vooral in 2002, heeft IFB evenmin alle facturen betaald. De NMBS lijkt dat te hebben geduld. De totale waarde van de facturen van de NMBS die niet door IFB werden betaald, bedroeg eind januari 2003 63 miljoen euro.
71. Als gevolg van de financiële moeilijkheden van IFB raakten zowel de raad van bestuur van IFB als de voornaamste aandeelhouder, de NMBS, er steeds meer van overtuigd dat voor het overleven van de groep IFB op lange termijn het beheer van de onderneming structureel moest worden veranderd.
72. Op 19 september 2002 heeft de gedelegeerd bestuurder van IFB aan twee accountants de opdracht gegeven een bijzonder rapport op te stellen over de financiële toestand van de onderneming. Op 24 december 2002 heeft de bijzondere algemene vergadering der aandeelhouders (BAV) van IFB er kennis van genomen dat de NMBS, naar aanleiding van de vergadering van de raad van bestuur van 20 december 2002, bereid was in te tekenen op een kapitaalverhoging ter verbetering van de financiële toestand van IFB ten belope van maximaal 80 miljoen euro, waarvan 20 miljoen euro bestemd was om tegemoet te komen aan de behoeften van IFB aan liquide middelen. De raden van bestuur van de NMBS en IFB hebben in principe hun goedkeuring gehecht aan twee kapitaalverhogingen — van 60 miljoen euro door omzetting van vorderingen van de NMBS op IFB en van 20 miljoen euro door terbeschikkingstelling aan IFB van liquide middelen -, te onderschrijven door de NMBS om de voortzetting van de activiteiten van IFB te waarborgen.
73. IFB en de NMBS hebben op 7 april 2003 een "kaderovereenkomst m.b.t. de herstructurering van IFB" gesloten, teneinde tot genoemde kapitaalverhogingen over te gaan. Deze overeenkomst, een privaatrechtelijke overeenkomst, bestaat uit twee delen: een deel "reddingsmaatregelen" en een deel "herstructureringsmaatregelen".
74. Gezien de omstandigheden heeft de raad van bestuur van IFB na overleg met de voornaamste aandeelhouder, de NMBS, besloten een bijzondere algemene vergadering der aandeelhouders samen te roepen, zoals artikel 633 van het Belgische wetboek van vennootschappen voorschrijft wanneer het verlies minstens de helft van het maatschappelijk kapitaal bedraagt. Op deze vergadering, die op 20 mei 2003 werd gehouden, konden de aandeelhouders van IFB kennis nemen van het bijzondere rapport van de raad van bestuur van IFB, waarin de kaderovereenkomst tussen de NMBS en IFB werd besproken, en werd voorgesteld om de activiteiten van IFB na een herstructurering voort te zetten. Op basis hiervan zijn de aandeelhouders van IFB akkoord gegaan met de voortzetting van de activiteiten van IFB.
2.2.3. De reactie van de particuliere schuldeisers van IFB
75. Particuliere zakenbanken hebben IFB leningen en bankgaranties toegestaan. Volgens de door de Belgische regering verstrekte gegevens hebben de financiële moeilijkheden van IFB geen enkele invloed gehad op de relaties tussen IFB en de banken: alle banken hebben de bij overeenkomst vastgelegde voorwaarden gehandhaafd zonder andere aanvullende garanties, waarborgen of zekerheden te eisen dan de gebruikelijke. Nog volgens de Belgische regering waren alle banken bereid nieuwe leningen toe te staan tegen concurrerende voorwaarden.
76. Op 31 december 2004 had IFB de volgende leningsovereenkomsten gesloten met particuliere banken:
Doel van de lening | Bank | Jaar | % | Bedrag (in EUR) | Situatie op 31.12.2004 (in EUR) |
[…] | […] | 1997 | [tussen 2 % en 6 %] | 328334,97 | […] |
[…] | […] | 1999 | [tussen 2 % en 6 %] | 1264930,18 | […] |
[…] | […] | 1999 | [tussen 2 % en 6 %] | 1611307,91 | […] |
[…] | […] | 2001 | [tussen 2 % en 6 %] | 4945476,00 | […] |
[…] | […] | 2003 | [tussen 2 % en 6 %] | 2000000,00 | […] |
TOTAAL | | | | 10150049,06 | 5550066,03 |
77. De laatste leningsovereenkomst werd gesloten in juli 2003, dus na het sluiten van de kaderovereenkomst tussen IFB en de NMBS en nadat de banken hadden gehoord van de financiële moeilijkheden van IFB.
78. Op 31 december 2004 beschikte IFB over de volgende bankgaranties:
Begunstigde van de bankgarantie | Bedrag (in euro) |
Federale overheidsdienst FINANCIËN Garantie douane en accijnzen | 2401220,64 |
Federale overheidsdienst FINANCIËN Garantie fiscaal geschil | 1772817,63 |
Federale overheidsdienst MOBILITEIT EN VERVOER Garantie expediteur | 111552,12 |
Andere garanties | 44767,12 |
79. Alle kredietlijnen in verband met deze garanties zijn gehandhaafd zonder wijziging van de bij overeenkomst vastgestelde voorwaarden.
2.3. De belangrijkste bepalingen van de "kaderovereenkomst tussen de NMBS en IFB m.b.t. de herstructurering van IFB"
80. Om het voortbestaan van IFB te waarborgen hebben de NMBS en IFB de reeds aangehaalde kaderovereenkomst gesloten. Daarin wordt bepaald dat de voorgestelde maatregelen in twee fasen worden uitgevoerd: in een eerste fase wordt een reeks reddingsmaatregelen ten behoeve van IFB genomen totdat een herstructureringsplan voor IFB kan worden uitgevoerd; in een tweede fase zouden in het kader van een herstructureringsplan voor IFB maatregelen worden uitgewerkt en bij die gelegenheid zouden de reddingsmaatregelen in kapitaal kunnen worden omgezet.
81. In de preambule van de overeenkomst bevestigt de NMBS haar voornemen om "haar goedkeuring te hechten aan een door de NMBS te onderschrijven kapitaalverhoging van IFB ten belope van ongeveer 60 miljoen euro door omzetting van vorderingen van de NMBS op IFB en om IFB eveneens een bijkomend bedrag van 20 miljoen euro ter beschikking te stellen, waarvan 5 miljoen euro onmiddellijk zou worden vrijgegeven."
82. Artikel 2 van de kaderovereenkomst tussen de NMBS en IFB voorziet in twee pakketten maatregelen, namelijk een pakket "reddingsmaatregelen" en een pakket "herstructureringsmaatregelen".
2.3.1. Modaliteiten en voorwaarden voor de reddingsmaatregelen
83. Het eerste deel van artikel 2 voorziet in een pakket van drie reddingsmaatregelen:
(1) een terugvorderbaar voorschot van 5 miljoen euro;
(2) het toekennen van een kredietfaciliteit van maximaal 15 miljoen euro, en
(3) het verlenen van een voorlopig uitstel van betaling voor alle schulden van IFB.
84. Artikel 3 van de kaderovereenkomst bepaalt dat de rentevoet op het terugvorderbare voorschot en op de opgenomen sommen van de kredietfaciliteit ten minste gelijk moet zijn aan de door de Commissie gehanteerde referentierentevoet voor overheidssteun [58]. Het bepaalt tevens dat de rente bij het kapitaal zal worden gevoegd. De betaling ervan zal plaatsvinden op het ogenblik waarop de nog uitstaande vorderingen worden betaald.
85. Het voorschot en de kredietfaciliteit worden voorlopig ter beschikking gesteld teneinde te voldoen aan de dringende financiële behoeften van IFB. Zij zullen in het kader van het nog op te stellen herstructureringsplan in kapitaal worden omgezet.
86. Wat met name de toekenning van een kredietfaciliteit van maximaal 15 miljoen euro betreft, mag IFB de schuldvorderingen van de NMBS op IFB vanaf 1 januari 2003 in mindering brengen, met uitzondering van een factuur van 31 januari 2003 ten belope van 8 miljoen euro.
87. Het voorlopige uitstel van betaling heeft betrekking op alle schulden van IFB die op 31 december 2002 waren gefactureerd, met inbegrip van een factuur van 31 januari 2003 ten belope van 8 miljoen euro, en van de schulden waarvan het bedrag op 31 december 2002 zeker en vaststaand was maar die in regel niet werden gefactureerd. Het aan de NMBS verschuldigde bedrag beliep in totaal 63 miljoen euro. Bovendien moet het betrokken bedrag worden verhoogd met de gebruikelijke rente op achterstallige betalingen van [tussen 1 en 2] per duizend per volledige periode van tien dagen [59], of met de wettelijk vastgestelde rente. De rente wordt bij het kapitaal gevoegd en wordt betaald op het ogenblik dat de hoofdvordering wordt betaald.
88. De door IFB aan de NMBS verschuldigde rente op de schuld en de kredietfaciliteit beliep 2,2 miljoen euro in 2002, 3,9 miljoen euro in 2003 en 4,7 miljoen euro in 2004. In de kaderovereenkomst is bepaald dat de rente wordt betaald op het ogenblik dat de vorderingen worden betaald.
89. IFB heeft tegenover de NMBS ook afstand gedaan van de verjaring van haar schulden. Al deze maatregelen zijn, met uitzondering van het terugvorderbaar voorschot, ten uitvoer gelegd van bij de ondertekening van het contract op 7 april 2003. Het uitstel van betaling van zijn kant was de facto al verleend voordat de kaderovereenkomst werd gesloten en is door de kaderovereenkomst geformaliseerd.
2.3.2. Modaliteiten en voorwaarden voor de herstructureringsmaatregelen
90. Het tweede deel van artikel 2 van de kaderovereenkomst bepaalt dat door de raden van bestuur van de NMBS en IFB herstructureringsmaatregelen zullen worden uitgewerkt en dat deze vervolgens ter goedkeuring aan de Belgische overheid zullen worden voorgelegd.
91. Artikel 4 van de kaderovereenkomst betreffende de modaliteiten voor de herstructureringsmaatregelen luidt als volgt:
"Partijen bevestigen hun voornemen om — indien en voor zover deze conform zijn met een herstructureringsplan dat is goedgekeurd door hun beider raden van bestuur, door de Belgische overheid, en voor zover vereist, door de EC, en onder voorbehoud van goedkeuring door de aandeelhouders van IFB — de volgende maatregelen ten uitvoer te leggen:
- de omzetting in kapitaal van het terugvorderbaar voorschot t.b.v. 5 miljoen euro;
- de omzetting in kapitaal van het opgenomen gedeelte van de kredietfaciliteit t.b.v. maximum 15 miljoen euro […];
- de omzetting in kapitaal van de schulden […] van 63 miljoen euro;
- eventueel, en op voorwaarde dat beide partijen daarover akkoord zijn, een bijkomende kapitaalverhoging […]".
92. De Belgische regering heeft de Commissie tijdens de bijeenkomsten van 12 december 2003 en 16 september 2005, alsmede bij brief van 13 januari 2004, 28 januari 2005, 25 maart 2005 en 30 juni 2005 in kennis gesteld van de bijzonderheden betreffende de herstructureringsmaatregelen, die ad-hocmaatregelen omvatten welke door IFB zijn getroffen ten aanzien van haar dochtermaatschappijen die in Frankrijk terminals exploiteren, alsmede van een herstructureringsplan voor IFB en van een kapitaalverhoging.
93. Op dit ogenblik is nog geen van deze maatregelen ten uitvoer gelegd.
2.3.2.1. Ad-hocmaatregelen die door IFB zijn getroffen ten aanzien van haar dochtermaatschappijen die in Frankrijk terminals exploiteren
94. Zoals hiervoor is uiteengezet, heeft IFB voor haar Franse dochtermaatschappijen een strategie van desinvestering gevolgd. Dit beleid is vrijwel voltooid (zie de beschrijving van de participaties hiervoor); voorts werden de patronaatsverklaringen ingetrokken.
2.3.2.2. Het herstructureringsplan
95. IFB en de NMBS hebben met adviesbureau McKinsey een herstructureringsplan voor IFB uitgewerkt dat de economische levensvatbaarheid van IFB op de lange termijn garandeert. Dit plan bestaat uit twee delen:
- Herstructurering van de activiteit "IFB Logistics"
- Herstructurering van de activiteit "IFB Terminals"
96. Met de uitvoering van het herstructureringsplan werd een begin gemaakt in 2003 en het zal worden voltooid in 2005. In het plan was voorzien dat IFB een exploitatiewinst van 0,5 miljoen euro in 2003 en van 0,8 miljoen euro in 2004 zou behalen, na in 2002 bedrijfsverliezen van 13,4 miljoen euro te hebben geleden. Onderstaande tabel laat de voor 2002-2004 verwachte verdeling zien van de winst en het verlies tussen de verschillende activiteiten:
| 2002 | 2003 | 2004 |
Dochtermaatschappijen | […] | […] | […] |
IFB Terminals | […] | […] | […] |
IFB Logistics | […] | […] | […] |
Totaal | - 13,4 | 0,5 | 0,8 |
97. De in 2003 behaalde resultaten bleven achter bij de verwachtingen, aangezien het bedrijfsresultaat –2,9 miljoen euro beliep. Dit was voornamelijk te wijten aan de verliezen van de dochterondernemingen (verliezen van […] miljoen euro in plaats van een winst van […] miljoen euro) en aan de geringe winst van IFB Logistics (winst van […] miljoen euro in plaats van een verwachte winst van […] miljoen euro).
98. De in 2004 behaalde resultaten overtroffen de verwachtingen, aangezien het bedrijfsresultaat een winst van 5,7 miljoen euro vertoonde. Hieraan werd door IFB Logistics voor […] miljoen euro, door IFB Terminals voor […] miljoen euro en door de dochterondernemingen voor […] miljoen euro bijgedragen.
99. In het herstructureringsplan wordt tevens de noodzaak aangedragen van nieuwe investeringen ten belope van […] miljoen euro. De voor de verschillende sectoren geplande herstructureringsmaatregelen alsook de behoefte aan nieuwe investeringen dienen meer in detail te worden gepresenteerd.
a) Herstructurering van de logistieke activiteit
100. Ten aanzien van de activiteit "IFB Logistics" was in het herstructureringsplan voor 2003 een exploitatiewinst van […] miljoen euro geraamd, na een verlies van […] miljoen euro in 2002. Ter verwezenlijking hiervan bevatte het plan in totaal negen maatregelen die een besparing van […] miljoen euro mogelijk zouden maken. Door de daling van het volume aan conventioneel vervoer, die naar verwachting een verlies van […] miljoen euro met zich zal meebrengen, zou de totale verbetering dus […] miljoen euro belopen. Onderstaande tabel bevat de negen maatregelen:
Maatregelen | Besparing |
1.Vermindering van de loonkosten | […] miljoen |
2.Advies en outsourcing | […] miljoen |
3.Waardevermindering en bijzondere afschrijvingen | […] miljoen |
4.Stopzetting van niet-rendabele afdelingen van het North European Network | […] miljoen |
5.Volumedaling van het conventioneel vervoer | […] miljoen |
6.Terugneming uit voorzieningen onderhoud wagons | […] miljoen |
7.Groei van het intermodaal vervoer | […] miljoen |
8.Herziening van de Railbarge-overeenkomst (verhoging van de prijzen en verwezenlijkte re-engineering) | […] miljoen |
9.Verhoging van de provisies van de vertegenwoordigers (agent) | […] miljoen |
10.Verlaging van de algemene kosten | […] miljoen |
101. De herstructureringsmaatregelen bestonden dus in hoofdzaak uit een prijsverhoging, gekoppeld aan een nieuw design van de producten, terugneming van voorzieningen en bijzondere afschrijvingen, vermindering van de loonkosten en de algemene kosten, en stopzetting van onrendabele activiteiten.
102. Voor de activiteit "IFB Logistics" zal de herstructurering volgens de planning dus tussen medio-2003 en medio-2004 zijn voltooid.
b) Herstructurering van de terminalactiviteit
103. De herstructurering van de activiteit "IFB Terminals" daarentegen zal waarschijnlijk drie jaar in beslag nemen. Volgens de verwachtingen zullen de operationele verliezen van deze activiteit van […] miljoen euro in 2002 dalen tot […] miljoen euro in 2003 en […] miljoen euro in 2004, alvorens 2005 af te sluiten met een exploitatiewinst van […] miljoen euro. Ter verwezenlijking hiervan bevatte het plan de volgende acht maatregelen:
Maatregelen | Besparing |
1.Mainhub:PersoneelsinkrimpingComputeraanpassingenVermindering van de afschrijvingen en terugneming van de voorzieningenUitbreiding van het aantal bewerkingen | […] miljoen |
2.CirkeldijckVermindering van de operaties op het terreinVerkoop van activaVerhuring van de terminalVermindering van het volumePersoneelsinkrimping | […] miljoen |
3.ZomerwegTransfer RailbargeVergroting van het volumeUitbreidingenInvesteringen | […] miljoen |
4.Dry port MuizenVermindering van personeelskosten dankzij het nieuwe bewakingssysteemVergroting van het volume | […] miljoen |
5.SchijnpoortVergroting van het volumeVermindering van de exploitatiekosten | […] miljoen |
6.RenoryVerkoop van een stackerStopzetting financiële solidariteit van IFB | […] miljoen |
7.Bressoux: Sluiting van de terminal | […] miljoen |
104. De belangrijkste maatregelen hebben dus betrekking op de terminals Mainhub, Cirkeldijck en Zomerweg. In onderstaande paragrafen worden zij meer gedetailleerd uiteengezet.
105. Mainhub. Mainhub zal tussen medio 2003 en eind 2005 volledig worden gereorganiseerd, hetgeen — met name dankzij omvangrijke computeraanpassingen — personeelsinkrimping in combinatie met een verhoging van het aantal bewerkingen mogelijk zal maken. Daardoor kan worden gezorgd voor een betere capaciteitsbezetting van de terminal, die in 2002 slechts voor […] % is gebruikt.
106. Cirkeldijck. In de Cirkeldijck-terminal zal IFB haar samenwerking met Hesse NoordNatie (HNN) verstevigen. HNN zal de operaties op het terrein overnemen, terwijl IFB de planning en het laden van het spoorvervoer behoudt. […].
107. Zomerweg. De Zomerweg-terminal zal van bimodale terminal tot een trimodale terminal worden omgevormd, waarbij alle Railbarge-vervoer naar deze terminal wordt overgebracht. In deze context worden het terrein en het perron uitgebreid, worden het terrein, de ingang en de wegen aangepast en zullen investeringen in materieel vereist zijn.
c) Noodzaak van investeringen
108. Voor de herstructurering van Mainhub en de herstructurering van Zomerweg zijn nieuwe investeringen, elk ten belope van […] miljoen euro, vereist. Terzelfder tijd kan het benodigde bedrag door de verkoop van de portaalkraan van de Cirkeldijck-terminal worden verlaagd tot in totaal […] miljoen euro.
2.3.2.3. Kapitaalverhoging
109. Bij schrijven van 28 januari 2005 heeft de Belgische regering de Commissie ervan in kennis gesteld dat het leidinggevend personeel van zowel IFB als de NMBS van oordeel is dat het herstructureringsplan vergezeld moet gaan van een verhoging van het kapitaal van IFB, zoals in de kaderovereenkomst was vastgelegd. Het benodigde bedrag, ten opzichte van de ramingen van de kaderovereenkomst iets naar boven bijgesteld, zou 96,5 miljoen euro bedragen.
110. De kapitaalverhoging zal als volgt verlopen: eerst worden de schulden van IFB jegens de NMBS, die 78 miljoen euro belopen, en de rente over die schulden, die eind 2005 13,5 miljoen euro zal belopen, in kapitaal omgezet. De oorsprong van deze schulden ligt in reddingsmaatregelen 1 en 2, dat wil zeggen het uitstel van betaling en de kredietfaciliteit. Vervolgens zal de NMBS de rest, dat wil zeggen 5 miljoen euro, in natura inbrengen. De procedure komt dus overeen met de in artikel 4 van de kaderovereenkomst vastgelegde procedure.
111. De inbreng in natura bestaat uit de participatie van de NMBS in TRW. Deze deelneming beloopt, zoals hierboven is uiteengezet, 47 %; IFB bezit al een participatie van 0,9 % in de onderneming. TRW exploiteert terminals in Antwerpen, Zeebrugge, Oostende, Charleroi, Luik, Brussel, Etge, Genk en Muizen, en biedt vrachttreinen aan voor 11 EU-landen.
112. De kapitaalverhoging bedraagt meer dan bij het afsluiten van de kaderovereenkomst tussen IFB en de NMBS was bepaald — hierin was namelijk een kapitaalverhoging van 80 miljoen euro vastgesteld — maar minder dan het voorstel van adviesbureau McKinsey, dat in het herstructureringsplan uitging van een kapitaalverhoging van 120 miljoen euro.
113. De Belgische regering is van mening dat IFB met deze kapitaalverhoging, na de aftrek van kapitaal om de overgedragen verliezen te dekken, een eigen vermogen van 23,9 miljoen euro zou hebben, wat een gezonde kapitaalstructuur zou zijn met een aan de activiteiten van IFB aangepaste verhouding tussen de financiering met eigen vermogen en de schulden.
114. De solvabiliteitscoëfficiënt, dat wil zeggen de verhouding tussen eigen vermogen en passiva, van IFB voor en na de kapitaalverhoging wordt door onderstaande tabel verduidelijkt:
| Situatie op 30.06.2005 | Voorgestelde verhoging | Situatie na verhoging |
Eigen vermogen | - 72,6 | 96,5 | 23,9 |
Voorzieningen en belastinglatenties | 14,3 | | 14,3 |
Schulden | 125,6 | - 91,5 | 34,1 |
Totaal passiva | 67,3 | | 72,3 |
Solvabiliteits-coëfficiënt | | | 33 % [60] |
115. De kapitaalverhoging is voorzien voor het tweede halfjaar 2005, na goedkeuring door de Europese Commissie en de Raad van Bestuur van de NMBS.
116. In tegenstelling tot hetgeen in artikel 4 van de kaderovereenkomst is bepaald, is het plan voor de kapitaalverhoging niet ter goedkeuring aan de Belgische regering voorgelegd. De Belgische regering is van mening dat een dergelijke goedkeuring niet vereist is omdat het een louter commerciële beslissing van de NMBS betreft, die deze onderneming zonder goedkeuring van de staat kan nemen.
2.4. Financiële ontwikkeling van IFB sinds de sluiting van de kaderovereenkomst
117. De economisch-financiële situatie van IFB is sedert de sluiting van de kaderovereenkomst in april 2003 aanmerkelijk verbeterd. Zo vertoonde het bedrijfsresultaat een positieve ontwikkeling van -47,36 miljoen euro in 2002 tot 5,74 miljoen euro in 2004. Het resultaat van het boekjaar voor aftrek van belastingen steeg van -109,76 miljoen euro in 2002 naar 13,21 miljoen euro in 2004.
118. Onderstaande tabel bevat een kort overzicht van de ontwikkeling van de belangrijkste economische en financiële indicatoren van IFB:
Tabel: Economisch-financiële situatie van IFB (in 000 euro)
| 31.12.2002 (aan audit onder-worpen) | 30.09.2003 | 31.12.2003 (aan audit onder-worpen) | 30.09.2004 | 31.12.2004 (aan audit onder-worpen) |
Verkopen en verrichtingen | 65377 | 43184 | 59091 | 61369 | 85751 |
Waarvan omzet | 63669 | 42445 | 58079 | 59903 | 83343 |
Kosten van verkopen en verrichtingen | 112734 | 43781 | 62051 | 58759 | 80011 |
Bedrijfsresultaat | (47357) | (1336) | (2960) | 2610 | 5740 |
Financieel resultaat | (3034) | — | (4458) | (3247) | (3303) |
Uitzonderlijk resultaat | (59369) | — | 7342 | 6754 | 10773 |
Resultaat van het boekjaar voor aftrek van belastingen | (109760) | (1200) | (76) | 6117 | 13210 |
Cash Flow | | (101) | | | |
Eigen vermogen | (84068) | (85277) | (83941) | (77775) | (74850) |
119. De verbetering van de economisch-financiële situatie is enerzijds te danken aan de uitvoering van het herstructureringsplan en anderzijds aan de strategie van afsplitsing ten aanzien van de participaties.
120. Ook in het eerste halfjaar 2005 boekte IFB winst: het bedrijfsresultaat beliep 1,6 miljoen euro en het resultaat voor aftrek van belastingen was 2,2 miljoen euro.
2.4.1. Uitvoering van het herstructureringsplan
121. Voor de tenuitvoerlegging van het herstructureringsplan moet een onderscheid worden gemaakt tussen de maatregelen die gevolgen hebben voor alle activiteiten van IFB en de specifieke maatregelen voor IFB Logistics en IFB Terminals.
2.4.1.1. Maatregelen die gevolgen hebben voor alle activiteiten van IFB
122. Door de sluiting van een nieuwe arbeidsovereenkomst op het niveau van de onderneming en de wijziging van het arbeidsreglement kon een hogere participatiegraad (het aantal dagen dat per jaar moet worden gewerkt is toegenomen) tegen geringere kosten (de vergoeding voor weekendwerk en ploegenarbeid is verlaagd). De administratieve en commerciële diensten zijn centraal in Berchem ondergebracht, waardoor de vestiging in Gent kon worden gesloten en de capaciteit van die in Zeebrugge kon worden teruggebracht.
123. Deze maatregelen hebben bijgedragen tot vermindering van het benodigde personeel en verlaging van de algemene kosten.
2.4.1.2. Specifieke maatregelen voor IFB Terminals
124. Naast de in het herstructureringsplan vervatte maatregelen zijn nog twee maatregelen genomen: Voor de terminal te Cirkeldijck is de prijs voor de afhandeling naar boven bijgesteld. Meer algemeen zijn de vervoersstromen geanalyseerd en vervolgens in onderling overleg met de klanten geheroriënteerd.
125. Dankzij al deze maatregelen, en door de groei van de behandelde hoeveelheden, kon IFB Terminals al in 2004 weer winstgevend worden, met een winst voor belastingaftrek van […] euro, na een verlies na belastingaftrek van […] miljoen euro in 2003. De doelstelling die in het herstructureringsplan was vastgelegd is dus ruimschoots gehaald (ter herinnering: in het herstructureringsplan was op een verlies van […] euro gerekend.)
2.4.1.3. Specifieke maatregelen voor IFB Logistics
126. Naast de in het herstructureringsplan vervatte maatregelen heeft IFB Logistics een diepgaande analyse verricht van zijn spoorvervoerproducten; hierbij zijn onrendabele producten aangetroffen, die IFB sindsdien niet meer produceert.
127. Voor andere producten heeft deze analyse de noodzaak van verbeteringen op technisch niveau aangetoond. Deze verbeteringen zijn aangebracht, met name voor de sector intermodaal containervervoer.
128. Dankzij al deze maatregelen kon IFB Logistics al in 2003 weer winstgevend worden met een winst voor belastingaftrek van […] euro. In 2004 waren de resultaten verder verbeterd tot […] miljoen euro. IFB Logistics heeft de doelstelling die voor 2003 in het herstructureringsplan was vastgelegd ([…] miljoen euro) dat jaar niet kunnen halen, maar wel in 2004 (het streefcijfer was […] miljoen euro).
2.5. Budget
129. Het geraamde totaalbedrag van de reddingsmaatregelen beloopt maximaal 78 miljoen euro [61].
130. Het totaalbedrag van de beoogde kapitaalverhoging beloopt 96,5 miljoen euro, waarvan 78 miljoen euro zal resulteren uit de omzetting van de bestaande schulden (63 miljoen) en van de reddingsmaatregelen (15 miljoen) in kapitaal, en 13,5 miljoen euro uit de omzetting van de gekapitaliseerde rente in kapitaal. Nog eens 5 miljoen euro zal door de NMBS in natura worden ingebracht, door overdracht van de deelneming van de NMBS in TRW aan IFB.
2.6. Terbeschikkingstelling van financiële middelen en looptijd
131. In haar brieven van 28 januari en 25 maart 2005 verklaart de Belgische regering dat de maatregelen 2 (kredietlijn van 15 miljoen euro) en 3 (uitstel van betaling voor de bestaande schulden van 63 miljoen euro) van het deel "reddingsmaatregelen" met ingang van 7 april 2003 door de NMBS en IFB ten uitvoer zijn gelegd. Daarentegen had IFB het in maatregel 1 vastgelegde terug te betalen voorschot niet nodig.
132. In de kaderovereenkomst is bepaald dat, behoudens omzetting in kapitaal in het kader van een goedgekeurd eventueel herstructureringsplan of enige andere overeengekomen maatregel van vergelijkbare strekking, alle bedragen vermeerderd met rente twaalf maanden nadat zij door de NMBS ter beschikking van IFB zijn gesteld dienen te worden terugbetaald. Aangezien het leidinggevend personeel van IFB en van de NMBS had ingestemd met het principe van een kapitaalverhoging, is volgens hen de leningovereenkomst stilzwijgend verlengd totdat de kapitaalverhoging plaatsvindt. IFB accumuleert intussen de in de kaderovereenkomst vastgelegde rente, te weten de gebruikelijke rente op achterstallige betalingen van [tussen 1 en 2]‰ per volledige periode van 10 dagen [62], of een wettelijk vastgestelde rentepercentage. De gemiddelde rente bedraagt [tussen 3,6 en 7,2] %. De volledige rente moet worden betaald op het ogenblik dat de schuld wordt voldaan of wordt omgezet in maatschappelijk kapitaal.
133. De kapitaalverhoging zal in het tweede halfjaar 2005 plaatsvinden, na goedkeuring ervan door de Commissie.
3. BEOORDELING
3.1. Beoordeling van het steunkarakter van de reddings- en herstructureringsmaatregelen
134. Overeenkomstig artikel 87, lid 1, van het Verdrag "zijn steunmaatregelen van de staten of in welke vorm ook met staatsmiddelen bekostigd, die de mededinging door begunstiging van bepaalde ondernemingen of bepaalde producties vervalsen of dreigen te vervalsen, onverenigbaar met de gemeenschappelijke markt, voorzover deze steun het handelsverkeer tussen de lidstaten ongunstig beïnvloedt".
3.1.1. Steunmaatregel van de staat of met staatsmiddelen bekostigd
135. Daarom rijst allereerst de vraag of het bij de financiële steun van de NMBS aan IFB om "steunmaatregelen van de staten of met staatsmiddelen bekostigd" gaat. Volgens de jurisprudentie van het Hof van Justitie in de zaak Stardust Marine [63] wordt aan dit criterium voldaan indien het om staatsmiddelen gaat en indien de beslissing om deze te verlenen aan de betrokken lidstaat, in casu België, kan worden toegerekend.
3.1.1.1. Staatsmiddelen
136. Wat het aspect "staatsmiddelen" betreft, constateert de Commissie dat de NMBS als een openbaar bedrijf in de zin van artikel 2 van Richtlijn 2000/52/EG [64] van de Commissie moet worden aangemerkt: de Belgische staat bezit 100 % van het geplaatst kapitaal van de NMBS en de Raad van Bestuur en de gedelegeerd bestuurder worden bij koninklijk besluit benoemd na overleg in de Raad van ministers. Derhalve is zowel aan criterium a) als aan criterium c) van de tweede alinea van artikel 2 van de richtlijn voldaan.
137. In dit verband "... volgt reeds uit de rechtspraak van het Hof dat artikel 87, lid 1, EG alle geldelijke middelen omvat die de overheid daadwerkelijk kan gebruiken om ondernemingen te steunen, ongeacht of deze middelen permanent deel uitmaken van het vermogen van de staat. Dus ook al zijn de bedragen die overeenkomen met de betrokken maatregel niet permanent in het bezit van de schatkist, dan nog volstaat het feit dat zij constant onder staatscontrole, en daarmee ter beschikking van de bevoegde nationale autoriteiten staan, om ze als staatsmiddelen aan te merken" [65].
138. Op grond hiervan is de Commissie van mening dat de ter beschikking van IFB gestelde bedragen als staatsmiddelen zijn aan te merken.
3.1.1.2. Toerekenbaarheid
3.1.1.3. Wat het criterium van de toerekenbaarheid van de maatregelen aan de betrokken staat betreft, bepaalt het arrest in de zaak Stardust Marine dat het feit "dat een openbaar bedrijf onder staatscontrole staat, op zich dus niet volstaat om door dit bedrijf genomen maatregelen, zoals de onderhavige financiële steunmaatregelen, aan de staat toe te rekenen. Daarnaast dient te worden nagegaan of de overheid op een of andere manier bij de vaststelling van de maatregelen was betrokken." [66]
139. Uit de jurisprudentie van het Hof blijkt dus dat het criterium van de toerekenbaarheid aan de staat van geval tot geval door de Commissie dient te worden onderzocht. Het Hof geeft toe dat het "…juist als gevolg van de bevoorrechte betrekkingen tussen de staat en openbare bedrijven voor derden" in de regel "zeer moeilijk" zal "zijn om in een concreet geval aan te tonen dat door dergelijke bedrijven genomen steunmaatregelen werkelijk in opdracht van de overheid zijn getroffen. Dienaangaande kan niet worden geëist dat op basis van een gedetailleerd onderzoek wordt aangetoond dat de overheid het openbare bedrijf er concreet toe heeft aangezet de betrokken steunmaatregelen te nemen." [67] Op deze gronden dient volgens hetzelfde arrest "... te worden aangenomen dat de toerekenbaarheid aan de staat van een door een openbaar bedrijf genomen steunmaatregel kan worden afgeleid uit een samenstel van aanwijzingen die blijken uit de omstandigheden van de zaak en de context waarin deze maatregel is genomen".
140. In het onderhavige geval moet, wat de toerekenbaarheid betreft, een onderscheid worden gemaakt tussen de periode vóór de sluiting van de kaderovereenkomst op 7 april 2003 en de periode daarna.
141. Wat de periode vóór de sluiting van de kaderovereenkomst betreft, rijst de vraag of het besluit van de NMBS om geen betaling te eisen voor de geleverde vervoerdiensten vanaf 2000 aan de Belgische staat is toe te rekenen.
142. De Commissie beschikt over geen gegevens met betrekking tot de vraag hoe en waarom de NMBS heeft besloten geen betaling van haar uitstaande facturen te eisen. Maar omdat deze facturen in de periode van eind 2000 tot begin 2003 systematisch niet blijken te zijn betaald, betwijfelt de Commissie toch of een dergelijk besluit door het middenkader van de onderneming kon worden genomen. Normaal moeten de auditors van de onderneming dit hebben geconstateerd en de bedrijfsleiding — en eventueel ook de met de NMBS belaste regeringscommissaris — hiervan in kennis hebben gesteld. De Commissie heeft in dit stadium dus vermoedens dat het besluit van de NMBS om vanaf eind 2000 geen betaling meer te eisen van haar facturen aan IFB, toerekenbaar is aan de Belgische staat en verzoekt de Belgische autoriteiten haar alle nuttige elementen te bezorgen om na te gaan hoe dit besluit tot stand is gekomen.
143. Wat de periode na de sluiting van de kaderovereenkomst betreft, resulteerde de analyse van het dossier door de Commissie in drie concrete aanwijzingen voor toerekenbaarheid van de reddings- en herstructureringsmaatregelen ten behoeve van IFB aan de Belgische staat:
- Het feit dat het herstructureringsplan ter goedkeuring aan de Belgische staat is voorgelegd
- De artikelen in de pers waaruit blijkt dat de Belgische regering gedurende 2003 een sterke invloed op de NMBS had
- Omvang, inhoud en voorwaarden van de kaderovereenkomst.
a) De goedkeuring door de overheid
144. In zijn arresten Van der Kooy [68], Italië/Commissie [69] en Commissie/Frankrijk [70], beschouwde het Hof de steun als staatssteun omdat hij toegekend werd met instemming van de overheid. Terwijl dit element in het arrest Van der Kooy volstaat om de steun als dusdanig te beoordelen, wordt in de arresten Italië/Commissie en Commissie/Frankrijk de goedkeuring gecombineerd met andere elementen die de invloed van de overheid aantonen [71]. De Commissie heeft in haar recente beschikking betreffende het Space Park Development GmbH, de eerste beschikking waarbij zij zich heeft gebaseerd op het Stardust Marine-arrest, geoordeeld dat de steun moest worden aangemerkt als staatssteun, omdat voor de toekenning van de betrokken lening toelating moest worden gegeven door de overheid van de deelstaat Bremen [72]. Daarom is het feit dat een maatregel ter goedkeuring aan de lidstaat wordt voorgelegd een aanwijzing van de toerekenbaarheid aan de staat.
145. In de onderhavige zaak zijn de Raden van Bestuur van de NMBS en IFB op grond van artikel 2 van de kaderovereenkomst verplicht het herstructureringsplan ter goedkeuring voor te leggen aan de Belgische staat. Dit vormt er een extra aanwijzing voor dat de besluiten van de NMBS in onderhavig geval aan de Belgische staat toe te rekenen zijn.
146. De Belgische regering heeft de Commissie inmiddels laten weten dat, in tegenstelling tot hetgeen in de kaderovereenkomst is vastgelegd, de NMBS en IFB geen herstructureringsplan ter goedkeuring aan de Belgische regering hebben voorgelegd, aangezien dit een inbreuk op de commerciële autonomie van de NMBS zou zijn geweest.
147. Volgens de Commissie blijft de indicatie van de toerekenbaarheid desondanks in stand: het lijkt uitgesloten dat de twee partijen bij de overeenkomst, de NMBS en IFB, een dergelijke bepaling in de overeenkomst zouden hebben opgenomen indien er geen invloed in deze zin was van de Belgische regering. Het feit dat de Belgische regering er niet op heeft aangedrongen om formeel over de uitvoering van de herstructurering te worden geraadpleegd volstaat daarom niet om informele beïnvloeding door de Belgische regering bij de voorbereiding van de kaderovereenkomst, waarin de reddings- en herstructureringsmaatregelen al in grote lijnen zijn vervat, uit te sluiten. In ieder geval betekent het feit dat de Belgische staat de controlemiddelen waarover hij beschikte niet heeft gebruikt, niet dat de maatregelen niet aan hem kunnen worden toegerekend.
b) Berichten in de pers
148. Aanwijzingen voor bemoeienis van de Belgische regering in deze zaak zijn tevens in de pers te vinden [73]. Zo wordt in een artikel dat in La libre Belgique van 19 mei 2003 is verschenen [74] de persdienst van de NMBS geciteerd, waarin het feit dat België de reddingsmaatregelen op 19 mei 2003 nog niet bij de Commissie had aangemeld, terwijl de kaderovereenkomst op 7 april 2003 was ondertekend, verklaard wordt door het feit dat de federale overheid zich er nog over moet [moest] uitspreken. In een artikel dat in maart 2003 is verschenen in www.cheminots.be wordt Karel Vinck, destijds gedelegeerd bestuurder van de NMBS, met betrekking tot de dossiers ABX en IFB als volgt geciteerd: "Hij verlangt een voldoende ruime manœuvreerruimte voor het management van de onderneming". Hieruit valt op te maken dat de bedrijfsleiding van de NMBS vond dat de staat zich teveel met deze zaken bemoeide.
c) Omvang, inhoud en voorwaarden van de kaderovereenkomst
149. Meer algemeen herinnert de Commissie eraan dat, volgens punt 56 van hogervermeld arrest-Stardust Marine "elke andere aanwijzing waaruit in het concrete geval blijkt dat de overheid bij de vaststelling van een maatregel is betrokken of dat het onwaarschijnlijk is dat zij hierbij niet betrokken is, mede gelet op de omvang van deze maatregel, op de inhoud ervan of op de eraan verbonden voorwaarden" in aanmerking moet worden genomen om de toerekenbaarheid van een maatregel aan de lidstaat in kwestie vast te stellen. Aangezien het hier omvangrijke herstructureringsmaatregelen betreft, waar de goedkeuring door de Belgische autoriteiten aan vooraf moet gaan, is de Commissie van mening dat de omvang, de inhoud en de voorwaarden van de kaderovereenkomst in dit concrete geval extra aanwijzingen voor de toerekenbaarheid vormen.
d) Conclusie
150. De Commissie is in deze fase dan ook van mening dat de financiële steun voor wat de periode na de sluiting van de kaderovereenkomst betreft, aan de staat is toe te rekenen. Er moet dus worden nagegaan of de steun de begunstigde een voordeel heeft opgeleverd dan wel of, integendeel, België heeft gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan.
3.1.2. Financiële steun aan bepaalde ondernemingen
151. Als blijkt dat het besluit van de NMBS om vanaf eind 2000 geen betaling van haar facturen aan IFB meer te eisen, aan de Belgische staat is toe te rekenen, moet worden nagegaan of deze steun ook door een particulier investeerder in een markteconomie zou zijn verleend.
152. Aangezien het besluit van de NMBS om de kaderovereenkomst met IFB te ondertekenen aan België valt toe te rekenen, moet daarna worden nagegaan of de NMBS, door IFB eerst reddingssteun en vervolgens herstructureringssteun te verlenen, dit bedrijf ten opzichte van andere bedrijven heeft bevoordeeld. Dit is niet het geval indien de NMBS zich tegenover IFB heeft opgesteld zoals een bedachtzaam investeerder/bedachtzaam kredietverlener in een markteconomie zou hebben gedaan. Om deze tweede beoordeling te kunnen maken, moet een onderscheid worden gemaakt tussen de reddingsmaatregelen en de herstructureringsmaatregelen.
3.1.2.1. Het niet betalen van de facturen van de NMBS door IFB tussen 2000 en 20033
153. Wat het niet betalen van de facturen van de NMBS door IFB betreft, moet worden nagegaan of een bedachtzaam schuldeiser in de plaats van de NMBS zou hebben aanvaard dat IFB zijn facturen niet betaalde, dan wel of een bedachtzaam schuldeiser zich in de plaats van de NMBS tot de rechter zou hebben gewend om de betaling van zijn facturen te verkrijgen.
154. In dit verband moet er allereerst op worden gewezen dat het een gangbare handelspraktijk is om aan een klant die tijdelijke liquiditeitsproblemen heeft, maar die voor het overige economisch gezond is, in afwachting van de betaling van de facturen veeleer een stilzwijgende termijn toe te kennen dan hem onmiddellijk voor het gerecht te dagen.
155. Kennelijk zijn de financiële moeilijkheden van de onderneming pas in de loop van 2002 zichtbaar geworden (zie onderstaande beschrijving van de financiële situatie). Het feit dat IFB in 2001 van de commerciële bank […] een lening van meer dan 4 miljoen euro tegen marktrente heeft gekregen, en dat het eigen vermogen van IFB eind 2001 28 miljoen euro beliep wijst eveneens in die richting.
156. Niettemin kan de Commissie in dit stadium niet uitsluiten dat de NMBS als moedermaatschappij van IFB had moeten inzien dat er in 2001 bij IFB verder stroomopwaarts problemen waren.
157. Pas op zijn vroegst vanaf 2001 had een particulier investeerder dus voorzichtiger kunnen handelen. Het valt moeilijk te zeggen vanaf wanneer een particulier schuldeiser zou hebben getracht terugbetaling van zijn vorderingen of aanvullende zekerheden te verkrijgen; momenteel is de Commissie van oordeel dat dit ogenblik uiterlijk op 19 september 2002 was aangebroken, toen de gedelegeerd bestuurder van IFB twee bedrijfsrevisoren ermee belastte een speciaal verslag over de financiële situatie van IFB op te stellen.
158. Deze gang van zaken heeft geleid tot de ontwikkeling van de kaderovereenkomst, waarin uitdrukkelijk reddings- en herstructureringsmaatregelen zijn vastgelegd. Door aan IFB diensten op het gebied van het spoorvervoer te blijven leveren heeft de NMBS op zijn vroegst in de loop van 2001 en uiterlijk sinds 19 september 2002 aan IFB economische voordelen verschaft, die als staatssteun moeten worden beschouwd. Door IFB niet uiterlijk vanaf dat ogenblik voor het gerecht te dagen ter verkrijging van de betaling van de facturen uit 2000 heeft de NMBS, ook wat het niet betalen van deze facturen betreft, IFB een voordeel verschaft.
159. De NMBS heeft derhalve op zijn vroegst sinds 2001 en uiterlijk sinds 19 september 2002 de facto steun verleend aan IFB; de kaderovereenkomst heeft deze steun alleen maar officieel gemaakt.
3.1.2.2. Reddingsmaatregelen
160. De reddingsmaatregelen zijn hierboven in deel 2 beschreven. Het ging om:
- Verlening van uitstel van betaling voor de schuld van 63 miljoen euro,
- Verlening van een kredietfaciliteit van 15 miljoen euro
- Verlening van een terugvorderbaar voorschot van 5 miljoen euro
161. Hierbij moet een onderscheid worden gemaakt tussen de maatregelen die de NMBS heeft getroffen als schuldeiser van IFB, te weten de verlening van uitstel van betaling voor de reeds bestaande schulden ten belope van 63 miljoen euro, en de maatregelen die de NMBS heeft getroffen als investeerder in IFB, namelijk verlening van een nieuwe kredietfaciliteit van 15 miljoen euro en verstrekking van een nieuw terug te betalen voorschot van 5 miljoen euro.
162. Zoals Advocaat-generaal Poiares Maduro verklaart, mag het criterium van de particuliere schuldeiser niet worden verward met dat […] van de particuliere investeerder. Waar een investeerder tracht winst te maken door zich bij de betrokken ondernemingen aan te bieden, tracht een schuldeiser van een debiteur in financiële moeilijkheden de terugbetaling te verkrijgen van aan hem verschuldigde bedragen. […] In dat geval is het doorslaggevende criterium niet of er een economisch voordeel is, maar of dit voordeel neerkomt op een behandeling die gunstiger is dan die welke onder soortgelijke omstandigheden door een particuliere schuldeiser zou worden verleend aan een onderneming die bij hem schulden heeft. [75]
163. Hieronder moet daarom worden nagegaan, eerst, of België ten aanzien van de verlening van uitstel van betaling heeft gehandeld als een bedachtzaam schuldeiser in een markteconomie, en vervolgens of België wat het verlenen van de kredietfaciliteit en het terugvorderbare voorschot betreft heeft gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan.
a) Heeft de NMBS door verlening van uitstel van betaling gehandeld zoals een bedachtzaam schuldeiser in een markteconomie zou hebben gedaan?
164. Volgens het Gerecht moet het gedrag van de staat worden vergeleken met dat van "een particuliere schuldeiser, die betaling tracht te verkrijgen van de bedragen die hem verschuldigd zijn door een schuldenaar in financiële moeilijkheden". [76] In dit geval moest schuldeiser NMBS dus beslissen of een bedachtzaam schuldeiser IFB geen uitstel van betaling zou hebben verleend en er de voorkeur aan zou hebben gegeven het bedrijf failliet te laten gaan.
165. De kaderovereenkomst is op 7 april 2003 ondertekend, maar het uitstel van betaling dat staatssteun zou kunnen zijn werd al in 2001 verleend. De analyse moet worden gemaakt uit het oogpunt van de feiten waarvan de NMBS destijds op de hoogte was [77].
166. Voor 2002 had IFB exploitatieverliezen geleden ten belope van 47,4 miljoen euro, waarvan 34 miljoen specifieke afschrijvingen waren die reeds bij de exploitatiekosten waren geconstateerd, en uitzonderlijke verliezen van 59,369 miljoen euro. De uitzonderlijke verliezen waren met name het gevolg van de waardevermindering in een aantal, hoofdzakelijk Franse, dochterondernemingen. Ten gevolge van deze verliezen had IFB aan het eind van boekjaar 2002 een negatief eigen vermogen van 84,07 miljoen euro.
167. In geval van faillissement zou de NMBS, die 89,03 % van het aandelenkapitaal van IFB in handen had, eventueel pas tot de resultaten van de liquidatie toegang hebben gehad nadat de schuldeisers waren voldaan. Bovendien hadden haar vorderingen die uit niet-betaalde facturen voortvloeiden waarschijnlijk slechts ten dele kunnen worden voldaan.
168. Dit was overigens de reden waarom de NMBS in haar jaarrekening van 2002 de waarde van deze aandelen en schuldvorderingen op nul had gesteld, [78] omdat, gelet op de financiële situatie van deze groep [d.i. IFB] en in afwachting van de voltooiing van het herstructureringsplan van deze groep binnen de vrachtsector van de NMBS, de commerciële schuldvorderingen en de lopende bestellingen die de NMBS heeft als twijfelachtig [moeten worden] geboekt. [79]
169. De NMBS was op dat ogenblik verreweg de grootste schuldeiser van IFB: volgens de jaarrekening 2003 van IFB had deze onderneming bij kredietinstellingen schulden ten belope van 12 miljoen euro, en schulden bij haar leveranciers, dus voornamelijk bij de NMBS, ten belope van 108 miljoen euro.
170. Bij een faillissement had de NMBS tevens 50 werknemers weer in de onderneming moeten opnemen die bij IFB waren gedetacheerd. Aangezien de NMBS het aantal werknemers juist tracht te verminderen, zou dat een extra nadeel voor de NMBS hebben opgeleverd.
171. Kortom: het faillissement van IFB zou voor de NMBS tot extra kosten hebben geleid, zonder dat de onderneming de zekerheid had dat de uitstaande schulden zouden worden vereffend.
172. Niettemin is het de vraag of de NMBS met het alternatief, namelijk het verlenen van uitstel van betaling, gecombineerd met de betaling van de vertragingsrente tegen de wettelijke rentevoet of tegen de marktrentevoet (naar gelang van de schulden, zie onderstaande beschrijving), de toezegging dat geen beroep zou worden gedaan op de verjaring van de schuldvorderingen en nieuwe investeringen, redelijkerwijs kon verwachten dat IFB voldoende winstgevend zou zijn om haar nieuwe investeringen te compenseren op een voor een particuliere investeerder in een markteconomie aanvaardbaar niveau en om de vooruitzichten op vereffening van de eerdere vorderingen op middellange of lange termijn te verbeteren.
173. In april 2003, op het tijdstip waarop de kaderovereenkomst werd afgesloten, had IFB een begin gemaakt met de herstructurering, die enerzijds een diepgaande herstructurering van de operaties van IFB zelf inhield en anderzijds een afsplitsingsstrategie om de exploitatieverliezen van de Franse dochterondernemingen op te vangen, zoals in deel 2.3.2 is beschreven.
174. Wat de kansen op hernieuwde rentabiliteit van IFB betreft, moet worden geconstateerd dat de financiële moeilijkheden met name het gevolg waren van de expansiestrategie in Frankrijk en slechts in mindere mate te wijten waren aan de structurele problemen van IFB Logistics en IFB Terminals.
175. Niettemin is in de kaderovereenkomst bepaald dat het uitstel van betaling gepaard zou gaan met een kredietfaciliteit van 15 miljoen en een terugvorderbaar voorschot van 5 miljoen euro. Daarom moest de NMBS, om redelijkerwijs te kunnen verwachten dat haar vorderingen zouden worden betaald, vers kapitaal investeren. Derhalve had een particuliere investeerder slechts uitstel van betaling verleend indien zijn aanvullende investering van 20 miljoen euro aan vers kapitaal een investering met een aanvaardbaar rendement was.
176. Het uitstel van betaling moet dan ook tezamen worden onderzocht met de door de NMBS in de kaderovereenkomst genomen investeringsbesluiten, aangezien de maatregelen, in de zin van de jurisprudentie in de zaak-BP Chemicals [80], een geheel vormen.
b) Heeft de NMBS door toekenning van een kredietfaciliteit en van een terugvorderbaar voorschot gehandeld zoals een bedachtzame investeerder in een markteconomie zou hebben gedaan?
177. Wat de toekenning van de kredietfaciliteit van 15 miljoen euro en de toekenning van het terugvorderbare voorschot van 5 miljoen euro betreft, had de NMBS, aangezien zij niet als investeerder optrad en dus geen schuldeiser van IFB was, de vrije keus om dit geld in IFB dan wel elders te investeren, en was zij dus een investeerder.
178. Derhalve moet worden nagegaan of de NMBS heeft gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan. Volgens de jurisprudentie van het Hof dient te worden beoordeeld of in soortgelijke omstandigheden een particulier investeerder die qua omvang vergelijkbaar is met de NMBS, ertoe zou kunnen worden gebracht een zo belangrijke kapitaalinbreng te doen. [81]
179. Het Hof heeft verduidelijkt dat een particulier investeerder, waarmee de deelneming van een publiek investeerder die doelstellingen van economisch beleid nastreeft, moet worden vergeleken, zich weliswaar niet noodzakelijkerwijs zal gedragen als een gewone investeerder die zijn kapitaal belegt om daaruit op min of meer korte termijn een rendement te halen, doch dat hij zich ten minste zal moeten gedragen als een particuliere holding of een particuliere groep ondernemingen met een algemene of sectoriële structuurpolitiek, die wordt geleid door het uitzicht op rendement op langere termijn [82]. Het Gerecht heeft de door de Commissie toe te passen beoordelingsmethode nauwkeuriger omschreven. Het heeft verduidelijkt dat de Commissie verplicht is "alle relevante elementen van de litigieuze transactie en haar context volledig te onderzoeken", teneinde te weten of de staat heeft gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan. [83]
180. In dit geval moet dus de rentabiliteit van het optreden van de NMBS worden vastgesteld, wat veronderstelt dat wordt nagegaan of de investering in IFB een normale winstmarge zou opleveren.
181. De NMBS heeft in april 2003, via reddingsmaatregelen, besloten 20 miljoen euro vrij te maken voor IFB in de vorm van een lening (kredietfaciliteit van 15 miljoen euro en terugvorderbaar voorschot van 5 miljoen euro).
182. De kaderovereenkomst, waarin reddingsmaatregelen waren vastgelegd, is op 7 april 2003 gesloten. De investering van 20 miljoen euro die op dat ogenblik bij wijze van reddingsmaatregel werd gedaan, moet worden geanalyseerd uit het oogpunt van de feiten waarvan de NMBS destijds op de hoogte was [84].
183. Bij het bepalen of de rentevoet voor een lening is afgestemd op de marktomstandigheden maakt de Commissie gewoonlijk een vergelijking met de referentierente die is vastgesteld voor de desbetreffende lidstaat op de desbetreffende datum [85]. Aangezien de leningen in kwestie tegen de marktrente worden vergoed, en ten dele zelfs tegen een hogere rentevoet dan de marktrente, lijkt deze op het eerste gezicht geen steunelement te bevatten. Niettemin moet worden geconstateerd dat IFB op het tijdstip waarop de leningen werden toegekend een onderneming met ernstige financiële moeilijkheden was. Het lijkt onwaarschijnlijk dat het bedrijf op de kapitaalmarkt een lening had kunnen krijgen tegen vergelijkbare voorwaarden als de door de NMBS geboden voorwaarden. Een bank had dus zeer waarschijnlijk een hogere rente verlangd dan de door de NMBS gevraagde rente of had zelfs geweigerd IFB een lening te geven. Het besluit van de NMBS om voor de bestaande schuldvorderingen uitstel van betaling te verlenen is trouwens een aanwijzing voor de moeilijkheden die IFB heeft moeten ondervinden om zich elders te herfinancieren.
184. De Belgische autoriteiten zijn van mening dat het feit dat IFB in juli 2003, dus na de sluiting van de kaderovereenkomst, een lening van 2 miljoen euro van de ING-bank heeft gekregen, aantoont dat particuliere banken geen vergoeding vroegen die hoger was dan de marktrentevoet.
185. Dit argument is om twee redenen niet overtuigend. Ten eerste is het bedrag van 2 miljoen euro zeer laag in vergelijking met de verbintenissen van de NMBS, die voorzagen in investeringen ten belope van 20 miljoen euro plus de mogelijkheid om de schuld van 63 miljoen euro om te zetten in kapitaal. Voorts heeft ING deze lening pas toegestaan nadat de NMBS, door de kaderovereenkomst te ondertekenen, zich ertoe verbonden had het voortbestaan van IFB te garanderen.
186. Geconstateerd moet daarom worden dat de NMBS door de toekenning van leningen tegen een lagere rente dan die welke voor de financiële situatie van IFB adequaat zou zijn geweest, niet heeft gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan.
187. De Belgische regering van haar kant is van mening dat de NMBS heeft gehandeld zoals iedere moedermaatschappij, waarvan een dochteronderneming in moeilijkheden verkeert, zou hebben gedaan, zonder dit standpunt nader toe te lichten. De Commissie merkt op dit punt op dat België dit standpunt niet heeft onderbouwd en met name niet heeft aangetoond dat de nieuwe investering noodzakelijk was om te kunnen verwachten er een hoger bedrag dan al haar bestaande en nieuwe vorderingen aan over te houden.
c) Conclusie ten aanzien van de reddingsmaatregelen
188. Bij wijze van conclusie is de Commissie in dit stadium van oordeel dat de NMBS, wat de toekenning van een kredietfaciliteit van 15 miljoen euro en de toekenning van een terugvorderbaar voorschot van 5 miljoen euro betreft, niet heeft gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan. Aangezien de verlening van uitstel van betaling voor een particuliere schuldeiser slechts redelijk was indien de investering dit eveneens was, volgt hieruit dat de NMBS, wat de verlening van uitstel van betaling aan IFB betreft, evenmin heeft gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan.
3.1.2.3. Herstructureringsmaatregelen
189. De herstructureringsmaatregelen zijn in deel 2 hierboven beschreven. Ter herinnering zij erop gewezen dat het gaat om:
- de omzetting van de schulden ten bedrage van 63 miljoen euro waarvoor uitstel van betaling is toegestaan, in maatschappelijk kapitaal;
- de omzetting van de kredietfaciliteit van 15 miljoen euro in maatschappelijk kapitaal;
- de omzetting van de gekapitaliseerde rente in verband met het uitstel van betaling ten bedrage van 11 miljoen euro in maatschappelijk kapitaal;
- de omzetting van de gekapitaliseerde rente op het terugvorderbare voorschot van 2,5 miljoen euro in maatschappelijk kapitaal;
- de injectie van 5 miljoen euro door de inbreng in natura van de participatie van de NMBS in TRW.
190. De kapitaalverhoging zal dus in totaal 96,5 miljoen euro bedragen. Daar IFB op dit ogenblik een negatief eigen vermogen van 72,6 miljoen euro heeft, zal het bedrijf door de kapitaalverhoging beschikken over 23,8 miljoen euro eigen kapitaal.
191. Bij deze maatregelen moet een onderscheid worden gemaakt tussen de maatregelen die de NMBS als schuldeiser van IFB heeft genomen, namelijk de omzetting van de bestaande schulden van 63 miljoen euro en van de bijbehorende rente van 11 miljoen euro in maatschappelijk kapitaal, en de maatregelen die de NMBS als investeerder in IFB heeft genomen, namelijk de omzetting van de kredietfaciliteit van 15 miljoen euro en van de bijbehorende rente van 2,5 miljoen euro in maatschappelijk kapitaal en de injectie van vers kapitaal van 5 miljoen euro.
192. Wat betreft de omzetting van de kredietfaciliteit van 15 miljoen euro in maatschappelijk kapitaal, zou kunnen worden aangevoerd dat de NMBS op het moment van de omzetting geen investeerder meer was, maar schuldeiser. Daarmee wordt echter het feit genegeerd dat in de kaderovereenkomst was bepaald dat de kredietfaciliteit eventueel in maatschappelijk kapitaal zou worden omgezet (zie de beschrijving in deel 2) en dat de kredietfaciliteit slechts een tijdelijke maatregel was. Bijgevolg moet worden aangenomen dat de omzetting van de kredietfaciliteit in maatschappelijk kapitaal te vergelijken is met een investering.
a) Heeft de NMBS gehandeld zoals een bedachtzaam schuldeiser in een markteconomie zou hebben gedaan, door haar schuldvorderingen van 63 miljoen euro en de bijbehorende rente van 11 miljoen euro om te zetten in maatschappelijk kapitaal?
193. Door haar schuldvorderingen van 63 miljoen euro en de bijbehorende rente van 11 miljoen euro om te zetten in maatschappelijk kapitaal, ziet de NMBS af van de terugbetaling van deze schulden. Daartegenover staat dat zij recht zal hebben op de dividenden die IFB aan zijn eigenaars zal uitkeren, en dat zij aandelen verwerft.
194. Zoals hierboven is aangetoond, dient in dit stadium te worden aangenomen dat een bedachtzaam particulier schuldeiser het door de NMBS toegekende uitstel van betaling niet zou hebben toegekend, maar het faillissement van IFB zou hebben aangevraagd en zou hebben getracht de betaling van de schuldvorderingen in het kader van de collectieve procedure te verkrijgen.
195. Bijgevolg zou een bedachtzaam particulier schuldeiser zijn vorderingen ook niet hebben omgezet in maatschappelijk kapitaal van een onderneming die slechts kon overleven indien hij tegelijkertijd ook vers kapitaal zou verstrekken. De NMBS heeft dus, door haar vorderingen in maatschappelijk kapitaal om te zetten, niet gehandeld zoals een particuliere schuldeiser in een markteconomie zou hebben gedaan.
b) Heeft de NMBS gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan, door de kredietfaciliteit van 15 miljoen euro en de bijbehorende rente van 2,5 miljoen euro om te zetten in maatschappelijk kapitaal en door 5 miljoen euro vers kapitaal te verstrekken?
196. Er moet worden nagegaan of de NMBS heeft gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan wat betreft de omzetting van de kredietfaciliteit van 15 miljoen euro en van de bijbehorende rente van 2,5 miljoen euro in maatschappelijk kapitaal, alsmede de kapitaalverhoging van IFB ten bedrage van 5 miljoen euro.
197. Volgens de jurisprudentie van het Hof dient te worden beoordeeld of in soortgelijke omstandigheden een particuliere investeerder die qua omvang vergelijkbaar is met de NMBS, ertoe zou kunnen worden gebracht een zo belangrijke kapitaalinbreng te doen [86].
198. Het Hof heeft verduidelijkt dat een particuliere investeerder, waarmee de deelneming van een publieke investeerder die doelstellingen van economisch beleid nastreeft, moet worden vergeleken, zich weliswaar niet noodzakelijkerwijs zal gedragen als een gewone investeerder die zijn kapitaal belegt om daaruit op min of meer korte termijn een rendement te halen, doch dat hij zich ten minste zal moeten gedragen als een particuliere holding of een particuliere groep ondernemingen met een algemene of sectoriële structuurpolitiek, die wordt geleid door het uitzicht op rendement op langere termijn [87]. Het Gerecht heeft de door de Commissie toe te passen beoordelingsmethode nauwkeuriger omschreven. Het heeft verduidelijkt dat de Commissie verplicht is "een volledig onderzoek uit te voeren van alle relevante elementen van de litigieuze transactie en haar context", teneinde te weten of de staat heeft gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan. [88]
199. In dit geval moet dus de rentabiliteit van het optreden van de NMBS worden vastgesteld, wat veronderstelt dat wordt aangetoond dat de investering in IFB een normale winstmarge zal opleveren.
200. Door haar beslissing om de kredietfaciliteit van 15 miljoen euro en de bijbehorende rente van 2,5 miljoen euro, die een tijdelijke reddingsmaatregel was, in een kapitaalverhoging om te zetten, zal de NMBS deze investering een duurzaam karakter geven.
201. Met haar beslissing aan deze kapitaalverhoging het bedrag van 5 miljoen euro toe te voegen, heeft zij een aanvullende investering van 5 miljoen verricht.
202. Over de omzetting van de kredietfaciliteit van 15 miljoen euro en van de bijbehorende rente van 2,5 miljoen euro in maatschappelijk kapitaal en het beginsel van de aanvullende kapitaalverhoging van 5 miljoen euro is in het voorjaar 2005 een beslissing genomen; bij het onderzoek ervan moet dus worden uitgegaan van de feiten waarvan de NMBS op dat ogenblik kennis had. [89]
203. Deze twee maatregelen moeten worden vergeleken met de beslissing van een particuliere investeerder om deel te nemen in een kapitaalverhoging van IFB.
204. De Commissie neemt in de eerste plaats nota van de afwezigheid van een particuliere investeerder die, met de NMBS, zou hebben deelgenomen in de kapitaalverhoging van IFB.
205. De Belgische regering is van oordeel dat de NMBS heeft gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan. Om dat aan te tonen, geeft zij het volgende voorbeeld: indien de NMBS op 1 januari 2004 nieuw kapitaal aan IFB had verstrekt door omzetting van de schulden van IFB ten aanzien van de NMBS (ca. 79 miljoen euro op dat ogenblik) en een aanvullende inbreng van ca. 21 miljoen euro, had IFB aan het begin van het boekjaar over ongeveer 16 miljoen euro eigen vermogen beschikt. Bovendien zou het bedrijf een bedrijfswinst van 5,74 miljoen euro (rendement van 36 % op eigen vermogen) en een lopende winst vóór belasting van meer dan 7,18 miljoen euro (45 % op eigen kapitaal) hebben gemaakt. De operationele winstmarge op de omzet zou dan ca. 7 % hebben bedragen in 2004. Aangezien het resultaat over 2004 sterk is beïnvloed door het gebruik en de overname van bepaalde in 2001 en 2002 gemaakte voorzieningen voor de verwachte verliezen van de Franse dochtermaatschappijen, stelt de Belgische regering voor deze buitengewone gebeurtenissen te neutraliseren, waardoor voor 2004 een operationele winstmarge op de omzet van 2,9 % overblijft. De Belgische regering heeft geen raming van de winst van IFB voor de volgende jaren verstrekt.
206. De Commissie is van oordeel dat de ontwikkeling van IFB sinds 2003 zeker aantoont dat het bedrijf economisch levensvatbaar is. De toets van de particuliere investeerder in een markteconomie heeft echter niet alleen betrekking op de economische levensvatbaarheid van een onderneming, maar ook op haar rentabiliteit. Volgens het Hof "moet worden beoordeeld of een particuliere aandeelhouder in gelijkaardige omstandigheden, op grond van de te verwachten rentabiliteit en afgezien van elke overweging van sociale aard of van regionaal of sectorieel beleid, een dergelijke kapitaalinbreng zou hebben gedaan" [90]. Deze mogelijkheid van rentabiliteit moet ten minste gelijk zijn aan die van "een particuliere holding of een particuliere groep ondernemingen met een algemene of sectoriële structuurpolitiek, die wordt geleid door het uitzicht op rendement op langere termijn". [91]
207. Bij de beoordeling van de normale vergoeding wordt met name rekening gehouden met de gemiddelde rentabiliteit van de concurrenten. In dit verband heeft de Belgische regering de Commissie meegedeeld dat de omzet en de rentabiliteit van de concurrenten van IFB als volgt waren (in miljoenen euro's):
| Omzet 2003 | Winst 2003 | Winst 2003 in % | Omzet 2004 | Winst 2004 | Winst 2004 in % |
CEMAT | 164,1 | 1,4 | 0,9 | 176,6 | 3,9 | 2,2 |
CNC | 193,5 | - 17,0 | - 8,8 | 164,4 | - 20,6 | - 12,5 |
HUPAC | 195,2 | 5,7 | 2,9 | 225,6 | 6,0 | 2,7 |
ICF | 276,5 | 0,5 | 0,2 | 261,1 | - 3,7 | - 1,4 |
Kombiverkehr | 289,2 | 0,8 | 0,3 | n.v.t. | n.v.t. | n.v.t. |
Novatrans | 109,0 | - 7,1 | - 6,5 | 102,5 | - 5,5 | - 5,4 |
208. Hierbij zij opgemerkt dat in deze tabel niet het rendement van de grote concurrenten Hesse-Noordnatie, Danzas, Ziegler, en Schenker wordt weergegeven en dat de meeste van de door de Belgische regering vermelde ondernemingen in 2004 verlies hebben geleden.
209. De door de Belgische regering verstrekte cijfers kunnen dus niet worden gebruikt om te beoordelen of het rendement van IFB een normaal rendement is. Bij gebrek aan een adequaat vergelijkingscijfer constateert de Commissie dat een rendement van 2,9 % een zeer laag rendement is, want het komt min of meer overeen met het rendement van overheidsobligaties. Aan een investering in IFB is echter een duidelijk hoger risico verbonden dan aan overheidsobligaties.
210. Bijgevolg is de Commissie van oordeel dat het rendement van een investering in IFB niet voldoende zou zijn om een bedachtzaam investeerder in een markteconomie ertoe over te halen een dergelijke investering te doen. Een bedachtzaam investeerder zou dus niet de investeringen hebben gedaan die de NMBS in IFB heeft gedaan.
c) Conclusie wat de herstructureringsmaatregelen betreft
211. De Commissie is bijgevolg in dit stadium van oordeel dat de NMBS niet heeft gehandeld zoals een particuliere schuldeiser in een markteconomie zou hebben gedaan, door de schulden van 63 miljoen euro en de bijbehorende rente van 11 miljoen om te zetten in maatschappelijk kapitaal. Zij is van oordeel dat de NMBS evenmin heeft gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan wat betreft de omzetting van de kredietfaciliteit van 15 miljoen euro en de bijbehorende rente van 2,5 miljoen euro in maatschappelijk kapitaal en wat betreft de injectie van 5 miljoen euro in IFB.
3.1.3 Vervalsing van de mededinging en ongunstige beïnvloeding van het handelsverkeer tussen de lidstaten
212. De Commissie moet een analyse maken van de situatie op de desbetreffende markt en van het marktaandeel van de begunstigde ondernemingen op deze markt, alsmede van het effect dat de financiële steun zal hebben op de concurrentiesituatie [92].
213. In dit geval is de financiële steun toegekend aan een onderneming die actief is op voor mededinging opengestelde markten en die zich met andere marktdeelnemers uit diverse lidstaten in een concurrentiesituatie bevindt, zoals hierboven in het deel "beschrijving" is aangetoond. De financiële steun vervalst dus de mededinging of dreigt die te vervalsen en beïnvloedt ongunstig het handelsverkeer tussen de lidstaten of dreigt dit ongunstig te beïnvloeden.
3.1.4. Conclusie: aanwezigheid van staatssteun
214. Bij wijze van conclusie is de Commissie in dit stadium van oordeel dat de NMBS niet heeft gehandeld zoals een bedachtzaam schuldeiser in een markteconomie zou hebben gedaan wat betreft het uitstel van betaling en de omzetting van de op 31 januari 2003 vervallen en niet betaalde schuldvorderingen ten bedrage van 63 miljoen euro, en dat zij niet heeft gehandeld zoals een bedachtzaam investeerder in een markteconomie zou hebben gedaan wat betreft de toekenning van een kredietfaciliteit van 15 miljoen euro, de toekenning van een terugvorderbaar voorschot van 5 miljoen euro, de omzetting van de kredietfaciliteit van 15 miljoen euro in maatschappelijk kapitaal, alsmede wat betreft de injectie van vers kapitaal ten bedrage van 5 miljoen euro.
3.2. Verenigbaarheid van de steun
215. In artikel 87, lid 3, onder c), van het EG-Verdrag is het volgende bepaald: "met de gemeenschappelijke markt zijn verenigbaar: steunmaatregelen om de ontwikkeling van bepaalde vormen van economische bedrijvigheid of van bepaalde regionale economieën te vergemakkelijken, mits de voorwaarden waaronder het handelsverkeer plaatsvindt daardoor niet zodanig worden veranderd dat het gemeenschappelijk belang wordt geschaad".
216. De door België via de NMBS toegekende steun zou met de gemeenschappelijke markt verenigbaar kunnen zijn op grond van artikel 87, lid 3, onder c), zoals door de Commissie geïnterpreteerd in haar Communautaire richtsnoeren voor reddings- en herstructureringssteun aan ondernemingen in moeilijkheden (hierna: de richtsnoeren) [93].
217. Om reddings- en herstructureringssteun te kunnen ontvangen, moet een onderneming om te beginnen in aanmerking komen voor de toepassing van de richtsnoeren. Om daarvoor in aanmerking te komen, mag de onderneming geen nieuw opgerichte onderneming zijn en moet het een onderneming in moeilijkheden zijn.
218. Geen nieuw opgerichte onderneming. In punt 12 van de richtsnoeren van 2004 wordt in dit verband het volgende bepaald (waarbij de richtsnoeren van 1999, punt 7, worden overgenomen en verduidelijkt):
Voor de toepassing van de onderhavige richtsnoeren komt een pas opgerichte onderneming niet voor reddings- of herstructureringssteun in aanmerking, zelfs niet wanneer haar aanvankelijke financiële positie onzeker is. Dit geldt bijvoorbeeld voor ondernemingen die uit de liquidatie van een bestaande onderneming ontstaan of die de activa van een dergelijke onderneming overnemen. Een onderneming wordt in beginsel als een nieuw opgerichte onderneming beschouwd gedurende de eerste drie jaar na de aanvang van activiteiten in de betrokken sector.
219. Om te beginnen rijst dus de vraag of IFB een nieuw opgerichte onderneming is. Zoals hierboven in deel 2 is beschreven, is IFB op 1 april 1998 opgericht door de fusie van drie andere maatschappijen, die respectievelijk in 1906, 1923 en 1967 waren opgericht.
220. Zoals hierboven in punt 3.1.2.1 is uitgelegd, was het eerste voordeel dat door de NMBS aan IFB werd toegekend, de stilzwijgende toekenning, ten vroegste vanaf 2001, van een uitstel van betaling voor de door de NMBS geleverde, maar door IFB niet betaalde diensten.
221. De onderneming IFB is op 1 april 1998 opgericht door de fusie van drie bestaande maatschappijen. In dit stadium is het niet duidelijk of de onderneming de rechtspersoonlijkheid van een van deze drie maatschappijen voortzet. Indien dit het geval zou zijn, zou IFB in 2001 duidelijk een onderneming van meer dan drie jaar oud zijn.
222. Indien IFB de rechtspersoonlijkheid van een van deze maatschappijen niet zou voortzetten, maar een op 1 april 1998 nieuw opgerichte onderneming zou zijn, zou zij op 1 april 2001 drie jaar oud zijn. In deze veronderstelling zou zij pas vanaf 1 april 2001 in aanmerking komen voor herstructureringssteun.
223. De Commissie uit dus twijfels over de vraag of IFB een onderneming is die in aanmerking komt voor herstructureringssteun, en verzoekt de Belgische autoriteiten haar alle nuttige informatie te verstrekken zodat zij kan nagaan of IFB in het licht van deze overwegingen een onderneming is die in aanmerking komt voor herstructureringssteun.
224. Onderneming in moeilijkheden Er is geen communautaire definitie van een onderneming in moeilijkheden. In de richtsnoeren wordt in punt 5 (versie van 1999), respectievelijk punt 10 (versie van 2004) aangenomen dat een vennootschap met beperkte aansprakelijkheid, zoals de maatschappij IFB, die een vennootschap op aandelen is, in elk geval als onderneming in moeilijkheden wordt beschouwd wanneer meer dan de helft van het maatschappelijk kapitaal verdwenen is en meer dan een kwart van dit kapitaal verloren is gegaan gedurende de afgelopen twaalf maanden. De jaarrekening over 2002 geeft een maatschappelijk kapitaal van 48 miljoen euro te zien en lopende verliezen vóór belasting van 50 miljoen euro. Bijgevolg was het maatschappelijk kapitaal verdwenen toen de NMBS in april 2003 besloot reddingssteun toe te kennen. Aangezien op dat ogenblik meer dan de helft van het maatschappelijk kapitaal verdwenen was, waarvan meer dan een kwart in de laatste twaalf maanden, is IFB een onderneming in moeilijkheden in de zin van de richtsnoeren.
225. De richtsnoeren zijn dus van toepassing. Er moet worden onderzocht of zij bij de toekenning van steun door de NMBS aan IFB zijn nageleefd. In dit verband moet in de eerste plaats worden onderzocht of het bij ten minste een deel van de steun ging om met de richtsnoeren verenigbare reddingssteun.
3.2.1. Verenigbaarheid als reddingssteun
226. Alleen maatregelen die bestaan in kassteun, zouden als reddingssteun verenigbaar kunnen zijn. In het onderhavige geval bestaat de kassteun in de toekenning van een stilzwijgend uitstel van betaling, ten vroegste in 2001, ten laatste op 19 september 2002, dat op 7 april 2003 uitdrukkelijk uitstel van betaling is geworden, de kredietfaciliteit en het terugvorderbare voorschot.
227. In de eerste plaats rijst de vraag welke versie van de richtsnoeren van toepassing is. De recentste versie van deze richtsnoeren is op 10 oktober 2004 in werking getreden. Daarin wordt in punt 7 "Datum van toepassing en duur" bepaald:
102. De Commissie zal deze richtsnoeren toepassen met ingang van 10 oktober 2004 tot 9 oktober 2009.
103. Aanmeldingen die door de Commissie vóór 10 oktober 2004 zijn geregistreerd, zullen worden getoetst aan de criteria die gelden op het tijdstip van de aanmelding.
104. De Commissie zal onderzoeken of reddings- of herstructureringssteun die zonder haar toestemming — en dus in strijd met artikel 88, lid 3, van het Verdrag — is toegekend, verenigbaar is met de gemeenschappelijke markt op basis van de onderhavige richtsnoeren wanneer die steun geheel of gedeeltelijk na de bekendmaking van deze richtsnoeren in het Publicatieblad van de Europese Unie is toegekend. In alle overige gevallen zal zij het onderzoek verrichten op basis van de op het tijdstip van de toekenning van de steun geldende richtsnoeren.
228. De kassteun is ten vroegste in 2001 of in de loop van 2002 en in zijn geheel op 7 april 2003 toegekend zonder voorafgaande kennisgeving aan de Commissie en dus in strijd met artikel 88, lid 3, van het EG-Verdrag. De vraag of hij als reddingssteun verenigbaar is, waarbij de andere, als herstructureringssteun aan te merken maatregelen buiten beschouwing worden gelaten, zal dus worden beoordeeld op basis van de richtsnoeren van 1999.
229. In punt 23 van de richtsnoeren van 1999, die van toepassing zijn op de reddingssteun die de NMBS mogelijkerwijs in 2001, zeker in 2002 en 2003, aan IFB heeft toegekend, worden de vijf voorwaarden bepaald waaraan reddingssteun moet voldoen om met de gemeenschappelijke markt verenigbaar te zijn. Deze vijf voorwaarden zijn:
a) bestaan in kassteun in de vorm van leninggaranties of leningen. In beide gevallen moet de rente op zijn minst vergelijkbaar zijn met de rentepercentages die gelden voor leningen aan gezonde ondernemingen en met name aan de referentiepercentages die door de Commissie zijn vastgesteld;
b) gekoppeld zijn aan leningen die over een periode van ten hoogste twaalf maanden na de laatste storting aan de onderneming moeten worden terugbetaald; eventueel kan de terugbetaling van de lening die in het kader van de reddingssteun is verstrekt, worden gedekt door herstructureringssteun die in een later stadium door de Commissie is goedgekeurd;
c) worden gerechtvaardigd door dringende sociale omstandigheden en geen ernstig "spill-over"-effect naar andere lidstaten hebben;
d) bij de aanmelding ervan gepaard gaan met een toezegging van de lidstaat, de Commissie binnen zes maanden na de goedkeuring van de reddingssteun, ofwel een herstructureringsplan, ofwel een liquidatieplan voor te leggen, dan wel aan te tonen dat de lening volledig is afgelost en/of dat de garantie is ingetrokken;
e) zich wat het bedrag betreft beperken tot hetgeen noodzakelijk is voor de exploitatie van de onderneming gedurende de periode waarvoor de steun is goedgekeurd (bijvoorbeeld dekking van de loonkosten, lopende leveringen).
3.2.1.1. Steun die bestaat in kassteun
230. Er zij aan herinnerd dat de reddingsmaatregelen bestaan in een uitstel van betaling voor schuldvorderingen voor een totaal bedrag van 63 miljoen euro, een terugvorderbaar voorschot van 5 miljoen euro, dat is toegekend, maar niet door IFB is gebruikt, en een kredietfaciliteit van 15 miljoen euro.
231. Bijgevolg bestaat de steun in kassteun, die bestaat uit een uitstel van betaling, een terugvorderbaar voorschot en een kredietfaciliteit.
3.2.1.2. Steun die gekoppeld is aan leningen die over een periode van ten hoogste twaalf maanden na de laatste storting aan de onderneming moeten worden terugbetaald
232. De in de kaderovereenkomst vastgestelde terugbetalingsperiode is twaalf maanden. De Belgische regering heeft de Commissie echter meegedeeld dat deze periode stilzwijgend is verlengd tot het tijdstip waarop de kapitaalverhoging plaatsvindt.
233. Bovendien is het voordeel dat voortvloeit uit het uitstel van betaling, reeds ten vroegste in de loop van 2001, ten laatste op 19 december 2002, toegekend. De Commissie is bijgevolg van oordeel dat aan dit criterium niet wordt voldaan en dat de kassteun niet als reddingssteun kan worden goedgekeurd.
3.2.1.3. Conclusie
234. Bij wijze van conclusie is de Commissie in dit stadium van oordeel dat de kassteun die de NMBS aan IFB heeft toegekend, als reddingssteun niet met de gemeenschappelijke markt verenigbaar is op grond van artikel 87, lid 3, onder c), van het Verdrag. Hij zou als herstructureringssteun echter wel met de gemeenschappelijke markt verenigbaar kunnen zijn.
3.2.2. Verenigbaarheid van de herstructureringssteun
235. Opnieuw rijst de vraag welke versie van de richtsnoeren van toepassing is. Er zij aan herinnerd dat de recentste versie van deze richtsnoeren op 10 oktober 2004 in werking is getreden. Daarin wordt in punt 7 "Datum van toepassing en duur" bepaald:
102. De Commissie zal deze richtsnoeren toepassen met ingang van 10 oktober 2004 tot 9 oktober 2009.
103. Aanmeldingen die door de Commissie vóór 10 oktober 2004 zijn geregistreerd, zullen worden getoetst aan de criteria die gelden op het tijdstip van de aanmelding.
104. De Commissie zal onderzoeken of reddings- of herstructureringssteun die zonder haar toestemming — en dus in strijd met artikel 88, lid 3, van het Verdrag — is toegekend, verenigbaar is met de gemeenschappelijke markt op basis van de onderhavige richtsnoeren wanneer die steun geheel of gedeeltelijk na de bekendmaking van deze richtsnoeren in het Publicatieblad van de Europese Unie is toegekend. In alle overige gevallen zal zij het onderzoek verrichten op basis van de op het tijdstip van de toekenning van de steun geldende richtsnoeren.
236. De kassteun is gedeeltelijk ten vroegste in de loop van 2001, ten laatste op 19 september 2002, en in zijn geheel op 7 april 2003 toegekend zonder voorafgaande kennisgeving aan de Commissie en dus in strijd met artikel 88, lid 3, van het EG-Verdrag. De omzetting ervan in kapitaal was gepland sinds de sluiting van de kaderovereenkomst op 7 april 2003, maar heeft tot op heden niet plaatsgevonden.
237. Aangezien de NMBS de kassteun zonder voorafgaande goedkeuring van de Commissie heeft verleend, moet punt 104 van de richtsnoeren van 2004 worden toegepast om te bepalen welke richtsnoeren op dit geval van toepassing zijn. De kassteun is gedeeltelijk ten vroegste in de loop van 2001, ten laatste op 19 september 2002, en voor de rest op 7 april 2003 toegekend, dat wil zeggen vóór de publicatie van de richtsnoeren van 2004 in het Publicatieblad. Indien de steun beperkt zou blijven tot kassteun, zouden dus de richtsnoeren van 1999 moeten worden toegepast, want de toekenning van de steun zou vóór de publicatie van de richtsnoeren van 2004 hebben plaatsgevonden.
238. De omzetting van de vorderingen in kapitaal is echter een latere maatregel, waardoor de aard van de voordien aan IFB toegekende voordelen wordt gewijzigd. In dit verband wordt in de kaderovereenkomst melding gemaakt van het voornemen van de partijen om over te gaan tot deze omzetting, evenwel onder voorbehoud van met name de goedkeuring van het herstructureringsplan door beide raden van bestuur en door de Belgische staat, alsmede onder voorbehoud van goedkeuring door de aandeelhouders van IFB. In dit stadium is dus niet aangetoond dat de maatregel definitief is toegekend vóór de publicatie van de richtsnoeren van 2004, in die zin dat de bevoegde autoriteit zich er door een juridisch bindend document toe heeft verbonden de steun vóór die datum toe te kennen [94]. Indien dit niet het geval was, en aangezien de omzetting van de vorderingen in kapitaal niet vóór 10 oktober 2004 ter kennis is gebracht, zouden de richtsnoeren van 2004 van toepassing zijn.
239. De Belgische autoriteiten hebben de Commissie er per brief van 28 januari 2005 van in kennis gesteld dat de NMBS in 2005 of 2006 een nieuw voordeel van 5 miljoen euro zou toekennen in de vorm van een kapitaalverhoging door inbreng in natura. In dat geval zou na 10 oktober 2004 kennisgeving zijn gedaan van steun. Krachtens punt 103 van de richtsnoeren van 2004 zouden dan de richtsnoeren van 2004 op die nieuwe kennisgeving moeten worden toegepast.
240. De Commissie moet zich uitspreken over alle maatregelen waarvan haar kennisgeving is gedaan; zij baseert dus haar juridische beoordeling op de richtsnoeren van 2004. Zij vestigt echter de aandacht van de Belgische regering en van belanghebbende derden op het feit dat, indien de NMBS besluit geen nieuw voordeel aan IFB toe te kennen, en indien het bewijs zou worden geleverd dat de NMBS zich ertoe verbonden had haar vorderingen vóór de publicatie van de richtsnoeren van 2004 in kapitaal om te zetten, de Commissie de door de NMBS aan IFB toegekende steun in haar eindbesluit zou moeten onderzoeken op basis van de richtsnoeren van 1999. De hierna op basis van de tekst van 2004 geuite twijfels gelden, mutatis mutandis, ook voor de tekst van 1999.
241. In punt 3.2.2 van de richtsnoeren van 2004 worden de voorwaarden voor de goedkeuring van herstructureringssteun omschreven. De voorwaarden zijn als volgt:
- Het herstructureringsplan dient binnen een redelijk tijdsbestek de levensvatbaarheid op lange termijn van de onderneming te herstellen.
- Er moeten maatregelen worden genomen om de nadelige gevolgen voor de concurrenten zoveel mogelijk te beperken.
- De steun moet worden beperkt tot het strikt noodzakelijke minimum om de herstructurering mogelijk te maken.
- De Commissie moet in staat worden gesteld zich aan de hand van regelmatige en gedetailleerde verslagen ervan te vergewissen dat het herstructureringsplan naar behoren wordt uitgevoerd.
- Er mag slechts eenmaal herstructureringssteun worden toegekend.
3.2.2.1. Herstructureringsplan
242. Voor de toekenning van herstructureringssteun geldt als voorwaarde dat een herstructureringsplan ten uitvoer wordt gelegd dat binnen een redelijk tijdsbestek de levensvatbaarheid op lange termijn van de onderneming dient te herstellen op grond van realistische veronderstellingen betreffende de toekomstige bedrijfsomstandigheden.
243. In de punten 32 tot en met 34 van de richtsnoeren worden de minimumvoorwaarden voor de goedkeuring van een herstructureringsplan door de Commissie bepaald. Het herstructureringsplan moet met name de volgende elementen bevatten:
- een marktstudie;
- een beschrijving van de omstandigheden die tot de moeilijkheden van de onderneming hebben geleid, zodat kan worden beoordeeld of de in het plan voorgestelde maatregelen passend zijn om de levensvatbaarheid van de onderneming te herstellen;
- een beschrijving van de voorgenomen veranderingen die ervoor moeten zorgen dat de onderneming, wanneer de herstructurering voltooid is, in staat is alle kosten, met inbegrip van aflossingen en financiële lasten, te dekken, en op eigen kracht op de markt te concurreren.
244. De Belgische regering heeft in december 2003 een herstructureringsplan voor IFB voorgelegd en heeft dit plan naderhand gedetailleerd. Het bevat de genoemde elementen en wordt in detail beschreven in deel 2 van deze beschikking.
245. Dit plan bevat een analyse van de logistiekmarkt en van de overslagmarkt, alsmede van de positie van IFB op die markten. In het plan worden de oorzaken van de moeilijkheden van IFB beschreven. Ze vinden met name hun oorsprong in een slecht aangepakt expansiebeleid in Frankrijk en in het slechte beheer van de activiteiten "IFB Terminals" en "IFB Logistics".
246. Ten slotte worden in dit plan de voorgenomen veranderingen beschreven die ervoor moeten zorgen dat de onderneming, wanneer de herstructurering voltooid is, in staat is op eigen kracht al haar kosten te dekken. De voorgenomen veranderingen zijn met name de opheffing van de Franse dochterondernemingen, alsmede een herstructurering van de activiteiten "IFB Logistics" en "IFB Terminals". Deze herstructureringen impliceren met name concentratie op rentabele onderdelen van het aanbod, een nieuwe collectieve overeenkomst en een reorganisatie van de terminals.
247. De tenuitvoerlegging van dit herstructureringsplan is in 2005 met succes voltooid.
3.2.2.2. Economische levensvatbaarheid van de onderneming
248. Het herstructureringsplan bevat de door IFB geplande maatregelen om zijn economische levensvatbaarheid te herstellen. Zoals hierboven werd beschreven, heeft IFB in 2003 zijn financiële doelstellingen niet kunnen verwezenlijken. Vanaf het boekjaar 2004 heeft de onderneming echter de in het herstructureringsplan geformuleerde doelstellingen kunnen bereiken en heeft zij zelfs een hogere winst gerealiseerd dan werd beoogd. Deze goede ontwikkeling heeft zich in 2005 voortgezet.
249. IFB is erin geslaagd om het vervoerde vrachtvolume sinds de aanvang van het herstructureringsprogramma aanzienlijk te vergroten (zie de beschrijving hierboven in deel 2). Dat verklaart ook de groei van zijn omzet van 58 miljoen euro in 2003 tot 83 miljoen euro in 2004.
250. De onderneming IFB heeft dus haar economische levensvatbaarheid kunnen aantonen, zowel in haar herstructureringsplan, dat in 2003 is voorgelegd, als in de sindsdien geboekte resultaten.
3.2.2.3. Maatregelen om de nadelige gevolgen van de steun voor de concurrenten zoveel mogelijk te beperken
251. Er moeten compenserende maatregelen worden genomen om de nadelige gevolgen van de steun voor de concurrenten zoveel mogelijk te beperken. Anders zou de staatssteun als "in strijd met het gemeenschappelijk belang" en derhalve als onverenigbaar met de gemeenschappelijke markt moeten worden beschouwd.
252. De Belgische autoriteiten leggen uit dat IFB twee maatregelen heeft genomen om de nadelige gevolgen van de steun voor de concurrenten zoveel mogelijk te beperken:
- de stopzetting van zijn overslagactiviteiten in Frankrijk;
- de sluiting van de terminal van Bressoux in België en de verkoop van de participaties in de terminals in Brussel en Zeebrugge in België.
253. Als gevolg van deze twee maatregelen is de omzet van IFB gedaald van 62 miljoen euro in 2002 tot 58 miljoen euro in 2003. In 2004 echter lag de omzet van de onderneming met 83 miljoen euro reeds boven die van 2002.
254. De Commissie vestigt evenwel de aandacht van België op punt 40 van de richtsnoeren van 2004, waarin het volgende staat:
Afschrijvingen en sluiting van verliesgevende activiteiten die in ieder geval nodig zijn om de levensvatbaarheid te herstellen, worden bij de beoordeling van de compenserende maatregelen niet als inkrimping van capaciteit of aanwezigheid op de markt beschouwd.
255. Volgens de informatie die de Belgische regering aan de Commissie heeft verstrekt, lijken de terugtrekking uit de Franse markt en de sluiting van de terminals in België betrekking te hebben op verliesgevende activiteiten.
256. Teneinde uit te maken of deze twee maatregelen toereikend zijn om de nadelige gevolgen van de steun voor de concurrenten zoveel mogelijk te beperken, dient te worden herinnerd aan de voornaamste ontwikkelingen van de twee markten waarop IFB actief is, namelijk de logistiekmarkt en de overslagmarkt. Vervolgens moet worden onderzocht of de voorgestelde maatregelen de nadelige gevolgen van de steun voor de concurrenten zoveel mogelijk beperken.
a) De logistiekmarkt en de steun voor IFB
257. Zoals in deel 2 van deze beschikking werd uitgelegd, is de logistiekmarkt een markt in volle verandering als gevolg van de openstelling van de markten van het spoorwegvervoer en het betreden van de markt door spoorweg- en postbedrijven, met tegelijkertijd een groot aantal kleine gespecialiseerde spelers en grote geïntegreerde spelers.
258. De Commissie stelt vast dat de voorgestelde maatregelen geen betrekking hebben op de logistiekmarkt. Zoals uit de tabel in punt 16 van deze beschikking blijkt, heeft IFB zijn volume op deze markt in 2004 aanzienlijk weten te verhogen (in vergelijking met 2003). België heeft geen enkele verbintenis voorgelegd waardoor de aanwezigheid van IFB op deze markt tijdens de herstructureringsperiode zou zijn beperkt.
259. De Commissie is bijgevolg van oordeel dat de afwezigheid van voorgestelde maatregelen voor de logistiekmarkt, alsmede de feiten dat de markt in volle verandering is en dat IFB zijn volume aanzienlijk heeft weten te verhogen, twijfels doen rijzen over de vraag of België de nadelige gevolgen voor de concurrentie zoveel mogelijk heeft beperkt wat de logistiekactiviteiten van IFB betreft.
b) De overslagmarkt en de steun voor IFB
260. De twee voorgestelde maatregelen hebben betrekking op de overslagmarkt. IFB heeft zijn activiteiten in Frankrijk zo goed als stopgezet, en heeft een terminal in België gesloten en zijn participaties in twee andere terminals verkocht.
261. De enige markt waarvoor de steun negatieve gevolgen voor de concurrentie kan hebben, is dus de Belgische markt. Op deze markt heeft IFB een marktaandeel van minder dan 7 % (zie de beschrijving van de markten in deel 2 van deze beschikking).
262. Om de negatieve gevolgen van de steun op de Belgische markt te beperken, heeft IFB een terminal gesloten en zijn participaties in twee andere terminals verkocht. De Commissie stelt echter enerzijds vast dat de sluiting de kleinste van deze terminals betrof en in de eerste plaats diende om de verliezen van IFB Terminals te verminderen, en anderzijds dat IFB opnieuw de twee terminals zal exploiteren die de onderneming na de kapitaalverhoging heeft verkocht, want de maatschappij TRW, waarvan de NMBS 47 % van de aandelen in IFB zal inbrengen, bezit aanzienlijke participaties in de terminals van Brussel en Zeebrugge.
263. Vervolgens stelt de Commissie vast dat IFB minderheidsparticipaties in een aantal belangrijke Belgische terminals bezit.
264. Bijgevolg heeft de Commissie twijfels over de vraag of de door IFB voorgestelde maatregelen om de nadelige gevolgen van de steun voor de concurrentie op de overslagmarkt zoveel mogelijk te beperken, toereikend zijn.
3.2.2.4. Beperking van de steun tot het strikte minimum en bijdrage van de begunstigde onderneming
265. Teneinde aan te tonen dat de steun tot het strikte minimum beperkt blijft, legt de Belgische regering uit dat de kapitaalverhoging ertoe beperkt blijft het maatschappelijk kapitaal van IFB, dat als gevolg van de in 2001 en 2002 geboekte verliezen negatief was geworden, in zoverre te herstellen dat de onderneming haar economische levensvatbaarheid kan terugvinden. Zoals hierboven in deel 2 is uitgelegd, zal de solvabiliteitsratio, d.w.z. de verhouding eigen vermogen/passiva, van IFB na de kapitaalverhoging 33 % bedragen.
266. België heeft de Commissie de solvabiliteitsratio's van de voornaamste concurrenten van IFB meegedeeld. Deze zijn als volgt:
Terminalexploitanten | |
ABP Ports | 59,60 |
Hesse-Noord Natie | 58,19 |
Katoennatie Terminals | 54,97 |
Schelde Container Terminal Noord | 53,33 |
Sea-Ro-Terminal | 43,75 |
RSC | 74,24 |
Gemiddelde | 57,35 |
| |
Transportondernemingen | |
DHL Freight (weg) | 34,60 |
ECS European Containers (weg) | 14,27 |
Gefco Benelux (spoor) | 39,92 |
Henri Essers (weg) | 15,71 |
Rhinecontainer (binnenvaart) | 18,63 |
TRW (spoor) | 20,74 |
Ziegler (weg) | 20,42 |
Gemiddelde | 23,47 |
| |
Ondernemingen met gemengde activiteiten | |
Gosselin | 38,92 |
Hupac | 34,90 |
Gemiddelde | 36,91 |
| |
Algemeen gemiddelde | 39,24 |
267. De Commissie neemt er nota van dat de voor IFB beoogde solvabiliteitsratio lager is dan die van de terminalexploitanten en ook, ofschoon in mindere mate, lager dan die van de ondernemingen met gemengde activiteiten. Het cijfer is echter wel hoger dan het gemiddelde van de solvabiliteitsratio's voor de transportondernemingen. Voorts ligt de kapitaalverhoging ook 20 miljoen euro onder het bedrag dat de consultant McKinsey in het herstructureringsplan had aanbevolen. De Commissie beschikt evenwel in dit stadium niet over voldoende elementen om definitief te concluderen dat de steun tot het strikte minimum is beperkt.
268. De Commissie vestigt de aandacht van de Belgische regering op de bepalingen van punt 42 en volgende van de richtsnoeren van 2004, die luiden als volgt:
Van de steun ontvangende ondernemingen wordt verwacht dat zij uit eigen middelen, zo nodig door de verkoop van activa die voor het voortbestaan van de onderneming niet onontbeerlijk zijn of door externe financiering tegen marktvoorwaarden, een belangrijke bijdrage aan het herstructureringsplan leveren. Deze bijdrage is een teken dat de markten er vertrouwen in hebben dat een herstel van de levensvatbaarheid haalbaar is. Zij moet reëel — dus actueel — zijn, onder uitsluiting van alle voor de toekomst verwachte winst en kasstromen, en zij moet zo hoog mogelijk zijn.
In de regel beschouwt de Commissie de volgende bijdragen aan de herstructurering als passend: minstens 25 % in het geval van kleine ondernemingen, minstens 40 % in het geval van middelgrote en minstens 50 % in het geval van grote ondernemingen. In uitzonderlijke omstandigheden en in geval van een door de lidstaat aan te tonen bijzondere noodsituatie kan de Commissie een lagere bijdrage accepteren.
Om de mededingingsverstorende effecten te beperken, moet de omvang van de steun of de vorm waarin hij wordt verleend zodanig zijn dat de onderneming niet de beschikking krijgt over extra kasmiddelen die kunnen worden gebruikt voor agressieve, marktverstorende activiteiten welke met het herstructureringsproces geen verband houden. Daartoe onderzoekt de Commissie de omvang van de passiva van de onderneming na de herstructurering, evenals de situatie na uitstel van betaling of vermindering van haar schulden, met name in het kader van de voortzetting van haar activiteiten na een collectieve insolventieprocedure volgens het nationale recht. De steun mag noch geheel noch gedeeltelijk worden gebruikt voor de financiering van nieuwe investeringen die voor het herstel van de levensvatbaarheid van de onderneming niet onmisbaar zijn.
269. De Commissie stelt vast dat IFB volgens het herstructureringsplan geen eigen bijdrage tot zijn herstructurering lijkt te leveren. De Commissie heeft dan ook twijfels over de vraag of IFB, zoals in de richtsnoeren van 2004 wordt geëist, op voldoende wijze aan zijn herstructureringssteun bijdraagt.
3.2.2.5. Jaarverslag en "one time, last time"
270. De Belgische regering heeft ermee ingestemd een jaarverslag bij de Commissie in te dienen zodat de Commissie kan beoordelen of het herstructureringsplan ten uitvoer wordt gelegd overeenkomstig de door de Belgische autoriteiten aangegane verbintenissen.
271. Ten slotte dient te worden nagegaan of in verband met de herstructureringssteun het beginsel "one time, last time" is nageleefd. Volgens de door de Belgische autoriteiten verstrekte informatie heeft IFB voordien geen herstructureringssteun ontvangen. De Commissie heeft voordien geen besluit betreffende IFB genomen. Zij is dus van oordeel dat aan het criterium "one time, last time" is voldaan.
3.3. CONCLUSIE
272. De Commissie is in dit stadium van oordeel dat de toekenning van een uitstel van betaling voor de bestaande schulden van 63 miljoen euro en de omzetting daarvan en van de bijbehorende rente van 11 miljoen euro in maatschappelijk kapitaal staatssteun vormen, omdat de NMBS niet heeft gehandeld zoals een particuliere investeerder in een markteconomie zou hebben gedaan.
273. Vormen evenzo staatssteun de toekenning van een terugvorderbaar voorschot van 5 miljoen euro en de toekenning van een kredietfaciliteit van 15 miljoen euro, de omzetting van de kredietfaciliteit van 15 miljoen euro en van de bijbehorende rente van 2,5 miljoen euro in maatschappelijk kapitaal, alsmede de inbreng in natura van 5 miljoen euro nieuw maatschappelijk kapitaal.
274. In zoverre deze steun kassteun vormt, kan hij als herstructureringssteun niet verenigbaar met de gemeenschappelijke markt worden verklaard, omdat hij voor een periode van langer dan 12 maanden is toegekend.
275. De Commissie heeft twijfels over de vraag of de steun in zijn geheel als herstructureringssteun verenigbaar met de gemeenschappelijke markt kan worden verklaard.
276. Haar twijfels hebben betrekking op de toerekenbaarheid van een deel van de steun aan de Belgische staat, de toereikendheid van de maatregelen die zijn genomen om de nadelige gevolgen van de steun voor de concurrenten zoveel mogelijk te beperken, alsmede op de beperking van de steun tot het strikte minimum en op de toereikendheid van de eigen bijdrage van de onderneming IFB aan de herstructureringssteun.
4. BESCHIKKING
De Commissie heeft besloten de reddingsmaatregelen en de herstructureringsmaatregelen ten gunste van IFB in dit stadium te beschouwen als staatssteun als bedoeld in artikel 87, lid 1, van het EG-Verdrag.
Zij uit twijfels over de vraag of deze steun op grond van de richtsnoeren voor herstructureringssteun verenigbaar met de gemeenschappelijke markt kan worden verklaard, en leidt bijgevolg voor dit deel van de zaak de bij artikel 88, lid 2, van het EG-Verdrag vastgestelde procedure in.
Gelet op de bovenstaande overwegingen verzoekt de Commissie België in het kader van de procedure van artikel 88, lid 2, van het EG-Verdrag binnen een maand vanaf de datum van ontvangst van dit schrijven zijn opmerkingen te maken en alle dienstige inlichtingen te verstrekken voor de beoordeling van de steunmaatregel. Zij verzoekt uw autoriteiten onverwijld een afschrift van deze brief aan de potentiële begunstigde van de steunmaatregel te doen toekomen.
De Commissie wijst België op de schorsende werking van artikel 88, lid 3, van het EG-Verdrag. Zij verwijst naar artikel 14 van Verordening (EG) nr. 659/1999, volgens hetwelk elke onrechtmatige steun van de begunstigde kan worden teruggevorderd.
Voorts deelt de Commissie België mee, dat zij de belanghebbenden door de bekendmaking van dit schrijven en van een samenvatting ervan in het Publicatieblad van de Europese Unie in kennis zal stellen. Tevens zal zij de belanghebbenden in de lidstaten van de EVA die partij zijn bij de EER-Overeenkomst door de bekendmaking van een mededeling in het EER-Supplement van het Publicatieblad in kennis stellen, alsmede de Toezichthoudende Autoriteit van de EVA door haar een afschrift van dit schrijven toe te zenden. Alle bovengenoemde belanghebbenden zal worden verzocht hun opmerkingen te maken binnen een maand vanaf de datum van deze bekendmaking."
[1] Secret d'affaires
[2] […]
[3] […]
[4] […]
[5] Essentiellement des produits chimiques, des granulats, du charbon et des marchandises générales.
[6] TEU est l'abréviation pour twenty foot equivalent unit, c'est-à-dire un container de vingt pied de longueur. Un container de cette taille est le standard pour décrire les volumes transportés en transport combiné.
[7] Moniteur Belge du 24 juillet 1926.
[8] Date de l'entrée en vigueur de l'arrêté royal du 30 septembre 1992 portant approbation du premier contrat de gestion de la Société nationale des chemins de fer belges et fixant les mesures relatives à cette société, Moniteur Belge du 14 octobre 1992.
[9] Tel que définies dans la loi du 21 mars 1991 portant réforme de certaines entreprises publiques économiques, Moniteur belge du 27 mars 1991.
[10] Moniteur Belge du 4 août 1966.
[11] A titre d'information: depuis le 1 janvier 2004, ce taux est fixé à 4,43 % sur une base annuelle.
[12] Ce qui équivaut au minimum à un taux annuel de [entre 3,6 et 7,2 %].
[13] 23,9/72,3 = 0,33
[14] EUR 15 millions (mesure 2) + EUR 63 millions. (mesure 3) = EUR 78 millions, les EUR 5 millions (mesure 1) n'ayant pas été utilisés.
[15] Ce qui équivaut au minimum à un taux annuel de 5,4 %.
[16] Arrêt de la Cour du 16 mai 2002, C-482/99, France/Commission, Affaire dite "Stardust Marine", considérant 37.
[17] Directive de la Commission 2000/52/CE du 26 juillet 2000, JO L 193 du 29.07.2000, qui modifie la Directive 80/723/CEE du 25 juin 1980 relative à la transparence des relations financières entre les Etats membres et les entreprises publiques, JO L 195 du 29.7.1980.
[18] Arrêt de la Cour du 16 mai 2002, C-482/99, précité, considérant 37.
[19] Arrêt de la Cour du 16 mai 2002, C-482/99, précité, considérants 52 et 55.
[20] Arrêt de la Cour du 16 mai 2002, C-482/99, précité, considérants 53 et 54.
[21] Arrêt de la Cour du 2 février 1988, C-67, 68 et 70/85.
[22] Arrêts de la Cour du 21 mars 1991, C-303/88 et C-305/89.
[23] Arrêt de la Cour du 30 janvier 1985, 290/83.
[24] À savoir la nomination des dirigeants par l'Etat pour les arrêts Commission/Italie; le financement par un établissement public, les modalités d'octroi qui correspondent à celles d'une aide étatique ordinaire, la présentation par le gouvernement de l'aide comme faisant partie d'un ensemble de mesures étatiques pour l'arrêt Commission/France.
[25] Décision de la Commission du 17 septembre 2003 relative à l'aide d'Etat accordée par l'Allemagne en faveur de Space Park Development GmbH, JO L 61 du 27.2.2004, p. 66, considérant 30.
[26] Des articles de presse peuvent constituer un indice d'imputabilité, cf. décisions ABX Logistics, JO C 9 du 14.1.2004, p. 32; Sniace SA, JO L 108 du 30.4.2003, p. 35.
[27] "Inter Ferry Boats coupée en 2 branches", mise en ligne le 19/05/2003 sur le site www.lalibre.be
[28] Conclusions dans le cas C-276/2002 Espagne contre Commission, 1er avril 2004.
[29] Arrêt du TPI du 8 juillet 2004, T-198/01, Technische Glaswerke Ilmenau, considérant 99.
[30] Cf. l'arrêt de la Cour du 16 mai 2002, C-482/99, précité, considérant 70
[31] Cf. rapport annuel de la SNCB pour 2002, p. 8.
[32] Idem, p. 7.
[33] Arrêt du Tribunal du 15 septembre 1998, T-11/95, points 70 et suivants.
[34] Arrêt du 21 mars 1991, Italie/Commission, C-305/89, point 19 et 20; cf. aussi Arrêt du Tribunal du 6 mars 2003, affaire T-228/99, WestLB/Commission, point 245.
[35] Arrêt du 21 mars 1991, Italie/Commission, C-305/89, point 19 et 20.
[36] Cf. Arrêt du 6 mars 2003, WestLB Girozentrale/Commission, T-228/99 et T-233/99, point 2251.
[37] Cf. Arrêt du 6 mars 2003, WestLB Girozentrale/Commission, T-228/99 et T-233/99, point 246.
[38] Pratique constante de la Commission, cf. Décision de la Commission du 30 avril 1996 concernant des aides d'Etat en faveur de La Seda de Barcelona, JO L 298, 22.11.1996, p. 14. Le taux de référence est publié au JOUE, cf. JOUE C 88 du 12 avril 2005, p. 5.
[39] Arrêt du 21 mars 1991, Italie/Commission, C-305/89, point 19 et 20.
[40] Arrêt du 21 mars 1991, Italie/Commission, C-305/89, point 19 et 20.
[41] Cf. Arrêt du 6 mars 2003, WestLB Girozentrale/Commission, T-228/99 et T-233/99, point 2251.
[42] Cf. Arrêt du 6 mars 2003, WestLB Girozentrale/Commission, T-228/99 et T-233/99, point 246.
[43] Arrêt du 10 juillet 1986, Belgique/Commission, 234/84, point 14.
[44] Arrêt du 21 mars 1991, Italie/Commission, C-305/89, point 19 et 20.
[45] Arrêt de la Cour du 13 mars 1985, affaires jointes 296 et 318/82, Royaume des Pays-Bas et Leeuwarder Papierwarenfabriek/Commission, point 24.
[46] JO C 289 du 9.10.1999, p. 2, et JO C 244 du 1.10.2004, p. 2.
[47] V., à cet égard, l'arrêt du 14 janvier 2004, Fleuren Compost/Commission (T-109/01, non encore publié au Rec., point 74 ).
[48] Zakengeheim
[49] […]
[50] […]
[51] […]
[52] Hoofdzakelijk chemische producten, granulaat, steenkool en algemeen goederenvervoer.
[53] TEU is de afkorting van twenty foot equivalent unit, d.w.z. een container met een lengte van 20 voet. Een container van die grootte is de standaard om de volumes te beschrijven die via gecombineerd vervoer worden getransporteerd.
[54] Belgisch Staatsblad van 24 juli 1926.
[55] Datum van inwerkingtreding van het Koninklijk Besluit van 30 september 1992 houdende goedkeuring van het eerste beheerscontract van de NMBS en vaststelling van de maatregelen betreffende deze maatschappij, Belgisch Staatsblad van 14 oktober 1992.
[56] Zoals omschreven in de wet van 21 maart 1991 houdende hervorming van sommige economische overheidsbedrijven, Belgisch Staatsblad van 27 maart 1991.
[57] Belgisch Staatsblad van 4 augustus 1966.
[58] Ter informatie: deze rentevoet is sinds 1 januari 2004 vastgesteld op 4,43 % op jaarbasis.
[59] Hetgeen overeenkomt met een jaarrente van minstens [tussen 3,6 en 7,2] %.
[60] 23,9/72,3 = 0,33
[61] 15 miljoen euro (maatregel 2) + 63 miljoen euro (maatregel 3) = 78 miljoen euro, aangezien de 5 miljoen euro (maatregel 1) niet waren gebruikt.
[62] Hetgeen overeenkomt met een jaarrente van minstens 5,4 %.
[63] Arrest van het Hof van 16 mei 2002, C-482/99, Frankrijk/Commissie, in de zaak "Stardust Marine", punt 37.
[64] Richtlijn 2000/52/EG van de Commissie van 26 juli 2000 (PB L 193 van 29.7.2000) tot wijziging van Richtlijn 80/723/EEG betreffende de doorzichtigheid in de financiële betrekkingen tussen lidstaten en openbare bedrijven (PB L 195 van 29.7.1980).
[65] Arrest van het Hof van 16 mei 2002, C-482/99, reeds aangehaald, punt 37.
[66] Arrest van het Hof van 16 mei 2002, C-482/99, reeds aangehaald, punten 52 en 55.
[67] Arrest van het Hof van 16 mei 2002, C-482/99, reeds aangehaald, punten 53 en 54.
[68] Arrest van het Hof van 2 februari 1988, C-67, 68 en 70/85.
[69] Arresten van het Hof van 21 maart 1991, C-303/88 en C-305/89.
[70] Arrest van het Hof van 30 januari 1985, 290/83.
[71] Namelijk: de benoeming van de bestuurders door de staat voor de arresten Commissie/Italië; de financiering door een publieke instantie, de toekenningsmodaliteiten die identiek zijn bij gewone staatssteun, het feit dat de regering de steun als onderdeel van een pakket overheidsmaatregelen voostelde voor het arrest Commissie/Frankrijk.
[72] Beschikking van de Commissie van 17 september 2003 betreffende de staatssteun die Duitsland aan Space Park Development GmbH heeft verleend, PB L 61 van 27.2.2004, blz. 66, overweging 30.
[73] Berichten in de pers kunnen een aanwijzing voor betrokkenheid vormen, zie de zaken ABX Logistics, PB C 9 van 14.1.2004, blz. 32; Sniace SA, PB L 108 van 30.4.2003, blz. 35.
[74] "Inter Ferry Boats coupée en 2 branches verdeeld", op 19/05/2003 op internet gezet op de website www.lalibre.be.
[75] Conclusies in zaak C-276/2002, Spanje tegen Commissie, 1 april 2004.
[76] Arrest van het Gerecht van eerste aanleg van 8 juli 2004, T-198/01, Technische Glaswerke Ilmenau, punt 99.
[77] Arrest van het Hof van 16 mei 2002, C-482/99, reeds aangehaald, punt 70.
[78] Zie jaarverslag 2002 van de NMBS, blz. 8.
[79] Idem, blz. 7.
[80] Arrest van het Gerecht van eerste aanleg van 15 september 1998, T-11/95, punten 70 e.v.
[81] Arrest van 21 maart 1991, Italië/Commissie, C-305/89, punten 19 en 20; zie ook Arrest van het Gerecht van eerste aanleg van 6 maart 2003, zaak T-228/99, WestLB/Commissie, punt 245.
[82] Arrest van 21 maart 1991, Italië/Commissie, C-305/89, punten 19 en 20.
[83] Zie arrest van 6 maart 2003, WestLB Girozentrale/Commissie, T-228/99 en T-233/99, punt 251.
[84] Zie arrest van 6 maart 2003, WestLB Girozentrale/Commissie, T-228/99 en T-233/99, punt 246.
[85] Vaste praktijk van de Commissie, zie Beschikking van de Commissie van 30 april 1996 betreffende staatssteun voor La Seda de Barcelona SA, PB L 298 van 22.11.1996, blz. 14. De referentierente wordt gepubliceerd in het PBEU, zie PBEU C 88 van 12.4.2005, blz. 5.
[86] Arrest van 21 maart 1991, Italië/Commissie, C-305/89, punten 19 en 20.
[87] Arrest van 21 maart 1991, Italië/Commissie, C-305/89, punten 19 en 20.
[88] Zie arrest van 6 maart 2003, WestLB Girozentrale/Commissie, T-228/99 en T-233/99, punt 251.
[89] Zie arrest van 6 maart 2003, WestLB Girozentrale/Commissie, T-228/99 en T-233/99, punt 246.
[90] Arrest van 10 juli 1986, België/Commissie, 234/84, punt 14.
[91] Arrest van 21 maart 1991, Italië/Commissie, C-305/89, punten 19 en 20.
[92] Arrest van het Hof van 13 maart 1985, gevoegde zaken 296 en 318/82, Koninkrijk der Nederlanden en Leeuwarder Papierwarenfabriek/Commissie, punt 24.
[93] PB C 288 van 9.10.1999, blz. 2, en PB C 244 van 1.10.2004, blz. 2.
[94] Zie in dit verband het arrest van 14 januari 2004, Fleuren Compost/Commissie (T-109/01, nog niet in de Jurisprudentie gepubliceerd, punt 74).
--------------------------------------------------
Riktlinjer för beräkning av böter som döms ut enligt artikel 23.2 a i förordning nr 1/2003
(2006/C 210/02)
(Text av betydelse för EES)
INLEDNING
1. Enligt artikel 23.2 a i förordning nr 1/2003 [1] får kommissionen genom beslut ålägga företag och företagssammanslutningar böter, om de uppsåtligen eller av oaktsamhet överträder artikel 81 eller artikel 82 i fördraget.
2. Inom de gränser som fastställs i förordning nr 1/2003 har kommissionen stort utrymme för att göra egna bedömningar [2] när den ålägger företag sådana böter. Först och främst skall kommissionen beakta överträdelsens allvar och varaktighet. Böterna får inte överskrida de gränser som anges i artikel 23.2 andra och tredje stycket i förordning nr 1/2003.
3. För att garantera insyn och objektivitet i sina beslut offentliggjorde kommissionen den 14 januari 1998 riktlinjer för beräkning av böter [3]. Riktlinjerna har nu tillämpats i över åtta år och kommissionen har därför fått tillräcklig erfarenhet av tillämpningen för att kunna utveckla och finslipa sin politik i fråga om böter.
4. Kommissionen har fått behörighet att ålägga företag och företagssammanslutningar böter om de uppsåtligen eller av oaktsamhet överträder bestämmelserna i artikel 81 eller 82 i fördraget för att den skall kunna utföra det övervakningsuppdrag som den anförtros i fördraget. Övervakningsuppdraget innebär inte enbart att kommissionen skall undersöka och bestraffa individuella överträdelser, utan också att dess politik rent allmänt skall vara att i konkurrensfrågor tillämpa de principer som fastställs i fördraget och på så sätt styra företagens beteende [4]. I samband med detta måste kommissionen se till att dess åtgärder har tillräckligt avskräckande verkan [5]. När kommissionen finner att bestämmelserna i artikel 81 eller 82 i fördraget har överträtts, kan det därför bli nödvändigt att ålägga företag som har överträtt bestämmelserna böter. Böterna skall vara så stora att de är tillräckligt avskräckande, inte bara för att bestraffa de berörda företagen (specifik avskräckande verkan), utan också för att avskräcka andra företag från att agera på ett sätt som strider mot artiklarna 81 och 82 i fördraget (allmän avskräckande verkan).
5. För att nå dessa mål bör kommissionen fastställa böterna på grundval av försäljningsvärdet av de varor eller tjänster som överträdelsen avser. Överträdelsens varaktighet bör också spela en viktig roll vid fastställandet av bötesbeloppet. Varaktigheten har naturligtvis stor betydelse för i vilken utsträckning överträdelsen påverkar marknaden. Det är därför viktigt att böterna återspeglar hur många år företaget har deltagit i överträdelsen.
6. Kombinationen av försäljningsvärdet och varaktigheten är ett lämpligt beräkningstal för att värdera överträdelsens ekonomiska betydelse och omfattningen av varje företags delaktighet i överträdelsen. Dessa mått ger en god indikation om ett rimligt bötesbelopp, men de skall inte ses som en automatisk och aritmetisk grund för beräkningen av böterna.
7. I böterna bör det också ingå ett särskilt belopp som inte är beroende av överträdelsens varaktighet och som har till syfte att avskräcka företagen från att begå nya överträdelser.
8. I följande avsnitt beskrivs de principer som kommissionen följer när den fastställer böter enligt artikel 23.2 a i förordning nr 1/2003.
METOD FÖR ATT FASTSTÄLLA BÖTER
9. När kommissionen fastställer de böter som skall åläggas företag eller företagssammanslutningar använder den en tvåstegsmetod (följande beskrivning påverkar inte tillämpningen av punkt 37 nedan).
10. I det första steget fastställer kommissionen ett grundbelopp för varje företag eller företagssammanslutning (se avsnitt 1 nedan).
11. I det andra steget kan kommissionen höja eller sänka grundbeloppet (se avsnitt 2 nedan).
1) Grundbelopp
12. Grundbeloppet fastställs på grundval av försäljningsvärdet med hjälp av den metod som beskrivs nedan.
A. Fastställande av försäljningsvärdet
13. Kommissionen fastställer grundbeloppet genom att utgå från försäljningsvärdet från de varor eller tjänster som har ett direkt eller indirekt [6] samband med överträdelsen och som företaget sålt i det berörda geografiska området inom EES. Kommissionen utgår i regel ifrån företagets försäljning under det sista kompletta räkenskapsåret då det deltar i överträdelsen (nedan kallat "försäljningsvärdet").
14. Om det är en företagssammanslutning som begått överträdelsen och överträdelsen avser medlemmarnas verksamhet, utgår kommissionen i regel från medlemmarnas sammanlagda försäljningsvärde.
15. När kommissionen fastställer ett företags försäljningsvärde utgår den från de bästa uppgifter som finns tillgängliga för företaget.
16. Om ett företags uppgifter är ofullständiga eller otillförlitliga, kan kommissionen fastställa företagets försäljningsvärde på grundval av de ofullständiga uppgifterna och/eller alla andra uppgifter som den anser relevanta.
17. I försäljningsvärdet ingår inte moms eller andra skatter som är direkt knutna till försäljningen.
18. Om överträdelsen sträcker sig utanför EES (till exempel världsomfattande karteller) räcker det i vissa fall inte med att fastställa ett företags försäljning inom EES för att ge en korrekt bild av företagets delaktighet i överträdelsen. Det kan framför allt vara fallet vid världsomfattande avtal om uppdelning av marknaden.
I sådana fall kan kommissionen fastställa försäljningsvärdet inom EES och omfattningen av varje företags delaktighet i överträdelsen genom att uppskatta det sammanlagda försäljningsvärdet av de varor eller tjänster överträdelsen avser i det berörda geografiska området (större än EES), fastställa varje deltagande företags andel av försäljningen på denna marknad, och lägga denna andel till varje företags totala försäljning inom EES. Resultatet betraktas som företagets försäljningsvärde när kommissionen fastställer grundbeloppet för böterna.
B. Fastställande av grundbeloppet
19. Grundbeloppet för böterna kommer att vara knutet till en andel av försäljningsvärdet och grundas på överträdelsens allvar multiplicerat med antalet år som företaget deltagit i överträdelsen.
20. Överträdelsens allvar fastställs från fall till fall för varje typ av överträdelse med beaktande av alla relevanta omständigheter i ärendet.
21. Regelmässigt uppgår den andel av försäljningsvärdet som beaktas till högst 30 %.
22. När kommissionen fastställer om den andel av försäljningsvärdet som skall beaktas i ett visst fall skall ligga i nedre eller övre delen av denna skala, tar den hänsyn till en rad faktorer, bland annat överträdelsens art, de berörda parternas sammanlagda marknadsandel, överträdelsens geografiska omfattning och om överträdelsen har genomförts eller ej.
23. Horisontella avtal [7] om fastställande av priser, uppdelning av marknaden och produktionsbegränsningar, som i allmänhet är hemliga, hör till mest allvarliga konkurrensbegränsningarna. EU:s konkurrenspolitik innebär att sådana överträdelser bestraffas hårt. I regel kommer därför den andel av försäljningsvärdet som skall beaktas vid sådana överträdelser att bestämmas i den övre delen av skalan.
24. För att överträdelsens varaktighet skall beaktas fullt ut för varje enskilt företag multipliceras det belopp som fastställs på grundval av försäljningsvärdet (se punkterna 20-23 ovan) med antalet år som företaget deltagit i överträdelsen. Perioder under sex månader räknas som ett halvår, medan perioder över sex månader, men kortare än ett år, räknas som ett helt år.
25. Dessutom skall kommissionen, oavsett varaktigheten av företagets överträdelse, höja grundbeloppet med ett belopp på mellan 15 och 25 % av försäljningsvärdet (se definitionen i avsnitt A ovan) för att avskräcka företagen från att över huvud taget delta i horisontella avtal om fastställande av priser, uppdelning av marknaden och produktionsbegränsningar. Kommissionen kan lägga till ett sådant belopp även vid andra typer av överträdelser. När kommissionen fastställer hur stor andel av försäljningsvärdet som skall beaktas i ett enskilt ärende tar den hänsyn till en rad faktorer, särskilt de som anges i punkt 22 ovan.
26. Om flera företag som deltagit i överträdelsen har ett försäljningsvärde som är nästan identisk, men inte helt, kan kommissionen ändå fastställa samma grundbelopp för vart och ett av företagen. Kommissionen avrundar dessutom siffrorna när den fastställer grundbeloppet för böterna.
2) Justering av grundbeloppet
27. När kommissionen fastställer böterna kan den beroende på omständigheterna höja eller sänka böterna på det sätt som beskrivs i avsnitt 1 ovan. Kommissionen beslutar om böterna skall höjas eller sänkas på grundval av en helhetsbedömning där den tar hänsyn till alla relevanta omständigheter.
A. Försvårande omständigheter
28. Grundbeloppet kan höjas om kommissionen konstaterar att det finns försvårande omständigheter, till exempel följande:
- Ett företag fortsätter med eller upprepar en identisk eller liknande överträdelse efter det att kommissionen eller en nationell konkurrensmyndighet har konstaterat att företaget har överträtt bestämmelserna i artikel 81 eller artikel 82 i fördraget. Grundbeloppet höjs med upp till 100 % för varje överträdelse som fastställs.
- Företaget vägrar att samarbeta eller hindrar kommissionens undersökning.
- Företaget har haft en ledande roll, eller initiativet, vid överträdelsen. Kommissionen riktar också särskild uppmärksamhet mot alla åtgärder som vidtas för att tvinga andra företag att delta i överträdelsen och/eller alla vedergällningsåtgärder som vidtas mot andra företag för att få dem hålla sig till det beteende som utgör överträdelsen.
B. Förmildrande omständigheter
29. Grundbeloppet kan sänkas om kommissionen konstaterar att det finns förmildrande omständigheter, till exempel följande:
- Det berörda företaget kan visa att det upphörde med överträdelsen omedelbart efter kommissionens första åtgärder. Detta gäller dock inte hemliga avtal eller åtgärder (särskilt karteller).
- Det berörda företaget kan visa att överträdelsen har begåtts av oaktsamhet.
- Det berörda företaget kan visa att dess deltagande i överträdelsen har varit mycket begränsat, eftersom företaget under den tid då det var det var bundet av de otillåtna avtalen i realiteten undvek att tillämpa dem genom att bete sig på ett konkurrensinriktat sätt på marknaden. Att ett företag har deltagit i en överträdelse under en kortare period än de andra företagen betraktas inte som någon förmildrande omständighet, eftersom kommissionen redan tagit hänsyn till detta när den fastställt grundbeloppet.
- Företaget samarbetar med kommissionen i en omfattning som går utöver tillämpningsområdet för tillkännagivandet om befrielse från eller nedsättning av böter i kartellärenden, samt företagets lagstadgade skyldighet att samarbeta.
- Företagets konkurrensbegränsande beteende har godkänts eller uppmuntrats av de offentliga myndigheterna eller lagstiftningen. [8]
C. Särskild höjning i avskräckande syfte
30. Kommissionen fäster särskild vikt vid att böterna har en tillräckligt avskräckande effekt. Därför kan kommissionen höja böterna för företag som har en särskilt stor omsättning som härrör från försäljningen av andra varor eller tjänster än de som berörs av överträdelsen.
31. Kommissionen anser det också nödvändigt att höja böterna så att de är högre än de olagliga vinster som erhållits på grund av överträdelsen, om det är möjligt att uppskatta dessa vinster.
D. Högsta tillåtna bötesbelopp
32. Enligt artikel 23.2 i förordning nr 1/2003 får böterna för varje företag och företagssammanslutning som deltagit i överträdelsen inte överstiga 10 % av föregående räkenskapsårs sammanlagda omsättning.
33. Om en företagssammanslutnings överträdelse har samband med dess medlemmars verksamhet, får böterna inte överstiga 10 % av summan av den sammanlagda omsättningen hos varje medlem med verksamhet på den marknad som påverkas av sammanslutningens överträdelse.
E. Tillkännagivandet om förmånlig behandling
34. Kommissionen kan ge företag förmånlig behandling i enlighet med bestämmelserna i tillkännagivandet om befrielse från eller nedsättning av böter i kartellärenden.
F. Faktisk betalningskapacitet
35. I undantagsfall kan kommissionen på begäran beakta ett företags faktiska betalningskapacitet i en viss ekonomisk kontext och i ett samhällssammanhang. För att kommissionen skall sätta ned böterna med hänsyn till företagets faktiska betalningskapacitet räcker det inte med att ett företag har en ogynnsam ekonomisk situation eller går med förlust. Böterna kan sättas ned endast om det finns objektiva bevis för att böter som åläggs på de villkor som fastställs i riktlinjerna för beräkning av böter oåterkalleligen skulle äventyra det berörda företagets ekonomiska bärkraft och leda till att företagets tillgångar förlorade allt värde.
SLUTKOMMENTAR
36. Kommissionen kan i vissa fall ålägga symboliska böter. Skälen för sådana symboliska böter bör anges i beslutet.
37. I riktlinjerna för beräkning av böter beskrivs en allmän metod för att fastställa böter, men kommissionen har rätt att avvika från denna metod eller från de gränser som fastställs i punkt 21 om omständigheterna i ett enskilt ärende kräver det eller om det krävs för att uppnå en tillräcklig avskräckande effekt.
38. Dessa riktlinjer tillämpas i alla ärenden där kommissionen har utfärdat ett meddelande om invändningar efter det att riktlinjerna offentliggjordes i den Europeiska unionens officiella tidning, oavsett om böterna åläggs enligt artikel 23.2 i förordning nr 1/2003 eller enligt artikel 15.2 i förordning nr 17 [9].
[1] Rådets förordning (EG) nr 1/2003 av den 16 december 2002 om tillämpning av konkurrensreglerna i artiklarna 81 och 82 i fördraget, EGT L 1, 4.1.2003, s. 1.
[2] Se t.ex. domstolens dom i förenade målen C-189/02 P, C-202/02 P, C-205/02 P till C-208/02 P och C-213/02 P av den 28 juni 2005, Dansk Rørindustri A/S m.fl. mot kommissionen, REG 2005, s. I-5425, punkt 172.
[3] Riktlinjer för beräkning av böter som döms ut enligt artikel 15.2 i förordning nr 17 och artikel 65.5 i EKSG-fördraget, EGT C 9, 14.1.1998, s. 3.
[4] Se till exempel punkt 170 i domen i mål Dansk Rørindustri A/S m.fl. mot kommissionen, som det hänvisas till i fotnot 2.
[5] Se domstolens dom av den 7 juni 1983 i förenade målen 100-103/80, Musique Diffusion française m.fl. mot kommissionen, Rec. 1983, s. 1825, punkt 106.
[6] Så kan till exempel ske i samband med horisontella arrangemang om fastställande av priser för en viss produkt när priset på denna produkt tjänar som grund för priset på andra produkter av antingen lägre eller högre kvalitet.
[7] Med detta avses avtal, samordnade förfaranden och beslut av företagssammanslutningar i enlighet med artikel 81 i fördraget.
[8] Detta påverkar dock inte eventuella förfaranden som inleds mot den berörda medlemsstaten.
[9] Artikel 15.2 i förordning nr 17 av den 6 februari, Första förordningen om tillämpning av fördragets artiklar 85 och 86 [nu artikel 81 och 82] (EGT 13, 21.2.1962, s. 204).
--------------------------------------------------
Kommissionens meddelande inom ramen för genomförandet av Europaparlamentets och rådets direktiv 2001/16/EG av den 19 mars 2001 om driftskompatibiliteten hos det transeuropeiska järnvägssystemet för konventionella tåg
(2006/C 243/02)
(Text av betydelse för EES)
(Offentliggörande av titlar på och hänvisningar till harmoniserade standarder inom ramen för direktivet)
ESO [1] | Titel på och hänvisning till standarden (samt referensdokument) | Hänvisning till den ersatta standarden | Datum då standarden upphör att gälla Anm. 1 |
CEN | EN 13715:2006 Hjulsatser och boggier – Hjul – Fälgprofil | — | |
CEN | EN 14531-1:2005 Järnvägar – Metoder för beräkning av stoppsträcka och nedbromsningssträcka, samt hållbroms och parkeringsbroms – Del 1: Allmänna algoritmer | — | |
CEN | EN 14535-1:2005 Järnvägar – Bromsskivor för rullande materiel – Del 1: Pressade eller krympta bromsskivor på axel eller drivaxel – Mått och kvalitetskrav | — | |
CEN | EN 14601:2005 Järnvägar – Rak och vinklad kran för broms- och huvudledning | — | |
Anmärkning 1 Det datum då den ersatta standarden upphör att gälla är i allmänhet det datum då den upphävs av det europeiska standardiseringsorganet. Användare av dessa standarder bör dock vara medvetna om att det i vissa undantagsfall kan vara ett annat datum
Anmärkning 3 Om tillägg förekommer innefattar hänvisningen såväl standarden EN CCCCC:YYYY som eventuella tidigare tillägg och det nya, angivna, tillägget. Den ersatta standarden (kolumn 3) består därför av EN CCCCC:YYYY med eventuella tidigare tillägg, men utan det nya, angivna, tillägget. Vid angivet datum upphör den ersatta standarden att gälla
Anmärkning:
- Närmare upplysningar om standarderna kan erhållas från de europeiska och nationella standardiseringsorgan som anges i bilagan till Europaparlamentets och rådets direktiv 98/34/EG [2], ändrat genom direktiv 98/48/EG [3].
- Offentliggörandet av hänvisningarna i Europeiska unionens officiella tidning innebär inte att de aktuella standarderna är tillgängliga på alla gemenskapsspråken.
- Denna förteckning ersätter alla tidigare förteckningar som har publicerats i Europeiska unionens officiella tidning. Kommissionen skall fortlöpande uppdatera denna förteckning.
Mer information återfinns på Europa-servern på Internet:
http://europa.eu.int/comm/enterprise/newapproach/standardization/harmstds/
[1] ESO: Europeiskt standardiseringsorgan:
- CEN: rue de Stassart 36, B-1050 Bryssel, Tel. (32-2) 550 08 11; fax (32-2) 550 08 19 (http://www.cenorm.be)
- CENELEC: rue de Stassart 35, B-1050 Bryssel, Tel. (32-2) 519 68 71; fax (32-2) 519 69 19 (http://www.cenelec.org)
- ETSI: 650, route des Lucioles, F-06921 Sophia Antipolis, Tel. (33) 492 94 42 00; fax (33) 493 65 47 16 (http://www.etsi.org)
[2] EGT L 204, 21.7.1998, s. 37
[3] EGT L 217, 5.8.1998, s. 18.
--------------------------------------------------
Frankrikes ändringar av den allmänna trafikplikten för regelbunden lufttrafik mellan Strasbourg och Madrid
(2006/C 246/04)
(Text av betydelse för EES)
1. Frankrike har beslutat att från och med den 25 mars 2007 ändra de bestämmelser om allmän trafikplikt för regelbunden lufttrafik mellan Strasbourg och Madrid som offentliggjorts i Europeiska gemenskapernas officiella tidning C 348 av den 5 december 2000 i enlighet med artikel 4.1 a i rådets förordning (EEG) nr 2408/92 av den 23 juli 1992 om EG-lufttrafikföretags tillträde till flyglinjer inom gemenskapen
2. Följande regler gäller för den allmänna trafikplikten:
2.1. Lägsta antalet flygningar
Flyglinjen skall trafikeras, utan mellanlandning, mellan Strasbourg och Madrid, med minst en tur- och returresor per dag, från måndag till fredag hela året.
2.2. Flygplanstyp och minimikapacitet
Trafiken skall bedrivas med flygplan med turbojetmotorer och med minst 48 platser.
2.3. Tidtabell
Flygningen varje dag från Madrid skall möjliggöra anslutningar med flyg från iberiska halvön.
Tidtabellen skall anpassas till Europaparlaments möten, så att en ankomst i Strasbourg läggs så nära kl. 14.00 som möjligt, men inte senare, för att passa till möten som börjar kl. 15.00, och en avgång från Strasbourg läggs så nära kl. 17.00 som möjligt, dock inte tidigare, för att passa till mötenas slut.
2.4. Biljettförsäljning
Flygningarna skall saluföras med hjälp av ett datoriserat reservationssystem.
2.5. Trafikens kontinuitet
Med undantag för force majeure får antalet flygningar som inställs av skäl som direkt kan tillskrivas trafikföretaget ej överstiga 2 % av antalet planerade flygningar per IATA-säsong. Lufttrafikföretaget får endast avbryta trafiken med minst sex månaders varsel.
Gemenskapens lufttrafikföretag upplyses om att trafikering av linjerna som är oförenlig med ovan fastställda bestämmelser om allmän trafikplikt kan medföra administrativa eller rättsliga åtgärder
--------------------------------------------------
Uppgifter från medlemsstaterna om statligt stöd som beviljats enligt kommissionens förordning (EG) nr 70/2001 av den 12 januari 2001 om tillämpningen av artiklarna 87 och 88 i EG-fördraget på statligt stöd till små och medelstora företag
(2006/C 289/02)
(Text av betydelse för EES)
Stöd nummer | XS 79/06 |
Medlemsstat | Tyskland |
Region | Freie und Hansestadt Hamburg |
Namnet på stödordningen eller namnet på det företag som tar emot det enskilda stödet | Hodorff Qualitätslogistic GmbH Banksstraße 28 D-20097 Hamburg |
Rättslig grund | Einzelfallentscheidung der Kreditkommission gemäß dem Gesetz über die Kreditkommission vom 29.4.1997 (Hamburgisches Gesetz- und Verordnungsblatt 1997, Nr. 18, Seite 133). Verordnung (EG) Nr. 70/2001 der Kommission vom 12. Januar 2001 über die Anwendung der Artikel 87 und 88 EG-Vertrag auf staatliche Beihilfen an kleine und mittlere Unternehmen (Amtsblatt der Europäischen Gemeinschaften 13.1.2001 L 10/33) |
Stödordningens beräknade utgifter per år eller totalt belopp som beviljats företaget som enskilt stöd | Stödordning | Årligt totalbelopp | |
Garanterade lån | |
Enskilt stöd | Totalt stödbelopp | 27300 EUR |
Garanterade lån | 5,46 milj. EUR |
Högsta tillåtna stödnivå | Överensstämmer med artikel 4.2-4.6 och artikel 5 i förordningen | Ja |
Datum för genomförande | Fr.o.m. den 15 maj 2006 |
Stödordningens eller det enskilda stödets varaktighet | Inget stöd eller utbetalning då det gäller engångsgaranti |
Stödets syfte | Stöd till små och medelstora företag | Ja |
Sektor(er) av ekonomin som berörs | Begränsat till vissa sektorer | Ja |
Andra tjänster | Ja |
Den beviljande myndighetens namn och adress | Freie und Hansestadt Hamburg Behörde für Wirtschaft und Arbeit Referat Finanzierungshilfen |
Alter Steinweg 4 D-20459 Hamburg |
Beviljande av stora enskilda stöd | I överensstämmelse med artikel 6 i förordningen | Ja |
Stöd nummer | XS 90/06 |
Medlemsstat | Tyskland |
Namnet på stödordningen eller namnet på det företag som tar emot det enskilda stödet | Programm zur Innovationsförderung/Bundesministerium für Ernährung, Landwirtschaft und Verbraucherschutz |
Rättslig grund | Programm und zugehörige Bekanntmachungen sind unter www.ble.de (Link Innovationsförderung — dort unter 3. Download des Programms zur Innovationsförderung des Bundesministeriums für Ernährung, Landwirtschaft und Verbraucherschutz (PDF-Dokument) und 3.1 Download der Bekanntmachung einer Richtlinie über die Förderung innovativer Pflanzenschutzvorhaben zur Reduzierung der Anwendung von Pflanzenschutzmitteln im Rahmen des Programms zur Innovationsförderung (PDF-Dokument)) einsehbar |
Stödordningens beräknade utgifter per år eller totalt belopp som beviljats företaget som enskilt stöd | Stödordning | Årligt totalbelopp | 21,6 milj. EUR |
Garanterade lån | |
Enskilt stöd | Totalt stödbelopp | |
Garanterade lån | |
Högsta tillåtna stödnivå | Överensstämmer med artikel 4.2-4.6 och artikel 5 i förordningen | Ja |
Datum för genomförande | Programmet sätts i verket omedelbart; anslagen utbetalas allteftersom, efter tillkännagivande och ansökan |
Stödordningens eller det enskilda stödets varaktighet | Ej begränsad. Programmet kommer att anpassas om förordning (EG) 70/2001 ersätts och detta gör en anpassning nödvändig. |
Stödets syfte | Stöd till små och medelstora företag | Ja |
Sektor(er) av ekonomin som berörs | Alla sektorer som är berättigade till stöd till små och medelstora företag | Ja |
Den beviljande myndighetens namn och adress | Bundesanstalt für Landwirtschaft und Ernährung (BLE) Projektgruppe Innovationsförderung |
Deichmanns Aue 29 D-53179 Bonn |
Beviljande av stora enskilda stöd | I överensstämmelse med artikel 6 i förordningen | (Inte relevant) |
Stöd nummer | XS 112/06 |
Medlemsstat | Nederländerna |
Region | Provinsen Zuid-Holland |
Namnet på stödordningen eller namnet på det företag som tar emot det enskilda stödet | Bioception B.V. |
Rättslig grund | Artikel 12 van de Algemene subsidieverordening Zuid-Holland, 1 juni 2005 |
Stödordningens beräknade utgifter per år eller totalt belopp som beviljats företaget som enskilt stöd | Stödordning | Årligt totalbelopp | |
Garanterade lån | |
Enskilt stöd | Totalt stödbelopp | 139001 EUR |
Garanterade lån | |
Högsta tillåtna stödnivå: | Överensstämmer med artikel 4.2-4.6 och artikel 5 i förordningen | Ja, nivån på det statliga stödet är 45 % (konkurrensneutral forskning) |
Datum för genomförande | 13.6.2006. Villkorat, stödet beviljas efter offentliggörande. |
Stödordningens eller det enskilda stödets varaktighet | T.o.m. den 31 december 2007 Åtgärden kommer vid behov att anpassas till tillämpliga bestämmelser i förordning 70/2001 när denna har ändrats. Kommissionen kommer att underrättas om detta |
Stödets syfte | Stöd till små och medelstora företag | Ja Detta forsknings- och utvecklingsprojekt syftar till att öka kunskapen om och utveckla tekniken när det gäller den praktiska användningen av biologiska testmedier. Det ställs allt högre krav på kvalitet och hygien vid tillverkning av läkemedel och livsmedel (bl.a. HACCP). Resultatet blir att störande mätningar leder till en försämring av produkten. De instrument som använts måste rengöras efteråt. För att upprätthålla den föreskrivna sterilitetsgraden måste allt dyrare apparater införskaffas. Detta projekt innebär ett möjligt alternativ, genom forskning och utveckling av ny kunskap och teknik när det gäller engångsbehållare som är utrustade med möjligheter att samla in och överföra data. Under tillverkningen mäts processparametrarna online och skickas till ett centralt system för processtyrning. Det är nödvändigt med teknisk forskning för att få fram de fysiska komponenterna, som måste vara små och billiga. Universitetet i Delft sörjer för den vetenskapliga kunskapen och för utvecklingen av de remsor där sensorerna placeras |
Sektor(er) av ekonomin som berörs | Begränsat till vissa sektorer | Ja |
Annan tillverkning | Verksamhetsområde som levererar till flera olika sektorer |
Den beviljande myndighetens namn och adress | Provincie Zuid-Holland |
Postbus 90602 2509 LP Den Haag Nederland |
Beviljande av stora enskilda stöd | I överensstämmelse med artikel 6 i förordningen | Ja |
Stöd nummer | XS 118/06 |
Medlemsstat | Nederländerna |
Region | Provinsen Flevoland |
Namnet på stödordningen eller namnet på det företag som tar emot det enskilda stödet | Eenmanszaak Pitch %amp% Putt Swifterbant te Swifterbant |
Rättslig grund | Decentralisatie-convenant Rijk/Flevoland m.b.t. het Leader+ programma Regio Randstad 2000-2006 d.d. 11 april 2001.Leader+ overeenkomst tussen de provincie Flevoland en Pitch %amp% Putt Swifterbant. |
Stödordningens beräknade utgifter per år eller totalt belopp som beviljats företaget som enskilt stöd | Stödordning | Årligt totalbelopp | |
Garanterade lån | |
Enskilt stöd | Totalt stödbelopp | 155700 EUR |
Garanterade lån | |
Högsta tillåtna stödnivå | Överensstämmer med artikel 4.2-4.6 och artikel 5 i förordningen | Ja Stödnivån är 12,4 %. Detta överensstämmer med artikel 4.2 a i förordning (EG) nr 70/2001 |
Datum för genomförande | Beslutet träder i kraft när det har offentliggjorts i EUT |
Stödordningens eller det enskilda stödets varaktighet | T.o.m. den 30 november 2007. Åtgärden kommer vid behov att anpassas till tillämpliga bestämmelser i förordning 70/2001 när denna har ändrats. Kommissionen kommer att underrättas om detta |
Stödets syfte | Stöd till små och medelstora företag | Ja. Stöd beviljas för investeringar i materiella tillgångar (art. 4.1). Syftet med stödet är att bidra till företagarens investeringskostnader för att anlägga en pitch %amp% putt-bana med tillhörande klubbhus. Denna turistaktivitet utgör en ny inkomstkälla för f.d. jordbrukare |
Sektor(er) av ekonomin som berörs | Alla sektorer som är berättigade till stöd till små och medelstora företag | Ja |
Den beviljande myndighetens namn och adress | Provincie Flevoland |
Postbus 55 8200 AB Lelystad Nederland |
Beviljande av stora enskilda stöd | I överensstämmelse med artikel 6 i förordningen | Ja |
Stöd nummer | XS 121/06 |
Medlemsstat | Grekland |
Region | Hela landet |
Namnet på stödordningen eller namnet på det företag som tar emot det enskilda stödet | Initiativet för grekiska teknikcentra (Hellenic Technology Clusters Initiative – HTCI) är godkänt och drivs av det grekiska ministeriet för utvecklingsfrågor. Initiativet avser att inrätta och utveckla konkurrenskraftiga teknikcentra i kunskapsintensiva och exportorienterade sektorer. De teknikcentra som deltar består huvudsakligen av små och medelstora företag |
Rättslig grund | Νόμος 1514/85 όπως τροποποιήθηκε από το Νόμο 2919/01. Ο ρόλος του Ερευνητικού Κέντρου %quot%Αθηνά%quot% περιγράφεται στο Άρθρο 8 του Νόμου 2919/01 και το Προεδρικό Διάταγμα 145/03 όπως τροποποιήθηκαν από το άρθρο 9 του Νόμου 3438/06 και το άρθρο 15 του Νόμου 3460/06 |
Stödordningens beräknade utgifter per år eller totalt belopp som beviljats företaget som enskilt stöd | Årligt totalbelopp | 2006: 1310000 EUR 2007: 1310000 EUR 2008: 652000 EUR |
Totalt stödbelopp De faktiska siffrorna per år kan variera något, men totalbeloppet är fast. | 1514000 EUR |
Högsta tillåtna stödnivå | Den högsta tillåtna stödnivån kommer inte att överstiga 50 % och ligger alltså under det tak för regionalt investeringsstöd som kommissionen fastställt för varje medlemsland samt i förordning (EG) nr 70/2001, senast ändrad genom förordning (EG) nr 364/2004 |
Datum för genomförande | Den första förslagsomgången inleddes i augusti 2006 |
Stödordningens eller det enskilda stödets varaktighet | T.o.m. den 31 december 2008. Rättsliga åtaganden t.o.m. den 31 december 2006 |
Stödets syfte | HTCI-programmet skall stödja initiativ för teknikcentra genom bidrag som ges under en kort period (2006-2008). Bidragen får användas för investeringar (kontorsinredning och ombyggnad, inköp av hårdvara och utrustning, inköp av mjukvara och användarlicenser), konsulttjänster (som inte utgör en permanent eller regelbunden verksamhet och inte ingår i företagets sedvanliga driftskostnader), övriga tjänster och övrig verksamhet (deltagande i mässor och utställningar), samt bidrag som skall täcka kostnader för licenser och andra immateriella rättigheter (patent). Stödets syfte är att hjälpa deltagarna i teknikcentrumen att utvidga sitt verksamhetsområde, upprätta stabila kontaktnät, hantera innovations- och FoTU-frågor, underlätta teknik- och kunskapsdelningen mellan deltagarna, tillvarata personalens begåvningsreserv samt höja de deltagande små och medelstora företagens kompetens |
Sektor(er) av ekonomin som berörs | Mikroelektronik och inbyggda system, förutom företag med verksamhet som avser produktion, utveckling eller marknadsföring av sådana produkter som upptas i bilaga I till fördraget om upprättandet av Europeiska gemenskapen |
Den beviljande myndighetens namn och adress | Υπουργείο Ανάπτυξης, Γενική Γραμματεία Έρευνας και Τεχνολογίας, Ερευνητικό Κέντρο %quot%Αθηνά%quot%, Γ. Αναστασίου 13, GR-11527 Αθήνα (Ministeriet för utveckling, Generalsekretariatet för forskning och teknisk utveckling, Forskningscenter %quot%Aten%quot%, G. Anastasiou 13 – GR-11527 Aten) |
Övriga upplysningar | Stödet är förenligt med förordning (EG) nr 70/2001, senast ändrad genom förordning (EG) nr 364/2004. Stödet avser åtgärd 4.6.3 i programmet för företagens konkurrenskraft som samfinansieras av strukturfonderna |
Stöd nummer | XS 127/06 |
Medlemsstat | Nederländerna |
Region | Alla regioner som kan komma i fråga |
Namnet på stödordningen eller namnet på det företag som tar emot det enskilda stödet | Hållbarhetsundersökningar för forskning och utveckling för projektet Boegbeelden |
Rättslig grund | Kaderwet EZ-subsidies |
Stödordningens beräknade utgifter per år eller totalt belopp som beviljats företaget som enskilt stöd | Stödordning | Årligt totalbelopp | 1 milj. EUR |
Garanterade lån | |
Enskilt stöd | Totalt stödbelopp | |
Garanterade lån | |
Högsta tillåtna stödnivå | Överensstämmer med artikel 4.2-4.6 och artikel 5 i förordningen | För stöd till forskning och utveckling: Följer bestämmelserna om maximala stödnivåer |
Datum för genomförande | Fr.o.m. den 21 juni 2006 |
Stödordningens eller det enskilda stödets varaktighet | 4 år |
Stödets syfte | Stöd till små och medelstora företag | Ja |
Sektor(er) av ekonomin som berörs | Alla sektorer som är berättigade till stöd till små och medelstora företag | Ja |
Den beviljande myndighetens namn och adress | Ministerie van Economische Zaken |
Bezuidenhoutseweg 20 2500 EC Den Haag Nederland |
Beviljande av stora enskilda stöd | I överensstämmelse med artikel 6 i förordningen | Ja |
Stöd nummer | XS 132/06 |
Medlemsstat | Nederländerna |
Region | Provinsen Flevoland |
Namnet på stödordningen eller namnet på det företag som tar emot det enskilda stödet | Maatschap M.T.M.%amp% I. Daniëls-Bisschop |
Rättslig grund | Decentralisatie-convenant Rijk/Flevoland m.b.t. het Leader+ programma Regio Randstad 2000-2006 d.d 11 april 2001.Leader+ overeenkomst tussen de provincie Flevoland en Maatschap M.T.M.%amp% I. Daniëls-Bisschop |
Stödordningens beräknade utgifter per år eller totalt belopp som beviljats företaget som enskilt stöd | Stödordning | Årligt totalbelopp | |
Garanterade lån | |
Enskilt stöd | Totalt stödbelopp | 121446 EUR |
Garanterade lån | |
Högsta tillåtna stödnivå | Överensstämmer med artikel 4.2-4.6 och artikel 5 i förordningen | Ja. Stödnivån är 15 %. Det är förenligt med art. 4.2a i förordning nr 70/2001 |
Datum för genomförande | Beslutet träder i kraft när det har offentliggjorts i EUT |
Stödordningens eller det enskilda stödets varaktighet | T.o.m. den 1 september 2006 |
Stödets syfte | Stöd till små och medelstora företag | Ja. Ett stöd beviljas för investeringar i materiella tillgångar (art. 4.1). Stödets syfte är att bidra till företagets investeringar för att bygga ett pensionat för inkvartering av utländska arbetstagare som tillfälligt utför arbete för ett stort antal jordbrukare i Flevoland |
Sektor(er) av ekonomin som berörs | Alla sektorer som är berättigade till stöd till små och medelstora företag | Ja |
Den beviljande myndighetens namn och adress | Provincie Flevoland |
Postbus 55 8200 AB Lelystad Nederland |
Beviljande av stora enskilda stöd | I överensstämmelse med artikel 6 i förordningen | Ja |
Stöd nummer | XS 146/06 |
Medlemsstat | Nederländerna |
Region | Provincie Zuid-Holland |
Namnet på stödordningen eller namnet på det företag som tar emot det enskilda stödet | Företagets namn: Vastgoed Ontwikkelings Combinatie |
Rättslig grund | Algemene subsidieverordening (Asv), hoofdstuk 6, Milieu, onderdeel regeling stimulering duurzame energie |
Stödordningens beräknade utgifter per år eller totalt belopp som beviljats företaget i form av enskilt stöd | Stödordning | Årligt totalbelopp | |
Garanterade lån | |
Enskilt stöd | Totalt stödbelopp | 370837 EUR (0,9 % av de totala investeringskostnaderna för företaget Vastgoed Ontwikkelings Combinatie) |
Garanterade lån | |
Högsta tillåtna stödnivå | Överensstämmer med artikel 4.2-4.6 och artikel 5 i förordningen | Ja |
Datum för genomförande | Datum för beslutet är den 15 juni 2006. Stödet beviljas först efter anmälan till Europeiska kommissionen |
Stödordningens eller det enskilda stödets varaktighet | Till den 1 september 2007. Sökanden kan ansöka om förskott på högst 80 % av det belopp som kan förväntas. Om denna möjlighet inte utnyttjas utbetalas beloppet 13 veckor efter det att stödet har fastställts |
Stödets syfte | Stöd till små och medelstora företag | Ja |
Projektmål | Syftet är att åstadkomma temperaturreglering i de företagsbyggnader vid Zuidelijke Randweg i Middelharnis som skall byggas, genom värme- och kyllagring i akviferer i golvet kombinerat med värmepumpar. Företagsområdet består av sex skiften som skall anslutas till en central anläggning för produktion av värme och kyla. På grund av obalansen i efterfrågan på värme och kyla (60/40 %) kommer värme att utvinnas från asfalt genom road-energy-system (rörledningar i asfalten) Härigenom kommer utsläppen av koldioxid att minska med 473 ton per år |
Sektor(er) av ekonomin som berörs | Alla sektorer som är berättigade till stöd till små och medelstora företag | Ja |
Den beviljande myndighetens namn och adress | Provincie Zuid Holland |
Zuid-Hollandlaan 1 2596 AW Den Haag Nederland |
Beviljande av stora enskilda stöd | I överensstämmelse med artikel 6 i förordningen | Ja |
--------------------------------------------------
